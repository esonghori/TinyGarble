
module modexp_2N_NN_N1024_CC2097152 ( clk, rst, g_init, e_init, o );
  input [1023:0] g_init;
  input [2047:0] e_init;
  output [1023:0] o;
  input clk, rst;
  wire   first_one, mul_pow, n6, n8, \modmult_1/N2052 , \modmult_1/N2051 ,
         \modmult_1/N2050 , \modmult_1/N2049 , \modmult_1/N2048 ,
         \modmult_1/N2047 , \modmult_1/N2046 , \modmult_1/N2045 ,
         \modmult_1/N2044 , \modmult_1/N2043 , \modmult_1/N2042 ,
         \modmult_1/N2041 , \modmult_1/N2040 , \modmult_1/N2039 ,
         \modmult_1/N2038 , \modmult_1/N2037 , \modmult_1/N2036 ,
         \modmult_1/N2035 , \modmult_1/N2034 , \modmult_1/N2033 ,
         \modmult_1/N2032 , \modmult_1/N2031 , \modmult_1/N2030 ,
         \modmult_1/N2029 , \modmult_1/N2028 , \modmult_1/N2027 ,
         \modmult_1/N2026 , \modmult_1/N2025 , \modmult_1/N2024 ,
         \modmult_1/N2023 , \modmult_1/N2022 , \modmult_1/N2021 ,
         \modmult_1/N2020 , \modmult_1/N2019 , \modmult_1/N2018 ,
         \modmult_1/N2017 , \modmult_1/N2016 , \modmult_1/N2015 ,
         \modmult_1/N2014 , \modmult_1/N2013 , \modmult_1/N2012 ,
         \modmult_1/N2011 , \modmult_1/N2010 , \modmult_1/N2009 ,
         \modmult_1/N2008 , \modmult_1/N2007 , \modmult_1/N2006 ,
         \modmult_1/N2005 , \modmult_1/N2004 , \modmult_1/N2003 ,
         \modmult_1/N2002 , \modmult_1/N2001 , \modmult_1/N2000 ,
         \modmult_1/N1999 , \modmult_1/N1998 , \modmult_1/N1997 ,
         \modmult_1/N1996 , \modmult_1/N1995 , \modmult_1/N1994 ,
         \modmult_1/N1993 , \modmult_1/N1992 , \modmult_1/N1991 ,
         \modmult_1/N1990 , \modmult_1/N1989 , \modmult_1/N1988 ,
         \modmult_1/N1987 , \modmult_1/N1986 , \modmult_1/N1985 ,
         \modmult_1/N1984 , \modmult_1/N1983 , \modmult_1/N1982 ,
         \modmult_1/N1981 , \modmult_1/N1980 , \modmult_1/N1979 ,
         \modmult_1/N1978 , \modmult_1/N1977 , \modmult_1/N1976 ,
         \modmult_1/N1975 , \modmult_1/N1974 , \modmult_1/N1973 ,
         \modmult_1/N1972 , \modmult_1/N1971 , \modmult_1/N1970 ,
         \modmult_1/N1969 , \modmult_1/N1968 , \modmult_1/N1967 ,
         \modmult_1/N1966 , \modmult_1/N1965 , \modmult_1/N1964 ,
         \modmult_1/N1963 , \modmult_1/N1962 , \modmult_1/N1961 ,
         \modmult_1/N1960 , \modmult_1/N1959 , \modmult_1/N1958 ,
         \modmult_1/N1957 , \modmult_1/N1956 , \modmult_1/N1955 ,
         \modmult_1/N1954 , \modmult_1/N1953 , \modmult_1/N1952 ,
         \modmult_1/N1951 , \modmult_1/N1950 , \modmult_1/N1949 ,
         \modmult_1/N1948 , \modmult_1/N1947 , \modmult_1/N1946 ,
         \modmult_1/N1945 , \modmult_1/N1944 , \modmult_1/N1943 ,
         \modmult_1/N1942 , \modmult_1/N1941 , \modmult_1/N1940 ,
         \modmult_1/N1939 , \modmult_1/N1938 , \modmult_1/N1937 ,
         \modmult_1/N1936 , \modmult_1/N1935 , \modmult_1/N1934 ,
         \modmult_1/N1933 , \modmult_1/N1932 , \modmult_1/N1931 ,
         \modmult_1/N1930 , \modmult_1/N1929 , \modmult_1/N1928 ,
         \modmult_1/N1927 , \modmult_1/N1926 , \modmult_1/N1925 ,
         \modmult_1/N1924 , \modmult_1/N1923 , \modmult_1/N1922 ,
         \modmult_1/N1921 , \modmult_1/N1920 , \modmult_1/N1919 ,
         \modmult_1/N1918 , \modmult_1/N1917 , \modmult_1/N1916 ,
         \modmult_1/N1915 , \modmult_1/N1914 , \modmult_1/N1913 ,
         \modmult_1/N1912 , \modmult_1/N1911 , \modmult_1/N1910 ,
         \modmult_1/N1909 , \modmult_1/N1908 , \modmult_1/N1907 ,
         \modmult_1/N1906 , \modmult_1/N1905 , \modmult_1/N1904 ,
         \modmult_1/N1903 , \modmult_1/N1902 , \modmult_1/N1901 ,
         \modmult_1/N1900 , \modmult_1/N1899 , \modmult_1/N1898 ,
         \modmult_1/N1897 , \modmult_1/N1896 , \modmult_1/N1895 ,
         \modmult_1/N1894 , \modmult_1/N1893 , \modmult_1/N1892 ,
         \modmult_1/N1891 , \modmult_1/N1890 , \modmult_1/N1889 ,
         \modmult_1/N1888 , \modmult_1/N1887 , \modmult_1/N1886 ,
         \modmult_1/N1885 , \modmult_1/N1884 , \modmult_1/N1883 ,
         \modmult_1/N1882 , \modmult_1/N1881 , \modmult_1/N1880 ,
         \modmult_1/N1879 , \modmult_1/N1878 , \modmult_1/N1877 ,
         \modmult_1/N1876 , \modmult_1/N1875 , \modmult_1/N1874 ,
         \modmult_1/N1873 , \modmult_1/N1872 , \modmult_1/N1871 ,
         \modmult_1/N1870 , \modmult_1/N1869 , \modmult_1/N1868 ,
         \modmult_1/N1867 , \modmult_1/N1866 , \modmult_1/N1865 ,
         \modmult_1/N1864 , \modmult_1/N1863 , \modmult_1/N1862 ,
         \modmult_1/N1861 , \modmult_1/N1860 , \modmult_1/N1859 ,
         \modmult_1/N1858 , \modmult_1/N1857 , \modmult_1/N1856 ,
         \modmult_1/N1855 , \modmult_1/N1854 , \modmult_1/N1853 ,
         \modmult_1/N1852 , \modmult_1/N1851 , \modmult_1/N1850 ,
         \modmult_1/N1849 , \modmult_1/N1848 , \modmult_1/N1847 ,
         \modmult_1/N1846 , \modmult_1/N1845 , \modmult_1/N1844 ,
         \modmult_1/N1843 , \modmult_1/N1842 , \modmult_1/N1841 ,
         \modmult_1/N1840 , \modmult_1/N1839 , \modmult_1/N1838 ,
         \modmult_1/N1837 , \modmult_1/N1836 , \modmult_1/N1835 ,
         \modmult_1/N1834 , \modmult_1/N1833 , \modmult_1/N1832 ,
         \modmult_1/N1831 , \modmult_1/N1830 , \modmult_1/N1829 ,
         \modmult_1/N1828 , \modmult_1/N1827 , \modmult_1/N1826 ,
         \modmult_1/N1825 , \modmult_1/N1824 , \modmult_1/N1823 ,
         \modmult_1/N1822 , \modmult_1/N1821 , \modmult_1/N1820 ,
         \modmult_1/N1819 , \modmult_1/N1818 , \modmult_1/N1817 ,
         \modmult_1/N1816 , \modmult_1/N1815 , \modmult_1/N1814 ,
         \modmult_1/N1813 , \modmult_1/N1812 , \modmult_1/N1811 ,
         \modmult_1/N1810 , \modmult_1/N1809 , \modmult_1/N1808 ,
         \modmult_1/N1807 , \modmult_1/N1806 , \modmult_1/N1805 ,
         \modmult_1/N1804 , \modmult_1/N1803 , \modmult_1/N1802 ,
         \modmult_1/N1801 , \modmult_1/N1800 , \modmult_1/N1799 ,
         \modmult_1/N1798 , \modmult_1/N1797 , \modmult_1/N1796 ,
         \modmult_1/N1795 , \modmult_1/N1794 , \modmult_1/N1793 ,
         \modmult_1/N1792 , \modmult_1/N1791 , \modmult_1/N1790 ,
         \modmult_1/N1789 , \modmult_1/N1788 , \modmult_1/N1787 ,
         \modmult_1/N1786 , \modmult_1/N1785 , \modmult_1/N1784 ,
         \modmult_1/N1783 , \modmult_1/N1782 , \modmult_1/N1781 ,
         \modmult_1/N1780 , \modmult_1/N1779 , \modmult_1/N1778 ,
         \modmult_1/N1777 , \modmult_1/N1776 , \modmult_1/N1775 ,
         \modmult_1/N1774 , \modmult_1/N1773 , \modmult_1/N1772 ,
         \modmult_1/N1771 , \modmult_1/N1770 , \modmult_1/N1769 ,
         \modmult_1/N1768 , \modmult_1/N1767 , \modmult_1/N1766 ,
         \modmult_1/N1765 , \modmult_1/N1764 , \modmult_1/N1763 ,
         \modmult_1/N1762 , \modmult_1/N1761 , \modmult_1/N1760 ,
         \modmult_1/N1759 , \modmult_1/N1758 , \modmult_1/N1757 ,
         \modmult_1/N1756 , \modmult_1/N1755 , \modmult_1/N1754 ,
         \modmult_1/N1753 , \modmult_1/N1752 , \modmult_1/N1751 ,
         \modmult_1/N1750 , \modmult_1/N1749 , \modmult_1/N1748 ,
         \modmult_1/N1747 , \modmult_1/N1746 , \modmult_1/N1745 ,
         \modmult_1/N1744 , \modmult_1/N1743 , \modmult_1/N1742 ,
         \modmult_1/N1741 , \modmult_1/N1740 , \modmult_1/N1739 ,
         \modmult_1/N1738 , \modmult_1/N1737 , \modmult_1/N1736 ,
         \modmult_1/N1735 , \modmult_1/N1734 , \modmult_1/N1733 ,
         \modmult_1/N1732 , \modmult_1/N1731 , \modmult_1/N1730 ,
         \modmult_1/N1729 , \modmult_1/N1728 , \modmult_1/N1727 ,
         \modmult_1/N1726 , \modmult_1/N1725 , \modmult_1/N1724 ,
         \modmult_1/N1723 , \modmult_1/N1722 , \modmult_1/N1721 ,
         \modmult_1/N1720 , \modmult_1/N1719 , \modmult_1/N1718 ,
         \modmult_1/N1717 , \modmult_1/N1716 , \modmult_1/N1715 ,
         \modmult_1/N1714 , \modmult_1/N1713 , \modmult_1/N1712 ,
         \modmult_1/N1711 , \modmult_1/N1710 , \modmult_1/N1709 ,
         \modmult_1/N1708 , \modmult_1/N1707 , \modmult_1/N1706 ,
         \modmult_1/N1705 , \modmult_1/N1704 , \modmult_1/N1703 ,
         \modmult_1/N1702 , \modmult_1/N1701 , \modmult_1/N1700 ,
         \modmult_1/N1699 , \modmult_1/N1698 , \modmult_1/N1697 ,
         \modmult_1/N1696 , \modmult_1/N1695 , \modmult_1/N1694 ,
         \modmult_1/N1693 , \modmult_1/N1692 , \modmult_1/N1691 ,
         \modmult_1/N1690 , \modmult_1/N1689 , \modmult_1/N1688 ,
         \modmult_1/N1687 , \modmult_1/N1686 , \modmult_1/N1685 ,
         \modmult_1/N1684 , \modmult_1/N1683 , \modmult_1/N1682 ,
         \modmult_1/N1681 , \modmult_1/N1680 , \modmult_1/N1679 ,
         \modmult_1/N1678 , \modmult_1/N1677 , \modmult_1/N1676 ,
         \modmult_1/N1675 , \modmult_1/N1674 , \modmult_1/N1673 ,
         \modmult_1/N1672 , \modmult_1/N1671 , \modmult_1/N1670 ,
         \modmult_1/N1669 , \modmult_1/N1668 , \modmult_1/N1667 ,
         \modmult_1/N1666 , \modmult_1/N1665 , \modmult_1/N1664 ,
         \modmult_1/N1663 , \modmult_1/N1662 , \modmult_1/N1661 ,
         \modmult_1/N1660 , \modmult_1/N1659 , \modmult_1/N1658 ,
         \modmult_1/N1657 , \modmult_1/N1656 , \modmult_1/N1655 ,
         \modmult_1/N1654 , \modmult_1/N1653 , \modmult_1/N1652 ,
         \modmult_1/N1651 , \modmult_1/N1650 , \modmult_1/N1649 ,
         \modmult_1/N1648 , \modmult_1/N1647 , \modmult_1/N1646 ,
         \modmult_1/N1645 , \modmult_1/N1644 , \modmult_1/N1643 ,
         \modmult_1/N1642 , \modmult_1/N1641 , \modmult_1/N1640 ,
         \modmult_1/N1639 , \modmult_1/N1638 , \modmult_1/N1637 ,
         \modmult_1/N1636 , \modmult_1/N1635 , \modmult_1/N1634 ,
         \modmult_1/N1633 , \modmult_1/N1632 , \modmult_1/N1631 ,
         \modmult_1/N1630 , \modmult_1/N1629 , \modmult_1/N1628 ,
         \modmult_1/N1627 , \modmult_1/N1626 , \modmult_1/N1625 ,
         \modmult_1/N1624 , \modmult_1/N1623 , \modmult_1/N1622 ,
         \modmult_1/N1621 , \modmult_1/N1620 , \modmult_1/N1619 ,
         \modmult_1/N1618 , \modmult_1/N1617 , \modmult_1/N1616 ,
         \modmult_1/N1615 , \modmult_1/N1614 , \modmult_1/N1613 ,
         \modmult_1/N1612 , \modmult_1/N1611 , \modmult_1/N1610 ,
         \modmult_1/N1609 , \modmult_1/N1608 , \modmult_1/N1607 ,
         \modmult_1/N1606 , \modmult_1/N1605 , \modmult_1/N1604 ,
         \modmult_1/N1603 , \modmult_1/N1602 , \modmult_1/N1601 ,
         \modmult_1/N1600 , \modmult_1/N1599 , \modmult_1/N1598 ,
         \modmult_1/N1597 , \modmult_1/N1596 , \modmult_1/N1595 ,
         \modmult_1/N1594 , \modmult_1/N1593 , \modmult_1/N1592 ,
         \modmult_1/N1591 , \modmult_1/N1590 , \modmult_1/N1589 ,
         \modmult_1/N1588 , \modmult_1/N1587 , \modmult_1/N1586 ,
         \modmult_1/N1585 , \modmult_1/N1584 , \modmult_1/N1583 ,
         \modmult_1/N1582 , \modmult_1/N1581 , \modmult_1/N1580 ,
         \modmult_1/N1579 , \modmult_1/N1578 , \modmult_1/N1577 ,
         \modmult_1/N1576 , \modmult_1/N1575 , \modmult_1/N1574 ,
         \modmult_1/N1573 , \modmult_1/N1572 , \modmult_1/N1571 ,
         \modmult_1/N1570 , \modmult_1/N1569 , \modmult_1/N1568 ,
         \modmult_1/N1567 , \modmult_1/N1566 , \modmult_1/N1565 ,
         \modmult_1/N1564 , \modmult_1/N1563 , \modmult_1/N1562 ,
         \modmult_1/N1561 , \modmult_1/N1560 , \modmult_1/N1559 ,
         \modmult_1/N1558 , \modmult_1/N1557 , \modmult_1/N1556 ,
         \modmult_1/N1555 , \modmult_1/N1554 , \modmult_1/N1553 ,
         \modmult_1/N1552 , \modmult_1/N1551 , \modmult_1/N1550 ,
         \modmult_1/N1549 , \modmult_1/N1548 , \modmult_1/N1547 ,
         \modmult_1/N1546 , \modmult_1/N1545 , \modmult_1/N1544 ,
         \modmult_1/N1543 , \modmult_1/N1542 , \modmult_1/N1541 ,
         \modmult_1/N1540 , \modmult_1/N1539 , \modmult_1/N1538 ,
         \modmult_1/N1537 , \modmult_1/N1536 , \modmult_1/N1535 ,
         \modmult_1/N1534 , \modmult_1/N1533 , \modmult_1/N1532 ,
         \modmult_1/N1531 , \modmult_1/N1530 , \modmult_1/N1529 ,
         \modmult_1/N1528 , \modmult_1/N1527 , \modmult_1/N1526 ,
         \modmult_1/N1525 , \modmult_1/N1524 , \modmult_1/N1523 ,
         \modmult_1/N1522 , \modmult_1/N1521 , \modmult_1/N1520 ,
         \modmult_1/N1519 , \modmult_1/N1518 , \modmult_1/N1517 ,
         \modmult_1/N1516 , \modmult_1/N1515 , \modmult_1/N1514 ,
         \modmult_1/N1513 , \modmult_1/N1512 , \modmult_1/N1511 ,
         \modmult_1/N1510 , \modmult_1/N1509 , \modmult_1/N1508 ,
         \modmult_1/N1507 , \modmult_1/N1506 , \modmult_1/N1505 ,
         \modmult_1/N1504 , \modmult_1/N1503 , \modmult_1/N1502 ,
         \modmult_1/N1501 , \modmult_1/N1500 , \modmult_1/N1499 ,
         \modmult_1/N1498 , \modmult_1/N1497 , \modmult_1/N1496 ,
         \modmult_1/N1495 , \modmult_1/N1494 , \modmult_1/N1493 ,
         \modmult_1/N1492 , \modmult_1/N1491 , \modmult_1/N1490 ,
         \modmult_1/N1489 , \modmult_1/N1488 , \modmult_1/N1487 ,
         \modmult_1/N1486 , \modmult_1/N1485 , \modmult_1/N1484 ,
         \modmult_1/N1483 , \modmult_1/N1482 , \modmult_1/N1481 ,
         \modmult_1/N1480 , \modmult_1/N1479 , \modmult_1/N1478 ,
         \modmult_1/N1477 , \modmult_1/N1476 , \modmult_1/N1475 ,
         \modmult_1/N1474 , \modmult_1/N1473 , \modmult_1/N1472 ,
         \modmult_1/N1471 , \modmult_1/N1470 , \modmult_1/N1469 ,
         \modmult_1/N1468 , \modmult_1/N1467 , \modmult_1/N1466 ,
         \modmult_1/N1465 , \modmult_1/N1464 , \modmult_1/N1463 ,
         \modmult_1/N1462 , \modmult_1/N1461 , \modmult_1/N1460 ,
         \modmult_1/N1459 , \modmult_1/N1458 , \modmult_1/N1457 ,
         \modmult_1/N1456 , \modmult_1/N1455 , \modmult_1/N1454 ,
         \modmult_1/N1453 , \modmult_1/N1452 , \modmult_1/N1451 ,
         \modmult_1/N1450 , \modmult_1/N1449 , \modmult_1/N1448 ,
         \modmult_1/N1447 , \modmult_1/N1446 , \modmult_1/N1445 ,
         \modmult_1/N1444 , \modmult_1/N1443 , \modmult_1/N1442 ,
         \modmult_1/N1441 , \modmult_1/N1440 , \modmult_1/N1439 ,
         \modmult_1/N1438 , \modmult_1/N1437 , \modmult_1/N1436 ,
         \modmult_1/N1435 , \modmult_1/N1434 , \modmult_1/N1433 ,
         \modmult_1/N1432 , \modmult_1/N1431 , \modmult_1/N1430 ,
         \modmult_1/N1429 , \modmult_1/N1428 , \modmult_1/N1427 ,
         \modmult_1/N1426 , \modmult_1/N1425 , \modmult_1/N1424 ,
         \modmult_1/N1423 , \modmult_1/N1422 , \modmult_1/N1421 ,
         \modmult_1/N1420 , \modmult_1/N1419 , \modmult_1/N1418 ,
         \modmult_1/N1417 , \modmult_1/N1416 , \modmult_1/N1415 ,
         \modmult_1/N1414 , \modmult_1/N1413 , \modmult_1/N1412 ,
         \modmult_1/N1411 , \modmult_1/N1410 , \modmult_1/N1409 ,
         \modmult_1/N1408 , \modmult_1/N1407 , \modmult_1/N1406 ,
         \modmult_1/N1405 , \modmult_1/N1404 , \modmult_1/N1403 ,
         \modmult_1/N1402 , \modmult_1/N1401 , \modmult_1/N1400 ,
         \modmult_1/N1399 , \modmult_1/N1398 , \modmult_1/N1397 ,
         \modmult_1/N1396 , \modmult_1/N1395 , \modmult_1/N1394 ,
         \modmult_1/N1393 , \modmult_1/N1392 , \modmult_1/N1391 ,
         \modmult_1/N1390 , \modmult_1/N1389 , \modmult_1/N1388 ,
         \modmult_1/N1387 , \modmult_1/N1386 , \modmult_1/N1385 ,
         \modmult_1/N1384 , \modmult_1/N1383 , \modmult_1/N1382 ,
         \modmult_1/N1381 , \modmult_1/N1380 , \modmult_1/N1379 ,
         \modmult_1/N1378 , \modmult_1/N1377 , \modmult_1/N1376 ,
         \modmult_1/N1375 , \modmult_1/N1374 , \modmult_1/N1373 ,
         \modmult_1/N1372 , \modmult_1/N1371 , \modmult_1/N1370 ,
         \modmult_1/N1369 , \modmult_1/N1368 , \modmult_1/N1367 ,
         \modmult_1/N1366 , \modmult_1/N1365 , \modmult_1/N1364 ,
         \modmult_1/N1363 , \modmult_1/N1362 , \modmult_1/N1361 ,
         \modmult_1/N1360 , \modmult_1/N1359 , \modmult_1/N1358 ,
         \modmult_1/N1357 , \modmult_1/N1356 , \modmult_1/N1355 ,
         \modmult_1/N1354 , \modmult_1/N1353 , \modmult_1/N1352 ,
         \modmult_1/N1351 , \modmult_1/N1350 , \modmult_1/N1349 ,
         \modmult_1/N1348 , \modmult_1/N1347 , \modmult_1/N1346 ,
         \modmult_1/N1345 , \modmult_1/N1344 , \modmult_1/N1343 ,
         \modmult_1/N1342 , \modmult_1/N1341 , \modmult_1/N1340 ,
         \modmult_1/N1339 , \modmult_1/N1338 , \modmult_1/N1337 ,
         \modmult_1/N1336 , \modmult_1/N1335 , \modmult_1/N1334 ,
         \modmult_1/N1333 , \modmult_1/N1332 , \modmult_1/N1331 ,
         \modmult_1/N1330 , \modmult_1/N1329 , \modmult_1/N1328 ,
         \modmult_1/N1327 , \modmult_1/N1326 , \modmult_1/N1325 ,
         \modmult_1/N1324 , \modmult_1/N1323 , \modmult_1/N1322 ,
         \modmult_1/N1321 , \modmult_1/N1320 , \modmult_1/N1319 ,
         \modmult_1/N1318 , \modmult_1/N1317 , \modmult_1/N1316 ,
         \modmult_1/N1315 , \modmult_1/N1314 , \modmult_1/N1313 ,
         \modmult_1/N1312 , \modmult_1/N1311 , \modmult_1/N1310 ,
         \modmult_1/N1309 , \modmult_1/N1308 , \modmult_1/N1307 ,
         \modmult_1/N1306 , \modmult_1/N1305 , \modmult_1/N1304 ,
         \modmult_1/N1303 , \modmult_1/N1302 , \modmult_1/N1301 ,
         \modmult_1/N1300 , \modmult_1/N1299 , \modmult_1/N1298 ,
         \modmult_1/N1297 , \modmult_1/N1296 , \modmult_1/N1295 ,
         \modmult_1/N1294 , \modmult_1/N1293 , \modmult_1/N1292 ,
         \modmult_1/N1291 , \modmult_1/N1290 , \modmult_1/N1289 ,
         \modmult_1/N1288 , \modmult_1/N1287 , \modmult_1/N1286 ,
         \modmult_1/N1285 , \modmult_1/N1284 , \modmult_1/N1283 ,
         \modmult_1/N1282 , \modmult_1/N1281 , \modmult_1/N1280 ,
         \modmult_1/N1279 , \modmult_1/N1278 , \modmult_1/N1277 ,
         \modmult_1/N1276 , \modmult_1/N1275 , \modmult_1/N1274 ,
         \modmult_1/N1273 , \modmult_1/N1272 , \modmult_1/N1271 ,
         \modmult_1/N1270 , \modmult_1/N1269 , \modmult_1/N1268 ,
         \modmult_1/N1267 , \modmult_1/N1266 , \modmult_1/N1265 ,
         \modmult_1/N1264 , \modmult_1/N1263 , \modmult_1/N1262 ,
         \modmult_1/N1261 , \modmult_1/N1260 , \modmult_1/N1259 ,
         \modmult_1/N1258 , \modmult_1/N1257 , \modmult_1/N1256 ,
         \modmult_1/N1255 , \modmult_1/N1254 , \modmult_1/N1253 ,
         \modmult_1/N1252 , \modmult_1/N1251 , \modmult_1/N1250 ,
         \modmult_1/N1249 , \modmult_1/N1248 , \modmult_1/N1247 ,
         \modmult_1/N1246 , \modmult_1/N1245 , \modmult_1/N1244 ,
         \modmult_1/N1243 , \modmult_1/N1242 , \modmult_1/N1241 ,
         \modmult_1/N1240 , \modmult_1/N1239 , \modmult_1/N1238 ,
         \modmult_1/N1237 , \modmult_1/N1236 , \modmult_1/N1235 ,
         \modmult_1/N1234 , \modmult_1/N1233 , \modmult_1/N1232 ,
         \modmult_1/N1231 , \modmult_1/N1230 , \modmult_1/N1229 ,
         \modmult_1/N1228 , \modmult_1/N1227 , \modmult_1/N1226 ,
         \modmult_1/N1225 , \modmult_1/N1224 , \modmult_1/N1223 ,
         \modmult_1/N1222 , \modmult_1/N1221 , \modmult_1/N1220 ,
         \modmult_1/N1219 , \modmult_1/N1218 , \modmult_1/N1217 ,
         \modmult_1/N1216 , \modmult_1/N1215 , \modmult_1/N1214 ,
         \modmult_1/N1213 , \modmult_1/N1212 , \modmult_1/N1211 ,
         \modmult_1/N1210 , \modmult_1/N1209 , \modmult_1/N1208 ,
         \modmult_1/N1207 , \modmult_1/N1206 , \modmult_1/N1205 ,
         \modmult_1/N1204 , \modmult_1/N1203 , \modmult_1/N1202 ,
         \modmult_1/N1201 , \modmult_1/N1200 , \modmult_1/N1199 ,
         \modmult_1/N1198 , \modmult_1/N1197 , \modmult_1/N1196 ,
         \modmult_1/N1195 , \modmult_1/N1194 , \modmult_1/N1193 ,
         \modmult_1/N1192 , \modmult_1/N1191 , \modmult_1/N1190 ,
         \modmult_1/N1189 , \modmult_1/N1188 , \modmult_1/N1187 ,
         \modmult_1/N1186 , \modmult_1/N1185 , \modmult_1/N1184 ,
         \modmult_1/N1183 , \modmult_1/N1182 , \modmult_1/N1181 ,
         \modmult_1/N1180 , \modmult_1/N1179 , \modmult_1/N1178 ,
         \modmult_1/N1177 , \modmult_1/N1176 , \modmult_1/N1175 ,
         \modmult_1/N1174 , \modmult_1/N1173 , \modmult_1/N1172 ,
         \modmult_1/N1171 , \modmult_1/N1170 , \modmult_1/N1169 ,
         \modmult_1/N1168 , \modmult_1/N1167 , \modmult_1/N1166 ,
         \modmult_1/N1165 , \modmult_1/N1164 , \modmult_1/N1163 ,
         \modmult_1/N1162 , \modmult_1/N1161 , \modmult_1/N1160 ,
         \modmult_1/N1159 , \modmult_1/N1158 , \modmult_1/N1157 ,
         \modmult_1/N1156 , \modmult_1/N1155 , \modmult_1/N1154 ,
         \modmult_1/N1153 , \modmult_1/N1152 , \modmult_1/N1151 ,
         \modmult_1/N1150 , \modmult_1/N1149 , \modmult_1/N1148 ,
         \modmult_1/N1147 , \modmult_1/N1146 , \modmult_1/N1145 ,
         \modmult_1/N1144 , \modmult_1/N1143 , \modmult_1/N1142 ,
         \modmult_1/N1141 , \modmult_1/N1140 , \modmult_1/N1139 ,
         \modmult_1/N1138 , \modmult_1/N1137 , \modmult_1/N1136 ,
         \modmult_1/N1135 , \modmult_1/N1134 , \modmult_1/N1133 ,
         \modmult_1/N1132 , \modmult_1/N1131 , \modmult_1/N1130 ,
         \modmult_1/N1129 , \modmult_1/N1128 , \modmult_1/N1127 ,
         \modmult_1/N1126 , \modmult_1/N1125 , \modmult_1/N1124 ,
         \modmult_1/N1123 , \modmult_1/N1122 , \modmult_1/N1121 ,
         \modmult_1/N1120 , \modmult_1/N1119 , \modmult_1/N1118 ,
         \modmult_1/N1117 , \modmult_1/N1116 , \modmult_1/N1115 ,
         \modmult_1/N1114 , \modmult_1/N1113 , \modmult_1/N1112 ,
         \modmult_1/N1111 , \modmult_1/N1110 , \modmult_1/N1109 ,
         \modmult_1/N1108 , \modmult_1/N1107 , \modmult_1/N1106 ,
         \modmult_1/N1105 , \modmult_1/N1104 , \modmult_1/N1103 ,
         \modmult_1/N1102 , \modmult_1/N1101 , \modmult_1/N1100 ,
         \modmult_1/N1099 , \modmult_1/N1098 , \modmult_1/N1097 ,
         \modmult_1/N1096 , \modmult_1/N1095 , \modmult_1/N1094 ,
         \modmult_1/N1093 , \modmult_1/N1092 , \modmult_1/N1091 ,
         \modmult_1/N1090 , \modmult_1/N1089 , \modmult_1/N1088 ,
         \modmult_1/N1087 , \modmult_1/N1086 , \modmult_1/N1085 ,
         \modmult_1/N1084 , \modmult_1/N1083 , \modmult_1/N1082 ,
         \modmult_1/N1081 , \modmult_1/N1080 , \modmult_1/N1079 ,
         \modmult_1/N1078 , \modmult_1/N1077 , \modmult_1/N1076 ,
         \modmult_1/N1075 , \modmult_1/N1074 , \modmult_1/N1073 ,
         \modmult_1/N1072 , \modmult_1/N1071 , \modmult_1/N1070 ,
         \modmult_1/N1069 , \modmult_1/N1068 , \modmult_1/N1067 ,
         \modmult_1/N1066 , \modmult_1/N1065 , \modmult_1/N1064 ,
         \modmult_1/N1063 , \modmult_1/N1062 , \modmult_1/N1061 ,
         \modmult_1/N1060 , \modmult_1/N1059 , \modmult_1/N1058 ,
         \modmult_1/N1057 , \modmult_1/N1056 , \modmult_1/N1055 ,
         \modmult_1/N1054 , \modmult_1/N1053 , \modmult_1/N1052 ,
         \modmult_1/N1051 , \modmult_1/N1050 , \modmult_1/N1049 ,
         \modmult_1/N1048 , \modmult_1/N1047 , \modmult_1/N1046 ,
         \modmult_1/N1045 , \modmult_1/N1044 , \modmult_1/N1043 ,
         \modmult_1/N1042 , \modmult_1/N1041 , \modmult_1/N1040 ,
         \modmult_1/N1039 , \modmult_1/N1038 , \modmult_1/N1037 ,
         \modmult_1/N1036 , \modmult_1/N1035 , \modmult_1/N1034 ,
         \modmult_1/N1033 , \modmult_1/N1032 , \modmult_1/N1031 ,
         \modmult_1/N1030 , \modmult_1/N1029 , \modmult_1/N1027 ,
         \modmult_1/N1026 , \modmult_1/N1025 , \modmult_1/N1024 ,
         \modmult_1/N1023 , \modmult_1/N1022 , \modmult_1/N1021 ,
         \modmult_1/N1020 , \modmult_1/N1019 , \modmult_1/N1018 ,
         \modmult_1/N1017 , \modmult_1/N1016 , \modmult_1/N1015 ,
         \modmult_1/N1014 , \modmult_1/N1013 , \modmult_1/N1012 ,
         \modmult_1/N1011 , \modmult_1/N1010 , \modmult_1/N1009 ,
         \modmult_1/N1008 , \modmult_1/N1007 , \modmult_1/N1006 ,
         \modmult_1/N1005 , \modmult_1/N1004 , \modmult_1/N1003 ,
         \modmult_1/N1002 , \modmult_1/N1001 , \modmult_1/N1000 ,
         \modmult_1/N999 , \modmult_1/N998 , \modmult_1/N997 ,
         \modmult_1/N996 , \modmult_1/N995 , \modmult_1/N994 ,
         \modmult_1/N993 , \modmult_1/N992 , \modmult_1/N991 ,
         \modmult_1/N990 , \modmult_1/N989 , \modmult_1/N988 ,
         \modmult_1/N987 , \modmult_1/N986 , \modmult_1/N985 ,
         \modmult_1/N984 , \modmult_1/N983 , \modmult_1/N982 ,
         \modmult_1/N981 , \modmult_1/N980 , \modmult_1/N979 ,
         \modmult_1/N978 , \modmult_1/N977 , \modmult_1/N976 ,
         \modmult_1/N975 , \modmult_1/N974 , \modmult_1/N973 ,
         \modmult_1/N972 , \modmult_1/N971 , \modmult_1/N970 ,
         \modmult_1/N969 , \modmult_1/N968 , \modmult_1/N967 ,
         \modmult_1/N966 , \modmult_1/N965 , \modmult_1/N964 ,
         \modmult_1/N963 , \modmult_1/N962 , \modmult_1/N961 ,
         \modmult_1/N960 , \modmult_1/N959 , \modmult_1/N958 ,
         \modmult_1/N957 , \modmult_1/N956 , \modmult_1/N955 ,
         \modmult_1/N954 , \modmult_1/N953 , \modmult_1/N952 ,
         \modmult_1/N951 , \modmult_1/N950 , \modmult_1/N949 ,
         \modmult_1/N948 , \modmult_1/N947 , \modmult_1/N946 ,
         \modmult_1/N945 , \modmult_1/N944 , \modmult_1/N943 ,
         \modmult_1/N942 , \modmult_1/N941 , \modmult_1/N940 ,
         \modmult_1/N939 , \modmult_1/N938 , \modmult_1/N937 ,
         \modmult_1/N936 , \modmult_1/N935 , \modmult_1/N934 ,
         \modmult_1/N933 , \modmult_1/N932 , \modmult_1/N931 ,
         \modmult_1/N930 , \modmult_1/N929 , \modmult_1/N928 ,
         \modmult_1/N927 , \modmult_1/N926 , \modmult_1/N925 ,
         \modmult_1/N924 , \modmult_1/N923 , \modmult_1/N922 ,
         \modmult_1/N921 , \modmult_1/N920 , \modmult_1/N919 ,
         \modmult_1/N918 , \modmult_1/N917 , \modmult_1/N916 ,
         \modmult_1/N915 , \modmult_1/N914 , \modmult_1/N913 ,
         \modmult_1/N912 , \modmult_1/N911 , \modmult_1/N910 ,
         \modmult_1/N909 , \modmult_1/N908 , \modmult_1/N907 ,
         \modmult_1/N906 , \modmult_1/N905 , \modmult_1/N904 ,
         \modmult_1/N903 , \modmult_1/N902 , \modmult_1/N901 ,
         \modmult_1/N900 , \modmult_1/N899 , \modmult_1/N898 ,
         \modmult_1/N897 , \modmult_1/N896 , \modmult_1/N895 ,
         \modmult_1/N894 , \modmult_1/N893 , \modmult_1/N892 ,
         \modmult_1/N891 , \modmult_1/N890 , \modmult_1/N889 ,
         \modmult_1/N888 , \modmult_1/N887 , \modmult_1/N886 ,
         \modmult_1/N885 , \modmult_1/N884 , \modmult_1/N883 ,
         \modmult_1/N882 , \modmult_1/N881 , \modmult_1/N880 ,
         \modmult_1/N879 , \modmult_1/N878 , \modmult_1/N877 ,
         \modmult_1/N876 , \modmult_1/N875 , \modmult_1/N874 ,
         \modmult_1/N873 , \modmult_1/N872 , \modmult_1/N871 ,
         \modmult_1/N870 , \modmult_1/N869 , \modmult_1/N868 ,
         \modmult_1/N867 , \modmult_1/N866 , \modmult_1/N865 ,
         \modmult_1/N864 , \modmult_1/N863 , \modmult_1/N862 ,
         \modmult_1/N861 , \modmult_1/N860 , \modmult_1/N859 ,
         \modmult_1/N858 , \modmult_1/N857 , \modmult_1/N856 ,
         \modmult_1/N855 , \modmult_1/N854 , \modmult_1/N853 ,
         \modmult_1/N852 , \modmult_1/N851 , \modmult_1/N850 ,
         \modmult_1/N849 , \modmult_1/N848 , \modmult_1/N847 ,
         \modmult_1/N846 , \modmult_1/N845 , \modmult_1/N844 ,
         \modmult_1/N843 , \modmult_1/N842 , \modmult_1/N841 ,
         \modmult_1/N840 , \modmult_1/N839 , \modmult_1/N838 ,
         \modmult_1/N837 , \modmult_1/N836 , \modmult_1/N835 ,
         \modmult_1/N834 , \modmult_1/N833 , \modmult_1/N832 ,
         \modmult_1/N831 , \modmult_1/N830 , \modmult_1/N829 ,
         \modmult_1/N828 , \modmult_1/N827 , \modmult_1/N826 ,
         \modmult_1/N825 , \modmult_1/N824 , \modmult_1/N823 ,
         \modmult_1/N822 , \modmult_1/N821 , \modmult_1/N820 ,
         \modmult_1/N819 , \modmult_1/N818 , \modmult_1/N817 ,
         \modmult_1/N816 , \modmult_1/N815 , \modmult_1/N814 ,
         \modmult_1/N813 , \modmult_1/N812 , \modmult_1/N811 ,
         \modmult_1/N810 , \modmult_1/N809 , \modmult_1/N808 ,
         \modmult_1/N807 , \modmult_1/N806 , \modmult_1/N805 ,
         \modmult_1/N804 , \modmult_1/N803 , \modmult_1/N802 ,
         \modmult_1/N801 , \modmult_1/N800 , \modmult_1/N799 ,
         \modmult_1/N798 , \modmult_1/N797 , \modmult_1/N796 ,
         \modmult_1/N795 , \modmult_1/N794 , \modmult_1/N793 ,
         \modmult_1/N792 , \modmult_1/N791 , \modmult_1/N790 ,
         \modmult_1/N789 , \modmult_1/N788 , \modmult_1/N787 ,
         \modmult_1/N786 , \modmult_1/N785 , \modmult_1/N784 ,
         \modmult_1/N783 , \modmult_1/N782 , \modmult_1/N781 ,
         \modmult_1/N780 , \modmult_1/N779 , \modmult_1/N778 ,
         \modmult_1/N777 , \modmult_1/N776 , \modmult_1/N775 ,
         \modmult_1/N774 , \modmult_1/N773 , \modmult_1/N772 ,
         \modmult_1/N771 , \modmult_1/N770 , \modmult_1/N769 ,
         \modmult_1/N768 , \modmult_1/N767 , \modmult_1/N766 ,
         \modmult_1/N765 , \modmult_1/N764 , \modmult_1/N763 ,
         \modmult_1/N762 , \modmult_1/N761 , \modmult_1/N760 ,
         \modmult_1/N759 , \modmult_1/N758 , \modmult_1/N757 ,
         \modmult_1/N756 , \modmult_1/N755 , \modmult_1/N754 ,
         \modmult_1/N753 , \modmult_1/N752 , \modmult_1/N751 ,
         \modmult_1/N750 , \modmult_1/N749 , \modmult_1/N748 ,
         \modmult_1/N747 , \modmult_1/N746 , \modmult_1/N745 ,
         \modmult_1/N744 , \modmult_1/N743 , \modmult_1/N742 ,
         \modmult_1/N741 , \modmult_1/N740 , \modmult_1/N739 ,
         \modmult_1/N738 , \modmult_1/N737 , \modmult_1/N736 ,
         \modmult_1/N735 , \modmult_1/N734 , \modmult_1/N733 ,
         \modmult_1/N732 , \modmult_1/N731 , \modmult_1/N730 ,
         \modmult_1/N729 , \modmult_1/N728 , \modmult_1/N727 ,
         \modmult_1/N726 , \modmult_1/N725 , \modmult_1/N724 ,
         \modmult_1/N723 , \modmult_1/N722 , \modmult_1/N721 ,
         \modmult_1/N720 , \modmult_1/N719 , \modmult_1/N718 ,
         \modmult_1/N717 , \modmult_1/N716 , \modmult_1/N715 ,
         \modmult_1/N714 , \modmult_1/N713 , \modmult_1/N712 ,
         \modmult_1/N711 , \modmult_1/N710 , \modmult_1/N709 ,
         \modmult_1/N708 , \modmult_1/N707 , \modmult_1/N706 ,
         \modmult_1/N705 , \modmult_1/N704 , \modmult_1/N703 ,
         \modmult_1/N702 , \modmult_1/N701 , \modmult_1/N700 ,
         \modmult_1/N699 , \modmult_1/N698 , \modmult_1/N697 ,
         \modmult_1/N696 , \modmult_1/N695 , \modmult_1/N694 ,
         \modmult_1/N693 , \modmult_1/N692 , \modmult_1/N691 ,
         \modmult_1/N690 , \modmult_1/N689 , \modmult_1/N688 ,
         \modmult_1/N687 , \modmult_1/N686 , \modmult_1/N685 ,
         \modmult_1/N684 , \modmult_1/N683 , \modmult_1/N682 ,
         \modmult_1/N681 , \modmult_1/N680 , \modmult_1/N679 ,
         \modmult_1/N678 , \modmult_1/N677 , \modmult_1/N676 ,
         \modmult_1/N675 , \modmult_1/N674 , \modmult_1/N673 ,
         \modmult_1/N672 , \modmult_1/N671 , \modmult_1/N670 ,
         \modmult_1/N669 , \modmult_1/N668 , \modmult_1/N667 ,
         \modmult_1/N666 , \modmult_1/N665 , \modmult_1/N664 ,
         \modmult_1/N663 , \modmult_1/N662 , \modmult_1/N661 ,
         \modmult_1/N660 , \modmult_1/N659 , \modmult_1/N658 ,
         \modmult_1/N657 , \modmult_1/N656 , \modmult_1/N655 ,
         \modmult_1/N654 , \modmult_1/N653 , \modmult_1/N652 ,
         \modmult_1/N651 , \modmult_1/N650 , \modmult_1/N649 ,
         \modmult_1/N648 , \modmult_1/N647 , \modmult_1/N646 ,
         \modmult_1/N645 , \modmult_1/N644 , \modmult_1/N643 ,
         \modmult_1/N642 , \modmult_1/N641 , \modmult_1/N640 ,
         \modmult_1/N639 , \modmult_1/N638 , \modmult_1/N637 ,
         \modmult_1/N636 , \modmult_1/N635 , \modmult_1/N634 ,
         \modmult_1/N633 , \modmult_1/N632 , \modmult_1/N631 ,
         \modmult_1/N630 , \modmult_1/N629 , \modmult_1/N628 ,
         \modmult_1/N627 , \modmult_1/N626 , \modmult_1/N625 ,
         \modmult_1/N624 , \modmult_1/N623 , \modmult_1/N622 ,
         \modmult_1/N621 , \modmult_1/N620 , \modmult_1/N619 ,
         \modmult_1/N618 , \modmult_1/N617 , \modmult_1/N616 ,
         \modmult_1/N615 , \modmult_1/N614 , \modmult_1/N613 ,
         \modmult_1/N612 , \modmult_1/N611 , \modmult_1/N610 ,
         \modmult_1/N609 , \modmult_1/N608 , \modmult_1/N607 ,
         \modmult_1/N606 , \modmult_1/N605 , \modmult_1/N604 ,
         \modmult_1/N603 , \modmult_1/N602 , \modmult_1/N601 ,
         \modmult_1/N600 , \modmult_1/N599 , \modmult_1/N598 ,
         \modmult_1/N597 , \modmult_1/N596 , \modmult_1/N595 ,
         \modmult_1/N594 , \modmult_1/N593 , \modmult_1/N592 ,
         \modmult_1/N591 , \modmult_1/N590 , \modmult_1/N589 ,
         \modmult_1/N588 , \modmult_1/N587 , \modmult_1/N586 ,
         \modmult_1/N585 , \modmult_1/N584 , \modmult_1/N583 ,
         \modmult_1/N582 , \modmult_1/N581 , \modmult_1/N580 ,
         \modmult_1/N579 , \modmult_1/N578 , \modmult_1/N577 ,
         \modmult_1/N576 , \modmult_1/N575 , \modmult_1/N574 ,
         \modmult_1/N573 , \modmult_1/N572 , \modmult_1/N571 ,
         \modmult_1/N570 , \modmult_1/N569 , \modmult_1/N568 ,
         \modmult_1/N567 , \modmult_1/N566 , \modmult_1/N565 ,
         \modmult_1/N564 , \modmult_1/N563 , \modmult_1/N562 ,
         \modmult_1/N561 , \modmult_1/N560 , \modmult_1/N559 ,
         \modmult_1/N558 , \modmult_1/N557 , \modmult_1/N556 ,
         \modmult_1/N555 , \modmult_1/N554 , \modmult_1/N553 ,
         \modmult_1/N552 , \modmult_1/N551 , \modmult_1/N550 ,
         \modmult_1/N549 , \modmult_1/N548 , \modmult_1/N547 ,
         \modmult_1/N546 , \modmult_1/N545 , \modmult_1/N544 ,
         \modmult_1/N543 , \modmult_1/N542 , \modmult_1/N541 ,
         \modmult_1/N540 , \modmult_1/N539 , \modmult_1/N538 ,
         \modmult_1/N537 , \modmult_1/N536 , \modmult_1/N535 ,
         \modmult_1/N534 , \modmult_1/N533 , \modmult_1/N532 ,
         \modmult_1/N531 , \modmult_1/N530 , \modmult_1/N529 ,
         \modmult_1/N528 , \modmult_1/N527 , \modmult_1/N526 ,
         \modmult_1/N525 , \modmult_1/N524 , \modmult_1/N523 ,
         \modmult_1/N522 , \modmult_1/N521 , \modmult_1/N520 ,
         \modmult_1/N519 , \modmult_1/N518 , \modmult_1/N517 ,
         \modmult_1/N516 , \modmult_1/N515 , \modmult_1/N514 ,
         \modmult_1/N513 , \modmult_1/N512 , \modmult_1/N511 ,
         \modmult_1/N510 , \modmult_1/N509 , \modmult_1/N508 ,
         \modmult_1/N507 , \modmult_1/N506 , \modmult_1/N505 ,
         \modmult_1/N504 , \modmult_1/N503 , \modmult_1/N502 ,
         \modmult_1/N501 , \modmult_1/N500 , \modmult_1/N499 ,
         \modmult_1/N498 , \modmult_1/N497 , \modmult_1/N496 ,
         \modmult_1/N495 , \modmult_1/N494 , \modmult_1/N493 ,
         \modmult_1/N492 , \modmult_1/N491 , \modmult_1/N490 ,
         \modmult_1/N489 , \modmult_1/N488 , \modmult_1/N487 ,
         \modmult_1/N486 , \modmult_1/N485 , \modmult_1/N484 ,
         \modmult_1/N483 , \modmult_1/N482 , \modmult_1/N481 ,
         \modmult_1/N480 , \modmult_1/N479 , \modmult_1/N478 ,
         \modmult_1/N477 , \modmult_1/N476 , \modmult_1/N475 ,
         \modmult_1/N474 , \modmult_1/N473 , \modmult_1/N472 ,
         \modmult_1/N471 , \modmult_1/N470 , \modmult_1/N469 ,
         \modmult_1/N468 , \modmult_1/N467 , \modmult_1/N466 ,
         \modmult_1/N465 , \modmult_1/N464 , \modmult_1/N463 ,
         \modmult_1/N462 , \modmult_1/N461 , \modmult_1/N460 ,
         \modmult_1/N459 , \modmult_1/N458 , \modmult_1/N457 ,
         \modmult_1/N456 , \modmult_1/N455 , \modmult_1/N454 ,
         \modmult_1/N453 , \modmult_1/N452 , \modmult_1/N451 ,
         \modmult_1/N450 , \modmult_1/N449 , \modmult_1/N448 ,
         \modmult_1/N447 , \modmult_1/N446 , \modmult_1/N445 ,
         \modmult_1/N444 , \modmult_1/N443 , \modmult_1/N442 ,
         \modmult_1/N441 , \modmult_1/N440 , \modmult_1/N439 ,
         \modmult_1/N438 , \modmult_1/N437 , \modmult_1/N436 ,
         \modmult_1/N435 , \modmult_1/N434 , \modmult_1/N433 ,
         \modmult_1/N432 , \modmult_1/N431 , \modmult_1/N430 ,
         \modmult_1/N429 , \modmult_1/N428 , \modmult_1/N427 ,
         \modmult_1/N426 , \modmult_1/N425 , \modmult_1/N424 ,
         \modmult_1/N423 , \modmult_1/N422 , \modmult_1/N421 ,
         \modmult_1/N420 , \modmult_1/N419 , \modmult_1/N418 ,
         \modmult_1/N417 , \modmult_1/N416 , \modmult_1/N415 ,
         \modmult_1/N414 , \modmult_1/N413 , \modmult_1/N412 ,
         \modmult_1/N411 , \modmult_1/N410 , \modmult_1/N409 ,
         \modmult_1/N408 , \modmult_1/N407 , \modmult_1/N406 ,
         \modmult_1/N405 , \modmult_1/N404 , \modmult_1/N403 ,
         \modmult_1/N402 , \modmult_1/N401 , \modmult_1/N400 ,
         \modmult_1/N399 , \modmult_1/N398 , \modmult_1/N397 ,
         \modmult_1/N396 , \modmult_1/N395 , \modmult_1/N394 ,
         \modmult_1/N393 , \modmult_1/N392 , \modmult_1/N391 ,
         \modmult_1/N390 , \modmult_1/N389 , \modmult_1/N388 ,
         \modmult_1/N387 , \modmult_1/N386 , \modmult_1/N385 ,
         \modmult_1/N384 , \modmult_1/N383 , \modmult_1/N382 ,
         \modmult_1/N381 , \modmult_1/N380 , \modmult_1/N379 ,
         \modmult_1/N378 , \modmult_1/N377 , \modmult_1/N376 ,
         \modmult_1/N375 , \modmult_1/N374 , \modmult_1/N373 ,
         \modmult_1/N372 , \modmult_1/N371 , \modmult_1/N370 ,
         \modmult_1/N369 , \modmult_1/N368 , \modmult_1/N367 ,
         \modmult_1/N366 , \modmult_1/N365 , \modmult_1/N364 ,
         \modmult_1/N363 , \modmult_1/N362 , \modmult_1/N361 ,
         \modmult_1/N360 , \modmult_1/N359 , \modmult_1/N358 ,
         \modmult_1/N357 , \modmult_1/N356 , \modmult_1/N355 ,
         \modmult_1/N354 , \modmult_1/N353 , \modmult_1/N352 ,
         \modmult_1/N351 , \modmult_1/N350 , \modmult_1/N349 ,
         \modmult_1/N348 , \modmult_1/N347 , \modmult_1/N346 ,
         \modmult_1/N345 , \modmult_1/N344 , \modmult_1/N343 ,
         \modmult_1/N342 , \modmult_1/N341 , \modmult_1/N340 ,
         \modmult_1/N339 , \modmult_1/N338 , \modmult_1/N337 ,
         \modmult_1/N336 , \modmult_1/N335 , \modmult_1/N334 ,
         \modmult_1/N333 , \modmult_1/N332 , \modmult_1/N331 ,
         \modmult_1/N330 , \modmult_1/N329 , \modmult_1/N328 ,
         \modmult_1/N327 , \modmult_1/N326 , \modmult_1/N325 ,
         \modmult_1/N324 , \modmult_1/N323 , \modmult_1/N322 ,
         \modmult_1/N321 , \modmult_1/N320 , \modmult_1/N319 ,
         \modmult_1/N318 , \modmult_1/N317 , \modmult_1/N316 ,
         \modmult_1/N315 , \modmult_1/N314 , \modmult_1/N313 ,
         \modmult_1/N312 , \modmult_1/N311 , \modmult_1/N310 ,
         \modmult_1/N309 , \modmult_1/N308 , \modmult_1/N307 ,
         \modmult_1/N306 , \modmult_1/N305 , \modmult_1/N304 ,
         \modmult_1/N303 , \modmult_1/N302 , \modmult_1/N301 ,
         \modmult_1/N300 , \modmult_1/N299 , \modmult_1/N298 ,
         \modmult_1/N297 , \modmult_1/N296 , \modmult_1/N295 ,
         \modmult_1/N294 , \modmult_1/N293 , \modmult_1/N292 ,
         \modmult_1/N291 , \modmult_1/N290 , \modmult_1/N289 ,
         \modmult_1/N288 , \modmult_1/N287 , \modmult_1/N286 ,
         \modmult_1/N285 , \modmult_1/N284 , \modmult_1/N283 ,
         \modmult_1/N282 , \modmult_1/N281 , \modmult_1/N280 ,
         \modmult_1/N279 , \modmult_1/N278 , \modmult_1/N277 ,
         \modmult_1/N276 , \modmult_1/N275 , \modmult_1/N274 ,
         \modmult_1/N273 , \modmult_1/N272 , \modmult_1/N271 ,
         \modmult_1/N270 , \modmult_1/N269 , \modmult_1/N268 ,
         \modmult_1/N267 , \modmult_1/N266 , \modmult_1/N265 ,
         \modmult_1/N264 , \modmult_1/N263 , \modmult_1/N262 ,
         \modmult_1/N261 , \modmult_1/N260 , \modmult_1/N259 ,
         \modmult_1/N258 , \modmult_1/N257 , \modmult_1/N256 ,
         \modmult_1/N255 , \modmult_1/N254 , \modmult_1/N253 ,
         \modmult_1/N252 , \modmult_1/N251 , \modmult_1/N250 ,
         \modmult_1/N249 , \modmult_1/N248 , \modmult_1/N247 ,
         \modmult_1/N246 , \modmult_1/N245 , \modmult_1/N244 ,
         \modmult_1/N243 , \modmult_1/N242 , \modmult_1/N241 ,
         \modmult_1/N240 , \modmult_1/N239 , \modmult_1/N238 ,
         \modmult_1/N237 , \modmult_1/N236 , \modmult_1/N235 ,
         \modmult_1/N234 , \modmult_1/N233 , \modmult_1/N232 ,
         \modmult_1/N231 , \modmult_1/N230 , \modmult_1/N229 ,
         \modmult_1/N228 , \modmult_1/N227 , \modmult_1/N226 ,
         \modmult_1/N225 , \modmult_1/N224 , \modmult_1/N223 ,
         \modmult_1/N222 , \modmult_1/N221 , \modmult_1/N220 ,
         \modmult_1/N219 , \modmult_1/N218 , \modmult_1/N217 ,
         \modmult_1/N216 , \modmult_1/N215 , \modmult_1/N214 ,
         \modmult_1/N213 , \modmult_1/N212 , \modmult_1/N211 ,
         \modmult_1/N210 , \modmult_1/N209 , \modmult_1/N208 ,
         \modmult_1/N207 , \modmult_1/N206 , \modmult_1/N205 ,
         \modmult_1/N204 , \modmult_1/N203 , \modmult_1/N202 ,
         \modmult_1/N201 , \modmult_1/N200 , \modmult_1/N199 ,
         \modmult_1/N198 , \modmult_1/N197 , \modmult_1/N196 ,
         \modmult_1/N195 , \modmult_1/N194 , \modmult_1/N193 ,
         \modmult_1/N192 , \modmult_1/N191 , \modmult_1/N190 ,
         \modmult_1/N189 , \modmult_1/N188 , \modmult_1/N187 ,
         \modmult_1/N186 , \modmult_1/N185 , \modmult_1/N184 ,
         \modmult_1/N183 , \modmult_1/N182 , \modmult_1/N181 ,
         \modmult_1/N180 , \modmult_1/N179 , \modmult_1/N178 ,
         \modmult_1/N177 , \modmult_1/N176 , \modmult_1/N175 ,
         \modmult_1/N174 , \modmult_1/N173 , \modmult_1/N172 ,
         \modmult_1/N171 , \modmult_1/N170 , \modmult_1/N169 ,
         \modmult_1/N168 , \modmult_1/N167 , \modmult_1/N166 ,
         \modmult_1/N165 , \modmult_1/N164 , \modmult_1/N163 ,
         \modmult_1/N162 , \modmult_1/N161 , \modmult_1/N160 ,
         \modmult_1/N159 , \modmult_1/N158 , \modmult_1/N157 ,
         \modmult_1/N156 , \modmult_1/N155 , \modmult_1/N154 ,
         \modmult_1/N153 , \modmult_1/N152 , \modmult_1/N151 ,
         \modmult_1/N150 , \modmult_1/N149 , \modmult_1/N148 ,
         \modmult_1/N147 , \modmult_1/N146 , \modmult_1/N145 ,
         \modmult_1/N144 , \modmult_1/N143 , \modmult_1/N142 ,
         \modmult_1/N141 , \modmult_1/N140 , \modmult_1/N139 ,
         \modmult_1/N138 , \modmult_1/N137 , \modmult_1/N136 ,
         \modmult_1/N135 , \modmult_1/N134 , \modmult_1/N133 ,
         \modmult_1/N132 , \modmult_1/N131 , \modmult_1/N130 ,
         \modmult_1/N129 , \modmult_1/N128 , \modmult_1/N127 ,
         \modmult_1/N126 , \modmult_1/N125 , \modmult_1/N124 ,
         \modmult_1/N123 , \modmult_1/N122 , \modmult_1/N121 ,
         \modmult_1/N120 , \modmult_1/N119 , \modmult_1/N118 ,
         \modmult_1/N117 , \modmult_1/N116 , \modmult_1/N115 ,
         \modmult_1/N114 , \modmult_1/N113 , \modmult_1/N112 ,
         \modmult_1/N111 , \modmult_1/N110 , \modmult_1/N109 ,
         \modmult_1/N108 , \modmult_1/N107 , \modmult_1/N106 ,
         \modmult_1/N105 , \modmult_1/N104 , \modmult_1/N103 ,
         \modmult_1/N102 , \modmult_1/N101 , \modmult_1/N100 , \modmult_1/N99 ,
         \modmult_1/N98 , \modmult_1/N97 , \modmult_1/N96 , \modmult_1/N95 ,
         \modmult_1/N94 , \modmult_1/N93 , \modmult_1/N92 , \modmult_1/N91 ,
         \modmult_1/N90 , \modmult_1/N89 , \modmult_1/N88 , \modmult_1/N87 ,
         \modmult_1/N86 , \modmult_1/N85 , \modmult_1/N84 , \modmult_1/N83 ,
         \modmult_1/N82 , \modmult_1/N81 , \modmult_1/N80 , \modmult_1/N79 ,
         \modmult_1/N78 , \modmult_1/N77 , \modmult_1/N76 , \modmult_1/N75 ,
         \modmult_1/N74 , \modmult_1/N73 , \modmult_1/N72 , \modmult_1/N71 ,
         \modmult_1/N70 , \modmult_1/N69 , \modmult_1/N68 , \modmult_1/N67 ,
         \modmult_1/N66 , \modmult_1/N65 , \modmult_1/N64 , \modmult_1/N63 ,
         \modmult_1/N62 , \modmult_1/N61 , \modmult_1/N60 , \modmult_1/N59 ,
         \modmult_1/N58 , \modmult_1/N57 , \modmult_1/N56 , \modmult_1/N55 ,
         \modmult_1/N54 , \modmult_1/N53 , \modmult_1/N52 , \modmult_1/N51 ,
         \modmult_1/N50 , \modmult_1/N49 , \modmult_1/N48 , \modmult_1/N47 ,
         \modmult_1/N46 , \modmult_1/N45 , \modmult_1/N44 , \modmult_1/N43 ,
         \modmult_1/N42 , \modmult_1/N41 , \modmult_1/N40 , \modmult_1/N39 ,
         \modmult_1/N38 , \modmult_1/N37 , \modmult_1/N36 , \modmult_1/N35 ,
         \modmult_1/N34 , \modmult_1/N33 , \modmult_1/N32 , \modmult_1/N31 ,
         \modmult_1/N30 , \modmult_1/N29 , \modmult_1/N28 , \modmult_1/N27 ,
         \modmult_1/N26 , \modmult_1/N25 , \modmult_1/N24 , \modmult_1/N23 ,
         \modmult_1/N22 , \modmult_1/N21 , \modmult_1/N20 , \modmult_1/N19 ,
         \modmult_1/N18 , \modmult_1/N17 , \modmult_1/N16 , \modmult_1/N15 ,
         \modmult_1/N14 , \modmult_1/N13 , \modmult_1/N12 , \modmult_1/N11 ,
         \modmult_1/N10 , \modmult_1/N9 , \modmult_1/N8 , \modmult_1/N7 ,
         \modmult_1/N6 , \modmult_1/N5 , \modmult_1/N4 , \modmult_1/N3 ,
         \modmult_1/xin[1023] , \modmult_1/xin[1022] , \modmult_1/xin[1021] ,
         \modmult_1/xin[1020] , \modmult_1/xin[1019] , \modmult_1/xin[1018] ,
         \modmult_1/xin[1017] , \modmult_1/xin[1016] , \modmult_1/xin[1015] ,
         \modmult_1/xin[1014] , \modmult_1/xin[1013] , \modmult_1/xin[1012] ,
         \modmult_1/xin[1011] , \modmult_1/xin[1010] , \modmult_1/xin[1009] ,
         \modmult_1/xin[1008] , \modmult_1/xin[1007] , \modmult_1/xin[1006] ,
         \modmult_1/xin[1005] , \modmult_1/xin[1004] , \modmult_1/xin[1003] ,
         \modmult_1/xin[1002] , \modmult_1/xin[1001] , \modmult_1/xin[1000] ,
         \modmult_1/xin[999] , \modmult_1/xin[998] , \modmult_1/xin[997] ,
         \modmult_1/xin[996] , \modmult_1/xin[995] , \modmult_1/xin[994] ,
         \modmult_1/xin[993] , \modmult_1/xin[992] , \modmult_1/xin[991] ,
         \modmult_1/xin[990] , \modmult_1/xin[989] , \modmult_1/xin[988] ,
         \modmult_1/xin[987] , \modmult_1/xin[986] , \modmult_1/xin[985] ,
         \modmult_1/xin[984] , \modmult_1/xin[983] , \modmult_1/xin[982] ,
         \modmult_1/xin[981] , \modmult_1/xin[980] , \modmult_1/xin[979] ,
         \modmult_1/xin[978] , \modmult_1/xin[977] , \modmult_1/xin[976] ,
         \modmult_1/xin[975] , \modmult_1/xin[974] , \modmult_1/xin[973] ,
         \modmult_1/xin[972] , \modmult_1/xin[971] , \modmult_1/xin[970] ,
         \modmult_1/xin[969] , \modmult_1/xin[968] , \modmult_1/xin[967] ,
         \modmult_1/xin[966] , \modmult_1/xin[965] , \modmult_1/xin[964] ,
         \modmult_1/xin[963] , \modmult_1/xin[962] , \modmult_1/xin[961] ,
         \modmult_1/xin[960] , \modmult_1/xin[959] , \modmult_1/xin[958] ,
         \modmult_1/xin[957] , \modmult_1/xin[956] , \modmult_1/xin[955] ,
         \modmult_1/xin[954] , \modmult_1/xin[953] , \modmult_1/xin[952] ,
         \modmult_1/xin[951] , \modmult_1/xin[950] , \modmult_1/xin[949] ,
         \modmult_1/xin[948] , \modmult_1/xin[947] , \modmult_1/xin[946] ,
         \modmult_1/xin[945] , \modmult_1/xin[944] , \modmult_1/xin[943] ,
         \modmult_1/xin[942] , \modmult_1/xin[941] , \modmult_1/xin[940] ,
         \modmult_1/xin[939] , \modmult_1/xin[938] , \modmult_1/xin[937] ,
         \modmult_1/xin[936] , \modmult_1/xin[935] , \modmult_1/xin[934] ,
         \modmult_1/xin[933] , \modmult_1/xin[932] , \modmult_1/xin[931] ,
         \modmult_1/xin[930] , \modmult_1/xin[929] , \modmult_1/xin[928] ,
         \modmult_1/xin[927] , \modmult_1/xin[926] , \modmult_1/xin[925] ,
         \modmult_1/xin[924] , \modmult_1/xin[923] , \modmult_1/xin[922] ,
         \modmult_1/xin[921] , \modmult_1/xin[920] , \modmult_1/xin[919] ,
         \modmult_1/xin[918] , \modmult_1/xin[917] , \modmult_1/xin[916] ,
         \modmult_1/xin[915] , \modmult_1/xin[914] , \modmult_1/xin[913] ,
         \modmult_1/xin[912] , \modmult_1/xin[911] , \modmult_1/xin[910] ,
         \modmult_1/xin[909] , \modmult_1/xin[908] , \modmult_1/xin[907] ,
         \modmult_1/xin[906] , \modmult_1/xin[905] , \modmult_1/xin[904] ,
         \modmult_1/xin[903] , \modmult_1/xin[902] , \modmult_1/xin[901] ,
         \modmult_1/xin[900] , \modmult_1/xin[899] , \modmult_1/xin[898] ,
         \modmult_1/xin[897] , \modmult_1/xin[896] , \modmult_1/xin[895] ,
         \modmult_1/xin[894] , \modmult_1/xin[893] , \modmult_1/xin[892] ,
         \modmult_1/xin[891] , \modmult_1/xin[890] , \modmult_1/xin[889] ,
         \modmult_1/xin[888] , \modmult_1/xin[887] , \modmult_1/xin[886] ,
         \modmult_1/xin[885] , \modmult_1/xin[884] , \modmult_1/xin[883] ,
         \modmult_1/xin[882] , \modmult_1/xin[881] , \modmult_1/xin[880] ,
         \modmult_1/xin[879] , \modmult_1/xin[878] , \modmult_1/xin[877] ,
         \modmult_1/xin[876] , \modmult_1/xin[875] , \modmult_1/xin[874] ,
         \modmult_1/xin[873] , \modmult_1/xin[872] , \modmult_1/xin[871] ,
         \modmult_1/xin[870] , \modmult_1/xin[869] , \modmult_1/xin[868] ,
         \modmult_1/xin[867] , \modmult_1/xin[866] , \modmult_1/xin[865] ,
         \modmult_1/xin[864] , \modmult_1/xin[863] , \modmult_1/xin[862] ,
         \modmult_1/xin[861] , \modmult_1/xin[860] , \modmult_1/xin[859] ,
         \modmult_1/xin[858] , \modmult_1/xin[857] , \modmult_1/xin[856] ,
         \modmult_1/xin[855] , \modmult_1/xin[854] , \modmult_1/xin[853] ,
         \modmult_1/xin[852] , \modmult_1/xin[851] , \modmult_1/xin[850] ,
         \modmult_1/xin[849] , \modmult_1/xin[848] , \modmult_1/xin[847] ,
         \modmult_1/xin[846] , \modmult_1/xin[845] , \modmult_1/xin[844] ,
         \modmult_1/xin[843] , \modmult_1/xin[842] , \modmult_1/xin[841] ,
         \modmult_1/xin[840] , \modmult_1/xin[839] , \modmult_1/xin[838] ,
         \modmult_1/xin[837] , \modmult_1/xin[836] , \modmult_1/xin[835] ,
         \modmult_1/xin[834] , \modmult_1/xin[833] , \modmult_1/xin[832] ,
         \modmult_1/xin[831] , \modmult_1/xin[830] , \modmult_1/xin[829] ,
         \modmult_1/xin[828] , \modmult_1/xin[827] , \modmult_1/xin[826] ,
         \modmult_1/xin[825] , \modmult_1/xin[824] , \modmult_1/xin[823] ,
         \modmult_1/xin[822] , \modmult_1/xin[821] , \modmult_1/xin[820] ,
         \modmult_1/xin[819] , \modmult_1/xin[818] , \modmult_1/xin[817] ,
         \modmult_1/xin[816] , \modmult_1/xin[815] , \modmult_1/xin[814] ,
         \modmult_1/xin[813] , \modmult_1/xin[812] , \modmult_1/xin[811] ,
         \modmult_1/xin[810] , \modmult_1/xin[809] , \modmult_1/xin[808] ,
         \modmult_1/xin[807] , \modmult_1/xin[806] , \modmult_1/xin[805] ,
         \modmult_1/xin[804] , \modmult_1/xin[803] , \modmult_1/xin[802] ,
         \modmult_1/xin[801] , \modmult_1/xin[800] , \modmult_1/xin[799] ,
         \modmult_1/xin[798] , \modmult_1/xin[797] , \modmult_1/xin[796] ,
         \modmult_1/xin[795] , \modmult_1/xin[794] , \modmult_1/xin[793] ,
         \modmult_1/xin[792] , \modmult_1/xin[791] , \modmult_1/xin[790] ,
         \modmult_1/xin[789] , \modmult_1/xin[788] , \modmult_1/xin[787] ,
         \modmult_1/xin[786] , \modmult_1/xin[785] , \modmult_1/xin[784] ,
         \modmult_1/xin[783] , \modmult_1/xin[782] , \modmult_1/xin[781] ,
         \modmult_1/xin[780] , \modmult_1/xin[779] , \modmult_1/xin[778] ,
         \modmult_1/xin[777] , \modmult_1/xin[776] , \modmult_1/xin[775] ,
         \modmult_1/xin[774] , \modmult_1/xin[773] , \modmult_1/xin[772] ,
         \modmult_1/xin[771] , \modmult_1/xin[770] , \modmult_1/xin[769] ,
         \modmult_1/xin[768] , \modmult_1/xin[767] , \modmult_1/xin[766] ,
         \modmult_1/xin[765] , \modmult_1/xin[764] , \modmult_1/xin[763] ,
         \modmult_1/xin[762] , \modmult_1/xin[761] , \modmult_1/xin[760] ,
         \modmult_1/xin[759] , \modmult_1/xin[758] , \modmult_1/xin[757] ,
         \modmult_1/xin[756] , \modmult_1/xin[755] , \modmult_1/xin[754] ,
         \modmult_1/xin[753] , \modmult_1/xin[752] , \modmult_1/xin[751] ,
         \modmult_1/xin[750] , \modmult_1/xin[749] , \modmult_1/xin[748] ,
         \modmult_1/xin[747] , \modmult_1/xin[746] , \modmult_1/xin[745] ,
         \modmult_1/xin[744] , \modmult_1/xin[743] , \modmult_1/xin[742] ,
         \modmult_1/xin[741] , \modmult_1/xin[740] , \modmult_1/xin[739] ,
         \modmult_1/xin[738] , \modmult_1/xin[737] , \modmult_1/xin[736] ,
         \modmult_1/xin[735] , \modmult_1/xin[734] , \modmult_1/xin[733] ,
         \modmult_1/xin[732] , \modmult_1/xin[731] , \modmult_1/xin[730] ,
         \modmult_1/xin[729] , \modmult_1/xin[728] , \modmult_1/xin[727] ,
         \modmult_1/xin[726] , \modmult_1/xin[725] , \modmult_1/xin[724] ,
         \modmult_1/xin[723] , \modmult_1/xin[722] , \modmult_1/xin[721] ,
         \modmult_1/xin[720] , \modmult_1/xin[719] , \modmult_1/xin[718] ,
         \modmult_1/xin[717] , \modmult_1/xin[716] , \modmult_1/xin[715] ,
         \modmult_1/xin[714] , \modmult_1/xin[713] , \modmult_1/xin[712] ,
         \modmult_1/xin[711] , \modmult_1/xin[710] , \modmult_1/xin[709] ,
         \modmult_1/xin[708] , \modmult_1/xin[707] , \modmult_1/xin[706] ,
         \modmult_1/xin[705] , \modmult_1/xin[704] , \modmult_1/xin[703] ,
         \modmult_1/xin[702] , \modmult_1/xin[701] , \modmult_1/xin[700] ,
         \modmult_1/xin[699] , \modmult_1/xin[698] , \modmult_1/xin[697] ,
         \modmult_1/xin[696] , \modmult_1/xin[695] , \modmult_1/xin[694] ,
         \modmult_1/xin[693] , \modmult_1/xin[692] , \modmult_1/xin[691] ,
         \modmult_1/xin[690] , \modmult_1/xin[689] , \modmult_1/xin[688] ,
         \modmult_1/xin[687] , \modmult_1/xin[686] , \modmult_1/xin[685] ,
         \modmult_1/xin[684] , \modmult_1/xin[683] , \modmult_1/xin[682] ,
         \modmult_1/xin[681] , \modmult_1/xin[680] , \modmult_1/xin[679] ,
         \modmult_1/xin[678] , \modmult_1/xin[677] , \modmult_1/xin[676] ,
         \modmult_1/xin[675] , \modmult_1/xin[674] , \modmult_1/xin[673] ,
         \modmult_1/xin[672] , \modmult_1/xin[671] , \modmult_1/xin[670] ,
         \modmult_1/xin[669] , \modmult_1/xin[668] , \modmult_1/xin[667] ,
         \modmult_1/xin[666] , \modmult_1/xin[665] , \modmult_1/xin[664] ,
         \modmult_1/xin[663] , \modmult_1/xin[662] , \modmult_1/xin[661] ,
         \modmult_1/xin[660] , \modmult_1/xin[659] , \modmult_1/xin[658] ,
         \modmult_1/xin[657] , \modmult_1/xin[656] , \modmult_1/xin[655] ,
         \modmult_1/xin[654] , \modmult_1/xin[653] , \modmult_1/xin[652] ,
         \modmult_1/xin[651] , \modmult_1/xin[650] , \modmult_1/xin[649] ,
         \modmult_1/xin[648] , \modmult_1/xin[647] , \modmult_1/xin[646] ,
         \modmult_1/xin[645] , \modmult_1/xin[644] , \modmult_1/xin[643] ,
         \modmult_1/xin[642] , \modmult_1/xin[641] , \modmult_1/xin[640] ,
         \modmult_1/xin[639] , \modmult_1/xin[638] , \modmult_1/xin[637] ,
         \modmult_1/xin[636] , \modmult_1/xin[635] , \modmult_1/xin[634] ,
         \modmult_1/xin[633] , \modmult_1/xin[632] , \modmult_1/xin[631] ,
         \modmult_1/xin[630] , \modmult_1/xin[629] , \modmult_1/xin[628] ,
         \modmult_1/xin[627] , \modmult_1/xin[626] , \modmult_1/xin[625] ,
         \modmult_1/xin[624] , \modmult_1/xin[623] , \modmult_1/xin[622] ,
         \modmult_1/xin[621] , \modmult_1/xin[620] , \modmult_1/xin[619] ,
         \modmult_1/xin[618] , \modmult_1/xin[617] , \modmult_1/xin[616] ,
         \modmult_1/xin[615] , \modmult_1/xin[614] , \modmult_1/xin[613] ,
         \modmult_1/xin[612] , \modmult_1/xin[611] , \modmult_1/xin[610] ,
         \modmult_1/xin[609] , \modmult_1/xin[608] , \modmult_1/xin[607] ,
         \modmult_1/xin[606] , \modmult_1/xin[605] , \modmult_1/xin[604] ,
         \modmult_1/xin[603] , \modmult_1/xin[602] , \modmult_1/xin[601] ,
         \modmult_1/xin[600] , \modmult_1/xin[599] , \modmult_1/xin[598] ,
         \modmult_1/xin[597] , \modmult_1/xin[596] , \modmult_1/xin[595] ,
         \modmult_1/xin[594] , \modmult_1/xin[593] , \modmult_1/xin[592] ,
         \modmult_1/xin[591] , \modmult_1/xin[590] , \modmult_1/xin[589] ,
         \modmult_1/xin[588] , \modmult_1/xin[587] , \modmult_1/xin[586] ,
         \modmult_1/xin[585] , \modmult_1/xin[584] , \modmult_1/xin[583] ,
         \modmult_1/xin[582] , \modmult_1/xin[581] , \modmult_1/xin[580] ,
         \modmult_1/xin[579] , \modmult_1/xin[578] , \modmult_1/xin[577] ,
         \modmult_1/xin[576] , \modmult_1/xin[575] , \modmult_1/xin[574] ,
         \modmult_1/xin[573] , \modmult_1/xin[572] , \modmult_1/xin[571] ,
         \modmult_1/xin[570] , \modmult_1/xin[569] , \modmult_1/xin[568] ,
         \modmult_1/xin[567] , \modmult_1/xin[566] , \modmult_1/xin[565] ,
         \modmult_1/xin[564] , \modmult_1/xin[563] , \modmult_1/xin[562] ,
         \modmult_1/xin[561] , \modmult_1/xin[560] , \modmult_1/xin[559] ,
         \modmult_1/xin[558] , \modmult_1/xin[557] , \modmult_1/xin[556] ,
         \modmult_1/xin[555] , \modmult_1/xin[554] , \modmult_1/xin[553] ,
         \modmult_1/xin[552] , \modmult_1/xin[551] , \modmult_1/xin[550] ,
         \modmult_1/xin[549] , \modmult_1/xin[548] , \modmult_1/xin[547] ,
         \modmult_1/xin[546] , \modmult_1/xin[545] , \modmult_1/xin[544] ,
         \modmult_1/xin[543] , \modmult_1/xin[542] , \modmult_1/xin[541] ,
         \modmult_1/xin[540] , \modmult_1/xin[539] , \modmult_1/xin[538] ,
         \modmult_1/xin[537] , \modmult_1/xin[536] , \modmult_1/xin[535] ,
         \modmult_1/xin[534] , \modmult_1/xin[533] , \modmult_1/xin[532] ,
         \modmult_1/xin[531] , \modmult_1/xin[530] , \modmult_1/xin[529] ,
         \modmult_1/xin[528] , \modmult_1/xin[527] , \modmult_1/xin[526] ,
         \modmult_1/xin[525] , \modmult_1/xin[524] , \modmult_1/xin[523] ,
         \modmult_1/xin[522] , \modmult_1/xin[521] , \modmult_1/xin[520] ,
         \modmult_1/xin[519] , \modmult_1/xin[518] , \modmult_1/xin[517] ,
         \modmult_1/xin[516] , \modmult_1/xin[515] , \modmult_1/xin[514] ,
         \modmult_1/xin[513] , \modmult_1/xin[512] , \modmult_1/xin[511] ,
         \modmult_1/xin[510] , \modmult_1/xin[509] , \modmult_1/xin[508] ,
         \modmult_1/xin[507] , \modmult_1/xin[506] , \modmult_1/xin[505] ,
         \modmult_1/xin[504] , \modmult_1/xin[503] , \modmult_1/xin[502] ,
         \modmult_1/xin[501] , \modmult_1/xin[500] , \modmult_1/xin[499] ,
         \modmult_1/xin[498] , \modmult_1/xin[497] , \modmult_1/xin[496] ,
         \modmult_1/xin[495] , \modmult_1/xin[494] , \modmult_1/xin[493] ,
         \modmult_1/xin[492] , \modmult_1/xin[491] , \modmult_1/xin[490] ,
         \modmult_1/xin[489] , \modmult_1/xin[488] , \modmult_1/xin[487] ,
         \modmult_1/xin[486] , \modmult_1/xin[485] , \modmult_1/xin[484] ,
         \modmult_1/xin[483] , \modmult_1/xin[482] , \modmult_1/xin[481] ,
         \modmult_1/xin[480] , \modmult_1/xin[479] , \modmult_1/xin[478] ,
         \modmult_1/xin[477] , \modmult_1/xin[476] , \modmult_1/xin[475] ,
         \modmult_1/xin[474] , \modmult_1/xin[473] , \modmult_1/xin[472] ,
         \modmult_1/xin[471] , \modmult_1/xin[470] , \modmult_1/xin[469] ,
         \modmult_1/xin[468] , \modmult_1/xin[467] , \modmult_1/xin[466] ,
         \modmult_1/xin[465] , \modmult_1/xin[464] , \modmult_1/xin[463] ,
         \modmult_1/xin[462] , \modmult_1/xin[461] , \modmult_1/xin[460] ,
         \modmult_1/xin[459] , \modmult_1/xin[458] , \modmult_1/xin[457] ,
         \modmult_1/xin[456] , \modmult_1/xin[455] , \modmult_1/xin[454] ,
         \modmult_1/xin[453] , \modmult_1/xin[452] , \modmult_1/xin[451] ,
         \modmult_1/xin[450] , \modmult_1/xin[449] , \modmult_1/xin[448] ,
         \modmult_1/xin[447] , \modmult_1/xin[446] , \modmult_1/xin[445] ,
         \modmult_1/xin[444] , \modmult_1/xin[443] , \modmult_1/xin[442] ,
         \modmult_1/xin[441] , \modmult_1/xin[440] , \modmult_1/xin[439] ,
         \modmult_1/xin[438] , \modmult_1/xin[437] , \modmult_1/xin[436] ,
         \modmult_1/xin[435] , \modmult_1/xin[434] , \modmult_1/xin[433] ,
         \modmult_1/xin[432] , \modmult_1/xin[431] , \modmult_1/xin[430] ,
         \modmult_1/xin[429] , \modmult_1/xin[428] , \modmult_1/xin[427] ,
         \modmult_1/xin[426] , \modmult_1/xin[425] , \modmult_1/xin[424] ,
         \modmult_1/xin[423] , \modmult_1/xin[422] , \modmult_1/xin[421] ,
         \modmult_1/xin[420] , \modmult_1/xin[419] , \modmult_1/xin[418] ,
         \modmult_1/xin[417] , \modmult_1/xin[416] , \modmult_1/xin[415] ,
         \modmult_1/xin[414] , \modmult_1/xin[413] , \modmult_1/xin[412] ,
         \modmult_1/xin[411] , \modmult_1/xin[410] , \modmult_1/xin[409] ,
         \modmult_1/xin[408] , \modmult_1/xin[407] , \modmult_1/xin[406] ,
         \modmult_1/xin[405] , \modmult_1/xin[404] , \modmult_1/xin[403] ,
         \modmult_1/xin[402] , \modmult_1/xin[401] , \modmult_1/xin[400] ,
         \modmult_1/xin[399] , \modmult_1/xin[398] , \modmult_1/xin[397] ,
         \modmult_1/xin[396] , \modmult_1/xin[395] , \modmult_1/xin[394] ,
         \modmult_1/xin[393] , \modmult_1/xin[392] , \modmult_1/xin[391] ,
         \modmult_1/xin[390] , \modmult_1/xin[389] , \modmult_1/xin[388] ,
         \modmult_1/xin[387] , \modmult_1/xin[386] , \modmult_1/xin[385] ,
         \modmult_1/xin[384] , \modmult_1/xin[383] , \modmult_1/xin[382] ,
         \modmult_1/xin[381] , \modmult_1/xin[380] , \modmult_1/xin[379] ,
         \modmult_1/xin[378] , \modmult_1/xin[377] , \modmult_1/xin[376] ,
         \modmult_1/xin[375] , \modmult_1/xin[374] , \modmult_1/xin[373] ,
         \modmult_1/xin[372] , \modmult_1/xin[371] , \modmult_1/xin[370] ,
         \modmult_1/xin[369] , \modmult_1/xin[368] , \modmult_1/xin[367] ,
         \modmult_1/xin[366] , \modmult_1/xin[365] , \modmult_1/xin[364] ,
         \modmult_1/xin[363] , \modmult_1/xin[362] , \modmult_1/xin[361] ,
         \modmult_1/xin[360] , \modmult_1/xin[359] , \modmult_1/xin[358] ,
         \modmult_1/xin[357] , \modmult_1/xin[356] , \modmult_1/xin[355] ,
         \modmult_1/xin[354] , \modmult_1/xin[353] , \modmult_1/xin[352] ,
         \modmult_1/xin[351] , \modmult_1/xin[350] , \modmult_1/xin[349] ,
         \modmult_1/xin[348] , \modmult_1/xin[347] , \modmult_1/xin[346] ,
         \modmult_1/xin[345] , \modmult_1/xin[344] , \modmult_1/xin[343] ,
         \modmult_1/xin[342] , \modmult_1/xin[341] , \modmult_1/xin[340] ,
         \modmult_1/xin[339] , \modmult_1/xin[338] , \modmult_1/xin[337] ,
         \modmult_1/xin[336] , \modmult_1/xin[335] , \modmult_1/xin[334] ,
         \modmult_1/xin[333] , \modmult_1/xin[332] , \modmult_1/xin[331] ,
         \modmult_1/xin[330] , \modmult_1/xin[329] , \modmult_1/xin[328] ,
         \modmult_1/xin[327] , \modmult_1/xin[326] , \modmult_1/xin[325] ,
         \modmult_1/xin[324] , \modmult_1/xin[323] , \modmult_1/xin[322] ,
         \modmult_1/xin[321] , \modmult_1/xin[320] , \modmult_1/xin[319] ,
         \modmult_1/xin[318] , \modmult_1/xin[317] , \modmult_1/xin[316] ,
         \modmult_1/xin[315] , \modmult_1/xin[314] , \modmult_1/xin[313] ,
         \modmult_1/xin[312] , \modmult_1/xin[311] , \modmult_1/xin[310] ,
         \modmult_1/xin[309] , \modmult_1/xin[308] , \modmult_1/xin[307] ,
         \modmult_1/xin[306] , \modmult_1/xin[305] , \modmult_1/xin[304] ,
         \modmult_1/xin[303] , \modmult_1/xin[302] , \modmult_1/xin[301] ,
         \modmult_1/xin[300] , \modmult_1/xin[299] , \modmult_1/xin[298] ,
         \modmult_1/xin[297] , \modmult_1/xin[296] , \modmult_1/xin[295] ,
         \modmult_1/xin[294] , \modmult_1/xin[293] , \modmult_1/xin[292] ,
         \modmult_1/xin[291] , \modmult_1/xin[290] , \modmult_1/xin[289] ,
         \modmult_1/xin[288] , \modmult_1/xin[287] , \modmult_1/xin[286] ,
         \modmult_1/xin[285] , \modmult_1/xin[284] , \modmult_1/xin[283] ,
         \modmult_1/xin[282] , \modmult_1/xin[281] , \modmult_1/xin[280] ,
         \modmult_1/xin[279] , \modmult_1/xin[278] , \modmult_1/xin[277] ,
         \modmult_1/xin[276] , \modmult_1/xin[275] , \modmult_1/xin[274] ,
         \modmult_1/xin[273] , \modmult_1/xin[272] , \modmult_1/xin[271] ,
         \modmult_1/xin[270] , \modmult_1/xin[269] , \modmult_1/xin[268] ,
         \modmult_1/xin[267] , \modmult_1/xin[266] , \modmult_1/xin[265] ,
         \modmult_1/xin[264] , \modmult_1/xin[263] , \modmult_1/xin[262] ,
         \modmult_1/xin[261] , \modmult_1/xin[260] , \modmult_1/xin[259] ,
         \modmult_1/xin[258] , \modmult_1/xin[257] , \modmult_1/xin[256] ,
         \modmult_1/xin[255] , \modmult_1/xin[254] , \modmult_1/xin[253] ,
         \modmult_1/xin[252] , \modmult_1/xin[251] , \modmult_1/xin[250] ,
         \modmult_1/xin[249] , \modmult_1/xin[248] , \modmult_1/xin[247] ,
         \modmult_1/xin[246] , \modmult_1/xin[245] , \modmult_1/xin[244] ,
         \modmult_1/xin[243] , \modmult_1/xin[242] , \modmult_1/xin[241] ,
         \modmult_1/xin[240] , \modmult_1/xin[239] , \modmult_1/xin[238] ,
         \modmult_1/xin[237] , \modmult_1/xin[236] , \modmult_1/xin[235] ,
         \modmult_1/xin[234] , \modmult_1/xin[233] , \modmult_1/xin[232] ,
         \modmult_1/xin[231] , \modmult_1/xin[230] , \modmult_1/xin[229] ,
         \modmult_1/xin[228] , \modmult_1/xin[227] , \modmult_1/xin[226] ,
         \modmult_1/xin[225] , \modmult_1/xin[224] , \modmult_1/xin[223] ,
         \modmult_1/xin[222] , \modmult_1/xin[221] , \modmult_1/xin[220] ,
         \modmult_1/xin[219] , \modmult_1/xin[218] , \modmult_1/xin[217] ,
         \modmult_1/xin[216] , \modmult_1/xin[215] , \modmult_1/xin[214] ,
         \modmult_1/xin[213] , \modmult_1/xin[212] , \modmult_1/xin[211] ,
         \modmult_1/xin[210] , \modmult_1/xin[209] , \modmult_1/xin[208] ,
         \modmult_1/xin[207] , \modmult_1/xin[206] , \modmult_1/xin[205] ,
         \modmult_1/xin[204] , \modmult_1/xin[203] , \modmult_1/xin[202] ,
         \modmult_1/xin[201] , \modmult_1/xin[200] , \modmult_1/xin[199] ,
         \modmult_1/xin[198] , \modmult_1/xin[197] , \modmult_1/xin[196] ,
         \modmult_1/xin[195] , \modmult_1/xin[194] , \modmult_1/xin[193] ,
         \modmult_1/xin[192] , \modmult_1/xin[191] , \modmult_1/xin[190] ,
         \modmult_1/xin[189] , \modmult_1/xin[188] , \modmult_1/xin[187] ,
         \modmult_1/xin[186] , \modmult_1/xin[185] , \modmult_1/xin[184] ,
         \modmult_1/xin[183] , \modmult_1/xin[182] , \modmult_1/xin[181] ,
         \modmult_1/xin[180] , \modmult_1/xin[179] , \modmult_1/xin[178] ,
         \modmult_1/xin[177] , \modmult_1/xin[176] , \modmult_1/xin[175] ,
         \modmult_1/xin[174] , \modmult_1/xin[173] , \modmult_1/xin[172] ,
         \modmult_1/xin[171] , \modmult_1/xin[170] , \modmult_1/xin[169] ,
         \modmult_1/xin[168] , \modmult_1/xin[167] , \modmult_1/xin[166] ,
         \modmult_1/xin[165] , \modmult_1/xin[164] , \modmult_1/xin[163] ,
         \modmult_1/xin[162] , \modmult_1/xin[161] , \modmult_1/xin[160] ,
         \modmult_1/xin[159] , \modmult_1/xin[158] , \modmult_1/xin[157] ,
         \modmult_1/xin[156] , \modmult_1/xin[155] , \modmult_1/xin[154] ,
         \modmult_1/xin[153] , \modmult_1/xin[152] , \modmult_1/xin[151] ,
         \modmult_1/xin[150] , \modmult_1/xin[149] , \modmult_1/xin[148] ,
         \modmult_1/xin[147] , \modmult_1/xin[146] , \modmult_1/xin[145] ,
         \modmult_1/xin[144] , \modmult_1/xin[143] , \modmult_1/xin[142] ,
         \modmult_1/xin[141] , \modmult_1/xin[140] , \modmult_1/xin[139] ,
         \modmult_1/xin[138] , \modmult_1/xin[137] , \modmult_1/xin[136] ,
         \modmult_1/xin[135] , \modmult_1/xin[134] , \modmult_1/xin[133] ,
         \modmult_1/xin[132] , \modmult_1/xin[131] , \modmult_1/xin[130] ,
         \modmult_1/xin[129] , \modmult_1/xin[128] , \modmult_1/xin[127] ,
         \modmult_1/xin[126] , \modmult_1/xin[125] , \modmult_1/xin[124] ,
         \modmult_1/xin[123] , \modmult_1/xin[122] , \modmult_1/xin[121] ,
         \modmult_1/xin[120] , \modmult_1/xin[119] , \modmult_1/xin[118] ,
         \modmult_1/xin[117] , \modmult_1/xin[116] , \modmult_1/xin[115] ,
         \modmult_1/xin[114] , \modmult_1/xin[113] , \modmult_1/xin[112] ,
         \modmult_1/xin[111] , \modmult_1/xin[110] , \modmult_1/xin[109] ,
         \modmult_1/xin[108] , \modmult_1/xin[107] , \modmult_1/xin[106] ,
         \modmult_1/xin[105] , \modmult_1/xin[104] , \modmult_1/xin[103] ,
         \modmult_1/xin[102] , \modmult_1/xin[101] , \modmult_1/xin[100] ,
         \modmult_1/xin[99] , \modmult_1/xin[98] , \modmult_1/xin[97] ,
         \modmult_1/xin[96] , \modmult_1/xin[95] , \modmult_1/xin[94] ,
         \modmult_1/xin[93] , \modmult_1/xin[92] , \modmult_1/xin[91] ,
         \modmult_1/xin[90] , \modmult_1/xin[89] , \modmult_1/xin[88] ,
         \modmult_1/xin[87] , \modmult_1/xin[86] , \modmult_1/xin[85] ,
         \modmult_1/xin[84] , \modmult_1/xin[83] , \modmult_1/xin[82] ,
         \modmult_1/xin[81] , \modmult_1/xin[80] , \modmult_1/xin[79] ,
         \modmult_1/xin[78] , \modmult_1/xin[77] , \modmult_1/xin[76] ,
         \modmult_1/xin[75] , \modmult_1/xin[74] , \modmult_1/xin[73] ,
         \modmult_1/xin[72] , \modmult_1/xin[71] , \modmult_1/xin[70] ,
         \modmult_1/xin[69] , \modmult_1/xin[68] , \modmult_1/xin[67] ,
         \modmult_1/xin[66] , \modmult_1/xin[65] , \modmult_1/xin[64] ,
         \modmult_1/xin[63] , \modmult_1/xin[62] , \modmult_1/xin[61] ,
         \modmult_1/xin[60] , \modmult_1/xin[59] , \modmult_1/xin[58] ,
         \modmult_1/xin[57] , \modmult_1/xin[56] , \modmult_1/xin[55] ,
         \modmult_1/xin[54] , \modmult_1/xin[53] , \modmult_1/xin[52] ,
         \modmult_1/xin[51] , \modmult_1/xin[50] , \modmult_1/xin[49] ,
         \modmult_1/xin[48] , \modmult_1/xin[47] , \modmult_1/xin[46] ,
         \modmult_1/xin[45] , \modmult_1/xin[44] , \modmult_1/xin[43] ,
         \modmult_1/xin[42] , \modmult_1/xin[41] , \modmult_1/xin[40] ,
         \modmult_1/xin[39] , \modmult_1/xin[38] , \modmult_1/xin[37] ,
         \modmult_1/xin[36] , \modmult_1/xin[35] , \modmult_1/xin[34] ,
         \modmult_1/xin[33] , \modmult_1/xin[32] , \modmult_1/xin[31] ,
         \modmult_1/xin[30] , \modmult_1/xin[29] , \modmult_1/xin[28] ,
         \modmult_1/xin[27] , \modmult_1/xin[26] , \modmult_1/xin[25] ,
         \modmult_1/xin[24] , \modmult_1/xin[23] , \modmult_1/xin[22] ,
         \modmult_1/xin[21] , \modmult_1/xin[20] , \modmult_1/xin[19] ,
         \modmult_1/xin[18] , \modmult_1/xin[17] , \modmult_1/xin[16] ,
         \modmult_1/xin[15] , \modmult_1/xin[14] , \modmult_1/xin[13] ,
         \modmult_1/xin[12] , \modmult_1/xin[11] , \modmult_1/xin[10] ,
         \modmult_1/xin[9] , \modmult_1/xin[8] , \modmult_1/xin[7] ,
         \modmult_1/xin[6] , \modmult_1/xin[5] , \modmult_1/xin[4] ,
         \modmult_1/xin[3] , \modmult_1/xin[2] , \modmult_1/xin[1] ,
         \modmult_1/xin[0] , \modmult_1/zin[0][1024] ,
         \modmult_1/zin[0][1023] , \modmult_1/zin[0][1022] ,
         \modmult_1/zin[0][1021] , \modmult_1/zin[0][1020] ,
         \modmult_1/zin[0][1019] , \modmult_1/zin[0][1018] ,
         \modmult_1/zin[0][1017] , \modmult_1/zin[0][1016] ,
         \modmult_1/zin[0][1015] , \modmult_1/zin[0][1014] ,
         \modmult_1/zin[0][1013] , \modmult_1/zin[0][1012] ,
         \modmult_1/zin[0][1011] , \modmult_1/zin[0][1010] ,
         \modmult_1/zin[0][1009] , \modmult_1/zin[0][1008] ,
         \modmult_1/zin[0][1007] , \modmult_1/zin[0][1006] ,
         \modmult_1/zin[0][1005] , \modmult_1/zin[0][1004] ,
         \modmult_1/zin[0][1003] , \modmult_1/zin[0][1002] ,
         \modmult_1/zin[0][1001] , \modmult_1/zin[0][1000] ,
         \modmult_1/zin[0][999] , \modmult_1/zin[0][998] ,
         \modmult_1/zin[0][997] , \modmult_1/zin[0][996] ,
         \modmult_1/zin[0][995] , \modmult_1/zin[0][994] ,
         \modmult_1/zin[0][993] , \modmult_1/zin[0][992] ,
         \modmult_1/zin[0][991] , \modmult_1/zin[0][990] ,
         \modmult_1/zin[0][989] , \modmult_1/zin[0][988] ,
         \modmult_1/zin[0][987] , \modmult_1/zin[0][986] ,
         \modmult_1/zin[0][985] , \modmult_1/zin[0][984] ,
         \modmult_1/zin[0][983] , \modmult_1/zin[0][982] ,
         \modmult_1/zin[0][981] , \modmult_1/zin[0][980] ,
         \modmult_1/zin[0][979] , \modmult_1/zin[0][978] ,
         \modmult_1/zin[0][977] , \modmult_1/zin[0][976] ,
         \modmult_1/zin[0][975] , \modmult_1/zin[0][974] ,
         \modmult_1/zin[0][973] , \modmult_1/zin[0][972] ,
         \modmult_1/zin[0][971] , \modmult_1/zin[0][970] ,
         \modmult_1/zin[0][969] , \modmult_1/zin[0][968] ,
         \modmult_1/zin[0][967] , \modmult_1/zin[0][966] ,
         \modmult_1/zin[0][965] , \modmult_1/zin[0][964] ,
         \modmult_1/zin[0][963] , \modmult_1/zin[0][962] ,
         \modmult_1/zin[0][961] , \modmult_1/zin[0][960] ,
         \modmult_1/zin[0][959] , \modmult_1/zin[0][958] ,
         \modmult_1/zin[0][957] , \modmult_1/zin[0][956] ,
         \modmult_1/zin[0][955] , \modmult_1/zin[0][954] ,
         \modmult_1/zin[0][953] , \modmult_1/zin[0][952] ,
         \modmult_1/zin[0][951] , \modmult_1/zin[0][950] ,
         \modmult_1/zin[0][949] , \modmult_1/zin[0][948] ,
         \modmult_1/zin[0][947] , \modmult_1/zin[0][946] ,
         \modmult_1/zin[0][945] , \modmult_1/zin[0][944] ,
         \modmult_1/zin[0][943] , \modmult_1/zin[0][942] ,
         \modmult_1/zin[0][941] , \modmult_1/zin[0][940] ,
         \modmult_1/zin[0][939] , \modmult_1/zin[0][938] ,
         \modmult_1/zin[0][937] , \modmult_1/zin[0][936] ,
         \modmult_1/zin[0][935] , \modmult_1/zin[0][934] ,
         \modmult_1/zin[0][933] , \modmult_1/zin[0][932] ,
         \modmult_1/zin[0][931] , \modmult_1/zin[0][930] ,
         \modmult_1/zin[0][929] , \modmult_1/zin[0][928] ,
         \modmult_1/zin[0][927] , \modmult_1/zin[0][926] ,
         \modmult_1/zin[0][925] , \modmult_1/zin[0][924] ,
         \modmult_1/zin[0][923] , \modmult_1/zin[0][922] ,
         \modmult_1/zin[0][921] , \modmult_1/zin[0][920] ,
         \modmult_1/zin[0][919] , \modmult_1/zin[0][918] ,
         \modmult_1/zin[0][917] , \modmult_1/zin[0][916] ,
         \modmult_1/zin[0][915] , \modmult_1/zin[0][914] ,
         \modmult_1/zin[0][913] , \modmult_1/zin[0][912] ,
         \modmult_1/zin[0][911] , \modmult_1/zin[0][910] ,
         \modmult_1/zin[0][909] , \modmult_1/zin[0][908] ,
         \modmult_1/zin[0][907] , \modmult_1/zin[0][906] ,
         \modmult_1/zin[0][905] , \modmult_1/zin[0][904] ,
         \modmult_1/zin[0][903] , \modmult_1/zin[0][902] ,
         \modmult_1/zin[0][901] , \modmult_1/zin[0][900] ,
         \modmult_1/zin[0][899] , \modmult_1/zin[0][898] ,
         \modmult_1/zin[0][897] , \modmult_1/zin[0][896] ,
         \modmult_1/zin[0][895] , \modmult_1/zin[0][894] ,
         \modmult_1/zin[0][893] , \modmult_1/zin[0][892] ,
         \modmult_1/zin[0][891] , \modmult_1/zin[0][890] ,
         \modmult_1/zin[0][889] , \modmult_1/zin[0][888] ,
         \modmult_1/zin[0][887] , \modmult_1/zin[0][886] ,
         \modmult_1/zin[0][885] , \modmult_1/zin[0][884] ,
         \modmult_1/zin[0][883] , \modmult_1/zin[0][882] ,
         \modmult_1/zin[0][881] , \modmult_1/zin[0][880] ,
         \modmult_1/zin[0][879] , \modmult_1/zin[0][878] ,
         \modmult_1/zin[0][877] , \modmult_1/zin[0][876] ,
         \modmult_1/zin[0][875] , \modmult_1/zin[0][874] ,
         \modmult_1/zin[0][873] , \modmult_1/zin[0][872] ,
         \modmult_1/zin[0][871] , \modmult_1/zin[0][870] ,
         \modmult_1/zin[0][869] , \modmult_1/zin[0][868] ,
         \modmult_1/zin[0][867] , \modmult_1/zin[0][866] ,
         \modmult_1/zin[0][865] , \modmult_1/zin[0][864] ,
         \modmult_1/zin[0][863] , \modmult_1/zin[0][862] ,
         \modmult_1/zin[0][861] , \modmult_1/zin[0][860] ,
         \modmult_1/zin[0][859] , \modmult_1/zin[0][858] ,
         \modmult_1/zin[0][857] , \modmult_1/zin[0][856] ,
         \modmult_1/zin[0][855] , \modmult_1/zin[0][854] ,
         \modmult_1/zin[0][853] , \modmult_1/zin[0][852] ,
         \modmult_1/zin[0][851] , \modmult_1/zin[0][850] ,
         \modmult_1/zin[0][849] , \modmult_1/zin[0][848] ,
         \modmult_1/zin[0][847] , \modmult_1/zin[0][846] ,
         \modmult_1/zin[0][845] , \modmult_1/zin[0][844] ,
         \modmult_1/zin[0][843] , \modmult_1/zin[0][842] ,
         \modmult_1/zin[0][841] , \modmult_1/zin[0][840] ,
         \modmult_1/zin[0][839] , \modmult_1/zin[0][838] ,
         \modmult_1/zin[0][837] , \modmult_1/zin[0][836] ,
         \modmult_1/zin[0][835] , \modmult_1/zin[0][834] ,
         \modmult_1/zin[0][833] , \modmult_1/zin[0][832] ,
         \modmult_1/zin[0][831] , \modmult_1/zin[0][830] ,
         \modmult_1/zin[0][829] , \modmult_1/zin[0][828] ,
         \modmult_1/zin[0][827] , \modmult_1/zin[0][826] ,
         \modmult_1/zin[0][825] , \modmult_1/zin[0][824] ,
         \modmult_1/zin[0][823] , \modmult_1/zin[0][822] ,
         \modmult_1/zin[0][821] , \modmult_1/zin[0][820] ,
         \modmult_1/zin[0][819] , \modmult_1/zin[0][818] ,
         \modmult_1/zin[0][817] , \modmult_1/zin[0][816] ,
         \modmult_1/zin[0][815] , \modmult_1/zin[0][814] ,
         \modmult_1/zin[0][813] , \modmult_1/zin[0][812] ,
         \modmult_1/zin[0][811] , \modmult_1/zin[0][810] ,
         \modmult_1/zin[0][809] , \modmult_1/zin[0][808] ,
         \modmult_1/zin[0][807] , \modmult_1/zin[0][806] ,
         \modmult_1/zin[0][805] , \modmult_1/zin[0][804] ,
         \modmult_1/zin[0][803] , \modmult_1/zin[0][802] ,
         \modmult_1/zin[0][801] , \modmult_1/zin[0][800] ,
         \modmult_1/zin[0][799] , \modmult_1/zin[0][798] ,
         \modmult_1/zin[0][797] , \modmult_1/zin[0][796] ,
         \modmult_1/zin[0][795] , \modmult_1/zin[0][794] ,
         \modmult_1/zin[0][793] , \modmult_1/zin[0][792] ,
         \modmult_1/zin[0][791] , \modmult_1/zin[0][790] ,
         \modmult_1/zin[0][789] , \modmult_1/zin[0][788] ,
         \modmult_1/zin[0][787] , \modmult_1/zin[0][786] ,
         \modmult_1/zin[0][785] , \modmult_1/zin[0][784] ,
         \modmult_1/zin[0][783] , \modmult_1/zin[0][782] ,
         \modmult_1/zin[0][781] , \modmult_1/zin[0][780] ,
         \modmult_1/zin[0][779] , \modmult_1/zin[0][778] ,
         \modmult_1/zin[0][777] , \modmult_1/zin[0][776] ,
         \modmult_1/zin[0][775] , \modmult_1/zin[0][774] ,
         \modmult_1/zin[0][773] , \modmult_1/zin[0][772] ,
         \modmult_1/zin[0][771] , \modmult_1/zin[0][770] ,
         \modmult_1/zin[0][769] , \modmult_1/zin[0][768] ,
         \modmult_1/zin[0][767] , \modmult_1/zin[0][766] ,
         \modmult_1/zin[0][765] , \modmult_1/zin[0][764] ,
         \modmult_1/zin[0][763] , \modmult_1/zin[0][762] ,
         \modmult_1/zin[0][761] , \modmult_1/zin[0][760] ,
         \modmult_1/zin[0][759] , \modmult_1/zin[0][758] ,
         \modmult_1/zin[0][757] , \modmult_1/zin[0][756] ,
         \modmult_1/zin[0][755] , \modmult_1/zin[0][754] ,
         \modmult_1/zin[0][753] , \modmult_1/zin[0][752] ,
         \modmult_1/zin[0][751] , \modmult_1/zin[0][750] ,
         \modmult_1/zin[0][749] , \modmult_1/zin[0][748] ,
         \modmult_1/zin[0][747] , \modmult_1/zin[0][746] ,
         \modmult_1/zin[0][745] , \modmult_1/zin[0][744] ,
         \modmult_1/zin[0][743] , \modmult_1/zin[0][742] ,
         \modmult_1/zin[0][741] , \modmult_1/zin[0][740] ,
         \modmult_1/zin[0][739] , \modmult_1/zin[0][738] ,
         \modmult_1/zin[0][737] , \modmult_1/zin[0][736] ,
         \modmult_1/zin[0][735] , \modmult_1/zin[0][734] ,
         \modmult_1/zin[0][733] , \modmult_1/zin[0][732] ,
         \modmult_1/zin[0][731] , \modmult_1/zin[0][730] ,
         \modmult_1/zin[0][729] , \modmult_1/zin[0][728] ,
         \modmult_1/zin[0][727] , \modmult_1/zin[0][726] ,
         \modmult_1/zin[0][725] , \modmult_1/zin[0][724] ,
         \modmult_1/zin[0][723] , \modmult_1/zin[0][722] ,
         \modmult_1/zin[0][721] , \modmult_1/zin[0][720] ,
         \modmult_1/zin[0][719] , \modmult_1/zin[0][718] ,
         \modmult_1/zin[0][717] , \modmult_1/zin[0][716] ,
         \modmult_1/zin[0][715] , \modmult_1/zin[0][714] ,
         \modmult_1/zin[0][713] , \modmult_1/zin[0][712] ,
         \modmult_1/zin[0][711] , \modmult_1/zin[0][710] ,
         \modmult_1/zin[0][709] , \modmult_1/zin[0][708] ,
         \modmult_1/zin[0][707] , \modmult_1/zin[0][706] ,
         \modmult_1/zin[0][705] , \modmult_1/zin[0][704] ,
         \modmult_1/zin[0][703] , \modmult_1/zin[0][702] ,
         \modmult_1/zin[0][701] , \modmult_1/zin[0][700] ,
         \modmult_1/zin[0][699] , \modmult_1/zin[0][698] ,
         \modmult_1/zin[0][697] , \modmult_1/zin[0][696] ,
         \modmult_1/zin[0][695] , \modmult_1/zin[0][694] ,
         \modmult_1/zin[0][693] , \modmult_1/zin[0][692] ,
         \modmult_1/zin[0][691] , \modmult_1/zin[0][690] ,
         \modmult_1/zin[0][689] , \modmult_1/zin[0][688] ,
         \modmult_1/zin[0][687] , \modmult_1/zin[0][686] ,
         \modmult_1/zin[0][685] , \modmult_1/zin[0][684] ,
         \modmult_1/zin[0][683] , \modmult_1/zin[0][682] ,
         \modmult_1/zin[0][681] , \modmult_1/zin[0][680] ,
         \modmult_1/zin[0][679] , \modmult_1/zin[0][678] ,
         \modmult_1/zin[0][677] , \modmult_1/zin[0][676] ,
         \modmult_1/zin[0][675] , \modmult_1/zin[0][674] ,
         \modmult_1/zin[0][673] , \modmult_1/zin[0][672] ,
         \modmult_1/zin[0][671] , \modmult_1/zin[0][670] ,
         \modmult_1/zin[0][669] , \modmult_1/zin[0][668] ,
         \modmult_1/zin[0][667] , \modmult_1/zin[0][666] ,
         \modmult_1/zin[0][665] , \modmult_1/zin[0][664] ,
         \modmult_1/zin[0][663] , \modmult_1/zin[0][662] ,
         \modmult_1/zin[0][661] , \modmult_1/zin[0][660] ,
         \modmult_1/zin[0][659] , \modmult_1/zin[0][658] ,
         \modmult_1/zin[0][657] , \modmult_1/zin[0][656] ,
         \modmult_1/zin[0][655] , \modmult_1/zin[0][654] ,
         \modmult_1/zin[0][653] , \modmult_1/zin[0][652] ,
         \modmult_1/zin[0][651] , \modmult_1/zin[0][650] ,
         \modmult_1/zin[0][649] , \modmult_1/zin[0][648] ,
         \modmult_1/zin[0][647] , \modmult_1/zin[0][646] ,
         \modmult_1/zin[0][645] , \modmult_1/zin[0][644] ,
         \modmult_1/zin[0][643] , \modmult_1/zin[0][642] ,
         \modmult_1/zin[0][641] , \modmult_1/zin[0][640] ,
         \modmult_1/zin[0][639] , \modmult_1/zin[0][638] ,
         \modmult_1/zin[0][637] , \modmult_1/zin[0][636] ,
         \modmult_1/zin[0][635] , \modmult_1/zin[0][634] ,
         \modmult_1/zin[0][633] , \modmult_1/zin[0][632] ,
         \modmult_1/zin[0][631] , \modmult_1/zin[0][630] ,
         \modmult_1/zin[0][629] , \modmult_1/zin[0][628] ,
         \modmult_1/zin[0][627] , \modmult_1/zin[0][626] ,
         \modmult_1/zin[0][625] , \modmult_1/zin[0][624] ,
         \modmult_1/zin[0][623] , \modmult_1/zin[0][622] ,
         \modmult_1/zin[0][621] , \modmult_1/zin[0][620] ,
         \modmult_1/zin[0][619] , \modmult_1/zin[0][618] ,
         \modmult_1/zin[0][617] , \modmult_1/zin[0][616] ,
         \modmult_1/zin[0][615] , \modmult_1/zin[0][614] ,
         \modmult_1/zin[0][613] , \modmult_1/zin[0][612] ,
         \modmult_1/zin[0][611] , \modmult_1/zin[0][610] ,
         \modmult_1/zin[0][609] , \modmult_1/zin[0][608] ,
         \modmult_1/zin[0][607] , \modmult_1/zin[0][606] ,
         \modmult_1/zin[0][605] , \modmult_1/zin[0][604] ,
         \modmult_1/zin[0][603] , \modmult_1/zin[0][602] ,
         \modmult_1/zin[0][601] , \modmult_1/zin[0][600] ,
         \modmult_1/zin[0][599] , \modmult_1/zin[0][598] ,
         \modmult_1/zin[0][597] , \modmult_1/zin[0][596] ,
         \modmult_1/zin[0][595] , \modmult_1/zin[0][594] ,
         \modmult_1/zin[0][593] , \modmult_1/zin[0][592] ,
         \modmult_1/zin[0][591] , \modmult_1/zin[0][590] ,
         \modmult_1/zin[0][589] , \modmult_1/zin[0][588] ,
         \modmult_1/zin[0][587] , \modmult_1/zin[0][586] ,
         \modmult_1/zin[0][585] , \modmult_1/zin[0][584] ,
         \modmult_1/zin[0][583] , \modmult_1/zin[0][582] ,
         \modmult_1/zin[0][581] , \modmult_1/zin[0][580] ,
         \modmult_1/zin[0][579] , \modmult_1/zin[0][578] ,
         \modmult_1/zin[0][577] , \modmult_1/zin[0][576] ,
         \modmult_1/zin[0][575] , \modmult_1/zin[0][574] ,
         \modmult_1/zin[0][573] , \modmult_1/zin[0][572] ,
         \modmult_1/zin[0][571] , \modmult_1/zin[0][570] ,
         \modmult_1/zin[0][569] , \modmult_1/zin[0][568] ,
         \modmult_1/zin[0][567] , \modmult_1/zin[0][566] ,
         \modmult_1/zin[0][565] , \modmult_1/zin[0][564] ,
         \modmult_1/zin[0][563] , \modmult_1/zin[0][562] ,
         \modmult_1/zin[0][561] , \modmult_1/zin[0][560] ,
         \modmult_1/zin[0][559] , \modmult_1/zin[0][558] ,
         \modmult_1/zin[0][557] , \modmult_1/zin[0][556] ,
         \modmult_1/zin[0][555] , \modmult_1/zin[0][554] ,
         \modmult_1/zin[0][553] , \modmult_1/zin[0][552] ,
         \modmult_1/zin[0][551] , \modmult_1/zin[0][550] ,
         \modmult_1/zin[0][549] , \modmult_1/zin[0][548] ,
         \modmult_1/zin[0][547] , \modmult_1/zin[0][546] ,
         \modmult_1/zin[0][545] , \modmult_1/zin[0][544] ,
         \modmult_1/zin[0][543] , \modmult_1/zin[0][542] ,
         \modmult_1/zin[0][541] , \modmult_1/zin[0][540] ,
         \modmult_1/zin[0][539] , \modmult_1/zin[0][538] ,
         \modmult_1/zin[0][537] , \modmult_1/zin[0][536] ,
         \modmult_1/zin[0][535] , \modmult_1/zin[0][534] ,
         \modmult_1/zin[0][533] , \modmult_1/zin[0][532] ,
         \modmult_1/zin[0][531] , \modmult_1/zin[0][530] ,
         \modmult_1/zin[0][529] , \modmult_1/zin[0][528] ,
         \modmult_1/zin[0][527] , \modmult_1/zin[0][526] ,
         \modmult_1/zin[0][525] , \modmult_1/zin[0][524] ,
         \modmult_1/zin[0][523] , \modmult_1/zin[0][522] ,
         \modmult_1/zin[0][521] , \modmult_1/zin[0][520] ,
         \modmult_1/zin[0][519] , \modmult_1/zin[0][518] ,
         \modmult_1/zin[0][517] , \modmult_1/zin[0][516] ,
         \modmult_1/zin[0][515] , \modmult_1/zin[0][514] ,
         \modmult_1/zin[0][513] , \modmult_1/zin[0][512] ,
         \modmult_1/zin[0][511] , \modmult_1/zin[0][510] ,
         \modmult_1/zin[0][509] , \modmult_1/zin[0][508] ,
         \modmult_1/zin[0][507] , \modmult_1/zin[0][506] ,
         \modmult_1/zin[0][505] , \modmult_1/zin[0][504] ,
         \modmult_1/zin[0][503] , \modmult_1/zin[0][502] ,
         \modmult_1/zin[0][501] , \modmult_1/zin[0][500] ,
         \modmult_1/zin[0][499] , \modmult_1/zin[0][498] ,
         \modmult_1/zin[0][497] , \modmult_1/zin[0][496] ,
         \modmult_1/zin[0][495] , \modmult_1/zin[0][494] ,
         \modmult_1/zin[0][493] , \modmult_1/zin[0][492] ,
         \modmult_1/zin[0][491] , \modmult_1/zin[0][490] ,
         \modmult_1/zin[0][489] , \modmult_1/zin[0][488] ,
         \modmult_1/zin[0][487] , \modmult_1/zin[0][486] ,
         \modmult_1/zin[0][485] , \modmult_1/zin[0][484] ,
         \modmult_1/zin[0][483] , \modmult_1/zin[0][482] ,
         \modmult_1/zin[0][481] , \modmult_1/zin[0][480] ,
         \modmult_1/zin[0][479] , \modmult_1/zin[0][478] ,
         \modmult_1/zin[0][477] , \modmult_1/zin[0][476] ,
         \modmult_1/zin[0][475] , \modmult_1/zin[0][474] ,
         \modmult_1/zin[0][473] , \modmult_1/zin[0][472] ,
         \modmult_1/zin[0][471] , \modmult_1/zin[0][470] ,
         \modmult_1/zin[0][469] , \modmult_1/zin[0][468] ,
         \modmult_1/zin[0][467] , \modmult_1/zin[0][466] ,
         \modmult_1/zin[0][465] , \modmult_1/zin[0][464] ,
         \modmult_1/zin[0][463] , \modmult_1/zin[0][462] ,
         \modmult_1/zin[0][461] , \modmult_1/zin[0][460] ,
         \modmult_1/zin[0][459] , \modmult_1/zin[0][458] ,
         \modmult_1/zin[0][457] , \modmult_1/zin[0][456] ,
         \modmult_1/zin[0][455] , \modmult_1/zin[0][454] ,
         \modmult_1/zin[0][453] , \modmult_1/zin[0][452] ,
         \modmult_1/zin[0][451] , \modmult_1/zin[0][450] ,
         \modmult_1/zin[0][449] , \modmult_1/zin[0][448] ,
         \modmult_1/zin[0][447] , \modmult_1/zin[0][446] ,
         \modmult_1/zin[0][445] , \modmult_1/zin[0][444] ,
         \modmult_1/zin[0][443] , \modmult_1/zin[0][442] ,
         \modmult_1/zin[0][441] , \modmult_1/zin[0][440] ,
         \modmult_1/zin[0][439] , \modmult_1/zin[0][438] ,
         \modmult_1/zin[0][437] , \modmult_1/zin[0][436] ,
         \modmult_1/zin[0][435] , \modmult_1/zin[0][434] ,
         \modmult_1/zin[0][433] , \modmult_1/zin[0][432] ,
         \modmult_1/zin[0][431] , \modmult_1/zin[0][430] ,
         \modmult_1/zin[0][429] , \modmult_1/zin[0][428] ,
         \modmult_1/zin[0][427] , \modmult_1/zin[0][426] ,
         \modmult_1/zin[0][425] , \modmult_1/zin[0][424] ,
         \modmult_1/zin[0][423] , \modmult_1/zin[0][422] ,
         \modmult_1/zin[0][421] , \modmult_1/zin[0][420] ,
         \modmult_1/zin[0][419] , \modmult_1/zin[0][418] ,
         \modmult_1/zin[0][417] , \modmult_1/zin[0][416] ,
         \modmult_1/zin[0][415] , \modmult_1/zin[0][414] ,
         \modmult_1/zin[0][413] , \modmult_1/zin[0][412] ,
         \modmult_1/zin[0][411] , \modmult_1/zin[0][410] ,
         \modmult_1/zin[0][409] , \modmult_1/zin[0][408] ,
         \modmult_1/zin[0][407] , \modmult_1/zin[0][406] ,
         \modmult_1/zin[0][405] , \modmult_1/zin[0][404] ,
         \modmult_1/zin[0][403] , \modmult_1/zin[0][402] ,
         \modmult_1/zin[0][401] , \modmult_1/zin[0][400] ,
         \modmult_1/zin[0][399] , \modmult_1/zin[0][398] ,
         \modmult_1/zin[0][397] , \modmult_1/zin[0][396] ,
         \modmult_1/zin[0][395] , \modmult_1/zin[0][394] ,
         \modmult_1/zin[0][393] , \modmult_1/zin[0][392] ,
         \modmult_1/zin[0][391] , \modmult_1/zin[0][390] ,
         \modmult_1/zin[0][389] , \modmult_1/zin[0][388] ,
         \modmult_1/zin[0][387] , \modmult_1/zin[0][386] ,
         \modmult_1/zin[0][385] , \modmult_1/zin[0][384] ,
         \modmult_1/zin[0][383] , \modmult_1/zin[0][382] ,
         \modmult_1/zin[0][381] , \modmult_1/zin[0][380] ,
         \modmult_1/zin[0][379] , \modmult_1/zin[0][378] ,
         \modmult_1/zin[0][377] , \modmult_1/zin[0][376] ,
         \modmult_1/zin[0][375] , \modmult_1/zin[0][374] ,
         \modmult_1/zin[0][373] , \modmult_1/zin[0][372] ,
         \modmult_1/zin[0][371] , \modmult_1/zin[0][370] ,
         \modmult_1/zin[0][369] , \modmult_1/zin[0][368] ,
         \modmult_1/zin[0][367] , \modmult_1/zin[0][366] ,
         \modmult_1/zin[0][365] , \modmult_1/zin[0][364] ,
         \modmult_1/zin[0][363] , \modmult_1/zin[0][362] ,
         \modmult_1/zin[0][361] , \modmult_1/zin[0][360] ,
         \modmult_1/zin[0][359] , \modmult_1/zin[0][358] ,
         \modmult_1/zin[0][357] , \modmult_1/zin[0][356] ,
         \modmult_1/zin[0][355] , \modmult_1/zin[0][354] ,
         \modmult_1/zin[0][353] , \modmult_1/zin[0][352] ,
         \modmult_1/zin[0][351] , \modmult_1/zin[0][350] ,
         \modmult_1/zin[0][349] , \modmult_1/zin[0][348] ,
         \modmult_1/zin[0][347] , \modmult_1/zin[0][346] ,
         \modmult_1/zin[0][345] , \modmult_1/zin[0][344] ,
         \modmult_1/zin[0][343] , \modmult_1/zin[0][342] ,
         \modmult_1/zin[0][341] , \modmult_1/zin[0][340] ,
         \modmult_1/zin[0][339] , \modmult_1/zin[0][338] ,
         \modmult_1/zin[0][337] , \modmult_1/zin[0][336] ,
         \modmult_1/zin[0][335] , \modmult_1/zin[0][334] ,
         \modmult_1/zin[0][333] , \modmult_1/zin[0][332] ,
         \modmult_1/zin[0][331] , \modmult_1/zin[0][330] ,
         \modmult_1/zin[0][329] , \modmult_1/zin[0][328] ,
         \modmult_1/zin[0][327] , \modmult_1/zin[0][326] ,
         \modmult_1/zin[0][325] , \modmult_1/zin[0][324] ,
         \modmult_1/zin[0][323] , \modmult_1/zin[0][322] ,
         \modmult_1/zin[0][321] , \modmult_1/zin[0][320] ,
         \modmult_1/zin[0][319] , \modmult_1/zin[0][318] ,
         \modmult_1/zin[0][317] , \modmult_1/zin[0][316] ,
         \modmult_1/zin[0][315] , \modmult_1/zin[0][314] ,
         \modmult_1/zin[0][313] , \modmult_1/zin[0][312] ,
         \modmult_1/zin[0][311] , \modmult_1/zin[0][310] ,
         \modmult_1/zin[0][309] , \modmult_1/zin[0][308] ,
         \modmult_1/zin[0][307] , \modmult_1/zin[0][306] ,
         \modmult_1/zin[0][305] , \modmult_1/zin[0][304] ,
         \modmult_1/zin[0][303] , \modmult_1/zin[0][302] ,
         \modmult_1/zin[0][301] , \modmult_1/zin[0][300] ,
         \modmult_1/zin[0][299] , \modmult_1/zin[0][298] ,
         \modmult_1/zin[0][297] , \modmult_1/zin[0][296] ,
         \modmult_1/zin[0][295] , \modmult_1/zin[0][294] ,
         \modmult_1/zin[0][293] , \modmult_1/zin[0][292] ,
         \modmult_1/zin[0][291] , \modmult_1/zin[0][290] ,
         \modmult_1/zin[0][289] , \modmult_1/zin[0][288] ,
         \modmult_1/zin[0][287] , \modmult_1/zin[0][286] ,
         \modmult_1/zin[0][285] , \modmult_1/zin[0][284] ,
         \modmult_1/zin[0][283] , \modmult_1/zin[0][282] ,
         \modmult_1/zin[0][281] , \modmult_1/zin[0][280] ,
         \modmult_1/zin[0][279] , \modmult_1/zin[0][278] ,
         \modmult_1/zin[0][277] , \modmult_1/zin[0][276] ,
         \modmult_1/zin[0][275] , \modmult_1/zin[0][274] ,
         \modmult_1/zin[0][273] , \modmult_1/zin[0][272] ,
         \modmult_1/zin[0][271] , \modmult_1/zin[0][270] ,
         \modmult_1/zin[0][269] , \modmult_1/zin[0][268] ,
         \modmult_1/zin[0][267] , \modmult_1/zin[0][266] ,
         \modmult_1/zin[0][265] , \modmult_1/zin[0][264] ,
         \modmult_1/zin[0][263] , \modmult_1/zin[0][262] ,
         \modmult_1/zin[0][261] , \modmult_1/zin[0][260] ,
         \modmult_1/zin[0][259] , \modmult_1/zin[0][258] ,
         \modmult_1/zin[0][257] , \modmult_1/zin[0][256] ,
         \modmult_1/zin[0][255] , \modmult_1/zin[0][254] ,
         \modmult_1/zin[0][253] , \modmult_1/zin[0][252] ,
         \modmult_1/zin[0][251] , \modmult_1/zin[0][250] ,
         \modmult_1/zin[0][249] , \modmult_1/zin[0][248] ,
         \modmult_1/zin[0][247] , \modmult_1/zin[0][246] ,
         \modmult_1/zin[0][245] , \modmult_1/zin[0][244] ,
         \modmult_1/zin[0][243] , \modmult_1/zin[0][242] ,
         \modmult_1/zin[0][241] , \modmult_1/zin[0][240] ,
         \modmult_1/zin[0][239] , \modmult_1/zin[0][238] ,
         \modmult_1/zin[0][237] , \modmult_1/zin[0][236] ,
         \modmult_1/zin[0][235] , \modmult_1/zin[0][234] ,
         \modmult_1/zin[0][233] , \modmult_1/zin[0][232] ,
         \modmult_1/zin[0][231] , \modmult_1/zin[0][230] ,
         \modmult_1/zin[0][229] , \modmult_1/zin[0][228] ,
         \modmult_1/zin[0][227] , \modmult_1/zin[0][226] ,
         \modmult_1/zin[0][225] , \modmult_1/zin[0][224] ,
         \modmult_1/zin[0][223] , \modmult_1/zin[0][222] ,
         \modmult_1/zin[0][221] , \modmult_1/zin[0][220] ,
         \modmult_1/zin[0][219] , \modmult_1/zin[0][218] ,
         \modmult_1/zin[0][217] , \modmult_1/zin[0][216] ,
         \modmult_1/zin[0][215] , \modmult_1/zin[0][214] ,
         \modmult_1/zin[0][213] , \modmult_1/zin[0][212] ,
         \modmult_1/zin[0][211] , \modmult_1/zin[0][210] ,
         \modmult_1/zin[0][209] , \modmult_1/zin[0][208] ,
         \modmult_1/zin[0][207] , \modmult_1/zin[0][206] ,
         \modmult_1/zin[0][205] , \modmult_1/zin[0][204] ,
         \modmult_1/zin[0][203] , \modmult_1/zin[0][202] ,
         \modmult_1/zin[0][201] , \modmult_1/zin[0][200] ,
         \modmult_1/zin[0][199] , \modmult_1/zin[0][198] ,
         \modmult_1/zin[0][197] , \modmult_1/zin[0][196] ,
         \modmult_1/zin[0][195] , \modmult_1/zin[0][194] ,
         \modmult_1/zin[0][193] , \modmult_1/zin[0][192] ,
         \modmult_1/zin[0][191] , \modmult_1/zin[0][190] ,
         \modmult_1/zin[0][189] , \modmult_1/zin[0][188] ,
         \modmult_1/zin[0][187] , \modmult_1/zin[0][186] ,
         \modmult_1/zin[0][185] , \modmult_1/zin[0][184] ,
         \modmult_1/zin[0][183] , \modmult_1/zin[0][182] ,
         \modmult_1/zin[0][181] , \modmult_1/zin[0][180] ,
         \modmult_1/zin[0][179] , \modmult_1/zin[0][178] ,
         \modmult_1/zin[0][177] , \modmult_1/zin[0][176] ,
         \modmult_1/zin[0][175] , \modmult_1/zin[0][174] ,
         \modmult_1/zin[0][173] , \modmult_1/zin[0][172] ,
         \modmult_1/zin[0][171] , \modmult_1/zin[0][170] ,
         \modmult_1/zin[0][169] , \modmult_1/zin[0][168] ,
         \modmult_1/zin[0][167] , \modmult_1/zin[0][166] ,
         \modmult_1/zin[0][165] , \modmult_1/zin[0][164] ,
         \modmult_1/zin[0][163] , \modmult_1/zin[0][162] ,
         \modmult_1/zin[0][161] , \modmult_1/zin[0][160] ,
         \modmult_1/zin[0][159] , \modmult_1/zin[0][158] ,
         \modmult_1/zin[0][157] , \modmult_1/zin[0][156] ,
         \modmult_1/zin[0][155] , \modmult_1/zin[0][154] ,
         \modmult_1/zin[0][153] , \modmult_1/zin[0][152] ,
         \modmult_1/zin[0][151] , \modmult_1/zin[0][150] ,
         \modmult_1/zin[0][149] , \modmult_1/zin[0][148] ,
         \modmult_1/zin[0][147] , \modmult_1/zin[0][146] ,
         \modmult_1/zin[0][145] , \modmult_1/zin[0][144] ,
         \modmult_1/zin[0][143] , \modmult_1/zin[0][142] ,
         \modmult_1/zin[0][141] , \modmult_1/zin[0][140] ,
         \modmult_1/zin[0][139] , \modmult_1/zin[0][138] ,
         \modmult_1/zin[0][137] , \modmult_1/zin[0][136] ,
         \modmult_1/zin[0][135] , \modmult_1/zin[0][134] ,
         \modmult_1/zin[0][133] , \modmult_1/zin[0][132] ,
         \modmult_1/zin[0][131] , \modmult_1/zin[0][130] ,
         \modmult_1/zin[0][129] , \modmult_1/zin[0][128] ,
         \modmult_1/zin[0][127] , \modmult_1/zin[0][126] ,
         \modmult_1/zin[0][125] , \modmult_1/zin[0][124] ,
         \modmult_1/zin[0][123] , \modmult_1/zin[0][122] ,
         \modmult_1/zin[0][121] , \modmult_1/zin[0][120] ,
         \modmult_1/zin[0][119] , \modmult_1/zin[0][118] ,
         \modmult_1/zin[0][117] , \modmult_1/zin[0][116] ,
         \modmult_1/zin[0][115] , \modmult_1/zin[0][114] ,
         \modmult_1/zin[0][113] , \modmult_1/zin[0][112] ,
         \modmult_1/zin[0][111] , \modmult_1/zin[0][110] ,
         \modmult_1/zin[0][109] , \modmult_1/zin[0][108] ,
         \modmult_1/zin[0][107] , \modmult_1/zin[0][106] ,
         \modmult_1/zin[0][105] , \modmult_1/zin[0][104] ,
         \modmult_1/zin[0][103] , \modmult_1/zin[0][102] ,
         \modmult_1/zin[0][101] , \modmult_1/zin[0][100] ,
         \modmult_1/zin[0][99] , \modmult_1/zin[0][98] ,
         \modmult_1/zin[0][97] , \modmult_1/zin[0][96] ,
         \modmult_1/zin[0][95] , \modmult_1/zin[0][94] ,
         \modmult_1/zin[0][93] , \modmult_1/zin[0][92] ,
         \modmult_1/zin[0][91] , \modmult_1/zin[0][90] ,
         \modmult_1/zin[0][89] , \modmult_1/zin[0][88] ,
         \modmult_1/zin[0][87] , \modmult_1/zin[0][86] ,
         \modmult_1/zin[0][85] , \modmult_1/zin[0][84] ,
         \modmult_1/zin[0][83] , \modmult_1/zin[0][82] ,
         \modmult_1/zin[0][81] , \modmult_1/zin[0][80] ,
         \modmult_1/zin[0][79] , \modmult_1/zin[0][78] ,
         \modmult_1/zin[0][77] , \modmult_1/zin[0][76] ,
         \modmult_1/zin[0][75] , \modmult_1/zin[0][74] ,
         \modmult_1/zin[0][73] , \modmult_1/zin[0][72] ,
         \modmult_1/zin[0][71] , \modmult_1/zin[0][70] ,
         \modmult_1/zin[0][69] , \modmult_1/zin[0][68] ,
         \modmult_1/zin[0][67] , \modmult_1/zin[0][66] ,
         \modmult_1/zin[0][65] , \modmult_1/zin[0][64] ,
         \modmult_1/zin[0][63] , \modmult_1/zin[0][62] ,
         \modmult_1/zin[0][61] , \modmult_1/zin[0][60] ,
         \modmult_1/zin[0][59] , \modmult_1/zin[0][58] ,
         \modmult_1/zin[0][57] , \modmult_1/zin[0][56] ,
         \modmult_1/zin[0][55] , \modmult_1/zin[0][54] ,
         \modmult_1/zin[0][53] , \modmult_1/zin[0][52] ,
         \modmult_1/zin[0][51] , \modmult_1/zin[0][50] ,
         \modmult_1/zin[0][49] , \modmult_1/zin[0][48] ,
         \modmult_1/zin[0][47] , \modmult_1/zin[0][46] ,
         \modmult_1/zin[0][45] , \modmult_1/zin[0][44] ,
         \modmult_1/zin[0][43] , \modmult_1/zin[0][42] ,
         \modmult_1/zin[0][41] , \modmult_1/zin[0][40] ,
         \modmult_1/zin[0][39] , \modmult_1/zin[0][38] ,
         \modmult_1/zin[0][37] , \modmult_1/zin[0][36] ,
         \modmult_1/zin[0][35] , \modmult_1/zin[0][34] ,
         \modmult_1/zin[0][33] , \modmult_1/zin[0][32] ,
         \modmult_1/zin[0][31] , \modmult_1/zin[0][30] ,
         \modmult_1/zin[0][29] , \modmult_1/zin[0][28] ,
         \modmult_1/zin[0][27] , \modmult_1/zin[0][26] ,
         \modmult_1/zin[0][25] , \modmult_1/zin[0][24] ,
         \modmult_1/zin[0][23] , \modmult_1/zin[0][22] ,
         \modmult_1/zin[0][21] , \modmult_1/zin[0][20] ,
         \modmult_1/zin[0][19] , \modmult_1/zin[0][18] ,
         \modmult_1/zin[0][17] , \modmult_1/zin[0][16] ,
         \modmult_1/zin[0][15] , \modmult_1/zin[0][14] ,
         \modmult_1/zin[0][13] , \modmult_1/zin[0][12] ,
         \modmult_1/zin[0][11] , \modmult_1/zin[0][10] , \modmult_1/zin[0][9] ,
         \modmult_1/zin[0][8] , \modmult_1/zin[0][7] , \modmult_1/zin[0][6] ,
         \modmult_1/zin[0][5] , \modmult_1/zin[0][4] , \modmult_1/zin[0][3] ,
         \modmult_1/zin[0][2] , \modmult_1/zin[0][1] , \modmult_1/zin[0][0] ,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
         n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313,
         n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
         n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
         n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337,
         n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
         n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
         n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361,
         n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369,
         n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
         n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
         n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
         n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
         n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
         n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
         n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
         n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433,
         n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441,
         n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
         n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
         n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
         n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473,
         n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481,
         n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489,
         n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497,
         n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505,
         n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513,
         n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529,
         n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537,
         n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545,
         n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553,
         n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561,
         n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569,
         n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577,
         n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585,
         n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
         n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601,
         n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609,
         n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617,
         n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625,
         n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633,
         n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641,
         n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649,
         n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657,
         n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665,
         n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673,
         n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681,
         n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689,
         n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697,
         n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705,
         n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713,
         n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721,
         n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729,
         n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737,
         n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745,
         n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753,
         n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761,
         n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769,
         n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777,
         n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785,
         n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793,
         n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801,
         n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
         n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817,
         n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825,
         n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833,
         n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841,
         n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849,
         n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857,
         n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865,
         n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873,
         n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881,
         n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889,
         n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897,
         n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905,
         n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913,
         n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921,
         n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929,
         n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937,
         n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945,
         n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953,
         n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961,
         n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969,
         n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977,
         n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985,
         n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993,
         n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001,
         n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009,
         n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017,
         n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025,
         n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033,
         n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
         n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049,
         n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057,
         n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065,
         n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073,
         n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081,
         n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089,
         n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097,
         n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105,
         n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113,
         n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121,
         n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129,
         n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137,
         n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145,
         n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153,
         n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161,
         n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169,
         n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177,
         n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185,
         n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193,
         n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201,
         n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209,
         n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217,
         n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225,
         n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233,
         n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241,
         n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249,
         n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257,
         n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265,
         n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273,
         n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281,
         n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289,
         n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297,
         n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305,
         n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
         n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321,
         n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329,
         n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337,
         n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345,
         n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353,
         n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361,
         n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369,
         n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377,
         n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385,
         n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393,
         n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401,
         n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409,
         n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417,
         n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425,
         n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433,
         n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441,
         n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449,
         n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457,
         n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465,
         n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473,
         n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481,
         n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489,
         n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497,
         n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505,
         n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513,
         n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521,
         n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529,
         n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537,
         n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545,
         n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553,
         n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561,
         n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569,
         n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577,
         n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585,
         n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593,
         n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601,
         n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609,
         n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617,
         n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625,
         n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633,
         n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641,
         n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649,
         n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657,
         n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665,
         n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673,
         n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681,
         n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689,
         n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697,
         n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705,
         n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713,
         n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721,
         n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729,
         n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737,
         n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745,
         n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753,
         n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761,
         n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769,
         n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777,
         n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785,
         n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793,
         n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801,
         n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809,
         n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817,
         n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825,
         n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833,
         n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841,
         n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849,
         n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857,
         n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865,
         n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873,
         n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881,
         n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889,
         n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897,
         n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905,
         n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913,
         n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921,
         n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929,
         n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937,
         n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945,
         n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953,
         n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961,
         n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969,
         n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977,
         n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985,
         n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993,
         n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001,
         n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009,
         n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017,
         n40018, n40019, n40020, n40021, n40022, n40023, n40024, n40025,
         n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033,
         n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041,
         n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049,
         n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057,
         n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065,
         n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073,
         n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081,
         n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089,
         n40090, n40091, n40092, n40093, n40094, n40095, n40096, n40097,
         n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105,
         n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113,
         n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121,
         n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129,
         n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137,
         n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145,
         n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153,
         n40154, n40155, n40156, n40157, n40158, n40159, n40160, n40161,
         n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169,
         n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177,
         n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185,
         n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
         n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201,
         n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209,
         n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217,
         n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225,
         n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233,
         n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241,
         n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249,
         n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257,
         n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265,
         n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273,
         n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281,
         n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289,
         n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297,
         n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305,
         n40306, n40307, n40308, n40309, n40310, n40311, n40312, n40313,
         n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321,
         n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329,
         n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337,
         n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345,
         n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353,
         n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361,
         n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369,
         n40370, n40371, n40372, n40373, n40374, n40375, n40376, n40377,
         n40378, n40379, n40380, n40381, n40382, n40383, n40384, n40385,
         n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393,
         n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401,
         n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409,
         n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417,
         n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425,
         n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433,
         n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441,
         n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449,
         n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457,
         n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465,
         n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473,
         n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481,
         n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489,
         n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497,
         n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505,
         n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513,
         n40514, n40515, n40516, n40517, n40518, n40519, n40520, n40521,
         n40522, n40523, n40524, n40525, n40526, n40527, n40528, n40529,
         n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537,
         n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545,
         n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553,
         n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561,
         n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569,
         n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577,
         n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585,
         n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593,
         n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601,
         n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609,
         n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617,
         n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625,
         n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633,
         n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641,
         n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649,
         n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657,
         n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665,
         n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673,
         n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681,
         n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689,
         n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697,
         n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705,
         n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713,
         n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721,
         n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729,
         n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737,
         n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745,
         n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753,
         n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761,
         n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769,
         n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777,
         n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785,
         n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793,
         n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801,
         n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809,
         n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817,
         n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825,
         n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833,
         n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841,
         n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849,
         n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857,
         n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865,
         n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873,
         n40874, n40875, n40876, n40877, n40878, n40879, n40880, n40881,
         n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889,
         n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897,
         n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905,
         n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913,
         n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921,
         n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929,
         n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937,
         n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945,
         n40946, n40947, n40948, n40949, n40950, n40951, n40952, n40953,
         n40954, n40955, n40956, n40957, n40958, n40959, n40960, n40961,
         n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969,
         n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977,
         n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985,
         n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993,
         n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001,
         n41002, n41003, n41004, n41005, n41006, n41007, n41008, n41009,
         n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41017,
         n41018, n41019, n41020, n41021, n41022, n41023, n41024, n41025,
         n41026, n41027, n41028, n41029, n41030, n41031, n41032, n41033,
         n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041,
         n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049,
         n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057,
         n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065,
         n41066, n41067, n41068, n41069, n41070, n41071, n41072, n41073,
         n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081,
         n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089,
         n41090, n41091, n41092, n41093, n41094, n41095, n41096, n41097,
         n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105,
         n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113,
         n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121,
         n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129,
         n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137,
         n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145,
         n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153,
         n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161,
         n41162, n41163, n41164, n41165, n41166, n41167, n41168, n41169,
         n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177,
         n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185,
         n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193,
         n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201,
         n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209,
         n41210, n41211, n41212, n41213, n41214, n41215, n41216, n41217,
         n41218, n41219, n41220, n41221, n41222, n41223, n41224, n41225,
         n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233,
         n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241,
         n41242, n41243, n41244, n41245, n41246, n41247, n41248, n41249,
         n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257,
         n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265,
         n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273,
         n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281,
         n41282, n41283, n41284, n41285, n41286, n41287, n41288, n41289,
         n41290, n41291, n41292, n41293, n41294, n41295, n41296, n41297,
         n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305,
         n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313,
         n41314, n41315, n41316, n41317, n41318, n41319, n41320, n41321,
         n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329,
         n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337,
         n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345,
         n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353,
         n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361,
         n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369,
         n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377,
         n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385,
         n41386, n41387, n41388, n41389, n41390, n41391, n41392, n41393,
         n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401,
         n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409,
         n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417,
         n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425,
         n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433,
         n41434, n41435, n41436, n41437, n41438, n41439, n41440, n41441,
         n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449,
         n41450, n41451, n41452, n41453, n41454, n41455, n41456, n41457,
         n41458, n41459, n41460, n41461, n41462, n41463, n41464, n41465,
         n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473,
         n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481,
         n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489,
         n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497,
         n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505,
         n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513,
         n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521,
         n41522, n41523, n41524, n41525, n41526, n41527, n41528, n41529,
         n41530, n41531, n41532, n41533, n41534, n41535, n41536, n41537,
         n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545,
         n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553,
         n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561,
         n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569,
         n41570, n41571, n41572, n41573, n41574, n41575, n41576, n41577,
         n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585,
         n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593,
         n41594, n41595, n41596, n41597, n41598, n41599, n41600, n41601,
         n41602, n41603, n41604, n41605, n41606, n41607, n41608, n41609,
         n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617,
         n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625,
         n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633,
         n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641,
         n41642, n41643, n41644, n41645, n41646, n41647, n41648, n41649,
         n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657,
         n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665,
         n41666, n41667, n41668, n41669, n41670, n41671, n41672, n41673,
         n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41681,
         n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689,
         n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697,
         n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705,
         n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713,
         n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721,
         n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729,
         n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737,
         n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745,
         n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753,
         n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761,
         n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769,
         n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777,
         n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785,
         n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793,
         n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801,
         n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809,
         n41810, n41811, n41812, n41813, n41814, n41815, n41816, n41817,
         n41818, n41819, n41820, n41821, n41822, n41823, n41824, n41825,
         n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833,
         n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841,
         n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849,
         n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857,
         n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865,
         n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873,
         n41874, n41875, n41876, n41877, n41878, n41879, n41880, n41881,
         n41882, n41883, n41884, n41885, n41886, n41887, n41888, n41889,
         n41890, n41891, n41892, n41893, n41894, n41895, n41896, n41897,
         n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905,
         n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913,
         n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921,
         n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929,
         n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937,
         n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945,
         n41946, n41947, n41948, n41949, n41950, n41951, n41952, n41953,
         n41954, n41955, n41956, n41957, n41958, n41959, n41960, n41961,
         n41962, n41963, n41964, n41965, n41966, n41967, n41968, n41969,
         n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977,
         n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985,
         n41986, n41987, n41988, n41989, n41990, n41991, n41992;
  wire   [1023:0] start_in;
  wire   [1023:0] ein;
  wire   [1023:0] creg;
  wire   [1023:0] ereg_next;
  wire   [1023:0] mreg;
  wire   [1023:0] nreg;

  DFF \start_reg_reg[0]  ( .D(start_in[1023]), .CLK(clk), .RST(rst), .I(1'b1), 
        .Q(start_in[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[127]) );
  DFF \start_reg_reg[128]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[128]) );
  DFF \start_reg_reg[129]  ( .D(start_in[128]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[129]) );
  DFF \start_reg_reg[130]  ( .D(start_in[129]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[130]) );
  DFF \start_reg_reg[131]  ( .D(start_in[130]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[131]) );
  DFF \start_reg_reg[132]  ( .D(start_in[131]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[132]) );
  DFF \start_reg_reg[133]  ( .D(start_in[132]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[133]) );
  DFF \start_reg_reg[134]  ( .D(start_in[133]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[134]) );
  DFF \start_reg_reg[135]  ( .D(start_in[134]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[135]) );
  DFF \start_reg_reg[136]  ( .D(start_in[135]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[136]) );
  DFF \start_reg_reg[137]  ( .D(start_in[136]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[137]) );
  DFF \start_reg_reg[138]  ( .D(start_in[137]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[138]) );
  DFF \start_reg_reg[139]  ( .D(start_in[138]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[139]) );
  DFF \start_reg_reg[140]  ( .D(start_in[139]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[140]) );
  DFF \start_reg_reg[141]  ( .D(start_in[140]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[141]) );
  DFF \start_reg_reg[142]  ( .D(start_in[141]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[142]) );
  DFF \start_reg_reg[143]  ( .D(start_in[142]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[143]) );
  DFF \start_reg_reg[144]  ( .D(start_in[143]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[144]) );
  DFF \start_reg_reg[145]  ( .D(start_in[144]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[145]) );
  DFF \start_reg_reg[146]  ( .D(start_in[145]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[146]) );
  DFF \start_reg_reg[147]  ( .D(start_in[146]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[147]) );
  DFF \start_reg_reg[148]  ( .D(start_in[147]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[148]) );
  DFF \start_reg_reg[149]  ( .D(start_in[148]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[149]) );
  DFF \start_reg_reg[150]  ( .D(start_in[149]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[150]) );
  DFF \start_reg_reg[151]  ( .D(start_in[150]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[151]) );
  DFF \start_reg_reg[152]  ( .D(start_in[151]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[152]) );
  DFF \start_reg_reg[153]  ( .D(start_in[152]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[153]) );
  DFF \start_reg_reg[154]  ( .D(start_in[153]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[154]) );
  DFF \start_reg_reg[155]  ( .D(start_in[154]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[155]) );
  DFF \start_reg_reg[156]  ( .D(start_in[155]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[156]) );
  DFF \start_reg_reg[157]  ( .D(start_in[156]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[157]) );
  DFF \start_reg_reg[158]  ( .D(start_in[157]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[158]) );
  DFF \start_reg_reg[159]  ( .D(start_in[158]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[159]) );
  DFF \start_reg_reg[160]  ( .D(start_in[159]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[160]) );
  DFF \start_reg_reg[161]  ( .D(start_in[160]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[161]) );
  DFF \start_reg_reg[162]  ( .D(start_in[161]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[162]) );
  DFF \start_reg_reg[163]  ( .D(start_in[162]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[163]) );
  DFF \start_reg_reg[164]  ( .D(start_in[163]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[164]) );
  DFF \start_reg_reg[165]  ( .D(start_in[164]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[165]) );
  DFF \start_reg_reg[166]  ( .D(start_in[165]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[166]) );
  DFF \start_reg_reg[167]  ( .D(start_in[166]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[167]) );
  DFF \start_reg_reg[168]  ( .D(start_in[167]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[168]) );
  DFF \start_reg_reg[169]  ( .D(start_in[168]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[169]) );
  DFF \start_reg_reg[170]  ( .D(start_in[169]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[170]) );
  DFF \start_reg_reg[171]  ( .D(start_in[170]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[171]) );
  DFF \start_reg_reg[172]  ( .D(start_in[171]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[172]) );
  DFF \start_reg_reg[173]  ( .D(start_in[172]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[173]) );
  DFF \start_reg_reg[174]  ( .D(start_in[173]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[174]) );
  DFF \start_reg_reg[175]  ( .D(start_in[174]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[175]) );
  DFF \start_reg_reg[176]  ( .D(start_in[175]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[176]) );
  DFF \start_reg_reg[177]  ( .D(start_in[176]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[177]) );
  DFF \start_reg_reg[178]  ( .D(start_in[177]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[178]) );
  DFF \start_reg_reg[179]  ( .D(start_in[178]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[179]) );
  DFF \start_reg_reg[180]  ( .D(start_in[179]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[180]) );
  DFF \start_reg_reg[181]  ( .D(start_in[180]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[181]) );
  DFF \start_reg_reg[182]  ( .D(start_in[181]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[182]) );
  DFF \start_reg_reg[183]  ( .D(start_in[182]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[183]) );
  DFF \start_reg_reg[184]  ( .D(start_in[183]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[184]) );
  DFF \start_reg_reg[185]  ( .D(start_in[184]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[185]) );
  DFF \start_reg_reg[186]  ( .D(start_in[185]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[186]) );
  DFF \start_reg_reg[187]  ( .D(start_in[186]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[187]) );
  DFF \start_reg_reg[188]  ( .D(start_in[187]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[188]) );
  DFF \start_reg_reg[189]  ( .D(start_in[188]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[189]) );
  DFF \start_reg_reg[190]  ( .D(start_in[189]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[190]) );
  DFF \start_reg_reg[191]  ( .D(start_in[190]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[191]) );
  DFF \start_reg_reg[192]  ( .D(start_in[191]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[192]) );
  DFF \start_reg_reg[193]  ( .D(start_in[192]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[193]) );
  DFF \start_reg_reg[194]  ( .D(start_in[193]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[194]) );
  DFF \start_reg_reg[195]  ( .D(start_in[194]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[195]) );
  DFF \start_reg_reg[196]  ( .D(start_in[195]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[196]) );
  DFF \start_reg_reg[197]  ( .D(start_in[196]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[197]) );
  DFF \start_reg_reg[198]  ( .D(start_in[197]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[198]) );
  DFF \start_reg_reg[199]  ( .D(start_in[198]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[199]) );
  DFF \start_reg_reg[200]  ( .D(start_in[199]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[200]) );
  DFF \start_reg_reg[201]  ( .D(start_in[200]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[201]) );
  DFF \start_reg_reg[202]  ( .D(start_in[201]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[202]) );
  DFF \start_reg_reg[203]  ( .D(start_in[202]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[203]) );
  DFF \start_reg_reg[204]  ( .D(start_in[203]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[204]) );
  DFF \start_reg_reg[205]  ( .D(start_in[204]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[205]) );
  DFF \start_reg_reg[206]  ( .D(start_in[205]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[206]) );
  DFF \start_reg_reg[207]  ( .D(start_in[206]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[207]) );
  DFF \start_reg_reg[208]  ( .D(start_in[207]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[208]) );
  DFF \start_reg_reg[209]  ( .D(start_in[208]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[209]) );
  DFF \start_reg_reg[210]  ( .D(start_in[209]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[210]) );
  DFF \start_reg_reg[211]  ( .D(start_in[210]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[211]) );
  DFF \start_reg_reg[212]  ( .D(start_in[211]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[212]) );
  DFF \start_reg_reg[213]  ( .D(start_in[212]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[213]) );
  DFF \start_reg_reg[214]  ( .D(start_in[213]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[214]) );
  DFF \start_reg_reg[215]  ( .D(start_in[214]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[215]) );
  DFF \start_reg_reg[216]  ( .D(start_in[215]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[216]) );
  DFF \start_reg_reg[217]  ( .D(start_in[216]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[217]) );
  DFF \start_reg_reg[218]  ( .D(start_in[217]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[218]) );
  DFF \start_reg_reg[219]  ( .D(start_in[218]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[219]) );
  DFF \start_reg_reg[220]  ( .D(start_in[219]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[220]) );
  DFF \start_reg_reg[221]  ( .D(start_in[220]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[221]) );
  DFF \start_reg_reg[222]  ( .D(start_in[221]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[222]) );
  DFF \start_reg_reg[223]  ( .D(start_in[222]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[223]) );
  DFF \start_reg_reg[224]  ( .D(start_in[223]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[224]) );
  DFF \start_reg_reg[225]  ( .D(start_in[224]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[225]) );
  DFF \start_reg_reg[226]  ( .D(start_in[225]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[226]) );
  DFF \start_reg_reg[227]  ( .D(start_in[226]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[227]) );
  DFF \start_reg_reg[228]  ( .D(start_in[227]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[228]) );
  DFF \start_reg_reg[229]  ( .D(start_in[228]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[229]) );
  DFF \start_reg_reg[230]  ( .D(start_in[229]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[230]) );
  DFF \start_reg_reg[231]  ( .D(start_in[230]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[231]) );
  DFF \start_reg_reg[232]  ( .D(start_in[231]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[232]) );
  DFF \start_reg_reg[233]  ( .D(start_in[232]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[233]) );
  DFF \start_reg_reg[234]  ( .D(start_in[233]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[234]) );
  DFF \start_reg_reg[235]  ( .D(start_in[234]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[235]) );
  DFF \start_reg_reg[236]  ( .D(start_in[235]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[236]) );
  DFF \start_reg_reg[237]  ( .D(start_in[236]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[237]) );
  DFF \start_reg_reg[238]  ( .D(start_in[237]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[238]) );
  DFF \start_reg_reg[239]  ( .D(start_in[238]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[239]) );
  DFF \start_reg_reg[240]  ( .D(start_in[239]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[240]) );
  DFF \start_reg_reg[241]  ( .D(start_in[240]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[241]) );
  DFF \start_reg_reg[242]  ( .D(start_in[241]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[242]) );
  DFF \start_reg_reg[243]  ( .D(start_in[242]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[243]) );
  DFF \start_reg_reg[244]  ( .D(start_in[243]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[244]) );
  DFF \start_reg_reg[245]  ( .D(start_in[244]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[245]) );
  DFF \start_reg_reg[246]  ( .D(start_in[245]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[246]) );
  DFF \start_reg_reg[247]  ( .D(start_in[246]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[247]) );
  DFF \start_reg_reg[248]  ( .D(start_in[247]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[248]) );
  DFF \start_reg_reg[249]  ( .D(start_in[248]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[249]) );
  DFF \start_reg_reg[250]  ( .D(start_in[249]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[250]) );
  DFF \start_reg_reg[251]  ( .D(start_in[250]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[251]) );
  DFF \start_reg_reg[252]  ( .D(start_in[251]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[252]) );
  DFF \start_reg_reg[253]  ( .D(start_in[252]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[253]) );
  DFF \start_reg_reg[254]  ( .D(start_in[253]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[254]) );
  DFF \start_reg_reg[255]  ( .D(start_in[254]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[255]) );
  DFF \start_reg_reg[256]  ( .D(start_in[255]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[256]) );
  DFF \start_reg_reg[257]  ( .D(start_in[256]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[257]) );
  DFF \start_reg_reg[258]  ( .D(start_in[257]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[258]) );
  DFF \start_reg_reg[259]  ( .D(start_in[258]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[259]) );
  DFF \start_reg_reg[260]  ( .D(start_in[259]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[260]) );
  DFF \start_reg_reg[261]  ( .D(start_in[260]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[261]) );
  DFF \start_reg_reg[262]  ( .D(start_in[261]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[262]) );
  DFF \start_reg_reg[263]  ( .D(start_in[262]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[263]) );
  DFF \start_reg_reg[264]  ( .D(start_in[263]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[264]) );
  DFF \start_reg_reg[265]  ( .D(start_in[264]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[265]) );
  DFF \start_reg_reg[266]  ( .D(start_in[265]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[266]) );
  DFF \start_reg_reg[267]  ( .D(start_in[266]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[267]) );
  DFF \start_reg_reg[268]  ( .D(start_in[267]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[268]) );
  DFF \start_reg_reg[269]  ( .D(start_in[268]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[269]) );
  DFF \start_reg_reg[270]  ( .D(start_in[269]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[270]) );
  DFF \start_reg_reg[271]  ( .D(start_in[270]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[271]) );
  DFF \start_reg_reg[272]  ( .D(start_in[271]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[272]) );
  DFF \start_reg_reg[273]  ( .D(start_in[272]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[273]) );
  DFF \start_reg_reg[274]  ( .D(start_in[273]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[274]) );
  DFF \start_reg_reg[275]  ( .D(start_in[274]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[275]) );
  DFF \start_reg_reg[276]  ( .D(start_in[275]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[276]) );
  DFF \start_reg_reg[277]  ( .D(start_in[276]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[277]) );
  DFF \start_reg_reg[278]  ( .D(start_in[277]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[278]) );
  DFF \start_reg_reg[279]  ( .D(start_in[278]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[279]) );
  DFF \start_reg_reg[280]  ( .D(start_in[279]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[280]) );
  DFF \start_reg_reg[281]  ( .D(start_in[280]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[281]) );
  DFF \start_reg_reg[282]  ( .D(start_in[281]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[282]) );
  DFF \start_reg_reg[283]  ( .D(start_in[282]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[283]) );
  DFF \start_reg_reg[284]  ( .D(start_in[283]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[284]) );
  DFF \start_reg_reg[285]  ( .D(start_in[284]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[285]) );
  DFF \start_reg_reg[286]  ( .D(start_in[285]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[286]) );
  DFF \start_reg_reg[287]  ( .D(start_in[286]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[287]) );
  DFF \start_reg_reg[288]  ( .D(start_in[287]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[288]) );
  DFF \start_reg_reg[289]  ( .D(start_in[288]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[289]) );
  DFF \start_reg_reg[290]  ( .D(start_in[289]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[290]) );
  DFF \start_reg_reg[291]  ( .D(start_in[290]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[291]) );
  DFF \start_reg_reg[292]  ( .D(start_in[291]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[292]) );
  DFF \start_reg_reg[293]  ( .D(start_in[292]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[293]) );
  DFF \start_reg_reg[294]  ( .D(start_in[293]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[294]) );
  DFF \start_reg_reg[295]  ( .D(start_in[294]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[295]) );
  DFF \start_reg_reg[296]  ( .D(start_in[295]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[296]) );
  DFF \start_reg_reg[297]  ( .D(start_in[296]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[297]) );
  DFF \start_reg_reg[298]  ( .D(start_in[297]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[298]) );
  DFF \start_reg_reg[299]  ( .D(start_in[298]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[299]) );
  DFF \start_reg_reg[300]  ( .D(start_in[299]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[300]) );
  DFF \start_reg_reg[301]  ( .D(start_in[300]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[301]) );
  DFF \start_reg_reg[302]  ( .D(start_in[301]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[302]) );
  DFF \start_reg_reg[303]  ( .D(start_in[302]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[303]) );
  DFF \start_reg_reg[304]  ( .D(start_in[303]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[304]) );
  DFF \start_reg_reg[305]  ( .D(start_in[304]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[305]) );
  DFF \start_reg_reg[306]  ( .D(start_in[305]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[306]) );
  DFF \start_reg_reg[307]  ( .D(start_in[306]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[307]) );
  DFF \start_reg_reg[308]  ( .D(start_in[307]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[308]) );
  DFF \start_reg_reg[309]  ( .D(start_in[308]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[309]) );
  DFF \start_reg_reg[310]  ( .D(start_in[309]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[310]) );
  DFF \start_reg_reg[311]  ( .D(start_in[310]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[311]) );
  DFF \start_reg_reg[312]  ( .D(start_in[311]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[312]) );
  DFF \start_reg_reg[313]  ( .D(start_in[312]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[313]) );
  DFF \start_reg_reg[314]  ( .D(start_in[313]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[314]) );
  DFF \start_reg_reg[315]  ( .D(start_in[314]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[315]) );
  DFF \start_reg_reg[316]  ( .D(start_in[315]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[316]) );
  DFF \start_reg_reg[317]  ( .D(start_in[316]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[317]) );
  DFF \start_reg_reg[318]  ( .D(start_in[317]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[318]) );
  DFF \start_reg_reg[319]  ( .D(start_in[318]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[319]) );
  DFF \start_reg_reg[320]  ( .D(start_in[319]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[320]) );
  DFF \start_reg_reg[321]  ( .D(start_in[320]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[321]) );
  DFF \start_reg_reg[322]  ( .D(start_in[321]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[322]) );
  DFF \start_reg_reg[323]  ( .D(start_in[322]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[323]) );
  DFF \start_reg_reg[324]  ( .D(start_in[323]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[324]) );
  DFF \start_reg_reg[325]  ( .D(start_in[324]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[325]) );
  DFF \start_reg_reg[326]  ( .D(start_in[325]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[326]) );
  DFF \start_reg_reg[327]  ( .D(start_in[326]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[327]) );
  DFF \start_reg_reg[328]  ( .D(start_in[327]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[328]) );
  DFF \start_reg_reg[329]  ( .D(start_in[328]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[329]) );
  DFF \start_reg_reg[330]  ( .D(start_in[329]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[330]) );
  DFF \start_reg_reg[331]  ( .D(start_in[330]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[331]) );
  DFF \start_reg_reg[332]  ( .D(start_in[331]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[332]) );
  DFF \start_reg_reg[333]  ( .D(start_in[332]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[333]) );
  DFF \start_reg_reg[334]  ( .D(start_in[333]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[334]) );
  DFF \start_reg_reg[335]  ( .D(start_in[334]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[335]) );
  DFF \start_reg_reg[336]  ( .D(start_in[335]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[336]) );
  DFF \start_reg_reg[337]  ( .D(start_in[336]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[337]) );
  DFF \start_reg_reg[338]  ( .D(start_in[337]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[338]) );
  DFF \start_reg_reg[339]  ( .D(start_in[338]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[339]) );
  DFF \start_reg_reg[340]  ( .D(start_in[339]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[340]) );
  DFF \start_reg_reg[341]  ( .D(start_in[340]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[341]) );
  DFF \start_reg_reg[342]  ( .D(start_in[341]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[342]) );
  DFF \start_reg_reg[343]  ( .D(start_in[342]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[343]) );
  DFF \start_reg_reg[344]  ( .D(start_in[343]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[344]) );
  DFF \start_reg_reg[345]  ( .D(start_in[344]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[345]) );
  DFF \start_reg_reg[346]  ( .D(start_in[345]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[346]) );
  DFF \start_reg_reg[347]  ( .D(start_in[346]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[347]) );
  DFF \start_reg_reg[348]  ( .D(start_in[347]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[348]) );
  DFF \start_reg_reg[349]  ( .D(start_in[348]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[349]) );
  DFF \start_reg_reg[350]  ( .D(start_in[349]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[350]) );
  DFF \start_reg_reg[351]  ( .D(start_in[350]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[351]) );
  DFF \start_reg_reg[352]  ( .D(start_in[351]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[352]) );
  DFF \start_reg_reg[353]  ( .D(start_in[352]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[353]) );
  DFF \start_reg_reg[354]  ( .D(start_in[353]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[354]) );
  DFF \start_reg_reg[355]  ( .D(start_in[354]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[355]) );
  DFF \start_reg_reg[356]  ( .D(start_in[355]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[356]) );
  DFF \start_reg_reg[357]  ( .D(start_in[356]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[357]) );
  DFF \start_reg_reg[358]  ( .D(start_in[357]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[358]) );
  DFF \start_reg_reg[359]  ( .D(start_in[358]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[359]) );
  DFF \start_reg_reg[360]  ( .D(start_in[359]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[360]) );
  DFF \start_reg_reg[361]  ( .D(start_in[360]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[361]) );
  DFF \start_reg_reg[362]  ( .D(start_in[361]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[362]) );
  DFF \start_reg_reg[363]  ( .D(start_in[362]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[363]) );
  DFF \start_reg_reg[364]  ( .D(start_in[363]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[364]) );
  DFF \start_reg_reg[365]  ( .D(start_in[364]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[365]) );
  DFF \start_reg_reg[366]  ( .D(start_in[365]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[366]) );
  DFF \start_reg_reg[367]  ( .D(start_in[366]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[367]) );
  DFF \start_reg_reg[368]  ( .D(start_in[367]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[368]) );
  DFF \start_reg_reg[369]  ( .D(start_in[368]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[369]) );
  DFF \start_reg_reg[370]  ( .D(start_in[369]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[370]) );
  DFF \start_reg_reg[371]  ( .D(start_in[370]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[371]) );
  DFF \start_reg_reg[372]  ( .D(start_in[371]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[372]) );
  DFF \start_reg_reg[373]  ( .D(start_in[372]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[373]) );
  DFF \start_reg_reg[374]  ( .D(start_in[373]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[374]) );
  DFF \start_reg_reg[375]  ( .D(start_in[374]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[375]) );
  DFF \start_reg_reg[376]  ( .D(start_in[375]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[376]) );
  DFF \start_reg_reg[377]  ( .D(start_in[376]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[377]) );
  DFF \start_reg_reg[378]  ( .D(start_in[377]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[378]) );
  DFF \start_reg_reg[379]  ( .D(start_in[378]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[379]) );
  DFF \start_reg_reg[380]  ( .D(start_in[379]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[380]) );
  DFF \start_reg_reg[381]  ( .D(start_in[380]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[381]) );
  DFF \start_reg_reg[382]  ( .D(start_in[381]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[382]) );
  DFF \start_reg_reg[383]  ( .D(start_in[382]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[383]) );
  DFF \start_reg_reg[384]  ( .D(start_in[383]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[384]) );
  DFF \start_reg_reg[385]  ( .D(start_in[384]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[385]) );
  DFF \start_reg_reg[386]  ( .D(start_in[385]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[386]) );
  DFF \start_reg_reg[387]  ( .D(start_in[386]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[387]) );
  DFF \start_reg_reg[388]  ( .D(start_in[387]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[388]) );
  DFF \start_reg_reg[389]  ( .D(start_in[388]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[389]) );
  DFF \start_reg_reg[390]  ( .D(start_in[389]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[390]) );
  DFF \start_reg_reg[391]  ( .D(start_in[390]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[391]) );
  DFF \start_reg_reg[392]  ( .D(start_in[391]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[392]) );
  DFF \start_reg_reg[393]  ( .D(start_in[392]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[393]) );
  DFF \start_reg_reg[394]  ( .D(start_in[393]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[394]) );
  DFF \start_reg_reg[395]  ( .D(start_in[394]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[395]) );
  DFF \start_reg_reg[396]  ( .D(start_in[395]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[396]) );
  DFF \start_reg_reg[397]  ( .D(start_in[396]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[397]) );
  DFF \start_reg_reg[398]  ( .D(start_in[397]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[398]) );
  DFF \start_reg_reg[399]  ( .D(start_in[398]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[399]) );
  DFF \start_reg_reg[400]  ( .D(start_in[399]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[400]) );
  DFF \start_reg_reg[401]  ( .D(start_in[400]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[401]) );
  DFF \start_reg_reg[402]  ( .D(start_in[401]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[402]) );
  DFF \start_reg_reg[403]  ( .D(start_in[402]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[403]) );
  DFF \start_reg_reg[404]  ( .D(start_in[403]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[404]) );
  DFF \start_reg_reg[405]  ( .D(start_in[404]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[405]) );
  DFF \start_reg_reg[406]  ( .D(start_in[405]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[406]) );
  DFF \start_reg_reg[407]  ( .D(start_in[406]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[407]) );
  DFF \start_reg_reg[408]  ( .D(start_in[407]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[408]) );
  DFF \start_reg_reg[409]  ( .D(start_in[408]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[409]) );
  DFF \start_reg_reg[410]  ( .D(start_in[409]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[410]) );
  DFF \start_reg_reg[411]  ( .D(start_in[410]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[411]) );
  DFF \start_reg_reg[412]  ( .D(start_in[411]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[412]) );
  DFF \start_reg_reg[413]  ( .D(start_in[412]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[413]) );
  DFF \start_reg_reg[414]  ( .D(start_in[413]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[414]) );
  DFF \start_reg_reg[415]  ( .D(start_in[414]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[415]) );
  DFF \start_reg_reg[416]  ( .D(start_in[415]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[416]) );
  DFF \start_reg_reg[417]  ( .D(start_in[416]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[417]) );
  DFF \start_reg_reg[418]  ( .D(start_in[417]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[418]) );
  DFF \start_reg_reg[419]  ( .D(start_in[418]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[419]) );
  DFF \start_reg_reg[420]  ( .D(start_in[419]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[420]) );
  DFF \start_reg_reg[421]  ( .D(start_in[420]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[421]) );
  DFF \start_reg_reg[422]  ( .D(start_in[421]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[422]) );
  DFF \start_reg_reg[423]  ( .D(start_in[422]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[423]) );
  DFF \start_reg_reg[424]  ( .D(start_in[423]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[424]) );
  DFF \start_reg_reg[425]  ( .D(start_in[424]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[425]) );
  DFF \start_reg_reg[426]  ( .D(start_in[425]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[426]) );
  DFF \start_reg_reg[427]  ( .D(start_in[426]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[427]) );
  DFF \start_reg_reg[428]  ( .D(start_in[427]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[428]) );
  DFF \start_reg_reg[429]  ( .D(start_in[428]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[429]) );
  DFF \start_reg_reg[430]  ( .D(start_in[429]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[430]) );
  DFF \start_reg_reg[431]  ( .D(start_in[430]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[431]) );
  DFF \start_reg_reg[432]  ( .D(start_in[431]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[432]) );
  DFF \start_reg_reg[433]  ( .D(start_in[432]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[433]) );
  DFF \start_reg_reg[434]  ( .D(start_in[433]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[434]) );
  DFF \start_reg_reg[435]  ( .D(start_in[434]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[435]) );
  DFF \start_reg_reg[436]  ( .D(start_in[435]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[436]) );
  DFF \start_reg_reg[437]  ( .D(start_in[436]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[437]) );
  DFF \start_reg_reg[438]  ( .D(start_in[437]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[438]) );
  DFF \start_reg_reg[439]  ( .D(start_in[438]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[439]) );
  DFF \start_reg_reg[440]  ( .D(start_in[439]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[440]) );
  DFF \start_reg_reg[441]  ( .D(start_in[440]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[441]) );
  DFF \start_reg_reg[442]  ( .D(start_in[441]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[442]) );
  DFF \start_reg_reg[443]  ( .D(start_in[442]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[443]) );
  DFF \start_reg_reg[444]  ( .D(start_in[443]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[444]) );
  DFF \start_reg_reg[445]  ( .D(start_in[444]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[445]) );
  DFF \start_reg_reg[446]  ( .D(start_in[445]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[446]) );
  DFF \start_reg_reg[447]  ( .D(start_in[446]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[447]) );
  DFF \start_reg_reg[448]  ( .D(start_in[447]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[448]) );
  DFF \start_reg_reg[449]  ( .D(start_in[448]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[449]) );
  DFF \start_reg_reg[450]  ( .D(start_in[449]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[450]) );
  DFF \start_reg_reg[451]  ( .D(start_in[450]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[451]) );
  DFF \start_reg_reg[452]  ( .D(start_in[451]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[452]) );
  DFF \start_reg_reg[453]  ( .D(start_in[452]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[453]) );
  DFF \start_reg_reg[454]  ( .D(start_in[453]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[454]) );
  DFF \start_reg_reg[455]  ( .D(start_in[454]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[455]) );
  DFF \start_reg_reg[456]  ( .D(start_in[455]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[456]) );
  DFF \start_reg_reg[457]  ( .D(start_in[456]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[457]) );
  DFF \start_reg_reg[458]  ( .D(start_in[457]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[458]) );
  DFF \start_reg_reg[459]  ( .D(start_in[458]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[459]) );
  DFF \start_reg_reg[460]  ( .D(start_in[459]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[460]) );
  DFF \start_reg_reg[461]  ( .D(start_in[460]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[461]) );
  DFF \start_reg_reg[462]  ( .D(start_in[461]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[462]) );
  DFF \start_reg_reg[463]  ( .D(start_in[462]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[463]) );
  DFF \start_reg_reg[464]  ( .D(start_in[463]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[464]) );
  DFF \start_reg_reg[465]  ( .D(start_in[464]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[465]) );
  DFF \start_reg_reg[466]  ( .D(start_in[465]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[466]) );
  DFF \start_reg_reg[467]  ( .D(start_in[466]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[467]) );
  DFF \start_reg_reg[468]  ( .D(start_in[467]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[468]) );
  DFF \start_reg_reg[469]  ( .D(start_in[468]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[469]) );
  DFF \start_reg_reg[470]  ( .D(start_in[469]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[470]) );
  DFF \start_reg_reg[471]  ( .D(start_in[470]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[471]) );
  DFF \start_reg_reg[472]  ( .D(start_in[471]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[472]) );
  DFF \start_reg_reg[473]  ( .D(start_in[472]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[473]) );
  DFF \start_reg_reg[474]  ( .D(start_in[473]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[474]) );
  DFF \start_reg_reg[475]  ( .D(start_in[474]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[475]) );
  DFF \start_reg_reg[476]  ( .D(start_in[475]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[476]) );
  DFF \start_reg_reg[477]  ( .D(start_in[476]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[477]) );
  DFF \start_reg_reg[478]  ( .D(start_in[477]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[478]) );
  DFF \start_reg_reg[479]  ( .D(start_in[478]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[479]) );
  DFF \start_reg_reg[480]  ( .D(start_in[479]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[480]) );
  DFF \start_reg_reg[481]  ( .D(start_in[480]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[481]) );
  DFF \start_reg_reg[482]  ( .D(start_in[481]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[482]) );
  DFF \start_reg_reg[483]  ( .D(start_in[482]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[483]) );
  DFF \start_reg_reg[484]  ( .D(start_in[483]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[484]) );
  DFF \start_reg_reg[485]  ( .D(start_in[484]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[485]) );
  DFF \start_reg_reg[486]  ( .D(start_in[485]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[486]) );
  DFF \start_reg_reg[487]  ( .D(start_in[486]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[487]) );
  DFF \start_reg_reg[488]  ( .D(start_in[487]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[488]) );
  DFF \start_reg_reg[489]  ( .D(start_in[488]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[489]) );
  DFF \start_reg_reg[490]  ( .D(start_in[489]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[490]) );
  DFF \start_reg_reg[491]  ( .D(start_in[490]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[491]) );
  DFF \start_reg_reg[492]  ( .D(start_in[491]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[492]) );
  DFF \start_reg_reg[493]  ( .D(start_in[492]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[493]) );
  DFF \start_reg_reg[494]  ( .D(start_in[493]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[494]) );
  DFF \start_reg_reg[495]  ( .D(start_in[494]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[495]) );
  DFF \start_reg_reg[496]  ( .D(start_in[495]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[496]) );
  DFF \start_reg_reg[497]  ( .D(start_in[496]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[497]) );
  DFF \start_reg_reg[498]  ( .D(start_in[497]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[498]) );
  DFF \start_reg_reg[499]  ( .D(start_in[498]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[499]) );
  DFF \start_reg_reg[500]  ( .D(start_in[499]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[500]) );
  DFF \start_reg_reg[501]  ( .D(start_in[500]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[501]) );
  DFF \start_reg_reg[502]  ( .D(start_in[501]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[502]) );
  DFF \start_reg_reg[503]  ( .D(start_in[502]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[503]) );
  DFF \start_reg_reg[504]  ( .D(start_in[503]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[504]) );
  DFF \start_reg_reg[505]  ( .D(start_in[504]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[505]) );
  DFF \start_reg_reg[506]  ( .D(start_in[505]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[506]) );
  DFF \start_reg_reg[507]  ( .D(start_in[506]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[507]) );
  DFF \start_reg_reg[508]  ( .D(start_in[507]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[508]) );
  DFF \start_reg_reg[509]  ( .D(start_in[508]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[509]) );
  DFF \start_reg_reg[510]  ( .D(start_in[509]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[510]) );
  DFF \start_reg_reg[511]  ( .D(start_in[510]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[511]) );
  DFF \start_reg_reg[512]  ( .D(start_in[511]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[512]) );
  DFF \start_reg_reg[513]  ( .D(start_in[512]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[513]) );
  DFF \start_reg_reg[514]  ( .D(start_in[513]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[514]) );
  DFF \start_reg_reg[515]  ( .D(start_in[514]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[515]) );
  DFF \start_reg_reg[516]  ( .D(start_in[515]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[516]) );
  DFF \start_reg_reg[517]  ( .D(start_in[516]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[517]) );
  DFF \start_reg_reg[518]  ( .D(start_in[517]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[518]) );
  DFF \start_reg_reg[519]  ( .D(start_in[518]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[519]) );
  DFF \start_reg_reg[520]  ( .D(start_in[519]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[520]) );
  DFF \start_reg_reg[521]  ( .D(start_in[520]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[521]) );
  DFF \start_reg_reg[522]  ( .D(start_in[521]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[522]) );
  DFF \start_reg_reg[523]  ( .D(start_in[522]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[523]) );
  DFF \start_reg_reg[524]  ( .D(start_in[523]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[524]) );
  DFF \start_reg_reg[525]  ( .D(start_in[524]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[525]) );
  DFF \start_reg_reg[526]  ( .D(start_in[525]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[526]) );
  DFF \start_reg_reg[527]  ( .D(start_in[526]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[527]) );
  DFF \start_reg_reg[528]  ( .D(start_in[527]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[528]) );
  DFF \start_reg_reg[529]  ( .D(start_in[528]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[529]) );
  DFF \start_reg_reg[530]  ( .D(start_in[529]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[530]) );
  DFF \start_reg_reg[531]  ( .D(start_in[530]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[531]) );
  DFF \start_reg_reg[532]  ( .D(start_in[531]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[532]) );
  DFF \start_reg_reg[533]  ( .D(start_in[532]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[533]) );
  DFF \start_reg_reg[534]  ( .D(start_in[533]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[534]) );
  DFF \start_reg_reg[535]  ( .D(start_in[534]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[535]) );
  DFF \start_reg_reg[536]  ( .D(start_in[535]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[536]) );
  DFF \start_reg_reg[537]  ( .D(start_in[536]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[537]) );
  DFF \start_reg_reg[538]  ( .D(start_in[537]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[538]) );
  DFF \start_reg_reg[539]  ( .D(start_in[538]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[539]) );
  DFF \start_reg_reg[540]  ( .D(start_in[539]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[540]) );
  DFF \start_reg_reg[541]  ( .D(start_in[540]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[541]) );
  DFF \start_reg_reg[542]  ( .D(start_in[541]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[542]) );
  DFF \start_reg_reg[543]  ( .D(start_in[542]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[543]) );
  DFF \start_reg_reg[544]  ( .D(start_in[543]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[544]) );
  DFF \start_reg_reg[545]  ( .D(start_in[544]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[545]) );
  DFF \start_reg_reg[546]  ( .D(start_in[545]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[546]) );
  DFF \start_reg_reg[547]  ( .D(start_in[546]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[547]) );
  DFF \start_reg_reg[548]  ( .D(start_in[547]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[548]) );
  DFF \start_reg_reg[549]  ( .D(start_in[548]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[549]) );
  DFF \start_reg_reg[550]  ( .D(start_in[549]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[550]) );
  DFF \start_reg_reg[551]  ( .D(start_in[550]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[551]) );
  DFF \start_reg_reg[552]  ( .D(start_in[551]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[552]) );
  DFF \start_reg_reg[553]  ( .D(start_in[552]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[553]) );
  DFF \start_reg_reg[554]  ( .D(start_in[553]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[554]) );
  DFF \start_reg_reg[555]  ( .D(start_in[554]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[555]) );
  DFF \start_reg_reg[556]  ( .D(start_in[555]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[556]) );
  DFF \start_reg_reg[557]  ( .D(start_in[556]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[557]) );
  DFF \start_reg_reg[558]  ( .D(start_in[557]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[558]) );
  DFF \start_reg_reg[559]  ( .D(start_in[558]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[559]) );
  DFF \start_reg_reg[560]  ( .D(start_in[559]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[560]) );
  DFF \start_reg_reg[561]  ( .D(start_in[560]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[561]) );
  DFF \start_reg_reg[562]  ( .D(start_in[561]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[562]) );
  DFF \start_reg_reg[563]  ( .D(start_in[562]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[563]) );
  DFF \start_reg_reg[564]  ( .D(start_in[563]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[564]) );
  DFF \start_reg_reg[565]  ( .D(start_in[564]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[565]) );
  DFF \start_reg_reg[566]  ( .D(start_in[565]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[566]) );
  DFF \start_reg_reg[567]  ( .D(start_in[566]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[567]) );
  DFF \start_reg_reg[568]  ( .D(start_in[567]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[568]) );
  DFF \start_reg_reg[569]  ( .D(start_in[568]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[569]) );
  DFF \start_reg_reg[570]  ( .D(start_in[569]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[570]) );
  DFF \start_reg_reg[571]  ( .D(start_in[570]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[571]) );
  DFF \start_reg_reg[572]  ( .D(start_in[571]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[572]) );
  DFF \start_reg_reg[573]  ( .D(start_in[572]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[573]) );
  DFF \start_reg_reg[574]  ( .D(start_in[573]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[574]) );
  DFF \start_reg_reg[575]  ( .D(start_in[574]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[575]) );
  DFF \start_reg_reg[576]  ( .D(start_in[575]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[576]) );
  DFF \start_reg_reg[577]  ( .D(start_in[576]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[577]) );
  DFF \start_reg_reg[578]  ( .D(start_in[577]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[578]) );
  DFF \start_reg_reg[579]  ( .D(start_in[578]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[579]) );
  DFF \start_reg_reg[580]  ( .D(start_in[579]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[580]) );
  DFF \start_reg_reg[581]  ( .D(start_in[580]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[581]) );
  DFF \start_reg_reg[582]  ( .D(start_in[581]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[582]) );
  DFF \start_reg_reg[583]  ( .D(start_in[582]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[583]) );
  DFF \start_reg_reg[584]  ( .D(start_in[583]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[584]) );
  DFF \start_reg_reg[585]  ( .D(start_in[584]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[585]) );
  DFF \start_reg_reg[586]  ( .D(start_in[585]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[586]) );
  DFF \start_reg_reg[587]  ( .D(start_in[586]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[587]) );
  DFF \start_reg_reg[588]  ( .D(start_in[587]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[588]) );
  DFF \start_reg_reg[589]  ( .D(start_in[588]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[589]) );
  DFF \start_reg_reg[590]  ( .D(start_in[589]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[590]) );
  DFF \start_reg_reg[591]  ( .D(start_in[590]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[591]) );
  DFF \start_reg_reg[592]  ( .D(start_in[591]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[592]) );
  DFF \start_reg_reg[593]  ( .D(start_in[592]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[593]) );
  DFF \start_reg_reg[594]  ( .D(start_in[593]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[594]) );
  DFF \start_reg_reg[595]  ( .D(start_in[594]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[595]) );
  DFF \start_reg_reg[596]  ( .D(start_in[595]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[596]) );
  DFF \start_reg_reg[597]  ( .D(start_in[596]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[597]) );
  DFF \start_reg_reg[598]  ( .D(start_in[597]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[598]) );
  DFF \start_reg_reg[599]  ( .D(start_in[598]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[599]) );
  DFF \start_reg_reg[600]  ( .D(start_in[599]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[600]) );
  DFF \start_reg_reg[601]  ( .D(start_in[600]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[601]) );
  DFF \start_reg_reg[602]  ( .D(start_in[601]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[602]) );
  DFF \start_reg_reg[603]  ( .D(start_in[602]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[603]) );
  DFF \start_reg_reg[604]  ( .D(start_in[603]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[604]) );
  DFF \start_reg_reg[605]  ( .D(start_in[604]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[605]) );
  DFF \start_reg_reg[606]  ( .D(start_in[605]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[606]) );
  DFF \start_reg_reg[607]  ( .D(start_in[606]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[607]) );
  DFF \start_reg_reg[608]  ( .D(start_in[607]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[608]) );
  DFF \start_reg_reg[609]  ( .D(start_in[608]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[609]) );
  DFF \start_reg_reg[610]  ( .D(start_in[609]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[610]) );
  DFF \start_reg_reg[611]  ( .D(start_in[610]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[611]) );
  DFF \start_reg_reg[612]  ( .D(start_in[611]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[612]) );
  DFF \start_reg_reg[613]  ( .D(start_in[612]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[613]) );
  DFF \start_reg_reg[614]  ( .D(start_in[613]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[614]) );
  DFF \start_reg_reg[615]  ( .D(start_in[614]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[615]) );
  DFF \start_reg_reg[616]  ( .D(start_in[615]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[616]) );
  DFF \start_reg_reg[617]  ( .D(start_in[616]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[617]) );
  DFF \start_reg_reg[618]  ( .D(start_in[617]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[618]) );
  DFF \start_reg_reg[619]  ( .D(start_in[618]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[619]) );
  DFF \start_reg_reg[620]  ( .D(start_in[619]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[620]) );
  DFF \start_reg_reg[621]  ( .D(start_in[620]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[621]) );
  DFF \start_reg_reg[622]  ( .D(start_in[621]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[622]) );
  DFF \start_reg_reg[623]  ( .D(start_in[622]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[623]) );
  DFF \start_reg_reg[624]  ( .D(start_in[623]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[624]) );
  DFF \start_reg_reg[625]  ( .D(start_in[624]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[625]) );
  DFF \start_reg_reg[626]  ( .D(start_in[625]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[626]) );
  DFF \start_reg_reg[627]  ( .D(start_in[626]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[627]) );
  DFF \start_reg_reg[628]  ( .D(start_in[627]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[628]) );
  DFF \start_reg_reg[629]  ( .D(start_in[628]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[629]) );
  DFF \start_reg_reg[630]  ( .D(start_in[629]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[630]) );
  DFF \start_reg_reg[631]  ( .D(start_in[630]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[631]) );
  DFF \start_reg_reg[632]  ( .D(start_in[631]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[632]) );
  DFF \start_reg_reg[633]  ( .D(start_in[632]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[633]) );
  DFF \start_reg_reg[634]  ( .D(start_in[633]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[634]) );
  DFF \start_reg_reg[635]  ( .D(start_in[634]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[635]) );
  DFF \start_reg_reg[636]  ( .D(start_in[635]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[636]) );
  DFF \start_reg_reg[637]  ( .D(start_in[636]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[637]) );
  DFF \start_reg_reg[638]  ( .D(start_in[637]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[638]) );
  DFF \start_reg_reg[639]  ( .D(start_in[638]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[639]) );
  DFF \start_reg_reg[640]  ( .D(start_in[639]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[640]) );
  DFF \start_reg_reg[641]  ( .D(start_in[640]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[641]) );
  DFF \start_reg_reg[642]  ( .D(start_in[641]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[642]) );
  DFF \start_reg_reg[643]  ( .D(start_in[642]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[643]) );
  DFF \start_reg_reg[644]  ( .D(start_in[643]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[644]) );
  DFF \start_reg_reg[645]  ( .D(start_in[644]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[645]) );
  DFF \start_reg_reg[646]  ( .D(start_in[645]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[646]) );
  DFF \start_reg_reg[647]  ( .D(start_in[646]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[647]) );
  DFF \start_reg_reg[648]  ( .D(start_in[647]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[648]) );
  DFF \start_reg_reg[649]  ( .D(start_in[648]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[649]) );
  DFF \start_reg_reg[650]  ( .D(start_in[649]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[650]) );
  DFF \start_reg_reg[651]  ( .D(start_in[650]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[651]) );
  DFF \start_reg_reg[652]  ( .D(start_in[651]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[652]) );
  DFF \start_reg_reg[653]  ( .D(start_in[652]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[653]) );
  DFF \start_reg_reg[654]  ( .D(start_in[653]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[654]) );
  DFF \start_reg_reg[655]  ( .D(start_in[654]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[655]) );
  DFF \start_reg_reg[656]  ( .D(start_in[655]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[656]) );
  DFF \start_reg_reg[657]  ( .D(start_in[656]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[657]) );
  DFF \start_reg_reg[658]  ( .D(start_in[657]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[658]) );
  DFF \start_reg_reg[659]  ( .D(start_in[658]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[659]) );
  DFF \start_reg_reg[660]  ( .D(start_in[659]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[660]) );
  DFF \start_reg_reg[661]  ( .D(start_in[660]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[661]) );
  DFF \start_reg_reg[662]  ( .D(start_in[661]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[662]) );
  DFF \start_reg_reg[663]  ( .D(start_in[662]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[663]) );
  DFF \start_reg_reg[664]  ( .D(start_in[663]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[664]) );
  DFF \start_reg_reg[665]  ( .D(start_in[664]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[665]) );
  DFF \start_reg_reg[666]  ( .D(start_in[665]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[666]) );
  DFF \start_reg_reg[667]  ( .D(start_in[666]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[667]) );
  DFF \start_reg_reg[668]  ( .D(start_in[667]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[668]) );
  DFF \start_reg_reg[669]  ( .D(start_in[668]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[669]) );
  DFF \start_reg_reg[670]  ( .D(start_in[669]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[670]) );
  DFF \start_reg_reg[671]  ( .D(start_in[670]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[671]) );
  DFF \start_reg_reg[672]  ( .D(start_in[671]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[672]) );
  DFF \start_reg_reg[673]  ( .D(start_in[672]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[673]) );
  DFF \start_reg_reg[674]  ( .D(start_in[673]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[674]) );
  DFF \start_reg_reg[675]  ( .D(start_in[674]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[675]) );
  DFF \start_reg_reg[676]  ( .D(start_in[675]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[676]) );
  DFF \start_reg_reg[677]  ( .D(start_in[676]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[677]) );
  DFF \start_reg_reg[678]  ( .D(start_in[677]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[678]) );
  DFF \start_reg_reg[679]  ( .D(start_in[678]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[679]) );
  DFF \start_reg_reg[680]  ( .D(start_in[679]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[680]) );
  DFF \start_reg_reg[681]  ( .D(start_in[680]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[681]) );
  DFF \start_reg_reg[682]  ( .D(start_in[681]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[682]) );
  DFF \start_reg_reg[683]  ( .D(start_in[682]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[683]) );
  DFF \start_reg_reg[684]  ( .D(start_in[683]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[684]) );
  DFF \start_reg_reg[685]  ( .D(start_in[684]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[685]) );
  DFF \start_reg_reg[686]  ( .D(start_in[685]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[686]) );
  DFF \start_reg_reg[687]  ( .D(start_in[686]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[687]) );
  DFF \start_reg_reg[688]  ( .D(start_in[687]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[688]) );
  DFF \start_reg_reg[689]  ( .D(start_in[688]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[689]) );
  DFF \start_reg_reg[690]  ( .D(start_in[689]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[690]) );
  DFF \start_reg_reg[691]  ( .D(start_in[690]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[691]) );
  DFF \start_reg_reg[692]  ( .D(start_in[691]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[692]) );
  DFF \start_reg_reg[693]  ( .D(start_in[692]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[693]) );
  DFF \start_reg_reg[694]  ( .D(start_in[693]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[694]) );
  DFF \start_reg_reg[695]  ( .D(start_in[694]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[695]) );
  DFF \start_reg_reg[696]  ( .D(start_in[695]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[696]) );
  DFF \start_reg_reg[697]  ( .D(start_in[696]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[697]) );
  DFF \start_reg_reg[698]  ( .D(start_in[697]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[698]) );
  DFF \start_reg_reg[699]  ( .D(start_in[698]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[699]) );
  DFF \start_reg_reg[700]  ( .D(start_in[699]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[700]) );
  DFF \start_reg_reg[701]  ( .D(start_in[700]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[701]) );
  DFF \start_reg_reg[702]  ( .D(start_in[701]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[702]) );
  DFF \start_reg_reg[703]  ( .D(start_in[702]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[703]) );
  DFF \start_reg_reg[704]  ( .D(start_in[703]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[704]) );
  DFF \start_reg_reg[705]  ( .D(start_in[704]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[705]) );
  DFF \start_reg_reg[706]  ( .D(start_in[705]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[706]) );
  DFF \start_reg_reg[707]  ( .D(start_in[706]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[707]) );
  DFF \start_reg_reg[708]  ( .D(start_in[707]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[708]) );
  DFF \start_reg_reg[709]  ( .D(start_in[708]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[709]) );
  DFF \start_reg_reg[710]  ( .D(start_in[709]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[710]) );
  DFF \start_reg_reg[711]  ( .D(start_in[710]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[711]) );
  DFF \start_reg_reg[712]  ( .D(start_in[711]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[712]) );
  DFF \start_reg_reg[713]  ( .D(start_in[712]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[713]) );
  DFF \start_reg_reg[714]  ( .D(start_in[713]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[714]) );
  DFF \start_reg_reg[715]  ( .D(start_in[714]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[715]) );
  DFF \start_reg_reg[716]  ( .D(start_in[715]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[716]) );
  DFF \start_reg_reg[717]  ( .D(start_in[716]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[717]) );
  DFF \start_reg_reg[718]  ( .D(start_in[717]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[718]) );
  DFF \start_reg_reg[719]  ( .D(start_in[718]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[719]) );
  DFF \start_reg_reg[720]  ( .D(start_in[719]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[720]) );
  DFF \start_reg_reg[721]  ( .D(start_in[720]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[721]) );
  DFF \start_reg_reg[722]  ( .D(start_in[721]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[722]) );
  DFF \start_reg_reg[723]  ( .D(start_in[722]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[723]) );
  DFF \start_reg_reg[724]  ( .D(start_in[723]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[724]) );
  DFF \start_reg_reg[725]  ( .D(start_in[724]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[725]) );
  DFF \start_reg_reg[726]  ( .D(start_in[725]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[726]) );
  DFF \start_reg_reg[727]  ( .D(start_in[726]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[727]) );
  DFF \start_reg_reg[728]  ( .D(start_in[727]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[728]) );
  DFF \start_reg_reg[729]  ( .D(start_in[728]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[729]) );
  DFF \start_reg_reg[730]  ( .D(start_in[729]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[730]) );
  DFF \start_reg_reg[731]  ( .D(start_in[730]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[731]) );
  DFF \start_reg_reg[732]  ( .D(start_in[731]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[732]) );
  DFF \start_reg_reg[733]  ( .D(start_in[732]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[733]) );
  DFF \start_reg_reg[734]  ( .D(start_in[733]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[734]) );
  DFF \start_reg_reg[735]  ( .D(start_in[734]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[735]) );
  DFF \start_reg_reg[736]  ( .D(start_in[735]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[736]) );
  DFF \start_reg_reg[737]  ( .D(start_in[736]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[737]) );
  DFF \start_reg_reg[738]  ( .D(start_in[737]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[738]) );
  DFF \start_reg_reg[739]  ( .D(start_in[738]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[739]) );
  DFF \start_reg_reg[740]  ( .D(start_in[739]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[740]) );
  DFF \start_reg_reg[741]  ( .D(start_in[740]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[741]) );
  DFF \start_reg_reg[742]  ( .D(start_in[741]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[742]) );
  DFF \start_reg_reg[743]  ( .D(start_in[742]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[743]) );
  DFF \start_reg_reg[744]  ( .D(start_in[743]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[744]) );
  DFF \start_reg_reg[745]  ( .D(start_in[744]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[745]) );
  DFF \start_reg_reg[746]  ( .D(start_in[745]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[746]) );
  DFF \start_reg_reg[747]  ( .D(start_in[746]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[747]) );
  DFF \start_reg_reg[748]  ( .D(start_in[747]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[748]) );
  DFF \start_reg_reg[749]  ( .D(start_in[748]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[749]) );
  DFF \start_reg_reg[750]  ( .D(start_in[749]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[750]) );
  DFF \start_reg_reg[751]  ( .D(start_in[750]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[751]) );
  DFF \start_reg_reg[752]  ( .D(start_in[751]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[752]) );
  DFF \start_reg_reg[753]  ( .D(start_in[752]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[753]) );
  DFF \start_reg_reg[754]  ( .D(start_in[753]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[754]) );
  DFF \start_reg_reg[755]  ( .D(start_in[754]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[755]) );
  DFF \start_reg_reg[756]  ( .D(start_in[755]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[756]) );
  DFF \start_reg_reg[757]  ( .D(start_in[756]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[757]) );
  DFF \start_reg_reg[758]  ( .D(start_in[757]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[758]) );
  DFF \start_reg_reg[759]  ( .D(start_in[758]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[759]) );
  DFF \start_reg_reg[760]  ( .D(start_in[759]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[760]) );
  DFF \start_reg_reg[761]  ( .D(start_in[760]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[761]) );
  DFF \start_reg_reg[762]  ( .D(start_in[761]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[762]) );
  DFF \start_reg_reg[763]  ( .D(start_in[762]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[763]) );
  DFF \start_reg_reg[764]  ( .D(start_in[763]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[764]) );
  DFF \start_reg_reg[765]  ( .D(start_in[764]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[765]) );
  DFF \start_reg_reg[766]  ( .D(start_in[765]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[766]) );
  DFF \start_reg_reg[767]  ( .D(start_in[766]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[767]) );
  DFF \start_reg_reg[768]  ( .D(start_in[767]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[768]) );
  DFF \start_reg_reg[769]  ( .D(start_in[768]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[769]) );
  DFF \start_reg_reg[770]  ( .D(start_in[769]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[770]) );
  DFF \start_reg_reg[771]  ( .D(start_in[770]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[771]) );
  DFF \start_reg_reg[772]  ( .D(start_in[771]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[772]) );
  DFF \start_reg_reg[773]  ( .D(start_in[772]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[773]) );
  DFF \start_reg_reg[774]  ( .D(start_in[773]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[774]) );
  DFF \start_reg_reg[775]  ( .D(start_in[774]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[775]) );
  DFF \start_reg_reg[776]  ( .D(start_in[775]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[776]) );
  DFF \start_reg_reg[777]  ( .D(start_in[776]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[777]) );
  DFF \start_reg_reg[778]  ( .D(start_in[777]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[778]) );
  DFF \start_reg_reg[779]  ( .D(start_in[778]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[779]) );
  DFF \start_reg_reg[780]  ( .D(start_in[779]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[780]) );
  DFF \start_reg_reg[781]  ( .D(start_in[780]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[781]) );
  DFF \start_reg_reg[782]  ( .D(start_in[781]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[782]) );
  DFF \start_reg_reg[783]  ( .D(start_in[782]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[783]) );
  DFF \start_reg_reg[784]  ( .D(start_in[783]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[784]) );
  DFF \start_reg_reg[785]  ( .D(start_in[784]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[785]) );
  DFF \start_reg_reg[786]  ( .D(start_in[785]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[786]) );
  DFF \start_reg_reg[787]  ( .D(start_in[786]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[787]) );
  DFF \start_reg_reg[788]  ( .D(start_in[787]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[788]) );
  DFF \start_reg_reg[789]  ( .D(start_in[788]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[789]) );
  DFF \start_reg_reg[790]  ( .D(start_in[789]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[790]) );
  DFF \start_reg_reg[791]  ( .D(start_in[790]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[791]) );
  DFF \start_reg_reg[792]  ( .D(start_in[791]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[792]) );
  DFF \start_reg_reg[793]  ( .D(start_in[792]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[793]) );
  DFF \start_reg_reg[794]  ( .D(start_in[793]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[794]) );
  DFF \start_reg_reg[795]  ( .D(start_in[794]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[795]) );
  DFF \start_reg_reg[796]  ( .D(start_in[795]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[796]) );
  DFF \start_reg_reg[797]  ( .D(start_in[796]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[797]) );
  DFF \start_reg_reg[798]  ( .D(start_in[797]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[798]) );
  DFF \start_reg_reg[799]  ( .D(start_in[798]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[799]) );
  DFF \start_reg_reg[800]  ( .D(start_in[799]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[800]) );
  DFF \start_reg_reg[801]  ( .D(start_in[800]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[801]) );
  DFF \start_reg_reg[802]  ( .D(start_in[801]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[802]) );
  DFF \start_reg_reg[803]  ( .D(start_in[802]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[803]) );
  DFF \start_reg_reg[804]  ( .D(start_in[803]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[804]) );
  DFF \start_reg_reg[805]  ( .D(start_in[804]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[805]) );
  DFF \start_reg_reg[806]  ( .D(start_in[805]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[806]) );
  DFF \start_reg_reg[807]  ( .D(start_in[806]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[807]) );
  DFF \start_reg_reg[808]  ( .D(start_in[807]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[808]) );
  DFF \start_reg_reg[809]  ( .D(start_in[808]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[809]) );
  DFF \start_reg_reg[810]  ( .D(start_in[809]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[810]) );
  DFF \start_reg_reg[811]  ( .D(start_in[810]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[811]) );
  DFF \start_reg_reg[812]  ( .D(start_in[811]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[812]) );
  DFF \start_reg_reg[813]  ( .D(start_in[812]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[813]) );
  DFF \start_reg_reg[814]  ( .D(start_in[813]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[814]) );
  DFF \start_reg_reg[815]  ( .D(start_in[814]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[815]) );
  DFF \start_reg_reg[816]  ( .D(start_in[815]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[816]) );
  DFF \start_reg_reg[817]  ( .D(start_in[816]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[817]) );
  DFF \start_reg_reg[818]  ( .D(start_in[817]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[818]) );
  DFF \start_reg_reg[819]  ( .D(start_in[818]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[819]) );
  DFF \start_reg_reg[820]  ( .D(start_in[819]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[820]) );
  DFF \start_reg_reg[821]  ( .D(start_in[820]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[821]) );
  DFF \start_reg_reg[822]  ( .D(start_in[821]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[822]) );
  DFF \start_reg_reg[823]  ( .D(start_in[822]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[823]) );
  DFF \start_reg_reg[824]  ( .D(start_in[823]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[824]) );
  DFF \start_reg_reg[825]  ( .D(start_in[824]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[825]) );
  DFF \start_reg_reg[826]  ( .D(start_in[825]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[826]) );
  DFF \start_reg_reg[827]  ( .D(start_in[826]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[827]) );
  DFF \start_reg_reg[828]  ( .D(start_in[827]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[828]) );
  DFF \start_reg_reg[829]  ( .D(start_in[828]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[829]) );
  DFF \start_reg_reg[830]  ( .D(start_in[829]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[830]) );
  DFF \start_reg_reg[831]  ( .D(start_in[830]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[831]) );
  DFF \start_reg_reg[832]  ( .D(start_in[831]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[832]) );
  DFF \start_reg_reg[833]  ( .D(start_in[832]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[833]) );
  DFF \start_reg_reg[834]  ( .D(start_in[833]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[834]) );
  DFF \start_reg_reg[835]  ( .D(start_in[834]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[835]) );
  DFF \start_reg_reg[836]  ( .D(start_in[835]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[836]) );
  DFF \start_reg_reg[837]  ( .D(start_in[836]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[837]) );
  DFF \start_reg_reg[838]  ( .D(start_in[837]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[838]) );
  DFF \start_reg_reg[839]  ( .D(start_in[838]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[839]) );
  DFF \start_reg_reg[840]  ( .D(start_in[839]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[840]) );
  DFF \start_reg_reg[841]  ( .D(start_in[840]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[841]) );
  DFF \start_reg_reg[842]  ( .D(start_in[841]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[842]) );
  DFF \start_reg_reg[843]  ( .D(start_in[842]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[843]) );
  DFF \start_reg_reg[844]  ( .D(start_in[843]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[844]) );
  DFF \start_reg_reg[845]  ( .D(start_in[844]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[845]) );
  DFF \start_reg_reg[846]  ( .D(start_in[845]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[846]) );
  DFF \start_reg_reg[847]  ( .D(start_in[846]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[847]) );
  DFF \start_reg_reg[848]  ( .D(start_in[847]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[848]) );
  DFF \start_reg_reg[849]  ( .D(start_in[848]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[849]) );
  DFF \start_reg_reg[850]  ( .D(start_in[849]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[850]) );
  DFF \start_reg_reg[851]  ( .D(start_in[850]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[851]) );
  DFF \start_reg_reg[852]  ( .D(start_in[851]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[852]) );
  DFF \start_reg_reg[853]  ( .D(start_in[852]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[853]) );
  DFF \start_reg_reg[854]  ( .D(start_in[853]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[854]) );
  DFF \start_reg_reg[855]  ( .D(start_in[854]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[855]) );
  DFF \start_reg_reg[856]  ( .D(start_in[855]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[856]) );
  DFF \start_reg_reg[857]  ( .D(start_in[856]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[857]) );
  DFF \start_reg_reg[858]  ( .D(start_in[857]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[858]) );
  DFF \start_reg_reg[859]  ( .D(start_in[858]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[859]) );
  DFF \start_reg_reg[860]  ( .D(start_in[859]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[860]) );
  DFF \start_reg_reg[861]  ( .D(start_in[860]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[861]) );
  DFF \start_reg_reg[862]  ( .D(start_in[861]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[862]) );
  DFF \start_reg_reg[863]  ( .D(start_in[862]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[863]) );
  DFF \start_reg_reg[864]  ( .D(start_in[863]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[864]) );
  DFF \start_reg_reg[865]  ( .D(start_in[864]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[865]) );
  DFF \start_reg_reg[866]  ( .D(start_in[865]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[866]) );
  DFF \start_reg_reg[867]  ( .D(start_in[866]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[867]) );
  DFF \start_reg_reg[868]  ( .D(start_in[867]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[868]) );
  DFF \start_reg_reg[869]  ( .D(start_in[868]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[869]) );
  DFF \start_reg_reg[870]  ( .D(start_in[869]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[870]) );
  DFF \start_reg_reg[871]  ( .D(start_in[870]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[871]) );
  DFF \start_reg_reg[872]  ( .D(start_in[871]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[872]) );
  DFF \start_reg_reg[873]  ( .D(start_in[872]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[873]) );
  DFF \start_reg_reg[874]  ( .D(start_in[873]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[874]) );
  DFF \start_reg_reg[875]  ( .D(start_in[874]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[875]) );
  DFF \start_reg_reg[876]  ( .D(start_in[875]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[876]) );
  DFF \start_reg_reg[877]  ( .D(start_in[876]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[877]) );
  DFF \start_reg_reg[878]  ( .D(start_in[877]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[878]) );
  DFF \start_reg_reg[879]  ( .D(start_in[878]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[879]) );
  DFF \start_reg_reg[880]  ( .D(start_in[879]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[880]) );
  DFF \start_reg_reg[881]  ( .D(start_in[880]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[881]) );
  DFF \start_reg_reg[882]  ( .D(start_in[881]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[882]) );
  DFF \start_reg_reg[883]  ( .D(start_in[882]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[883]) );
  DFF \start_reg_reg[884]  ( .D(start_in[883]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[884]) );
  DFF \start_reg_reg[885]  ( .D(start_in[884]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[885]) );
  DFF \start_reg_reg[886]  ( .D(start_in[885]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[886]) );
  DFF \start_reg_reg[887]  ( .D(start_in[886]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[887]) );
  DFF \start_reg_reg[888]  ( .D(start_in[887]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[888]) );
  DFF \start_reg_reg[889]  ( .D(start_in[888]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[889]) );
  DFF \start_reg_reg[890]  ( .D(start_in[889]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[890]) );
  DFF \start_reg_reg[891]  ( .D(start_in[890]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[891]) );
  DFF \start_reg_reg[892]  ( .D(start_in[891]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[892]) );
  DFF \start_reg_reg[893]  ( .D(start_in[892]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[893]) );
  DFF \start_reg_reg[894]  ( .D(start_in[893]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[894]) );
  DFF \start_reg_reg[895]  ( .D(start_in[894]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[895]) );
  DFF \start_reg_reg[896]  ( .D(start_in[895]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[896]) );
  DFF \start_reg_reg[897]  ( .D(start_in[896]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[897]) );
  DFF \start_reg_reg[898]  ( .D(start_in[897]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[898]) );
  DFF \start_reg_reg[899]  ( .D(start_in[898]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[899]) );
  DFF \start_reg_reg[900]  ( .D(start_in[899]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[900]) );
  DFF \start_reg_reg[901]  ( .D(start_in[900]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[901]) );
  DFF \start_reg_reg[902]  ( .D(start_in[901]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[902]) );
  DFF \start_reg_reg[903]  ( .D(start_in[902]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[903]) );
  DFF \start_reg_reg[904]  ( .D(start_in[903]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[904]) );
  DFF \start_reg_reg[905]  ( .D(start_in[904]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[905]) );
  DFF \start_reg_reg[906]  ( .D(start_in[905]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[906]) );
  DFF \start_reg_reg[907]  ( .D(start_in[906]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[907]) );
  DFF \start_reg_reg[908]  ( .D(start_in[907]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[908]) );
  DFF \start_reg_reg[909]  ( .D(start_in[908]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[909]) );
  DFF \start_reg_reg[910]  ( .D(start_in[909]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[910]) );
  DFF \start_reg_reg[911]  ( .D(start_in[910]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[911]) );
  DFF \start_reg_reg[912]  ( .D(start_in[911]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[912]) );
  DFF \start_reg_reg[913]  ( .D(start_in[912]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[913]) );
  DFF \start_reg_reg[914]  ( .D(start_in[913]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[914]) );
  DFF \start_reg_reg[915]  ( .D(start_in[914]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[915]) );
  DFF \start_reg_reg[916]  ( .D(start_in[915]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[916]) );
  DFF \start_reg_reg[917]  ( .D(start_in[916]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[917]) );
  DFF \start_reg_reg[918]  ( .D(start_in[917]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[918]) );
  DFF \start_reg_reg[919]  ( .D(start_in[918]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[919]) );
  DFF \start_reg_reg[920]  ( .D(start_in[919]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[920]) );
  DFF \start_reg_reg[921]  ( .D(start_in[920]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[921]) );
  DFF \start_reg_reg[922]  ( .D(start_in[921]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[922]) );
  DFF \start_reg_reg[923]  ( .D(start_in[922]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[923]) );
  DFF \start_reg_reg[924]  ( .D(start_in[923]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[924]) );
  DFF \start_reg_reg[925]  ( .D(start_in[924]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[925]) );
  DFF \start_reg_reg[926]  ( .D(start_in[925]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[926]) );
  DFF \start_reg_reg[927]  ( .D(start_in[926]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[927]) );
  DFF \start_reg_reg[928]  ( .D(start_in[927]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[928]) );
  DFF \start_reg_reg[929]  ( .D(start_in[928]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[929]) );
  DFF \start_reg_reg[930]  ( .D(start_in[929]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[930]) );
  DFF \start_reg_reg[931]  ( .D(start_in[930]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[931]) );
  DFF \start_reg_reg[932]  ( .D(start_in[931]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[932]) );
  DFF \start_reg_reg[933]  ( .D(start_in[932]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[933]) );
  DFF \start_reg_reg[934]  ( .D(start_in[933]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[934]) );
  DFF \start_reg_reg[935]  ( .D(start_in[934]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[935]) );
  DFF \start_reg_reg[936]  ( .D(start_in[935]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[936]) );
  DFF \start_reg_reg[937]  ( .D(start_in[936]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[937]) );
  DFF \start_reg_reg[938]  ( .D(start_in[937]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[938]) );
  DFF \start_reg_reg[939]  ( .D(start_in[938]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[939]) );
  DFF \start_reg_reg[940]  ( .D(start_in[939]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[940]) );
  DFF \start_reg_reg[941]  ( .D(start_in[940]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[941]) );
  DFF \start_reg_reg[942]  ( .D(start_in[941]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[942]) );
  DFF \start_reg_reg[943]  ( .D(start_in[942]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[943]) );
  DFF \start_reg_reg[944]  ( .D(start_in[943]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[944]) );
  DFF \start_reg_reg[945]  ( .D(start_in[944]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[945]) );
  DFF \start_reg_reg[946]  ( .D(start_in[945]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[946]) );
  DFF \start_reg_reg[947]  ( .D(start_in[946]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[947]) );
  DFF \start_reg_reg[948]  ( .D(start_in[947]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[948]) );
  DFF \start_reg_reg[949]  ( .D(start_in[948]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[949]) );
  DFF \start_reg_reg[950]  ( .D(start_in[949]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[950]) );
  DFF \start_reg_reg[951]  ( .D(start_in[950]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[951]) );
  DFF \start_reg_reg[952]  ( .D(start_in[951]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[952]) );
  DFF \start_reg_reg[953]  ( .D(start_in[952]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[953]) );
  DFF \start_reg_reg[954]  ( .D(start_in[953]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[954]) );
  DFF \start_reg_reg[955]  ( .D(start_in[954]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[955]) );
  DFF \start_reg_reg[956]  ( .D(start_in[955]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[956]) );
  DFF \start_reg_reg[957]  ( .D(start_in[956]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[957]) );
  DFF \start_reg_reg[958]  ( .D(start_in[957]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[958]) );
  DFF \start_reg_reg[959]  ( .D(start_in[958]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[959]) );
  DFF \start_reg_reg[960]  ( .D(start_in[959]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[960]) );
  DFF \start_reg_reg[961]  ( .D(start_in[960]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[961]) );
  DFF \start_reg_reg[962]  ( .D(start_in[961]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[962]) );
  DFF \start_reg_reg[963]  ( .D(start_in[962]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[963]) );
  DFF \start_reg_reg[964]  ( .D(start_in[963]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[964]) );
  DFF \start_reg_reg[965]  ( .D(start_in[964]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[965]) );
  DFF \start_reg_reg[966]  ( .D(start_in[965]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[966]) );
  DFF \start_reg_reg[967]  ( .D(start_in[966]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[967]) );
  DFF \start_reg_reg[968]  ( .D(start_in[967]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[968]) );
  DFF \start_reg_reg[969]  ( .D(start_in[968]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[969]) );
  DFF \start_reg_reg[970]  ( .D(start_in[969]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[970]) );
  DFF \start_reg_reg[971]  ( .D(start_in[970]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[971]) );
  DFF \start_reg_reg[972]  ( .D(start_in[971]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[972]) );
  DFF \start_reg_reg[973]  ( .D(start_in[972]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[973]) );
  DFF \start_reg_reg[974]  ( .D(start_in[973]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[974]) );
  DFF \start_reg_reg[975]  ( .D(start_in[974]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[975]) );
  DFF \start_reg_reg[976]  ( .D(start_in[975]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[976]) );
  DFF \start_reg_reg[977]  ( .D(start_in[976]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[977]) );
  DFF \start_reg_reg[978]  ( .D(start_in[977]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[978]) );
  DFF \start_reg_reg[979]  ( .D(start_in[978]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[979]) );
  DFF \start_reg_reg[980]  ( .D(start_in[979]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[980]) );
  DFF \start_reg_reg[981]  ( .D(start_in[980]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[981]) );
  DFF \start_reg_reg[982]  ( .D(start_in[981]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[982]) );
  DFF \start_reg_reg[983]  ( .D(start_in[982]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[983]) );
  DFF \start_reg_reg[984]  ( .D(start_in[983]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[984]) );
  DFF \start_reg_reg[985]  ( .D(start_in[984]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[985]) );
  DFF \start_reg_reg[986]  ( .D(start_in[985]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[986]) );
  DFF \start_reg_reg[987]  ( .D(start_in[986]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[987]) );
  DFF \start_reg_reg[988]  ( .D(start_in[987]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[988]) );
  DFF \start_reg_reg[989]  ( .D(start_in[988]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[989]) );
  DFF \start_reg_reg[990]  ( .D(start_in[989]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[990]) );
  DFF \start_reg_reg[991]  ( .D(start_in[990]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[991]) );
  DFF \start_reg_reg[992]  ( .D(start_in[991]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[992]) );
  DFF \start_reg_reg[993]  ( .D(start_in[992]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[993]) );
  DFF \start_reg_reg[994]  ( .D(start_in[993]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[994]) );
  DFF \start_reg_reg[995]  ( .D(start_in[994]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[995]) );
  DFF \start_reg_reg[996]  ( .D(start_in[995]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[996]) );
  DFF \start_reg_reg[997]  ( .D(start_in[996]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[997]) );
  DFF \start_reg_reg[998]  ( .D(start_in[997]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[998]) );
  DFF \start_reg_reg[999]  ( .D(start_in[998]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[999]) );
  DFF \start_reg_reg[1000]  ( .D(start_in[999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(start_in[1000]) );
  DFF \start_reg_reg[1001]  ( .D(start_in[1000]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1001]) );
  DFF \start_reg_reg[1002]  ( .D(start_in[1001]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1002]) );
  DFF \start_reg_reg[1003]  ( .D(start_in[1002]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1003]) );
  DFF \start_reg_reg[1004]  ( .D(start_in[1003]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1004]) );
  DFF \start_reg_reg[1005]  ( .D(start_in[1004]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1005]) );
  DFF \start_reg_reg[1006]  ( .D(start_in[1005]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1006]) );
  DFF \start_reg_reg[1007]  ( .D(start_in[1006]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1007]) );
  DFF \start_reg_reg[1008]  ( .D(start_in[1007]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1008]) );
  DFF \start_reg_reg[1009]  ( .D(start_in[1008]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1009]) );
  DFF \start_reg_reg[1010]  ( .D(start_in[1009]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1010]) );
  DFF \start_reg_reg[1011]  ( .D(start_in[1010]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1011]) );
  DFF \start_reg_reg[1012]  ( .D(start_in[1011]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1012]) );
  DFF \start_reg_reg[1013]  ( .D(start_in[1012]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1013]) );
  DFF \start_reg_reg[1014]  ( .D(start_in[1013]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1014]) );
  DFF \start_reg_reg[1015]  ( .D(start_in[1014]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1015]) );
  DFF \start_reg_reg[1016]  ( .D(start_in[1015]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1016]) );
  DFF \start_reg_reg[1017]  ( .D(start_in[1016]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1017]) );
  DFF \start_reg_reg[1018]  ( .D(start_in[1017]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1018]) );
  DFF \start_reg_reg[1019]  ( .D(start_in[1018]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1019]) );
  DFF \start_reg_reg[1020]  ( .D(start_in[1019]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1020]) );
  DFF \start_reg_reg[1021]  ( .D(start_in[1020]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1021]) );
  DFF \start_reg_reg[1022]  ( .D(start_in[1021]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1022]) );
  DFF \start_reg_reg[1023]  ( .D(start_in[1022]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1023]) );
  DFF \nreg_reg[1023]  ( .D(nreg[1023]), .CLK(clk), .RST(rst), .I(e_init[1023]), .Q(nreg[1023]) );
  DFF \nreg_reg[1022]  ( .D(nreg[1022]), .CLK(clk), .RST(rst), .I(e_init[1022]), .Q(nreg[1022]) );
  DFF \nreg_reg[1021]  ( .D(nreg[1021]), .CLK(clk), .RST(rst), .I(e_init[1021]), .Q(nreg[1021]) );
  DFF \nreg_reg[1020]  ( .D(nreg[1020]), .CLK(clk), .RST(rst), .I(e_init[1020]), .Q(nreg[1020]) );
  DFF \nreg_reg[1019]  ( .D(nreg[1019]), .CLK(clk), .RST(rst), .I(e_init[1019]), .Q(nreg[1019]) );
  DFF \nreg_reg[1018]  ( .D(nreg[1018]), .CLK(clk), .RST(rst), .I(e_init[1018]), .Q(nreg[1018]) );
  DFF \nreg_reg[1017]  ( .D(nreg[1017]), .CLK(clk), .RST(rst), .I(e_init[1017]), .Q(nreg[1017]) );
  DFF \nreg_reg[1016]  ( .D(nreg[1016]), .CLK(clk), .RST(rst), .I(e_init[1016]), .Q(nreg[1016]) );
  DFF \nreg_reg[1015]  ( .D(nreg[1015]), .CLK(clk), .RST(rst), .I(e_init[1015]), .Q(nreg[1015]) );
  DFF \nreg_reg[1014]  ( .D(nreg[1014]), .CLK(clk), .RST(rst), .I(e_init[1014]), .Q(nreg[1014]) );
  DFF \nreg_reg[1013]  ( .D(nreg[1013]), .CLK(clk), .RST(rst), .I(e_init[1013]), .Q(nreg[1013]) );
  DFF \nreg_reg[1012]  ( .D(nreg[1012]), .CLK(clk), .RST(rst), .I(e_init[1012]), .Q(nreg[1012]) );
  DFF \nreg_reg[1011]  ( .D(nreg[1011]), .CLK(clk), .RST(rst), .I(e_init[1011]), .Q(nreg[1011]) );
  DFF \nreg_reg[1010]  ( .D(nreg[1010]), .CLK(clk), .RST(rst), .I(e_init[1010]), .Q(nreg[1010]) );
  DFF \nreg_reg[1009]  ( .D(nreg[1009]), .CLK(clk), .RST(rst), .I(e_init[1009]), .Q(nreg[1009]) );
  DFF \nreg_reg[1008]  ( .D(nreg[1008]), .CLK(clk), .RST(rst), .I(e_init[1008]), .Q(nreg[1008]) );
  DFF \nreg_reg[1007]  ( .D(nreg[1007]), .CLK(clk), .RST(rst), .I(e_init[1007]), .Q(nreg[1007]) );
  DFF \nreg_reg[1006]  ( .D(nreg[1006]), .CLK(clk), .RST(rst), .I(e_init[1006]), .Q(nreg[1006]) );
  DFF \nreg_reg[1005]  ( .D(nreg[1005]), .CLK(clk), .RST(rst), .I(e_init[1005]), .Q(nreg[1005]) );
  DFF \nreg_reg[1004]  ( .D(nreg[1004]), .CLK(clk), .RST(rst), .I(e_init[1004]), .Q(nreg[1004]) );
  DFF \nreg_reg[1003]  ( .D(nreg[1003]), .CLK(clk), .RST(rst), .I(e_init[1003]), .Q(nreg[1003]) );
  DFF \nreg_reg[1002]  ( .D(nreg[1002]), .CLK(clk), .RST(rst), .I(e_init[1002]), .Q(nreg[1002]) );
  DFF \nreg_reg[1001]  ( .D(nreg[1001]), .CLK(clk), .RST(rst), .I(e_init[1001]), .Q(nreg[1001]) );
  DFF \nreg_reg[1000]  ( .D(nreg[1000]), .CLK(clk), .RST(rst), .I(e_init[1000]), .Q(nreg[1000]) );
  DFF \nreg_reg[999]  ( .D(nreg[999]), .CLK(clk), .RST(rst), .I(e_init[999]), 
        .Q(nreg[999]) );
  DFF \nreg_reg[998]  ( .D(nreg[998]), .CLK(clk), .RST(rst), .I(e_init[998]), 
        .Q(nreg[998]) );
  DFF \nreg_reg[997]  ( .D(nreg[997]), .CLK(clk), .RST(rst), .I(e_init[997]), 
        .Q(nreg[997]) );
  DFF \nreg_reg[996]  ( .D(nreg[996]), .CLK(clk), .RST(rst), .I(e_init[996]), 
        .Q(nreg[996]) );
  DFF \nreg_reg[995]  ( .D(nreg[995]), .CLK(clk), .RST(rst), .I(e_init[995]), 
        .Q(nreg[995]) );
  DFF \nreg_reg[994]  ( .D(nreg[994]), .CLK(clk), .RST(rst), .I(e_init[994]), 
        .Q(nreg[994]) );
  DFF \nreg_reg[993]  ( .D(nreg[993]), .CLK(clk), .RST(rst), .I(e_init[993]), 
        .Q(nreg[993]) );
  DFF \nreg_reg[992]  ( .D(nreg[992]), .CLK(clk), .RST(rst), .I(e_init[992]), 
        .Q(nreg[992]) );
  DFF \nreg_reg[991]  ( .D(nreg[991]), .CLK(clk), .RST(rst), .I(e_init[991]), 
        .Q(nreg[991]) );
  DFF \nreg_reg[990]  ( .D(nreg[990]), .CLK(clk), .RST(rst), .I(e_init[990]), 
        .Q(nreg[990]) );
  DFF \nreg_reg[989]  ( .D(nreg[989]), .CLK(clk), .RST(rst), .I(e_init[989]), 
        .Q(nreg[989]) );
  DFF \nreg_reg[988]  ( .D(nreg[988]), .CLK(clk), .RST(rst), .I(e_init[988]), 
        .Q(nreg[988]) );
  DFF \nreg_reg[987]  ( .D(nreg[987]), .CLK(clk), .RST(rst), .I(e_init[987]), 
        .Q(nreg[987]) );
  DFF \nreg_reg[986]  ( .D(nreg[986]), .CLK(clk), .RST(rst), .I(e_init[986]), 
        .Q(nreg[986]) );
  DFF \nreg_reg[985]  ( .D(nreg[985]), .CLK(clk), .RST(rst), .I(e_init[985]), 
        .Q(nreg[985]) );
  DFF \nreg_reg[984]  ( .D(nreg[984]), .CLK(clk), .RST(rst), .I(e_init[984]), 
        .Q(nreg[984]) );
  DFF \nreg_reg[983]  ( .D(nreg[983]), .CLK(clk), .RST(rst), .I(e_init[983]), 
        .Q(nreg[983]) );
  DFF \nreg_reg[982]  ( .D(nreg[982]), .CLK(clk), .RST(rst), .I(e_init[982]), 
        .Q(nreg[982]) );
  DFF \nreg_reg[981]  ( .D(nreg[981]), .CLK(clk), .RST(rst), .I(e_init[981]), 
        .Q(nreg[981]) );
  DFF \nreg_reg[980]  ( .D(nreg[980]), .CLK(clk), .RST(rst), .I(e_init[980]), 
        .Q(nreg[980]) );
  DFF \nreg_reg[979]  ( .D(nreg[979]), .CLK(clk), .RST(rst), .I(e_init[979]), 
        .Q(nreg[979]) );
  DFF \nreg_reg[978]  ( .D(nreg[978]), .CLK(clk), .RST(rst), .I(e_init[978]), 
        .Q(nreg[978]) );
  DFF \nreg_reg[977]  ( .D(nreg[977]), .CLK(clk), .RST(rst), .I(e_init[977]), 
        .Q(nreg[977]) );
  DFF \nreg_reg[976]  ( .D(nreg[976]), .CLK(clk), .RST(rst), .I(e_init[976]), 
        .Q(nreg[976]) );
  DFF \nreg_reg[975]  ( .D(nreg[975]), .CLK(clk), .RST(rst), .I(e_init[975]), 
        .Q(nreg[975]) );
  DFF \nreg_reg[974]  ( .D(nreg[974]), .CLK(clk), .RST(rst), .I(e_init[974]), 
        .Q(nreg[974]) );
  DFF \nreg_reg[973]  ( .D(nreg[973]), .CLK(clk), .RST(rst), .I(e_init[973]), 
        .Q(nreg[973]) );
  DFF \nreg_reg[972]  ( .D(nreg[972]), .CLK(clk), .RST(rst), .I(e_init[972]), 
        .Q(nreg[972]) );
  DFF \nreg_reg[971]  ( .D(nreg[971]), .CLK(clk), .RST(rst), .I(e_init[971]), 
        .Q(nreg[971]) );
  DFF \nreg_reg[970]  ( .D(nreg[970]), .CLK(clk), .RST(rst), .I(e_init[970]), 
        .Q(nreg[970]) );
  DFF \nreg_reg[969]  ( .D(nreg[969]), .CLK(clk), .RST(rst), .I(e_init[969]), 
        .Q(nreg[969]) );
  DFF \nreg_reg[968]  ( .D(nreg[968]), .CLK(clk), .RST(rst), .I(e_init[968]), 
        .Q(nreg[968]) );
  DFF \nreg_reg[967]  ( .D(nreg[967]), .CLK(clk), .RST(rst), .I(e_init[967]), 
        .Q(nreg[967]) );
  DFF \nreg_reg[966]  ( .D(nreg[966]), .CLK(clk), .RST(rst), .I(e_init[966]), 
        .Q(nreg[966]) );
  DFF \nreg_reg[965]  ( .D(nreg[965]), .CLK(clk), .RST(rst), .I(e_init[965]), 
        .Q(nreg[965]) );
  DFF \nreg_reg[964]  ( .D(nreg[964]), .CLK(clk), .RST(rst), .I(e_init[964]), 
        .Q(nreg[964]) );
  DFF \nreg_reg[963]  ( .D(nreg[963]), .CLK(clk), .RST(rst), .I(e_init[963]), 
        .Q(nreg[963]) );
  DFF \nreg_reg[962]  ( .D(nreg[962]), .CLK(clk), .RST(rst), .I(e_init[962]), 
        .Q(nreg[962]) );
  DFF \nreg_reg[961]  ( .D(nreg[961]), .CLK(clk), .RST(rst), .I(e_init[961]), 
        .Q(nreg[961]) );
  DFF \nreg_reg[960]  ( .D(nreg[960]), .CLK(clk), .RST(rst), .I(e_init[960]), 
        .Q(nreg[960]) );
  DFF \nreg_reg[959]  ( .D(nreg[959]), .CLK(clk), .RST(rst), .I(e_init[959]), 
        .Q(nreg[959]) );
  DFF \nreg_reg[958]  ( .D(nreg[958]), .CLK(clk), .RST(rst), .I(e_init[958]), 
        .Q(nreg[958]) );
  DFF \nreg_reg[957]  ( .D(nreg[957]), .CLK(clk), .RST(rst), .I(e_init[957]), 
        .Q(nreg[957]) );
  DFF \nreg_reg[956]  ( .D(nreg[956]), .CLK(clk), .RST(rst), .I(e_init[956]), 
        .Q(nreg[956]) );
  DFF \nreg_reg[955]  ( .D(nreg[955]), .CLK(clk), .RST(rst), .I(e_init[955]), 
        .Q(nreg[955]) );
  DFF \nreg_reg[954]  ( .D(nreg[954]), .CLK(clk), .RST(rst), .I(e_init[954]), 
        .Q(nreg[954]) );
  DFF \nreg_reg[953]  ( .D(nreg[953]), .CLK(clk), .RST(rst), .I(e_init[953]), 
        .Q(nreg[953]) );
  DFF \nreg_reg[952]  ( .D(nreg[952]), .CLK(clk), .RST(rst), .I(e_init[952]), 
        .Q(nreg[952]) );
  DFF \nreg_reg[951]  ( .D(nreg[951]), .CLK(clk), .RST(rst), .I(e_init[951]), 
        .Q(nreg[951]) );
  DFF \nreg_reg[950]  ( .D(nreg[950]), .CLK(clk), .RST(rst), .I(e_init[950]), 
        .Q(nreg[950]) );
  DFF \nreg_reg[949]  ( .D(nreg[949]), .CLK(clk), .RST(rst), .I(e_init[949]), 
        .Q(nreg[949]) );
  DFF \nreg_reg[948]  ( .D(nreg[948]), .CLK(clk), .RST(rst), .I(e_init[948]), 
        .Q(nreg[948]) );
  DFF \nreg_reg[947]  ( .D(nreg[947]), .CLK(clk), .RST(rst), .I(e_init[947]), 
        .Q(nreg[947]) );
  DFF \nreg_reg[946]  ( .D(nreg[946]), .CLK(clk), .RST(rst), .I(e_init[946]), 
        .Q(nreg[946]) );
  DFF \nreg_reg[945]  ( .D(nreg[945]), .CLK(clk), .RST(rst), .I(e_init[945]), 
        .Q(nreg[945]) );
  DFF \nreg_reg[944]  ( .D(nreg[944]), .CLK(clk), .RST(rst), .I(e_init[944]), 
        .Q(nreg[944]) );
  DFF \nreg_reg[943]  ( .D(nreg[943]), .CLK(clk), .RST(rst), .I(e_init[943]), 
        .Q(nreg[943]) );
  DFF \nreg_reg[942]  ( .D(nreg[942]), .CLK(clk), .RST(rst), .I(e_init[942]), 
        .Q(nreg[942]) );
  DFF \nreg_reg[941]  ( .D(nreg[941]), .CLK(clk), .RST(rst), .I(e_init[941]), 
        .Q(nreg[941]) );
  DFF \nreg_reg[940]  ( .D(nreg[940]), .CLK(clk), .RST(rst), .I(e_init[940]), 
        .Q(nreg[940]) );
  DFF \nreg_reg[939]  ( .D(nreg[939]), .CLK(clk), .RST(rst), .I(e_init[939]), 
        .Q(nreg[939]) );
  DFF \nreg_reg[938]  ( .D(nreg[938]), .CLK(clk), .RST(rst), .I(e_init[938]), 
        .Q(nreg[938]) );
  DFF \nreg_reg[937]  ( .D(nreg[937]), .CLK(clk), .RST(rst), .I(e_init[937]), 
        .Q(nreg[937]) );
  DFF \nreg_reg[936]  ( .D(nreg[936]), .CLK(clk), .RST(rst), .I(e_init[936]), 
        .Q(nreg[936]) );
  DFF \nreg_reg[935]  ( .D(nreg[935]), .CLK(clk), .RST(rst), .I(e_init[935]), 
        .Q(nreg[935]) );
  DFF \nreg_reg[934]  ( .D(nreg[934]), .CLK(clk), .RST(rst), .I(e_init[934]), 
        .Q(nreg[934]) );
  DFF \nreg_reg[933]  ( .D(nreg[933]), .CLK(clk), .RST(rst), .I(e_init[933]), 
        .Q(nreg[933]) );
  DFF \nreg_reg[932]  ( .D(nreg[932]), .CLK(clk), .RST(rst), .I(e_init[932]), 
        .Q(nreg[932]) );
  DFF \nreg_reg[931]  ( .D(nreg[931]), .CLK(clk), .RST(rst), .I(e_init[931]), 
        .Q(nreg[931]) );
  DFF \nreg_reg[930]  ( .D(nreg[930]), .CLK(clk), .RST(rst), .I(e_init[930]), 
        .Q(nreg[930]) );
  DFF \nreg_reg[929]  ( .D(nreg[929]), .CLK(clk), .RST(rst), .I(e_init[929]), 
        .Q(nreg[929]) );
  DFF \nreg_reg[928]  ( .D(nreg[928]), .CLK(clk), .RST(rst), .I(e_init[928]), 
        .Q(nreg[928]) );
  DFF \nreg_reg[927]  ( .D(nreg[927]), .CLK(clk), .RST(rst), .I(e_init[927]), 
        .Q(nreg[927]) );
  DFF \nreg_reg[926]  ( .D(nreg[926]), .CLK(clk), .RST(rst), .I(e_init[926]), 
        .Q(nreg[926]) );
  DFF \nreg_reg[925]  ( .D(nreg[925]), .CLK(clk), .RST(rst), .I(e_init[925]), 
        .Q(nreg[925]) );
  DFF \nreg_reg[924]  ( .D(nreg[924]), .CLK(clk), .RST(rst), .I(e_init[924]), 
        .Q(nreg[924]) );
  DFF \nreg_reg[923]  ( .D(nreg[923]), .CLK(clk), .RST(rst), .I(e_init[923]), 
        .Q(nreg[923]) );
  DFF \nreg_reg[922]  ( .D(nreg[922]), .CLK(clk), .RST(rst), .I(e_init[922]), 
        .Q(nreg[922]) );
  DFF \nreg_reg[921]  ( .D(nreg[921]), .CLK(clk), .RST(rst), .I(e_init[921]), 
        .Q(nreg[921]) );
  DFF \nreg_reg[920]  ( .D(nreg[920]), .CLK(clk), .RST(rst), .I(e_init[920]), 
        .Q(nreg[920]) );
  DFF \nreg_reg[919]  ( .D(nreg[919]), .CLK(clk), .RST(rst), .I(e_init[919]), 
        .Q(nreg[919]) );
  DFF \nreg_reg[918]  ( .D(nreg[918]), .CLK(clk), .RST(rst), .I(e_init[918]), 
        .Q(nreg[918]) );
  DFF \nreg_reg[917]  ( .D(nreg[917]), .CLK(clk), .RST(rst), .I(e_init[917]), 
        .Q(nreg[917]) );
  DFF \nreg_reg[916]  ( .D(nreg[916]), .CLK(clk), .RST(rst), .I(e_init[916]), 
        .Q(nreg[916]) );
  DFF \nreg_reg[915]  ( .D(nreg[915]), .CLK(clk), .RST(rst), .I(e_init[915]), 
        .Q(nreg[915]) );
  DFF \nreg_reg[914]  ( .D(nreg[914]), .CLK(clk), .RST(rst), .I(e_init[914]), 
        .Q(nreg[914]) );
  DFF \nreg_reg[913]  ( .D(nreg[913]), .CLK(clk), .RST(rst), .I(e_init[913]), 
        .Q(nreg[913]) );
  DFF \nreg_reg[912]  ( .D(nreg[912]), .CLK(clk), .RST(rst), .I(e_init[912]), 
        .Q(nreg[912]) );
  DFF \nreg_reg[911]  ( .D(nreg[911]), .CLK(clk), .RST(rst), .I(e_init[911]), 
        .Q(nreg[911]) );
  DFF \nreg_reg[910]  ( .D(nreg[910]), .CLK(clk), .RST(rst), .I(e_init[910]), 
        .Q(nreg[910]) );
  DFF \nreg_reg[909]  ( .D(nreg[909]), .CLK(clk), .RST(rst), .I(e_init[909]), 
        .Q(nreg[909]) );
  DFF \nreg_reg[908]  ( .D(nreg[908]), .CLK(clk), .RST(rst), .I(e_init[908]), 
        .Q(nreg[908]) );
  DFF \nreg_reg[907]  ( .D(nreg[907]), .CLK(clk), .RST(rst), .I(e_init[907]), 
        .Q(nreg[907]) );
  DFF \nreg_reg[906]  ( .D(nreg[906]), .CLK(clk), .RST(rst), .I(e_init[906]), 
        .Q(nreg[906]) );
  DFF \nreg_reg[905]  ( .D(nreg[905]), .CLK(clk), .RST(rst), .I(e_init[905]), 
        .Q(nreg[905]) );
  DFF \nreg_reg[904]  ( .D(nreg[904]), .CLK(clk), .RST(rst), .I(e_init[904]), 
        .Q(nreg[904]) );
  DFF \nreg_reg[903]  ( .D(nreg[903]), .CLK(clk), .RST(rst), .I(e_init[903]), 
        .Q(nreg[903]) );
  DFF \nreg_reg[902]  ( .D(nreg[902]), .CLK(clk), .RST(rst), .I(e_init[902]), 
        .Q(nreg[902]) );
  DFF \nreg_reg[901]  ( .D(nreg[901]), .CLK(clk), .RST(rst), .I(e_init[901]), 
        .Q(nreg[901]) );
  DFF \nreg_reg[900]  ( .D(nreg[900]), .CLK(clk), .RST(rst), .I(e_init[900]), 
        .Q(nreg[900]) );
  DFF \nreg_reg[899]  ( .D(nreg[899]), .CLK(clk), .RST(rst), .I(e_init[899]), 
        .Q(nreg[899]) );
  DFF \nreg_reg[898]  ( .D(nreg[898]), .CLK(clk), .RST(rst), .I(e_init[898]), 
        .Q(nreg[898]) );
  DFF \nreg_reg[897]  ( .D(nreg[897]), .CLK(clk), .RST(rst), .I(e_init[897]), 
        .Q(nreg[897]) );
  DFF \nreg_reg[896]  ( .D(nreg[896]), .CLK(clk), .RST(rst), .I(e_init[896]), 
        .Q(nreg[896]) );
  DFF \nreg_reg[895]  ( .D(nreg[895]), .CLK(clk), .RST(rst), .I(e_init[895]), 
        .Q(nreg[895]) );
  DFF \nreg_reg[894]  ( .D(nreg[894]), .CLK(clk), .RST(rst), .I(e_init[894]), 
        .Q(nreg[894]) );
  DFF \nreg_reg[893]  ( .D(nreg[893]), .CLK(clk), .RST(rst), .I(e_init[893]), 
        .Q(nreg[893]) );
  DFF \nreg_reg[892]  ( .D(nreg[892]), .CLK(clk), .RST(rst), .I(e_init[892]), 
        .Q(nreg[892]) );
  DFF \nreg_reg[891]  ( .D(nreg[891]), .CLK(clk), .RST(rst), .I(e_init[891]), 
        .Q(nreg[891]) );
  DFF \nreg_reg[890]  ( .D(nreg[890]), .CLK(clk), .RST(rst), .I(e_init[890]), 
        .Q(nreg[890]) );
  DFF \nreg_reg[889]  ( .D(nreg[889]), .CLK(clk), .RST(rst), .I(e_init[889]), 
        .Q(nreg[889]) );
  DFF \nreg_reg[888]  ( .D(nreg[888]), .CLK(clk), .RST(rst), .I(e_init[888]), 
        .Q(nreg[888]) );
  DFF \nreg_reg[887]  ( .D(nreg[887]), .CLK(clk), .RST(rst), .I(e_init[887]), 
        .Q(nreg[887]) );
  DFF \nreg_reg[886]  ( .D(nreg[886]), .CLK(clk), .RST(rst), .I(e_init[886]), 
        .Q(nreg[886]) );
  DFF \nreg_reg[885]  ( .D(nreg[885]), .CLK(clk), .RST(rst), .I(e_init[885]), 
        .Q(nreg[885]) );
  DFF \nreg_reg[884]  ( .D(nreg[884]), .CLK(clk), .RST(rst), .I(e_init[884]), 
        .Q(nreg[884]) );
  DFF \nreg_reg[883]  ( .D(nreg[883]), .CLK(clk), .RST(rst), .I(e_init[883]), 
        .Q(nreg[883]) );
  DFF \nreg_reg[882]  ( .D(nreg[882]), .CLK(clk), .RST(rst), .I(e_init[882]), 
        .Q(nreg[882]) );
  DFF \nreg_reg[881]  ( .D(nreg[881]), .CLK(clk), .RST(rst), .I(e_init[881]), 
        .Q(nreg[881]) );
  DFF \nreg_reg[880]  ( .D(nreg[880]), .CLK(clk), .RST(rst), .I(e_init[880]), 
        .Q(nreg[880]) );
  DFF \nreg_reg[879]  ( .D(nreg[879]), .CLK(clk), .RST(rst), .I(e_init[879]), 
        .Q(nreg[879]) );
  DFF \nreg_reg[878]  ( .D(nreg[878]), .CLK(clk), .RST(rst), .I(e_init[878]), 
        .Q(nreg[878]) );
  DFF \nreg_reg[877]  ( .D(nreg[877]), .CLK(clk), .RST(rst), .I(e_init[877]), 
        .Q(nreg[877]) );
  DFF \nreg_reg[876]  ( .D(nreg[876]), .CLK(clk), .RST(rst), .I(e_init[876]), 
        .Q(nreg[876]) );
  DFF \nreg_reg[875]  ( .D(nreg[875]), .CLK(clk), .RST(rst), .I(e_init[875]), 
        .Q(nreg[875]) );
  DFF \nreg_reg[874]  ( .D(nreg[874]), .CLK(clk), .RST(rst), .I(e_init[874]), 
        .Q(nreg[874]) );
  DFF \nreg_reg[873]  ( .D(nreg[873]), .CLK(clk), .RST(rst), .I(e_init[873]), 
        .Q(nreg[873]) );
  DFF \nreg_reg[872]  ( .D(nreg[872]), .CLK(clk), .RST(rst), .I(e_init[872]), 
        .Q(nreg[872]) );
  DFF \nreg_reg[871]  ( .D(nreg[871]), .CLK(clk), .RST(rst), .I(e_init[871]), 
        .Q(nreg[871]) );
  DFF \nreg_reg[870]  ( .D(nreg[870]), .CLK(clk), .RST(rst), .I(e_init[870]), 
        .Q(nreg[870]) );
  DFF \nreg_reg[869]  ( .D(nreg[869]), .CLK(clk), .RST(rst), .I(e_init[869]), 
        .Q(nreg[869]) );
  DFF \nreg_reg[868]  ( .D(nreg[868]), .CLK(clk), .RST(rst), .I(e_init[868]), 
        .Q(nreg[868]) );
  DFF \nreg_reg[867]  ( .D(nreg[867]), .CLK(clk), .RST(rst), .I(e_init[867]), 
        .Q(nreg[867]) );
  DFF \nreg_reg[866]  ( .D(nreg[866]), .CLK(clk), .RST(rst), .I(e_init[866]), 
        .Q(nreg[866]) );
  DFF \nreg_reg[865]  ( .D(nreg[865]), .CLK(clk), .RST(rst), .I(e_init[865]), 
        .Q(nreg[865]) );
  DFF \nreg_reg[864]  ( .D(nreg[864]), .CLK(clk), .RST(rst), .I(e_init[864]), 
        .Q(nreg[864]) );
  DFF \nreg_reg[863]  ( .D(nreg[863]), .CLK(clk), .RST(rst), .I(e_init[863]), 
        .Q(nreg[863]) );
  DFF \nreg_reg[862]  ( .D(nreg[862]), .CLK(clk), .RST(rst), .I(e_init[862]), 
        .Q(nreg[862]) );
  DFF \nreg_reg[861]  ( .D(nreg[861]), .CLK(clk), .RST(rst), .I(e_init[861]), 
        .Q(nreg[861]) );
  DFF \nreg_reg[860]  ( .D(nreg[860]), .CLK(clk), .RST(rst), .I(e_init[860]), 
        .Q(nreg[860]) );
  DFF \nreg_reg[859]  ( .D(nreg[859]), .CLK(clk), .RST(rst), .I(e_init[859]), 
        .Q(nreg[859]) );
  DFF \nreg_reg[858]  ( .D(nreg[858]), .CLK(clk), .RST(rst), .I(e_init[858]), 
        .Q(nreg[858]) );
  DFF \nreg_reg[857]  ( .D(nreg[857]), .CLK(clk), .RST(rst), .I(e_init[857]), 
        .Q(nreg[857]) );
  DFF \nreg_reg[856]  ( .D(nreg[856]), .CLK(clk), .RST(rst), .I(e_init[856]), 
        .Q(nreg[856]) );
  DFF \nreg_reg[855]  ( .D(nreg[855]), .CLK(clk), .RST(rst), .I(e_init[855]), 
        .Q(nreg[855]) );
  DFF \nreg_reg[854]  ( .D(nreg[854]), .CLK(clk), .RST(rst), .I(e_init[854]), 
        .Q(nreg[854]) );
  DFF \nreg_reg[853]  ( .D(nreg[853]), .CLK(clk), .RST(rst), .I(e_init[853]), 
        .Q(nreg[853]) );
  DFF \nreg_reg[852]  ( .D(nreg[852]), .CLK(clk), .RST(rst), .I(e_init[852]), 
        .Q(nreg[852]) );
  DFF \nreg_reg[851]  ( .D(nreg[851]), .CLK(clk), .RST(rst), .I(e_init[851]), 
        .Q(nreg[851]) );
  DFF \nreg_reg[850]  ( .D(nreg[850]), .CLK(clk), .RST(rst), .I(e_init[850]), 
        .Q(nreg[850]) );
  DFF \nreg_reg[849]  ( .D(nreg[849]), .CLK(clk), .RST(rst), .I(e_init[849]), 
        .Q(nreg[849]) );
  DFF \nreg_reg[848]  ( .D(nreg[848]), .CLK(clk), .RST(rst), .I(e_init[848]), 
        .Q(nreg[848]) );
  DFF \nreg_reg[847]  ( .D(nreg[847]), .CLK(clk), .RST(rst), .I(e_init[847]), 
        .Q(nreg[847]) );
  DFF \nreg_reg[846]  ( .D(nreg[846]), .CLK(clk), .RST(rst), .I(e_init[846]), 
        .Q(nreg[846]) );
  DFF \nreg_reg[845]  ( .D(nreg[845]), .CLK(clk), .RST(rst), .I(e_init[845]), 
        .Q(nreg[845]) );
  DFF \nreg_reg[844]  ( .D(nreg[844]), .CLK(clk), .RST(rst), .I(e_init[844]), 
        .Q(nreg[844]) );
  DFF \nreg_reg[843]  ( .D(nreg[843]), .CLK(clk), .RST(rst), .I(e_init[843]), 
        .Q(nreg[843]) );
  DFF \nreg_reg[842]  ( .D(nreg[842]), .CLK(clk), .RST(rst), .I(e_init[842]), 
        .Q(nreg[842]) );
  DFF \nreg_reg[841]  ( .D(nreg[841]), .CLK(clk), .RST(rst), .I(e_init[841]), 
        .Q(nreg[841]) );
  DFF \nreg_reg[840]  ( .D(nreg[840]), .CLK(clk), .RST(rst), .I(e_init[840]), 
        .Q(nreg[840]) );
  DFF \nreg_reg[839]  ( .D(nreg[839]), .CLK(clk), .RST(rst), .I(e_init[839]), 
        .Q(nreg[839]) );
  DFF \nreg_reg[838]  ( .D(nreg[838]), .CLK(clk), .RST(rst), .I(e_init[838]), 
        .Q(nreg[838]) );
  DFF \nreg_reg[837]  ( .D(nreg[837]), .CLK(clk), .RST(rst), .I(e_init[837]), 
        .Q(nreg[837]) );
  DFF \nreg_reg[836]  ( .D(nreg[836]), .CLK(clk), .RST(rst), .I(e_init[836]), 
        .Q(nreg[836]) );
  DFF \nreg_reg[835]  ( .D(nreg[835]), .CLK(clk), .RST(rst), .I(e_init[835]), 
        .Q(nreg[835]) );
  DFF \nreg_reg[834]  ( .D(nreg[834]), .CLK(clk), .RST(rst), .I(e_init[834]), 
        .Q(nreg[834]) );
  DFF \nreg_reg[833]  ( .D(nreg[833]), .CLK(clk), .RST(rst), .I(e_init[833]), 
        .Q(nreg[833]) );
  DFF \nreg_reg[832]  ( .D(nreg[832]), .CLK(clk), .RST(rst), .I(e_init[832]), 
        .Q(nreg[832]) );
  DFF \nreg_reg[831]  ( .D(nreg[831]), .CLK(clk), .RST(rst), .I(e_init[831]), 
        .Q(nreg[831]) );
  DFF \nreg_reg[830]  ( .D(nreg[830]), .CLK(clk), .RST(rst), .I(e_init[830]), 
        .Q(nreg[830]) );
  DFF \nreg_reg[829]  ( .D(nreg[829]), .CLK(clk), .RST(rst), .I(e_init[829]), 
        .Q(nreg[829]) );
  DFF \nreg_reg[828]  ( .D(nreg[828]), .CLK(clk), .RST(rst), .I(e_init[828]), 
        .Q(nreg[828]) );
  DFF \nreg_reg[827]  ( .D(nreg[827]), .CLK(clk), .RST(rst), .I(e_init[827]), 
        .Q(nreg[827]) );
  DFF \nreg_reg[826]  ( .D(nreg[826]), .CLK(clk), .RST(rst), .I(e_init[826]), 
        .Q(nreg[826]) );
  DFF \nreg_reg[825]  ( .D(nreg[825]), .CLK(clk), .RST(rst), .I(e_init[825]), 
        .Q(nreg[825]) );
  DFF \nreg_reg[824]  ( .D(nreg[824]), .CLK(clk), .RST(rst), .I(e_init[824]), 
        .Q(nreg[824]) );
  DFF \nreg_reg[823]  ( .D(nreg[823]), .CLK(clk), .RST(rst), .I(e_init[823]), 
        .Q(nreg[823]) );
  DFF \nreg_reg[822]  ( .D(nreg[822]), .CLK(clk), .RST(rst), .I(e_init[822]), 
        .Q(nreg[822]) );
  DFF \nreg_reg[821]  ( .D(nreg[821]), .CLK(clk), .RST(rst), .I(e_init[821]), 
        .Q(nreg[821]) );
  DFF \nreg_reg[820]  ( .D(nreg[820]), .CLK(clk), .RST(rst), .I(e_init[820]), 
        .Q(nreg[820]) );
  DFF \nreg_reg[819]  ( .D(nreg[819]), .CLK(clk), .RST(rst), .I(e_init[819]), 
        .Q(nreg[819]) );
  DFF \nreg_reg[818]  ( .D(nreg[818]), .CLK(clk), .RST(rst), .I(e_init[818]), 
        .Q(nreg[818]) );
  DFF \nreg_reg[817]  ( .D(nreg[817]), .CLK(clk), .RST(rst), .I(e_init[817]), 
        .Q(nreg[817]) );
  DFF \nreg_reg[816]  ( .D(nreg[816]), .CLK(clk), .RST(rst), .I(e_init[816]), 
        .Q(nreg[816]) );
  DFF \nreg_reg[815]  ( .D(nreg[815]), .CLK(clk), .RST(rst), .I(e_init[815]), 
        .Q(nreg[815]) );
  DFF \nreg_reg[814]  ( .D(nreg[814]), .CLK(clk), .RST(rst), .I(e_init[814]), 
        .Q(nreg[814]) );
  DFF \nreg_reg[813]  ( .D(nreg[813]), .CLK(clk), .RST(rst), .I(e_init[813]), 
        .Q(nreg[813]) );
  DFF \nreg_reg[812]  ( .D(nreg[812]), .CLK(clk), .RST(rst), .I(e_init[812]), 
        .Q(nreg[812]) );
  DFF \nreg_reg[811]  ( .D(nreg[811]), .CLK(clk), .RST(rst), .I(e_init[811]), 
        .Q(nreg[811]) );
  DFF \nreg_reg[810]  ( .D(nreg[810]), .CLK(clk), .RST(rst), .I(e_init[810]), 
        .Q(nreg[810]) );
  DFF \nreg_reg[809]  ( .D(nreg[809]), .CLK(clk), .RST(rst), .I(e_init[809]), 
        .Q(nreg[809]) );
  DFF \nreg_reg[808]  ( .D(nreg[808]), .CLK(clk), .RST(rst), .I(e_init[808]), 
        .Q(nreg[808]) );
  DFF \nreg_reg[807]  ( .D(nreg[807]), .CLK(clk), .RST(rst), .I(e_init[807]), 
        .Q(nreg[807]) );
  DFF \nreg_reg[806]  ( .D(nreg[806]), .CLK(clk), .RST(rst), .I(e_init[806]), 
        .Q(nreg[806]) );
  DFF \nreg_reg[805]  ( .D(nreg[805]), .CLK(clk), .RST(rst), .I(e_init[805]), 
        .Q(nreg[805]) );
  DFF \nreg_reg[804]  ( .D(nreg[804]), .CLK(clk), .RST(rst), .I(e_init[804]), 
        .Q(nreg[804]) );
  DFF \nreg_reg[803]  ( .D(nreg[803]), .CLK(clk), .RST(rst), .I(e_init[803]), 
        .Q(nreg[803]) );
  DFF \nreg_reg[802]  ( .D(nreg[802]), .CLK(clk), .RST(rst), .I(e_init[802]), 
        .Q(nreg[802]) );
  DFF \nreg_reg[801]  ( .D(nreg[801]), .CLK(clk), .RST(rst), .I(e_init[801]), 
        .Q(nreg[801]) );
  DFF \nreg_reg[800]  ( .D(nreg[800]), .CLK(clk), .RST(rst), .I(e_init[800]), 
        .Q(nreg[800]) );
  DFF \nreg_reg[799]  ( .D(nreg[799]), .CLK(clk), .RST(rst), .I(e_init[799]), 
        .Q(nreg[799]) );
  DFF \nreg_reg[798]  ( .D(nreg[798]), .CLK(clk), .RST(rst), .I(e_init[798]), 
        .Q(nreg[798]) );
  DFF \nreg_reg[797]  ( .D(nreg[797]), .CLK(clk), .RST(rst), .I(e_init[797]), 
        .Q(nreg[797]) );
  DFF \nreg_reg[796]  ( .D(nreg[796]), .CLK(clk), .RST(rst), .I(e_init[796]), 
        .Q(nreg[796]) );
  DFF \nreg_reg[795]  ( .D(nreg[795]), .CLK(clk), .RST(rst), .I(e_init[795]), 
        .Q(nreg[795]) );
  DFF \nreg_reg[794]  ( .D(nreg[794]), .CLK(clk), .RST(rst), .I(e_init[794]), 
        .Q(nreg[794]) );
  DFF \nreg_reg[793]  ( .D(nreg[793]), .CLK(clk), .RST(rst), .I(e_init[793]), 
        .Q(nreg[793]) );
  DFF \nreg_reg[792]  ( .D(nreg[792]), .CLK(clk), .RST(rst), .I(e_init[792]), 
        .Q(nreg[792]) );
  DFF \nreg_reg[791]  ( .D(nreg[791]), .CLK(clk), .RST(rst), .I(e_init[791]), 
        .Q(nreg[791]) );
  DFF \nreg_reg[790]  ( .D(nreg[790]), .CLK(clk), .RST(rst), .I(e_init[790]), 
        .Q(nreg[790]) );
  DFF \nreg_reg[789]  ( .D(nreg[789]), .CLK(clk), .RST(rst), .I(e_init[789]), 
        .Q(nreg[789]) );
  DFF \nreg_reg[788]  ( .D(nreg[788]), .CLK(clk), .RST(rst), .I(e_init[788]), 
        .Q(nreg[788]) );
  DFF \nreg_reg[787]  ( .D(nreg[787]), .CLK(clk), .RST(rst), .I(e_init[787]), 
        .Q(nreg[787]) );
  DFF \nreg_reg[786]  ( .D(nreg[786]), .CLK(clk), .RST(rst), .I(e_init[786]), 
        .Q(nreg[786]) );
  DFF \nreg_reg[785]  ( .D(nreg[785]), .CLK(clk), .RST(rst), .I(e_init[785]), 
        .Q(nreg[785]) );
  DFF \nreg_reg[784]  ( .D(nreg[784]), .CLK(clk), .RST(rst), .I(e_init[784]), 
        .Q(nreg[784]) );
  DFF \nreg_reg[783]  ( .D(nreg[783]), .CLK(clk), .RST(rst), .I(e_init[783]), 
        .Q(nreg[783]) );
  DFF \nreg_reg[782]  ( .D(nreg[782]), .CLK(clk), .RST(rst), .I(e_init[782]), 
        .Q(nreg[782]) );
  DFF \nreg_reg[781]  ( .D(nreg[781]), .CLK(clk), .RST(rst), .I(e_init[781]), 
        .Q(nreg[781]) );
  DFF \nreg_reg[780]  ( .D(nreg[780]), .CLK(clk), .RST(rst), .I(e_init[780]), 
        .Q(nreg[780]) );
  DFF \nreg_reg[779]  ( .D(nreg[779]), .CLK(clk), .RST(rst), .I(e_init[779]), 
        .Q(nreg[779]) );
  DFF \nreg_reg[778]  ( .D(nreg[778]), .CLK(clk), .RST(rst), .I(e_init[778]), 
        .Q(nreg[778]) );
  DFF \nreg_reg[777]  ( .D(nreg[777]), .CLK(clk), .RST(rst), .I(e_init[777]), 
        .Q(nreg[777]) );
  DFF \nreg_reg[776]  ( .D(nreg[776]), .CLK(clk), .RST(rst), .I(e_init[776]), 
        .Q(nreg[776]) );
  DFF \nreg_reg[775]  ( .D(nreg[775]), .CLK(clk), .RST(rst), .I(e_init[775]), 
        .Q(nreg[775]) );
  DFF \nreg_reg[774]  ( .D(nreg[774]), .CLK(clk), .RST(rst), .I(e_init[774]), 
        .Q(nreg[774]) );
  DFF \nreg_reg[773]  ( .D(nreg[773]), .CLK(clk), .RST(rst), .I(e_init[773]), 
        .Q(nreg[773]) );
  DFF \nreg_reg[772]  ( .D(nreg[772]), .CLK(clk), .RST(rst), .I(e_init[772]), 
        .Q(nreg[772]) );
  DFF \nreg_reg[771]  ( .D(nreg[771]), .CLK(clk), .RST(rst), .I(e_init[771]), 
        .Q(nreg[771]) );
  DFF \nreg_reg[770]  ( .D(nreg[770]), .CLK(clk), .RST(rst), .I(e_init[770]), 
        .Q(nreg[770]) );
  DFF \nreg_reg[769]  ( .D(nreg[769]), .CLK(clk), .RST(rst), .I(e_init[769]), 
        .Q(nreg[769]) );
  DFF \nreg_reg[768]  ( .D(nreg[768]), .CLK(clk), .RST(rst), .I(e_init[768]), 
        .Q(nreg[768]) );
  DFF \nreg_reg[767]  ( .D(nreg[767]), .CLK(clk), .RST(rst), .I(e_init[767]), 
        .Q(nreg[767]) );
  DFF \nreg_reg[766]  ( .D(nreg[766]), .CLK(clk), .RST(rst), .I(e_init[766]), 
        .Q(nreg[766]) );
  DFF \nreg_reg[765]  ( .D(nreg[765]), .CLK(clk), .RST(rst), .I(e_init[765]), 
        .Q(nreg[765]) );
  DFF \nreg_reg[764]  ( .D(nreg[764]), .CLK(clk), .RST(rst), .I(e_init[764]), 
        .Q(nreg[764]) );
  DFF \nreg_reg[763]  ( .D(nreg[763]), .CLK(clk), .RST(rst), .I(e_init[763]), 
        .Q(nreg[763]) );
  DFF \nreg_reg[762]  ( .D(nreg[762]), .CLK(clk), .RST(rst), .I(e_init[762]), 
        .Q(nreg[762]) );
  DFF \nreg_reg[761]  ( .D(nreg[761]), .CLK(clk), .RST(rst), .I(e_init[761]), 
        .Q(nreg[761]) );
  DFF \nreg_reg[760]  ( .D(nreg[760]), .CLK(clk), .RST(rst), .I(e_init[760]), 
        .Q(nreg[760]) );
  DFF \nreg_reg[759]  ( .D(nreg[759]), .CLK(clk), .RST(rst), .I(e_init[759]), 
        .Q(nreg[759]) );
  DFF \nreg_reg[758]  ( .D(nreg[758]), .CLK(clk), .RST(rst), .I(e_init[758]), 
        .Q(nreg[758]) );
  DFF \nreg_reg[757]  ( .D(nreg[757]), .CLK(clk), .RST(rst), .I(e_init[757]), 
        .Q(nreg[757]) );
  DFF \nreg_reg[756]  ( .D(nreg[756]), .CLK(clk), .RST(rst), .I(e_init[756]), 
        .Q(nreg[756]) );
  DFF \nreg_reg[755]  ( .D(nreg[755]), .CLK(clk), .RST(rst), .I(e_init[755]), 
        .Q(nreg[755]) );
  DFF \nreg_reg[754]  ( .D(nreg[754]), .CLK(clk), .RST(rst), .I(e_init[754]), 
        .Q(nreg[754]) );
  DFF \nreg_reg[753]  ( .D(nreg[753]), .CLK(clk), .RST(rst), .I(e_init[753]), 
        .Q(nreg[753]) );
  DFF \nreg_reg[752]  ( .D(nreg[752]), .CLK(clk), .RST(rst), .I(e_init[752]), 
        .Q(nreg[752]) );
  DFF \nreg_reg[751]  ( .D(nreg[751]), .CLK(clk), .RST(rst), .I(e_init[751]), 
        .Q(nreg[751]) );
  DFF \nreg_reg[750]  ( .D(nreg[750]), .CLK(clk), .RST(rst), .I(e_init[750]), 
        .Q(nreg[750]) );
  DFF \nreg_reg[749]  ( .D(nreg[749]), .CLK(clk), .RST(rst), .I(e_init[749]), 
        .Q(nreg[749]) );
  DFF \nreg_reg[748]  ( .D(nreg[748]), .CLK(clk), .RST(rst), .I(e_init[748]), 
        .Q(nreg[748]) );
  DFF \nreg_reg[747]  ( .D(nreg[747]), .CLK(clk), .RST(rst), .I(e_init[747]), 
        .Q(nreg[747]) );
  DFF \nreg_reg[746]  ( .D(nreg[746]), .CLK(clk), .RST(rst), .I(e_init[746]), 
        .Q(nreg[746]) );
  DFF \nreg_reg[745]  ( .D(nreg[745]), .CLK(clk), .RST(rst), .I(e_init[745]), 
        .Q(nreg[745]) );
  DFF \nreg_reg[744]  ( .D(nreg[744]), .CLK(clk), .RST(rst), .I(e_init[744]), 
        .Q(nreg[744]) );
  DFF \nreg_reg[743]  ( .D(nreg[743]), .CLK(clk), .RST(rst), .I(e_init[743]), 
        .Q(nreg[743]) );
  DFF \nreg_reg[742]  ( .D(nreg[742]), .CLK(clk), .RST(rst), .I(e_init[742]), 
        .Q(nreg[742]) );
  DFF \nreg_reg[741]  ( .D(nreg[741]), .CLK(clk), .RST(rst), .I(e_init[741]), 
        .Q(nreg[741]) );
  DFF \nreg_reg[740]  ( .D(nreg[740]), .CLK(clk), .RST(rst), .I(e_init[740]), 
        .Q(nreg[740]) );
  DFF \nreg_reg[739]  ( .D(nreg[739]), .CLK(clk), .RST(rst), .I(e_init[739]), 
        .Q(nreg[739]) );
  DFF \nreg_reg[738]  ( .D(nreg[738]), .CLK(clk), .RST(rst), .I(e_init[738]), 
        .Q(nreg[738]) );
  DFF \nreg_reg[737]  ( .D(nreg[737]), .CLK(clk), .RST(rst), .I(e_init[737]), 
        .Q(nreg[737]) );
  DFF \nreg_reg[736]  ( .D(nreg[736]), .CLK(clk), .RST(rst), .I(e_init[736]), 
        .Q(nreg[736]) );
  DFF \nreg_reg[735]  ( .D(nreg[735]), .CLK(clk), .RST(rst), .I(e_init[735]), 
        .Q(nreg[735]) );
  DFF \nreg_reg[734]  ( .D(nreg[734]), .CLK(clk), .RST(rst), .I(e_init[734]), 
        .Q(nreg[734]) );
  DFF \nreg_reg[733]  ( .D(nreg[733]), .CLK(clk), .RST(rst), .I(e_init[733]), 
        .Q(nreg[733]) );
  DFF \nreg_reg[732]  ( .D(nreg[732]), .CLK(clk), .RST(rst), .I(e_init[732]), 
        .Q(nreg[732]) );
  DFF \nreg_reg[731]  ( .D(nreg[731]), .CLK(clk), .RST(rst), .I(e_init[731]), 
        .Q(nreg[731]) );
  DFF \nreg_reg[730]  ( .D(nreg[730]), .CLK(clk), .RST(rst), .I(e_init[730]), 
        .Q(nreg[730]) );
  DFF \nreg_reg[729]  ( .D(nreg[729]), .CLK(clk), .RST(rst), .I(e_init[729]), 
        .Q(nreg[729]) );
  DFF \nreg_reg[728]  ( .D(nreg[728]), .CLK(clk), .RST(rst), .I(e_init[728]), 
        .Q(nreg[728]) );
  DFF \nreg_reg[727]  ( .D(nreg[727]), .CLK(clk), .RST(rst), .I(e_init[727]), 
        .Q(nreg[727]) );
  DFF \nreg_reg[726]  ( .D(nreg[726]), .CLK(clk), .RST(rst), .I(e_init[726]), 
        .Q(nreg[726]) );
  DFF \nreg_reg[725]  ( .D(nreg[725]), .CLK(clk), .RST(rst), .I(e_init[725]), 
        .Q(nreg[725]) );
  DFF \nreg_reg[724]  ( .D(nreg[724]), .CLK(clk), .RST(rst), .I(e_init[724]), 
        .Q(nreg[724]) );
  DFF \nreg_reg[723]  ( .D(nreg[723]), .CLK(clk), .RST(rst), .I(e_init[723]), 
        .Q(nreg[723]) );
  DFF \nreg_reg[722]  ( .D(nreg[722]), .CLK(clk), .RST(rst), .I(e_init[722]), 
        .Q(nreg[722]) );
  DFF \nreg_reg[721]  ( .D(nreg[721]), .CLK(clk), .RST(rst), .I(e_init[721]), 
        .Q(nreg[721]) );
  DFF \nreg_reg[720]  ( .D(nreg[720]), .CLK(clk), .RST(rst), .I(e_init[720]), 
        .Q(nreg[720]) );
  DFF \nreg_reg[719]  ( .D(nreg[719]), .CLK(clk), .RST(rst), .I(e_init[719]), 
        .Q(nreg[719]) );
  DFF \nreg_reg[718]  ( .D(nreg[718]), .CLK(clk), .RST(rst), .I(e_init[718]), 
        .Q(nreg[718]) );
  DFF \nreg_reg[717]  ( .D(nreg[717]), .CLK(clk), .RST(rst), .I(e_init[717]), 
        .Q(nreg[717]) );
  DFF \nreg_reg[716]  ( .D(nreg[716]), .CLK(clk), .RST(rst), .I(e_init[716]), 
        .Q(nreg[716]) );
  DFF \nreg_reg[715]  ( .D(nreg[715]), .CLK(clk), .RST(rst), .I(e_init[715]), 
        .Q(nreg[715]) );
  DFF \nreg_reg[714]  ( .D(nreg[714]), .CLK(clk), .RST(rst), .I(e_init[714]), 
        .Q(nreg[714]) );
  DFF \nreg_reg[713]  ( .D(nreg[713]), .CLK(clk), .RST(rst), .I(e_init[713]), 
        .Q(nreg[713]) );
  DFF \nreg_reg[712]  ( .D(nreg[712]), .CLK(clk), .RST(rst), .I(e_init[712]), 
        .Q(nreg[712]) );
  DFF \nreg_reg[711]  ( .D(nreg[711]), .CLK(clk), .RST(rst), .I(e_init[711]), 
        .Q(nreg[711]) );
  DFF \nreg_reg[710]  ( .D(nreg[710]), .CLK(clk), .RST(rst), .I(e_init[710]), 
        .Q(nreg[710]) );
  DFF \nreg_reg[709]  ( .D(nreg[709]), .CLK(clk), .RST(rst), .I(e_init[709]), 
        .Q(nreg[709]) );
  DFF \nreg_reg[708]  ( .D(nreg[708]), .CLK(clk), .RST(rst), .I(e_init[708]), 
        .Q(nreg[708]) );
  DFF \nreg_reg[707]  ( .D(nreg[707]), .CLK(clk), .RST(rst), .I(e_init[707]), 
        .Q(nreg[707]) );
  DFF \nreg_reg[706]  ( .D(nreg[706]), .CLK(clk), .RST(rst), .I(e_init[706]), 
        .Q(nreg[706]) );
  DFF \nreg_reg[705]  ( .D(nreg[705]), .CLK(clk), .RST(rst), .I(e_init[705]), 
        .Q(nreg[705]) );
  DFF \nreg_reg[704]  ( .D(nreg[704]), .CLK(clk), .RST(rst), .I(e_init[704]), 
        .Q(nreg[704]) );
  DFF \nreg_reg[703]  ( .D(nreg[703]), .CLK(clk), .RST(rst), .I(e_init[703]), 
        .Q(nreg[703]) );
  DFF \nreg_reg[702]  ( .D(nreg[702]), .CLK(clk), .RST(rst), .I(e_init[702]), 
        .Q(nreg[702]) );
  DFF \nreg_reg[701]  ( .D(nreg[701]), .CLK(clk), .RST(rst), .I(e_init[701]), 
        .Q(nreg[701]) );
  DFF \nreg_reg[700]  ( .D(nreg[700]), .CLK(clk), .RST(rst), .I(e_init[700]), 
        .Q(nreg[700]) );
  DFF \nreg_reg[699]  ( .D(nreg[699]), .CLK(clk), .RST(rst), .I(e_init[699]), 
        .Q(nreg[699]) );
  DFF \nreg_reg[698]  ( .D(nreg[698]), .CLK(clk), .RST(rst), .I(e_init[698]), 
        .Q(nreg[698]) );
  DFF \nreg_reg[697]  ( .D(nreg[697]), .CLK(clk), .RST(rst), .I(e_init[697]), 
        .Q(nreg[697]) );
  DFF \nreg_reg[696]  ( .D(nreg[696]), .CLK(clk), .RST(rst), .I(e_init[696]), 
        .Q(nreg[696]) );
  DFF \nreg_reg[695]  ( .D(nreg[695]), .CLK(clk), .RST(rst), .I(e_init[695]), 
        .Q(nreg[695]) );
  DFF \nreg_reg[694]  ( .D(nreg[694]), .CLK(clk), .RST(rst), .I(e_init[694]), 
        .Q(nreg[694]) );
  DFF \nreg_reg[693]  ( .D(nreg[693]), .CLK(clk), .RST(rst), .I(e_init[693]), 
        .Q(nreg[693]) );
  DFF \nreg_reg[692]  ( .D(nreg[692]), .CLK(clk), .RST(rst), .I(e_init[692]), 
        .Q(nreg[692]) );
  DFF \nreg_reg[691]  ( .D(nreg[691]), .CLK(clk), .RST(rst), .I(e_init[691]), 
        .Q(nreg[691]) );
  DFF \nreg_reg[690]  ( .D(nreg[690]), .CLK(clk), .RST(rst), .I(e_init[690]), 
        .Q(nreg[690]) );
  DFF \nreg_reg[689]  ( .D(nreg[689]), .CLK(clk), .RST(rst), .I(e_init[689]), 
        .Q(nreg[689]) );
  DFF \nreg_reg[688]  ( .D(nreg[688]), .CLK(clk), .RST(rst), .I(e_init[688]), 
        .Q(nreg[688]) );
  DFF \nreg_reg[687]  ( .D(nreg[687]), .CLK(clk), .RST(rst), .I(e_init[687]), 
        .Q(nreg[687]) );
  DFF \nreg_reg[686]  ( .D(nreg[686]), .CLK(clk), .RST(rst), .I(e_init[686]), 
        .Q(nreg[686]) );
  DFF \nreg_reg[685]  ( .D(nreg[685]), .CLK(clk), .RST(rst), .I(e_init[685]), 
        .Q(nreg[685]) );
  DFF \nreg_reg[684]  ( .D(nreg[684]), .CLK(clk), .RST(rst), .I(e_init[684]), 
        .Q(nreg[684]) );
  DFF \nreg_reg[683]  ( .D(nreg[683]), .CLK(clk), .RST(rst), .I(e_init[683]), 
        .Q(nreg[683]) );
  DFF \nreg_reg[682]  ( .D(nreg[682]), .CLK(clk), .RST(rst), .I(e_init[682]), 
        .Q(nreg[682]) );
  DFF \nreg_reg[681]  ( .D(nreg[681]), .CLK(clk), .RST(rst), .I(e_init[681]), 
        .Q(nreg[681]) );
  DFF \nreg_reg[680]  ( .D(nreg[680]), .CLK(clk), .RST(rst), .I(e_init[680]), 
        .Q(nreg[680]) );
  DFF \nreg_reg[679]  ( .D(nreg[679]), .CLK(clk), .RST(rst), .I(e_init[679]), 
        .Q(nreg[679]) );
  DFF \nreg_reg[678]  ( .D(nreg[678]), .CLK(clk), .RST(rst), .I(e_init[678]), 
        .Q(nreg[678]) );
  DFF \nreg_reg[677]  ( .D(nreg[677]), .CLK(clk), .RST(rst), .I(e_init[677]), 
        .Q(nreg[677]) );
  DFF \nreg_reg[676]  ( .D(nreg[676]), .CLK(clk), .RST(rst), .I(e_init[676]), 
        .Q(nreg[676]) );
  DFF \nreg_reg[675]  ( .D(nreg[675]), .CLK(clk), .RST(rst), .I(e_init[675]), 
        .Q(nreg[675]) );
  DFF \nreg_reg[674]  ( .D(nreg[674]), .CLK(clk), .RST(rst), .I(e_init[674]), 
        .Q(nreg[674]) );
  DFF \nreg_reg[673]  ( .D(nreg[673]), .CLK(clk), .RST(rst), .I(e_init[673]), 
        .Q(nreg[673]) );
  DFF \nreg_reg[672]  ( .D(nreg[672]), .CLK(clk), .RST(rst), .I(e_init[672]), 
        .Q(nreg[672]) );
  DFF \nreg_reg[671]  ( .D(nreg[671]), .CLK(clk), .RST(rst), .I(e_init[671]), 
        .Q(nreg[671]) );
  DFF \nreg_reg[670]  ( .D(nreg[670]), .CLK(clk), .RST(rst), .I(e_init[670]), 
        .Q(nreg[670]) );
  DFF \nreg_reg[669]  ( .D(nreg[669]), .CLK(clk), .RST(rst), .I(e_init[669]), 
        .Q(nreg[669]) );
  DFF \nreg_reg[668]  ( .D(nreg[668]), .CLK(clk), .RST(rst), .I(e_init[668]), 
        .Q(nreg[668]) );
  DFF \nreg_reg[667]  ( .D(nreg[667]), .CLK(clk), .RST(rst), .I(e_init[667]), 
        .Q(nreg[667]) );
  DFF \nreg_reg[666]  ( .D(nreg[666]), .CLK(clk), .RST(rst), .I(e_init[666]), 
        .Q(nreg[666]) );
  DFF \nreg_reg[665]  ( .D(nreg[665]), .CLK(clk), .RST(rst), .I(e_init[665]), 
        .Q(nreg[665]) );
  DFF \nreg_reg[664]  ( .D(nreg[664]), .CLK(clk), .RST(rst), .I(e_init[664]), 
        .Q(nreg[664]) );
  DFF \nreg_reg[663]  ( .D(nreg[663]), .CLK(clk), .RST(rst), .I(e_init[663]), 
        .Q(nreg[663]) );
  DFF \nreg_reg[662]  ( .D(nreg[662]), .CLK(clk), .RST(rst), .I(e_init[662]), 
        .Q(nreg[662]) );
  DFF \nreg_reg[661]  ( .D(nreg[661]), .CLK(clk), .RST(rst), .I(e_init[661]), 
        .Q(nreg[661]) );
  DFF \nreg_reg[660]  ( .D(nreg[660]), .CLK(clk), .RST(rst), .I(e_init[660]), 
        .Q(nreg[660]) );
  DFF \nreg_reg[659]  ( .D(nreg[659]), .CLK(clk), .RST(rst), .I(e_init[659]), 
        .Q(nreg[659]) );
  DFF \nreg_reg[658]  ( .D(nreg[658]), .CLK(clk), .RST(rst), .I(e_init[658]), 
        .Q(nreg[658]) );
  DFF \nreg_reg[657]  ( .D(nreg[657]), .CLK(clk), .RST(rst), .I(e_init[657]), 
        .Q(nreg[657]) );
  DFF \nreg_reg[656]  ( .D(nreg[656]), .CLK(clk), .RST(rst), .I(e_init[656]), 
        .Q(nreg[656]) );
  DFF \nreg_reg[655]  ( .D(nreg[655]), .CLK(clk), .RST(rst), .I(e_init[655]), 
        .Q(nreg[655]) );
  DFF \nreg_reg[654]  ( .D(nreg[654]), .CLK(clk), .RST(rst), .I(e_init[654]), 
        .Q(nreg[654]) );
  DFF \nreg_reg[653]  ( .D(nreg[653]), .CLK(clk), .RST(rst), .I(e_init[653]), 
        .Q(nreg[653]) );
  DFF \nreg_reg[652]  ( .D(nreg[652]), .CLK(clk), .RST(rst), .I(e_init[652]), 
        .Q(nreg[652]) );
  DFF \nreg_reg[651]  ( .D(nreg[651]), .CLK(clk), .RST(rst), .I(e_init[651]), 
        .Q(nreg[651]) );
  DFF \nreg_reg[650]  ( .D(nreg[650]), .CLK(clk), .RST(rst), .I(e_init[650]), 
        .Q(nreg[650]) );
  DFF \nreg_reg[649]  ( .D(nreg[649]), .CLK(clk), .RST(rst), .I(e_init[649]), 
        .Q(nreg[649]) );
  DFF \nreg_reg[648]  ( .D(nreg[648]), .CLK(clk), .RST(rst), .I(e_init[648]), 
        .Q(nreg[648]) );
  DFF \nreg_reg[647]  ( .D(nreg[647]), .CLK(clk), .RST(rst), .I(e_init[647]), 
        .Q(nreg[647]) );
  DFF \nreg_reg[646]  ( .D(nreg[646]), .CLK(clk), .RST(rst), .I(e_init[646]), 
        .Q(nreg[646]) );
  DFF \nreg_reg[645]  ( .D(nreg[645]), .CLK(clk), .RST(rst), .I(e_init[645]), 
        .Q(nreg[645]) );
  DFF \nreg_reg[644]  ( .D(nreg[644]), .CLK(clk), .RST(rst), .I(e_init[644]), 
        .Q(nreg[644]) );
  DFF \nreg_reg[643]  ( .D(nreg[643]), .CLK(clk), .RST(rst), .I(e_init[643]), 
        .Q(nreg[643]) );
  DFF \nreg_reg[642]  ( .D(nreg[642]), .CLK(clk), .RST(rst), .I(e_init[642]), 
        .Q(nreg[642]) );
  DFF \nreg_reg[641]  ( .D(nreg[641]), .CLK(clk), .RST(rst), .I(e_init[641]), 
        .Q(nreg[641]) );
  DFF \nreg_reg[640]  ( .D(nreg[640]), .CLK(clk), .RST(rst), .I(e_init[640]), 
        .Q(nreg[640]) );
  DFF \nreg_reg[639]  ( .D(nreg[639]), .CLK(clk), .RST(rst), .I(e_init[639]), 
        .Q(nreg[639]) );
  DFF \nreg_reg[638]  ( .D(nreg[638]), .CLK(clk), .RST(rst), .I(e_init[638]), 
        .Q(nreg[638]) );
  DFF \nreg_reg[637]  ( .D(nreg[637]), .CLK(clk), .RST(rst), .I(e_init[637]), 
        .Q(nreg[637]) );
  DFF \nreg_reg[636]  ( .D(nreg[636]), .CLK(clk), .RST(rst), .I(e_init[636]), 
        .Q(nreg[636]) );
  DFF \nreg_reg[635]  ( .D(nreg[635]), .CLK(clk), .RST(rst), .I(e_init[635]), 
        .Q(nreg[635]) );
  DFF \nreg_reg[634]  ( .D(nreg[634]), .CLK(clk), .RST(rst), .I(e_init[634]), 
        .Q(nreg[634]) );
  DFF \nreg_reg[633]  ( .D(nreg[633]), .CLK(clk), .RST(rst), .I(e_init[633]), 
        .Q(nreg[633]) );
  DFF \nreg_reg[632]  ( .D(nreg[632]), .CLK(clk), .RST(rst), .I(e_init[632]), 
        .Q(nreg[632]) );
  DFF \nreg_reg[631]  ( .D(nreg[631]), .CLK(clk), .RST(rst), .I(e_init[631]), 
        .Q(nreg[631]) );
  DFF \nreg_reg[630]  ( .D(nreg[630]), .CLK(clk), .RST(rst), .I(e_init[630]), 
        .Q(nreg[630]) );
  DFF \nreg_reg[629]  ( .D(nreg[629]), .CLK(clk), .RST(rst), .I(e_init[629]), 
        .Q(nreg[629]) );
  DFF \nreg_reg[628]  ( .D(nreg[628]), .CLK(clk), .RST(rst), .I(e_init[628]), 
        .Q(nreg[628]) );
  DFF \nreg_reg[627]  ( .D(nreg[627]), .CLK(clk), .RST(rst), .I(e_init[627]), 
        .Q(nreg[627]) );
  DFF \nreg_reg[626]  ( .D(nreg[626]), .CLK(clk), .RST(rst), .I(e_init[626]), 
        .Q(nreg[626]) );
  DFF \nreg_reg[625]  ( .D(nreg[625]), .CLK(clk), .RST(rst), .I(e_init[625]), 
        .Q(nreg[625]) );
  DFF \nreg_reg[624]  ( .D(nreg[624]), .CLK(clk), .RST(rst), .I(e_init[624]), 
        .Q(nreg[624]) );
  DFF \nreg_reg[623]  ( .D(nreg[623]), .CLK(clk), .RST(rst), .I(e_init[623]), 
        .Q(nreg[623]) );
  DFF \nreg_reg[622]  ( .D(nreg[622]), .CLK(clk), .RST(rst), .I(e_init[622]), 
        .Q(nreg[622]) );
  DFF \nreg_reg[621]  ( .D(nreg[621]), .CLK(clk), .RST(rst), .I(e_init[621]), 
        .Q(nreg[621]) );
  DFF \nreg_reg[620]  ( .D(nreg[620]), .CLK(clk), .RST(rst), .I(e_init[620]), 
        .Q(nreg[620]) );
  DFF \nreg_reg[619]  ( .D(nreg[619]), .CLK(clk), .RST(rst), .I(e_init[619]), 
        .Q(nreg[619]) );
  DFF \nreg_reg[618]  ( .D(nreg[618]), .CLK(clk), .RST(rst), .I(e_init[618]), 
        .Q(nreg[618]) );
  DFF \nreg_reg[617]  ( .D(nreg[617]), .CLK(clk), .RST(rst), .I(e_init[617]), 
        .Q(nreg[617]) );
  DFF \nreg_reg[616]  ( .D(nreg[616]), .CLK(clk), .RST(rst), .I(e_init[616]), 
        .Q(nreg[616]) );
  DFF \nreg_reg[615]  ( .D(nreg[615]), .CLK(clk), .RST(rst), .I(e_init[615]), 
        .Q(nreg[615]) );
  DFF \nreg_reg[614]  ( .D(nreg[614]), .CLK(clk), .RST(rst), .I(e_init[614]), 
        .Q(nreg[614]) );
  DFF \nreg_reg[613]  ( .D(nreg[613]), .CLK(clk), .RST(rst), .I(e_init[613]), 
        .Q(nreg[613]) );
  DFF \nreg_reg[612]  ( .D(nreg[612]), .CLK(clk), .RST(rst), .I(e_init[612]), 
        .Q(nreg[612]) );
  DFF \nreg_reg[611]  ( .D(nreg[611]), .CLK(clk), .RST(rst), .I(e_init[611]), 
        .Q(nreg[611]) );
  DFF \nreg_reg[610]  ( .D(nreg[610]), .CLK(clk), .RST(rst), .I(e_init[610]), 
        .Q(nreg[610]) );
  DFF \nreg_reg[609]  ( .D(nreg[609]), .CLK(clk), .RST(rst), .I(e_init[609]), 
        .Q(nreg[609]) );
  DFF \nreg_reg[608]  ( .D(nreg[608]), .CLK(clk), .RST(rst), .I(e_init[608]), 
        .Q(nreg[608]) );
  DFF \nreg_reg[607]  ( .D(nreg[607]), .CLK(clk), .RST(rst), .I(e_init[607]), 
        .Q(nreg[607]) );
  DFF \nreg_reg[606]  ( .D(nreg[606]), .CLK(clk), .RST(rst), .I(e_init[606]), 
        .Q(nreg[606]) );
  DFF \nreg_reg[605]  ( .D(nreg[605]), .CLK(clk), .RST(rst), .I(e_init[605]), 
        .Q(nreg[605]) );
  DFF \nreg_reg[604]  ( .D(nreg[604]), .CLK(clk), .RST(rst), .I(e_init[604]), 
        .Q(nreg[604]) );
  DFF \nreg_reg[603]  ( .D(nreg[603]), .CLK(clk), .RST(rst), .I(e_init[603]), 
        .Q(nreg[603]) );
  DFF \nreg_reg[602]  ( .D(nreg[602]), .CLK(clk), .RST(rst), .I(e_init[602]), 
        .Q(nreg[602]) );
  DFF \nreg_reg[601]  ( .D(nreg[601]), .CLK(clk), .RST(rst), .I(e_init[601]), 
        .Q(nreg[601]) );
  DFF \nreg_reg[600]  ( .D(nreg[600]), .CLK(clk), .RST(rst), .I(e_init[600]), 
        .Q(nreg[600]) );
  DFF \nreg_reg[599]  ( .D(nreg[599]), .CLK(clk), .RST(rst), .I(e_init[599]), 
        .Q(nreg[599]) );
  DFF \nreg_reg[598]  ( .D(nreg[598]), .CLK(clk), .RST(rst), .I(e_init[598]), 
        .Q(nreg[598]) );
  DFF \nreg_reg[597]  ( .D(nreg[597]), .CLK(clk), .RST(rst), .I(e_init[597]), 
        .Q(nreg[597]) );
  DFF \nreg_reg[596]  ( .D(nreg[596]), .CLK(clk), .RST(rst), .I(e_init[596]), 
        .Q(nreg[596]) );
  DFF \nreg_reg[595]  ( .D(nreg[595]), .CLK(clk), .RST(rst), .I(e_init[595]), 
        .Q(nreg[595]) );
  DFF \nreg_reg[594]  ( .D(nreg[594]), .CLK(clk), .RST(rst), .I(e_init[594]), 
        .Q(nreg[594]) );
  DFF \nreg_reg[593]  ( .D(nreg[593]), .CLK(clk), .RST(rst), .I(e_init[593]), 
        .Q(nreg[593]) );
  DFF \nreg_reg[592]  ( .D(nreg[592]), .CLK(clk), .RST(rst), .I(e_init[592]), 
        .Q(nreg[592]) );
  DFF \nreg_reg[591]  ( .D(nreg[591]), .CLK(clk), .RST(rst), .I(e_init[591]), 
        .Q(nreg[591]) );
  DFF \nreg_reg[590]  ( .D(nreg[590]), .CLK(clk), .RST(rst), .I(e_init[590]), 
        .Q(nreg[590]) );
  DFF \nreg_reg[589]  ( .D(nreg[589]), .CLK(clk), .RST(rst), .I(e_init[589]), 
        .Q(nreg[589]) );
  DFF \nreg_reg[588]  ( .D(nreg[588]), .CLK(clk), .RST(rst), .I(e_init[588]), 
        .Q(nreg[588]) );
  DFF \nreg_reg[587]  ( .D(nreg[587]), .CLK(clk), .RST(rst), .I(e_init[587]), 
        .Q(nreg[587]) );
  DFF \nreg_reg[586]  ( .D(nreg[586]), .CLK(clk), .RST(rst), .I(e_init[586]), 
        .Q(nreg[586]) );
  DFF \nreg_reg[585]  ( .D(nreg[585]), .CLK(clk), .RST(rst), .I(e_init[585]), 
        .Q(nreg[585]) );
  DFF \nreg_reg[584]  ( .D(nreg[584]), .CLK(clk), .RST(rst), .I(e_init[584]), 
        .Q(nreg[584]) );
  DFF \nreg_reg[583]  ( .D(nreg[583]), .CLK(clk), .RST(rst), .I(e_init[583]), 
        .Q(nreg[583]) );
  DFF \nreg_reg[582]  ( .D(nreg[582]), .CLK(clk), .RST(rst), .I(e_init[582]), 
        .Q(nreg[582]) );
  DFF \nreg_reg[581]  ( .D(nreg[581]), .CLK(clk), .RST(rst), .I(e_init[581]), 
        .Q(nreg[581]) );
  DFF \nreg_reg[580]  ( .D(nreg[580]), .CLK(clk), .RST(rst), .I(e_init[580]), 
        .Q(nreg[580]) );
  DFF \nreg_reg[579]  ( .D(nreg[579]), .CLK(clk), .RST(rst), .I(e_init[579]), 
        .Q(nreg[579]) );
  DFF \nreg_reg[578]  ( .D(nreg[578]), .CLK(clk), .RST(rst), .I(e_init[578]), 
        .Q(nreg[578]) );
  DFF \nreg_reg[577]  ( .D(nreg[577]), .CLK(clk), .RST(rst), .I(e_init[577]), 
        .Q(nreg[577]) );
  DFF \nreg_reg[576]  ( .D(nreg[576]), .CLK(clk), .RST(rst), .I(e_init[576]), 
        .Q(nreg[576]) );
  DFF \nreg_reg[575]  ( .D(nreg[575]), .CLK(clk), .RST(rst), .I(e_init[575]), 
        .Q(nreg[575]) );
  DFF \nreg_reg[574]  ( .D(nreg[574]), .CLK(clk), .RST(rst), .I(e_init[574]), 
        .Q(nreg[574]) );
  DFF \nreg_reg[573]  ( .D(nreg[573]), .CLK(clk), .RST(rst), .I(e_init[573]), 
        .Q(nreg[573]) );
  DFF \nreg_reg[572]  ( .D(nreg[572]), .CLK(clk), .RST(rst), .I(e_init[572]), 
        .Q(nreg[572]) );
  DFF \nreg_reg[571]  ( .D(nreg[571]), .CLK(clk), .RST(rst), .I(e_init[571]), 
        .Q(nreg[571]) );
  DFF \nreg_reg[570]  ( .D(nreg[570]), .CLK(clk), .RST(rst), .I(e_init[570]), 
        .Q(nreg[570]) );
  DFF \nreg_reg[569]  ( .D(nreg[569]), .CLK(clk), .RST(rst), .I(e_init[569]), 
        .Q(nreg[569]) );
  DFF \nreg_reg[568]  ( .D(nreg[568]), .CLK(clk), .RST(rst), .I(e_init[568]), 
        .Q(nreg[568]) );
  DFF \nreg_reg[567]  ( .D(nreg[567]), .CLK(clk), .RST(rst), .I(e_init[567]), 
        .Q(nreg[567]) );
  DFF \nreg_reg[566]  ( .D(nreg[566]), .CLK(clk), .RST(rst), .I(e_init[566]), 
        .Q(nreg[566]) );
  DFF \nreg_reg[565]  ( .D(nreg[565]), .CLK(clk), .RST(rst), .I(e_init[565]), 
        .Q(nreg[565]) );
  DFF \nreg_reg[564]  ( .D(nreg[564]), .CLK(clk), .RST(rst), .I(e_init[564]), 
        .Q(nreg[564]) );
  DFF \nreg_reg[563]  ( .D(nreg[563]), .CLK(clk), .RST(rst), .I(e_init[563]), 
        .Q(nreg[563]) );
  DFF \nreg_reg[562]  ( .D(nreg[562]), .CLK(clk), .RST(rst), .I(e_init[562]), 
        .Q(nreg[562]) );
  DFF \nreg_reg[561]  ( .D(nreg[561]), .CLK(clk), .RST(rst), .I(e_init[561]), 
        .Q(nreg[561]) );
  DFF \nreg_reg[560]  ( .D(nreg[560]), .CLK(clk), .RST(rst), .I(e_init[560]), 
        .Q(nreg[560]) );
  DFF \nreg_reg[559]  ( .D(nreg[559]), .CLK(clk), .RST(rst), .I(e_init[559]), 
        .Q(nreg[559]) );
  DFF \nreg_reg[558]  ( .D(nreg[558]), .CLK(clk), .RST(rst), .I(e_init[558]), 
        .Q(nreg[558]) );
  DFF \nreg_reg[557]  ( .D(nreg[557]), .CLK(clk), .RST(rst), .I(e_init[557]), 
        .Q(nreg[557]) );
  DFF \nreg_reg[556]  ( .D(nreg[556]), .CLK(clk), .RST(rst), .I(e_init[556]), 
        .Q(nreg[556]) );
  DFF \nreg_reg[555]  ( .D(nreg[555]), .CLK(clk), .RST(rst), .I(e_init[555]), 
        .Q(nreg[555]) );
  DFF \nreg_reg[554]  ( .D(nreg[554]), .CLK(clk), .RST(rst), .I(e_init[554]), 
        .Q(nreg[554]) );
  DFF \nreg_reg[553]  ( .D(nreg[553]), .CLK(clk), .RST(rst), .I(e_init[553]), 
        .Q(nreg[553]) );
  DFF \nreg_reg[552]  ( .D(nreg[552]), .CLK(clk), .RST(rst), .I(e_init[552]), 
        .Q(nreg[552]) );
  DFF \nreg_reg[551]  ( .D(nreg[551]), .CLK(clk), .RST(rst), .I(e_init[551]), 
        .Q(nreg[551]) );
  DFF \nreg_reg[550]  ( .D(nreg[550]), .CLK(clk), .RST(rst), .I(e_init[550]), 
        .Q(nreg[550]) );
  DFF \nreg_reg[549]  ( .D(nreg[549]), .CLK(clk), .RST(rst), .I(e_init[549]), 
        .Q(nreg[549]) );
  DFF \nreg_reg[548]  ( .D(nreg[548]), .CLK(clk), .RST(rst), .I(e_init[548]), 
        .Q(nreg[548]) );
  DFF \nreg_reg[547]  ( .D(nreg[547]), .CLK(clk), .RST(rst), .I(e_init[547]), 
        .Q(nreg[547]) );
  DFF \nreg_reg[546]  ( .D(nreg[546]), .CLK(clk), .RST(rst), .I(e_init[546]), 
        .Q(nreg[546]) );
  DFF \nreg_reg[545]  ( .D(nreg[545]), .CLK(clk), .RST(rst), .I(e_init[545]), 
        .Q(nreg[545]) );
  DFF \nreg_reg[544]  ( .D(nreg[544]), .CLK(clk), .RST(rst), .I(e_init[544]), 
        .Q(nreg[544]) );
  DFF \nreg_reg[543]  ( .D(nreg[543]), .CLK(clk), .RST(rst), .I(e_init[543]), 
        .Q(nreg[543]) );
  DFF \nreg_reg[542]  ( .D(nreg[542]), .CLK(clk), .RST(rst), .I(e_init[542]), 
        .Q(nreg[542]) );
  DFF \nreg_reg[541]  ( .D(nreg[541]), .CLK(clk), .RST(rst), .I(e_init[541]), 
        .Q(nreg[541]) );
  DFF \nreg_reg[540]  ( .D(nreg[540]), .CLK(clk), .RST(rst), .I(e_init[540]), 
        .Q(nreg[540]) );
  DFF \nreg_reg[539]  ( .D(nreg[539]), .CLK(clk), .RST(rst), .I(e_init[539]), 
        .Q(nreg[539]) );
  DFF \nreg_reg[538]  ( .D(nreg[538]), .CLK(clk), .RST(rst), .I(e_init[538]), 
        .Q(nreg[538]) );
  DFF \nreg_reg[537]  ( .D(nreg[537]), .CLK(clk), .RST(rst), .I(e_init[537]), 
        .Q(nreg[537]) );
  DFF \nreg_reg[536]  ( .D(nreg[536]), .CLK(clk), .RST(rst), .I(e_init[536]), 
        .Q(nreg[536]) );
  DFF \nreg_reg[535]  ( .D(nreg[535]), .CLK(clk), .RST(rst), .I(e_init[535]), 
        .Q(nreg[535]) );
  DFF \nreg_reg[534]  ( .D(nreg[534]), .CLK(clk), .RST(rst), .I(e_init[534]), 
        .Q(nreg[534]) );
  DFF \nreg_reg[533]  ( .D(nreg[533]), .CLK(clk), .RST(rst), .I(e_init[533]), 
        .Q(nreg[533]) );
  DFF \nreg_reg[532]  ( .D(nreg[532]), .CLK(clk), .RST(rst), .I(e_init[532]), 
        .Q(nreg[532]) );
  DFF \nreg_reg[531]  ( .D(nreg[531]), .CLK(clk), .RST(rst), .I(e_init[531]), 
        .Q(nreg[531]) );
  DFF \nreg_reg[530]  ( .D(nreg[530]), .CLK(clk), .RST(rst), .I(e_init[530]), 
        .Q(nreg[530]) );
  DFF \nreg_reg[529]  ( .D(nreg[529]), .CLK(clk), .RST(rst), .I(e_init[529]), 
        .Q(nreg[529]) );
  DFF \nreg_reg[528]  ( .D(nreg[528]), .CLK(clk), .RST(rst), .I(e_init[528]), 
        .Q(nreg[528]) );
  DFF \nreg_reg[527]  ( .D(nreg[527]), .CLK(clk), .RST(rst), .I(e_init[527]), 
        .Q(nreg[527]) );
  DFF \nreg_reg[526]  ( .D(nreg[526]), .CLK(clk), .RST(rst), .I(e_init[526]), 
        .Q(nreg[526]) );
  DFF \nreg_reg[525]  ( .D(nreg[525]), .CLK(clk), .RST(rst), .I(e_init[525]), 
        .Q(nreg[525]) );
  DFF \nreg_reg[524]  ( .D(nreg[524]), .CLK(clk), .RST(rst), .I(e_init[524]), 
        .Q(nreg[524]) );
  DFF \nreg_reg[523]  ( .D(nreg[523]), .CLK(clk), .RST(rst), .I(e_init[523]), 
        .Q(nreg[523]) );
  DFF \nreg_reg[522]  ( .D(nreg[522]), .CLK(clk), .RST(rst), .I(e_init[522]), 
        .Q(nreg[522]) );
  DFF \nreg_reg[521]  ( .D(nreg[521]), .CLK(clk), .RST(rst), .I(e_init[521]), 
        .Q(nreg[521]) );
  DFF \nreg_reg[520]  ( .D(nreg[520]), .CLK(clk), .RST(rst), .I(e_init[520]), 
        .Q(nreg[520]) );
  DFF \nreg_reg[519]  ( .D(nreg[519]), .CLK(clk), .RST(rst), .I(e_init[519]), 
        .Q(nreg[519]) );
  DFF \nreg_reg[518]  ( .D(nreg[518]), .CLK(clk), .RST(rst), .I(e_init[518]), 
        .Q(nreg[518]) );
  DFF \nreg_reg[517]  ( .D(nreg[517]), .CLK(clk), .RST(rst), .I(e_init[517]), 
        .Q(nreg[517]) );
  DFF \nreg_reg[516]  ( .D(nreg[516]), .CLK(clk), .RST(rst), .I(e_init[516]), 
        .Q(nreg[516]) );
  DFF \nreg_reg[515]  ( .D(nreg[515]), .CLK(clk), .RST(rst), .I(e_init[515]), 
        .Q(nreg[515]) );
  DFF \nreg_reg[514]  ( .D(nreg[514]), .CLK(clk), .RST(rst), .I(e_init[514]), 
        .Q(nreg[514]) );
  DFF \nreg_reg[513]  ( .D(nreg[513]), .CLK(clk), .RST(rst), .I(e_init[513]), 
        .Q(nreg[513]) );
  DFF \nreg_reg[512]  ( .D(nreg[512]), .CLK(clk), .RST(rst), .I(e_init[512]), 
        .Q(nreg[512]) );
  DFF \nreg_reg[511]  ( .D(nreg[511]), .CLK(clk), .RST(rst), .I(e_init[511]), 
        .Q(nreg[511]) );
  DFF \nreg_reg[510]  ( .D(nreg[510]), .CLK(clk), .RST(rst), .I(e_init[510]), 
        .Q(nreg[510]) );
  DFF \nreg_reg[509]  ( .D(nreg[509]), .CLK(clk), .RST(rst), .I(e_init[509]), 
        .Q(nreg[509]) );
  DFF \nreg_reg[508]  ( .D(nreg[508]), .CLK(clk), .RST(rst), .I(e_init[508]), 
        .Q(nreg[508]) );
  DFF \nreg_reg[507]  ( .D(nreg[507]), .CLK(clk), .RST(rst), .I(e_init[507]), 
        .Q(nreg[507]) );
  DFF \nreg_reg[506]  ( .D(nreg[506]), .CLK(clk), .RST(rst), .I(e_init[506]), 
        .Q(nreg[506]) );
  DFF \nreg_reg[505]  ( .D(nreg[505]), .CLK(clk), .RST(rst), .I(e_init[505]), 
        .Q(nreg[505]) );
  DFF \nreg_reg[504]  ( .D(nreg[504]), .CLK(clk), .RST(rst), .I(e_init[504]), 
        .Q(nreg[504]) );
  DFF \nreg_reg[503]  ( .D(nreg[503]), .CLK(clk), .RST(rst), .I(e_init[503]), 
        .Q(nreg[503]) );
  DFF \nreg_reg[502]  ( .D(nreg[502]), .CLK(clk), .RST(rst), .I(e_init[502]), 
        .Q(nreg[502]) );
  DFF \nreg_reg[501]  ( .D(nreg[501]), .CLK(clk), .RST(rst), .I(e_init[501]), 
        .Q(nreg[501]) );
  DFF \nreg_reg[500]  ( .D(nreg[500]), .CLK(clk), .RST(rst), .I(e_init[500]), 
        .Q(nreg[500]) );
  DFF \nreg_reg[499]  ( .D(nreg[499]), .CLK(clk), .RST(rst), .I(e_init[499]), 
        .Q(nreg[499]) );
  DFF \nreg_reg[498]  ( .D(nreg[498]), .CLK(clk), .RST(rst), .I(e_init[498]), 
        .Q(nreg[498]) );
  DFF \nreg_reg[497]  ( .D(nreg[497]), .CLK(clk), .RST(rst), .I(e_init[497]), 
        .Q(nreg[497]) );
  DFF \nreg_reg[496]  ( .D(nreg[496]), .CLK(clk), .RST(rst), .I(e_init[496]), 
        .Q(nreg[496]) );
  DFF \nreg_reg[495]  ( .D(nreg[495]), .CLK(clk), .RST(rst), .I(e_init[495]), 
        .Q(nreg[495]) );
  DFF \nreg_reg[494]  ( .D(nreg[494]), .CLK(clk), .RST(rst), .I(e_init[494]), 
        .Q(nreg[494]) );
  DFF \nreg_reg[493]  ( .D(nreg[493]), .CLK(clk), .RST(rst), .I(e_init[493]), 
        .Q(nreg[493]) );
  DFF \nreg_reg[492]  ( .D(nreg[492]), .CLK(clk), .RST(rst), .I(e_init[492]), 
        .Q(nreg[492]) );
  DFF \nreg_reg[491]  ( .D(nreg[491]), .CLK(clk), .RST(rst), .I(e_init[491]), 
        .Q(nreg[491]) );
  DFF \nreg_reg[490]  ( .D(nreg[490]), .CLK(clk), .RST(rst), .I(e_init[490]), 
        .Q(nreg[490]) );
  DFF \nreg_reg[489]  ( .D(nreg[489]), .CLK(clk), .RST(rst), .I(e_init[489]), 
        .Q(nreg[489]) );
  DFF \nreg_reg[488]  ( .D(nreg[488]), .CLK(clk), .RST(rst), .I(e_init[488]), 
        .Q(nreg[488]) );
  DFF \nreg_reg[487]  ( .D(nreg[487]), .CLK(clk), .RST(rst), .I(e_init[487]), 
        .Q(nreg[487]) );
  DFF \nreg_reg[486]  ( .D(nreg[486]), .CLK(clk), .RST(rst), .I(e_init[486]), 
        .Q(nreg[486]) );
  DFF \nreg_reg[485]  ( .D(nreg[485]), .CLK(clk), .RST(rst), .I(e_init[485]), 
        .Q(nreg[485]) );
  DFF \nreg_reg[484]  ( .D(nreg[484]), .CLK(clk), .RST(rst), .I(e_init[484]), 
        .Q(nreg[484]) );
  DFF \nreg_reg[483]  ( .D(nreg[483]), .CLK(clk), .RST(rst), .I(e_init[483]), 
        .Q(nreg[483]) );
  DFF \nreg_reg[482]  ( .D(nreg[482]), .CLK(clk), .RST(rst), .I(e_init[482]), 
        .Q(nreg[482]) );
  DFF \nreg_reg[481]  ( .D(nreg[481]), .CLK(clk), .RST(rst), .I(e_init[481]), 
        .Q(nreg[481]) );
  DFF \nreg_reg[480]  ( .D(nreg[480]), .CLK(clk), .RST(rst), .I(e_init[480]), 
        .Q(nreg[480]) );
  DFF \nreg_reg[479]  ( .D(nreg[479]), .CLK(clk), .RST(rst), .I(e_init[479]), 
        .Q(nreg[479]) );
  DFF \nreg_reg[478]  ( .D(nreg[478]), .CLK(clk), .RST(rst), .I(e_init[478]), 
        .Q(nreg[478]) );
  DFF \nreg_reg[477]  ( .D(nreg[477]), .CLK(clk), .RST(rst), .I(e_init[477]), 
        .Q(nreg[477]) );
  DFF \nreg_reg[476]  ( .D(nreg[476]), .CLK(clk), .RST(rst), .I(e_init[476]), 
        .Q(nreg[476]) );
  DFF \nreg_reg[475]  ( .D(nreg[475]), .CLK(clk), .RST(rst), .I(e_init[475]), 
        .Q(nreg[475]) );
  DFF \nreg_reg[474]  ( .D(nreg[474]), .CLK(clk), .RST(rst), .I(e_init[474]), 
        .Q(nreg[474]) );
  DFF \nreg_reg[473]  ( .D(nreg[473]), .CLK(clk), .RST(rst), .I(e_init[473]), 
        .Q(nreg[473]) );
  DFF \nreg_reg[472]  ( .D(nreg[472]), .CLK(clk), .RST(rst), .I(e_init[472]), 
        .Q(nreg[472]) );
  DFF \nreg_reg[471]  ( .D(nreg[471]), .CLK(clk), .RST(rst), .I(e_init[471]), 
        .Q(nreg[471]) );
  DFF \nreg_reg[470]  ( .D(nreg[470]), .CLK(clk), .RST(rst), .I(e_init[470]), 
        .Q(nreg[470]) );
  DFF \nreg_reg[469]  ( .D(nreg[469]), .CLK(clk), .RST(rst), .I(e_init[469]), 
        .Q(nreg[469]) );
  DFF \nreg_reg[468]  ( .D(nreg[468]), .CLK(clk), .RST(rst), .I(e_init[468]), 
        .Q(nreg[468]) );
  DFF \nreg_reg[467]  ( .D(nreg[467]), .CLK(clk), .RST(rst), .I(e_init[467]), 
        .Q(nreg[467]) );
  DFF \nreg_reg[466]  ( .D(nreg[466]), .CLK(clk), .RST(rst), .I(e_init[466]), 
        .Q(nreg[466]) );
  DFF \nreg_reg[465]  ( .D(nreg[465]), .CLK(clk), .RST(rst), .I(e_init[465]), 
        .Q(nreg[465]) );
  DFF \nreg_reg[464]  ( .D(nreg[464]), .CLK(clk), .RST(rst), .I(e_init[464]), 
        .Q(nreg[464]) );
  DFF \nreg_reg[463]  ( .D(nreg[463]), .CLK(clk), .RST(rst), .I(e_init[463]), 
        .Q(nreg[463]) );
  DFF \nreg_reg[462]  ( .D(nreg[462]), .CLK(clk), .RST(rst), .I(e_init[462]), 
        .Q(nreg[462]) );
  DFF \nreg_reg[461]  ( .D(nreg[461]), .CLK(clk), .RST(rst), .I(e_init[461]), 
        .Q(nreg[461]) );
  DFF \nreg_reg[460]  ( .D(nreg[460]), .CLK(clk), .RST(rst), .I(e_init[460]), 
        .Q(nreg[460]) );
  DFF \nreg_reg[459]  ( .D(nreg[459]), .CLK(clk), .RST(rst), .I(e_init[459]), 
        .Q(nreg[459]) );
  DFF \nreg_reg[458]  ( .D(nreg[458]), .CLK(clk), .RST(rst), .I(e_init[458]), 
        .Q(nreg[458]) );
  DFF \nreg_reg[457]  ( .D(nreg[457]), .CLK(clk), .RST(rst), .I(e_init[457]), 
        .Q(nreg[457]) );
  DFF \nreg_reg[456]  ( .D(nreg[456]), .CLK(clk), .RST(rst), .I(e_init[456]), 
        .Q(nreg[456]) );
  DFF \nreg_reg[455]  ( .D(nreg[455]), .CLK(clk), .RST(rst), .I(e_init[455]), 
        .Q(nreg[455]) );
  DFF \nreg_reg[454]  ( .D(nreg[454]), .CLK(clk), .RST(rst), .I(e_init[454]), 
        .Q(nreg[454]) );
  DFF \nreg_reg[453]  ( .D(nreg[453]), .CLK(clk), .RST(rst), .I(e_init[453]), 
        .Q(nreg[453]) );
  DFF \nreg_reg[452]  ( .D(nreg[452]), .CLK(clk), .RST(rst), .I(e_init[452]), 
        .Q(nreg[452]) );
  DFF \nreg_reg[451]  ( .D(nreg[451]), .CLK(clk), .RST(rst), .I(e_init[451]), 
        .Q(nreg[451]) );
  DFF \nreg_reg[450]  ( .D(nreg[450]), .CLK(clk), .RST(rst), .I(e_init[450]), 
        .Q(nreg[450]) );
  DFF \nreg_reg[449]  ( .D(nreg[449]), .CLK(clk), .RST(rst), .I(e_init[449]), 
        .Q(nreg[449]) );
  DFF \nreg_reg[448]  ( .D(nreg[448]), .CLK(clk), .RST(rst), .I(e_init[448]), 
        .Q(nreg[448]) );
  DFF \nreg_reg[447]  ( .D(nreg[447]), .CLK(clk), .RST(rst), .I(e_init[447]), 
        .Q(nreg[447]) );
  DFF \nreg_reg[446]  ( .D(nreg[446]), .CLK(clk), .RST(rst), .I(e_init[446]), 
        .Q(nreg[446]) );
  DFF \nreg_reg[445]  ( .D(nreg[445]), .CLK(clk), .RST(rst), .I(e_init[445]), 
        .Q(nreg[445]) );
  DFF \nreg_reg[444]  ( .D(nreg[444]), .CLK(clk), .RST(rst), .I(e_init[444]), 
        .Q(nreg[444]) );
  DFF \nreg_reg[443]  ( .D(nreg[443]), .CLK(clk), .RST(rst), .I(e_init[443]), 
        .Q(nreg[443]) );
  DFF \nreg_reg[442]  ( .D(nreg[442]), .CLK(clk), .RST(rst), .I(e_init[442]), 
        .Q(nreg[442]) );
  DFF \nreg_reg[441]  ( .D(nreg[441]), .CLK(clk), .RST(rst), .I(e_init[441]), 
        .Q(nreg[441]) );
  DFF \nreg_reg[440]  ( .D(nreg[440]), .CLK(clk), .RST(rst), .I(e_init[440]), 
        .Q(nreg[440]) );
  DFF \nreg_reg[439]  ( .D(nreg[439]), .CLK(clk), .RST(rst), .I(e_init[439]), 
        .Q(nreg[439]) );
  DFF \nreg_reg[438]  ( .D(nreg[438]), .CLK(clk), .RST(rst), .I(e_init[438]), 
        .Q(nreg[438]) );
  DFF \nreg_reg[437]  ( .D(nreg[437]), .CLK(clk), .RST(rst), .I(e_init[437]), 
        .Q(nreg[437]) );
  DFF \nreg_reg[436]  ( .D(nreg[436]), .CLK(clk), .RST(rst), .I(e_init[436]), 
        .Q(nreg[436]) );
  DFF \nreg_reg[435]  ( .D(nreg[435]), .CLK(clk), .RST(rst), .I(e_init[435]), 
        .Q(nreg[435]) );
  DFF \nreg_reg[434]  ( .D(nreg[434]), .CLK(clk), .RST(rst), .I(e_init[434]), 
        .Q(nreg[434]) );
  DFF \nreg_reg[433]  ( .D(nreg[433]), .CLK(clk), .RST(rst), .I(e_init[433]), 
        .Q(nreg[433]) );
  DFF \nreg_reg[432]  ( .D(nreg[432]), .CLK(clk), .RST(rst), .I(e_init[432]), 
        .Q(nreg[432]) );
  DFF \nreg_reg[431]  ( .D(nreg[431]), .CLK(clk), .RST(rst), .I(e_init[431]), 
        .Q(nreg[431]) );
  DFF \nreg_reg[430]  ( .D(nreg[430]), .CLK(clk), .RST(rst), .I(e_init[430]), 
        .Q(nreg[430]) );
  DFF \nreg_reg[429]  ( .D(nreg[429]), .CLK(clk), .RST(rst), .I(e_init[429]), 
        .Q(nreg[429]) );
  DFF \nreg_reg[428]  ( .D(nreg[428]), .CLK(clk), .RST(rst), .I(e_init[428]), 
        .Q(nreg[428]) );
  DFF \nreg_reg[427]  ( .D(nreg[427]), .CLK(clk), .RST(rst), .I(e_init[427]), 
        .Q(nreg[427]) );
  DFF \nreg_reg[426]  ( .D(nreg[426]), .CLK(clk), .RST(rst), .I(e_init[426]), 
        .Q(nreg[426]) );
  DFF \nreg_reg[425]  ( .D(nreg[425]), .CLK(clk), .RST(rst), .I(e_init[425]), 
        .Q(nreg[425]) );
  DFF \nreg_reg[424]  ( .D(nreg[424]), .CLK(clk), .RST(rst), .I(e_init[424]), 
        .Q(nreg[424]) );
  DFF \nreg_reg[423]  ( .D(nreg[423]), .CLK(clk), .RST(rst), .I(e_init[423]), 
        .Q(nreg[423]) );
  DFF \nreg_reg[422]  ( .D(nreg[422]), .CLK(clk), .RST(rst), .I(e_init[422]), 
        .Q(nreg[422]) );
  DFF \nreg_reg[421]  ( .D(nreg[421]), .CLK(clk), .RST(rst), .I(e_init[421]), 
        .Q(nreg[421]) );
  DFF \nreg_reg[420]  ( .D(nreg[420]), .CLK(clk), .RST(rst), .I(e_init[420]), 
        .Q(nreg[420]) );
  DFF \nreg_reg[419]  ( .D(nreg[419]), .CLK(clk), .RST(rst), .I(e_init[419]), 
        .Q(nreg[419]) );
  DFF \nreg_reg[418]  ( .D(nreg[418]), .CLK(clk), .RST(rst), .I(e_init[418]), 
        .Q(nreg[418]) );
  DFF \nreg_reg[417]  ( .D(nreg[417]), .CLK(clk), .RST(rst), .I(e_init[417]), 
        .Q(nreg[417]) );
  DFF \nreg_reg[416]  ( .D(nreg[416]), .CLK(clk), .RST(rst), .I(e_init[416]), 
        .Q(nreg[416]) );
  DFF \nreg_reg[415]  ( .D(nreg[415]), .CLK(clk), .RST(rst), .I(e_init[415]), 
        .Q(nreg[415]) );
  DFF \nreg_reg[414]  ( .D(nreg[414]), .CLK(clk), .RST(rst), .I(e_init[414]), 
        .Q(nreg[414]) );
  DFF \nreg_reg[413]  ( .D(nreg[413]), .CLK(clk), .RST(rst), .I(e_init[413]), 
        .Q(nreg[413]) );
  DFF \nreg_reg[412]  ( .D(nreg[412]), .CLK(clk), .RST(rst), .I(e_init[412]), 
        .Q(nreg[412]) );
  DFF \nreg_reg[411]  ( .D(nreg[411]), .CLK(clk), .RST(rst), .I(e_init[411]), 
        .Q(nreg[411]) );
  DFF \nreg_reg[410]  ( .D(nreg[410]), .CLK(clk), .RST(rst), .I(e_init[410]), 
        .Q(nreg[410]) );
  DFF \nreg_reg[409]  ( .D(nreg[409]), .CLK(clk), .RST(rst), .I(e_init[409]), 
        .Q(nreg[409]) );
  DFF \nreg_reg[408]  ( .D(nreg[408]), .CLK(clk), .RST(rst), .I(e_init[408]), 
        .Q(nreg[408]) );
  DFF \nreg_reg[407]  ( .D(nreg[407]), .CLK(clk), .RST(rst), .I(e_init[407]), 
        .Q(nreg[407]) );
  DFF \nreg_reg[406]  ( .D(nreg[406]), .CLK(clk), .RST(rst), .I(e_init[406]), 
        .Q(nreg[406]) );
  DFF \nreg_reg[405]  ( .D(nreg[405]), .CLK(clk), .RST(rst), .I(e_init[405]), 
        .Q(nreg[405]) );
  DFF \nreg_reg[404]  ( .D(nreg[404]), .CLK(clk), .RST(rst), .I(e_init[404]), 
        .Q(nreg[404]) );
  DFF \nreg_reg[403]  ( .D(nreg[403]), .CLK(clk), .RST(rst), .I(e_init[403]), 
        .Q(nreg[403]) );
  DFF \nreg_reg[402]  ( .D(nreg[402]), .CLK(clk), .RST(rst), .I(e_init[402]), 
        .Q(nreg[402]) );
  DFF \nreg_reg[401]  ( .D(nreg[401]), .CLK(clk), .RST(rst), .I(e_init[401]), 
        .Q(nreg[401]) );
  DFF \nreg_reg[400]  ( .D(nreg[400]), .CLK(clk), .RST(rst), .I(e_init[400]), 
        .Q(nreg[400]) );
  DFF \nreg_reg[399]  ( .D(nreg[399]), .CLK(clk), .RST(rst), .I(e_init[399]), 
        .Q(nreg[399]) );
  DFF \nreg_reg[398]  ( .D(nreg[398]), .CLK(clk), .RST(rst), .I(e_init[398]), 
        .Q(nreg[398]) );
  DFF \nreg_reg[397]  ( .D(nreg[397]), .CLK(clk), .RST(rst), .I(e_init[397]), 
        .Q(nreg[397]) );
  DFF \nreg_reg[396]  ( .D(nreg[396]), .CLK(clk), .RST(rst), .I(e_init[396]), 
        .Q(nreg[396]) );
  DFF \nreg_reg[395]  ( .D(nreg[395]), .CLK(clk), .RST(rst), .I(e_init[395]), 
        .Q(nreg[395]) );
  DFF \nreg_reg[394]  ( .D(nreg[394]), .CLK(clk), .RST(rst), .I(e_init[394]), 
        .Q(nreg[394]) );
  DFF \nreg_reg[393]  ( .D(nreg[393]), .CLK(clk), .RST(rst), .I(e_init[393]), 
        .Q(nreg[393]) );
  DFF \nreg_reg[392]  ( .D(nreg[392]), .CLK(clk), .RST(rst), .I(e_init[392]), 
        .Q(nreg[392]) );
  DFF \nreg_reg[391]  ( .D(nreg[391]), .CLK(clk), .RST(rst), .I(e_init[391]), 
        .Q(nreg[391]) );
  DFF \nreg_reg[390]  ( .D(nreg[390]), .CLK(clk), .RST(rst), .I(e_init[390]), 
        .Q(nreg[390]) );
  DFF \nreg_reg[389]  ( .D(nreg[389]), .CLK(clk), .RST(rst), .I(e_init[389]), 
        .Q(nreg[389]) );
  DFF \nreg_reg[388]  ( .D(nreg[388]), .CLK(clk), .RST(rst), .I(e_init[388]), 
        .Q(nreg[388]) );
  DFF \nreg_reg[387]  ( .D(nreg[387]), .CLK(clk), .RST(rst), .I(e_init[387]), 
        .Q(nreg[387]) );
  DFF \nreg_reg[386]  ( .D(nreg[386]), .CLK(clk), .RST(rst), .I(e_init[386]), 
        .Q(nreg[386]) );
  DFF \nreg_reg[385]  ( .D(nreg[385]), .CLK(clk), .RST(rst), .I(e_init[385]), 
        .Q(nreg[385]) );
  DFF \nreg_reg[384]  ( .D(nreg[384]), .CLK(clk), .RST(rst), .I(e_init[384]), 
        .Q(nreg[384]) );
  DFF \nreg_reg[383]  ( .D(nreg[383]), .CLK(clk), .RST(rst), .I(e_init[383]), 
        .Q(nreg[383]) );
  DFF \nreg_reg[382]  ( .D(nreg[382]), .CLK(clk), .RST(rst), .I(e_init[382]), 
        .Q(nreg[382]) );
  DFF \nreg_reg[381]  ( .D(nreg[381]), .CLK(clk), .RST(rst), .I(e_init[381]), 
        .Q(nreg[381]) );
  DFF \nreg_reg[380]  ( .D(nreg[380]), .CLK(clk), .RST(rst), .I(e_init[380]), 
        .Q(nreg[380]) );
  DFF \nreg_reg[379]  ( .D(nreg[379]), .CLK(clk), .RST(rst), .I(e_init[379]), 
        .Q(nreg[379]) );
  DFF \nreg_reg[378]  ( .D(nreg[378]), .CLK(clk), .RST(rst), .I(e_init[378]), 
        .Q(nreg[378]) );
  DFF \nreg_reg[377]  ( .D(nreg[377]), .CLK(clk), .RST(rst), .I(e_init[377]), 
        .Q(nreg[377]) );
  DFF \nreg_reg[376]  ( .D(nreg[376]), .CLK(clk), .RST(rst), .I(e_init[376]), 
        .Q(nreg[376]) );
  DFF \nreg_reg[375]  ( .D(nreg[375]), .CLK(clk), .RST(rst), .I(e_init[375]), 
        .Q(nreg[375]) );
  DFF \nreg_reg[374]  ( .D(nreg[374]), .CLK(clk), .RST(rst), .I(e_init[374]), 
        .Q(nreg[374]) );
  DFF \nreg_reg[373]  ( .D(nreg[373]), .CLK(clk), .RST(rst), .I(e_init[373]), 
        .Q(nreg[373]) );
  DFF \nreg_reg[372]  ( .D(nreg[372]), .CLK(clk), .RST(rst), .I(e_init[372]), 
        .Q(nreg[372]) );
  DFF \nreg_reg[371]  ( .D(nreg[371]), .CLK(clk), .RST(rst), .I(e_init[371]), 
        .Q(nreg[371]) );
  DFF \nreg_reg[370]  ( .D(nreg[370]), .CLK(clk), .RST(rst), .I(e_init[370]), 
        .Q(nreg[370]) );
  DFF \nreg_reg[369]  ( .D(nreg[369]), .CLK(clk), .RST(rst), .I(e_init[369]), 
        .Q(nreg[369]) );
  DFF \nreg_reg[368]  ( .D(nreg[368]), .CLK(clk), .RST(rst), .I(e_init[368]), 
        .Q(nreg[368]) );
  DFF \nreg_reg[367]  ( .D(nreg[367]), .CLK(clk), .RST(rst), .I(e_init[367]), 
        .Q(nreg[367]) );
  DFF \nreg_reg[366]  ( .D(nreg[366]), .CLK(clk), .RST(rst), .I(e_init[366]), 
        .Q(nreg[366]) );
  DFF \nreg_reg[365]  ( .D(nreg[365]), .CLK(clk), .RST(rst), .I(e_init[365]), 
        .Q(nreg[365]) );
  DFF \nreg_reg[364]  ( .D(nreg[364]), .CLK(clk), .RST(rst), .I(e_init[364]), 
        .Q(nreg[364]) );
  DFF \nreg_reg[363]  ( .D(nreg[363]), .CLK(clk), .RST(rst), .I(e_init[363]), 
        .Q(nreg[363]) );
  DFF \nreg_reg[362]  ( .D(nreg[362]), .CLK(clk), .RST(rst), .I(e_init[362]), 
        .Q(nreg[362]) );
  DFF \nreg_reg[361]  ( .D(nreg[361]), .CLK(clk), .RST(rst), .I(e_init[361]), 
        .Q(nreg[361]) );
  DFF \nreg_reg[360]  ( .D(nreg[360]), .CLK(clk), .RST(rst), .I(e_init[360]), 
        .Q(nreg[360]) );
  DFF \nreg_reg[359]  ( .D(nreg[359]), .CLK(clk), .RST(rst), .I(e_init[359]), 
        .Q(nreg[359]) );
  DFF \nreg_reg[358]  ( .D(nreg[358]), .CLK(clk), .RST(rst), .I(e_init[358]), 
        .Q(nreg[358]) );
  DFF \nreg_reg[357]  ( .D(nreg[357]), .CLK(clk), .RST(rst), .I(e_init[357]), 
        .Q(nreg[357]) );
  DFF \nreg_reg[356]  ( .D(nreg[356]), .CLK(clk), .RST(rst), .I(e_init[356]), 
        .Q(nreg[356]) );
  DFF \nreg_reg[355]  ( .D(nreg[355]), .CLK(clk), .RST(rst), .I(e_init[355]), 
        .Q(nreg[355]) );
  DFF \nreg_reg[354]  ( .D(nreg[354]), .CLK(clk), .RST(rst), .I(e_init[354]), 
        .Q(nreg[354]) );
  DFF \nreg_reg[353]  ( .D(nreg[353]), .CLK(clk), .RST(rst), .I(e_init[353]), 
        .Q(nreg[353]) );
  DFF \nreg_reg[352]  ( .D(nreg[352]), .CLK(clk), .RST(rst), .I(e_init[352]), 
        .Q(nreg[352]) );
  DFF \nreg_reg[351]  ( .D(nreg[351]), .CLK(clk), .RST(rst), .I(e_init[351]), 
        .Q(nreg[351]) );
  DFF \nreg_reg[350]  ( .D(nreg[350]), .CLK(clk), .RST(rst), .I(e_init[350]), 
        .Q(nreg[350]) );
  DFF \nreg_reg[349]  ( .D(nreg[349]), .CLK(clk), .RST(rst), .I(e_init[349]), 
        .Q(nreg[349]) );
  DFF \nreg_reg[348]  ( .D(nreg[348]), .CLK(clk), .RST(rst), .I(e_init[348]), 
        .Q(nreg[348]) );
  DFF \nreg_reg[347]  ( .D(nreg[347]), .CLK(clk), .RST(rst), .I(e_init[347]), 
        .Q(nreg[347]) );
  DFF \nreg_reg[346]  ( .D(nreg[346]), .CLK(clk), .RST(rst), .I(e_init[346]), 
        .Q(nreg[346]) );
  DFF \nreg_reg[345]  ( .D(nreg[345]), .CLK(clk), .RST(rst), .I(e_init[345]), 
        .Q(nreg[345]) );
  DFF \nreg_reg[344]  ( .D(nreg[344]), .CLK(clk), .RST(rst), .I(e_init[344]), 
        .Q(nreg[344]) );
  DFF \nreg_reg[343]  ( .D(nreg[343]), .CLK(clk), .RST(rst), .I(e_init[343]), 
        .Q(nreg[343]) );
  DFF \nreg_reg[342]  ( .D(nreg[342]), .CLK(clk), .RST(rst), .I(e_init[342]), 
        .Q(nreg[342]) );
  DFF \nreg_reg[341]  ( .D(nreg[341]), .CLK(clk), .RST(rst), .I(e_init[341]), 
        .Q(nreg[341]) );
  DFF \nreg_reg[340]  ( .D(nreg[340]), .CLK(clk), .RST(rst), .I(e_init[340]), 
        .Q(nreg[340]) );
  DFF \nreg_reg[339]  ( .D(nreg[339]), .CLK(clk), .RST(rst), .I(e_init[339]), 
        .Q(nreg[339]) );
  DFF \nreg_reg[338]  ( .D(nreg[338]), .CLK(clk), .RST(rst), .I(e_init[338]), 
        .Q(nreg[338]) );
  DFF \nreg_reg[337]  ( .D(nreg[337]), .CLK(clk), .RST(rst), .I(e_init[337]), 
        .Q(nreg[337]) );
  DFF \nreg_reg[336]  ( .D(nreg[336]), .CLK(clk), .RST(rst), .I(e_init[336]), 
        .Q(nreg[336]) );
  DFF \nreg_reg[335]  ( .D(nreg[335]), .CLK(clk), .RST(rst), .I(e_init[335]), 
        .Q(nreg[335]) );
  DFF \nreg_reg[334]  ( .D(nreg[334]), .CLK(clk), .RST(rst), .I(e_init[334]), 
        .Q(nreg[334]) );
  DFF \nreg_reg[333]  ( .D(nreg[333]), .CLK(clk), .RST(rst), .I(e_init[333]), 
        .Q(nreg[333]) );
  DFF \nreg_reg[332]  ( .D(nreg[332]), .CLK(clk), .RST(rst), .I(e_init[332]), 
        .Q(nreg[332]) );
  DFF \nreg_reg[331]  ( .D(nreg[331]), .CLK(clk), .RST(rst), .I(e_init[331]), 
        .Q(nreg[331]) );
  DFF \nreg_reg[330]  ( .D(nreg[330]), .CLK(clk), .RST(rst), .I(e_init[330]), 
        .Q(nreg[330]) );
  DFF \nreg_reg[329]  ( .D(nreg[329]), .CLK(clk), .RST(rst), .I(e_init[329]), 
        .Q(nreg[329]) );
  DFF \nreg_reg[328]  ( .D(nreg[328]), .CLK(clk), .RST(rst), .I(e_init[328]), 
        .Q(nreg[328]) );
  DFF \nreg_reg[327]  ( .D(nreg[327]), .CLK(clk), .RST(rst), .I(e_init[327]), 
        .Q(nreg[327]) );
  DFF \nreg_reg[326]  ( .D(nreg[326]), .CLK(clk), .RST(rst), .I(e_init[326]), 
        .Q(nreg[326]) );
  DFF \nreg_reg[325]  ( .D(nreg[325]), .CLK(clk), .RST(rst), .I(e_init[325]), 
        .Q(nreg[325]) );
  DFF \nreg_reg[324]  ( .D(nreg[324]), .CLK(clk), .RST(rst), .I(e_init[324]), 
        .Q(nreg[324]) );
  DFF \nreg_reg[323]  ( .D(nreg[323]), .CLK(clk), .RST(rst), .I(e_init[323]), 
        .Q(nreg[323]) );
  DFF \nreg_reg[322]  ( .D(nreg[322]), .CLK(clk), .RST(rst), .I(e_init[322]), 
        .Q(nreg[322]) );
  DFF \nreg_reg[321]  ( .D(nreg[321]), .CLK(clk), .RST(rst), .I(e_init[321]), 
        .Q(nreg[321]) );
  DFF \nreg_reg[320]  ( .D(nreg[320]), .CLK(clk), .RST(rst), .I(e_init[320]), 
        .Q(nreg[320]) );
  DFF \nreg_reg[319]  ( .D(nreg[319]), .CLK(clk), .RST(rst), .I(e_init[319]), 
        .Q(nreg[319]) );
  DFF \nreg_reg[318]  ( .D(nreg[318]), .CLK(clk), .RST(rst), .I(e_init[318]), 
        .Q(nreg[318]) );
  DFF \nreg_reg[317]  ( .D(nreg[317]), .CLK(clk), .RST(rst), .I(e_init[317]), 
        .Q(nreg[317]) );
  DFF \nreg_reg[316]  ( .D(nreg[316]), .CLK(clk), .RST(rst), .I(e_init[316]), 
        .Q(nreg[316]) );
  DFF \nreg_reg[315]  ( .D(nreg[315]), .CLK(clk), .RST(rst), .I(e_init[315]), 
        .Q(nreg[315]) );
  DFF \nreg_reg[314]  ( .D(nreg[314]), .CLK(clk), .RST(rst), .I(e_init[314]), 
        .Q(nreg[314]) );
  DFF \nreg_reg[313]  ( .D(nreg[313]), .CLK(clk), .RST(rst), .I(e_init[313]), 
        .Q(nreg[313]) );
  DFF \nreg_reg[312]  ( .D(nreg[312]), .CLK(clk), .RST(rst), .I(e_init[312]), 
        .Q(nreg[312]) );
  DFF \nreg_reg[311]  ( .D(nreg[311]), .CLK(clk), .RST(rst), .I(e_init[311]), 
        .Q(nreg[311]) );
  DFF \nreg_reg[310]  ( .D(nreg[310]), .CLK(clk), .RST(rst), .I(e_init[310]), 
        .Q(nreg[310]) );
  DFF \nreg_reg[309]  ( .D(nreg[309]), .CLK(clk), .RST(rst), .I(e_init[309]), 
        .Q(nreg[309]) );
  DFF \nreg_reg[308]  ( .D(nreg[308]), .CLK(clk), .RST(rst), .I(e_init[308]), 
        .Q(nreg[308]) );
  DFF \nreg_reg[307]  ( .D(nreg[307]), .CLK(clk), .RST(rst), .I(e_init[307]), 
        .Q(nreg[307]) );
  DFF \nreg_reg[306]  ( .D(nreg[306]), .CLK(clk), .RST(rst), .I(e_init[306]), 
        .Q(nreg[306]) );
  DFF \nreg_reg[305]  ( .D(nreg[305]), .CLK(clk), .RST(rst), .I(e_init[305]), 
        .Q(nreg[305]) );
  DFF \nreg_reg[304]  ( .D(nreg[304]), .CLK(clk), .RST(rst), .I(e_init[304]), 
        .Q(nreg[304]) );
  DFF \nreg_reg[303]  ( .D(nreg[303]), .CLK(clk), .RST(rst), .I(e_init[303]), 
        .Q(nreg[303]) );
  DFF \nreg_reg[302]  ( .D(nreg[302]), .CLK(clk), .RST(rst), .I(e_init[302]), 
        .Q(nreg[302]) );
  DFF \nreg_reg[301]  ( .D(nreg[301]), .CLK(clk), .RST(rst), .I(e_init[301]), 
        .Q(nreg[301]) );
  DFF \nreg_reg[300]  ( .D(nreg[300]), .CLK(clk), .RST(rst), .I(e_init[300]), 
        .Q(nreg[300]) );
  DFF \nreg_reg[299]  ( .D(nreg[299]), .CLK(clk), .RST(rst), .I(e_init[299]), 
        .Q(nreg[299]) );
  DFF \nreg_reg[298]  ( .D(nreg[298]), .CLK(clk), .RST(rst), .I(e_init[298]), 
        .Q(nreg[298]) );
  DFF \nreg_reg[297]  ( .D(nreg[297]), .CLK(clk), .RST(rst), .I(e_init[297]), 
        .Q(nreg[297]) );
  DFF \nreg_reg[296]  ( .D(nreg[296]), .CLK(clk), .RST(rst), .I(e_init[296]), 
        .Q(nreg[296]) );
  DFF \nreg_reg[295]  ( .D(nreg[295]), .CLK(clk), .RST(rst), .I(e_init[295]), 
        .Q(nreg[295]) );
  DFF \nreg_reg[294]  ( .D(nreg[294]), .CLK(clk), .RST(rst), .I(e_init[294]), 
        .Q(nreg[294]) );
  DFF \nreg_reg[293]  ( .D(nreg[293]), .CLK(clk), .RST(rst), .I(e_init[293]), 
        .Q(nreg[293]) );
  DFF \nreg_reg[292]  ( .D(nreg[292]), .CLK(clk), .RST(rst), .I(e_init[292]), 
        .Q(nreg[292]) );
  DFF \nreg_reg[291]  ( .D(nreg[291]), .CLK(clk), .RST(rst), .I(e_init[291]), 
        .Q(nreg[291]) );
  DFF \nreg_reg[290]  ( .D(nreg[290]), .CLK(clk), .RST(rst), .I(e_init[290]), 
        .Q(nreg[290]) );
  DFF \nreg_reg[289]  ( .D(nreg[289]), .CLK(clk), .RST(rst), .I(e_init[289]), 
        .Q(nreg[289]) );
  DFF \nreg_reg[288]  ( .D(nreg[288]), .CLK(clk), .RST(rst), .I(e_init[288]), 
        .Q(nreg[288]) );
  DFF \nreg_reg[287]  ( .D(nreg[287]), .CLK(clk), .RST(rst), .I(e_init[287]), 
        .Q(nreg[287]) );
  DFF \nreg_reg[286]  ( .D(nreg[286]), .CLK(clk), .RST(rst), .I(e_init[286]), 
        .Q(nreg[286]) );
  DFF \nreg_reg[285]  ( .D(nreg[285]), .CLK(clk), .RST(rst), .I(e_init[285]), 
        .Q(nreg[285]) );
  DFF \nreg_reg[284]  ( .D(nreg[284]), .CLK(clk), .RST(rst), .I(e_init[284]), 
        .Q(nreg[284]) );
  DFF \nreg_reg[283]  ( .D(nreg[283]), .CLK(clk), .RST(rst), .I(e_init[283]), 
        .Q(nreg[283]) );
  DFF \nreg_reg[282]  ( .D(nreg[282]), .CLK(clk), .RST(rst), .I(e_init[282]), 
        .Q(nreg[282]) );
  DFF \nreg_reg[281]  ( .D(nreg[281]), .CLK(clk), .RST(rst), .I(e_init[281]), 
        .Q(nreg[281]) );
  DFF \nreg_reg[280]  ( .D(nreg[280]), .CLK(clk), .RST(rst), .I(e_init[280]), 
        .Q(nreg[280]) );
  DFF \nreg_reg[279]  ( .D(nreg[279]), .CLK(clk), .RST(rst), .I(e_init[279]), 
        .Q(nreg[279]) );
  DFF \nreg_reg[278]  ( .D(nreg[278]), .CLK(clk), .RST(rst), .I(e_init[278]), 
        .Q(nreg[278]) );
  DFF \nreg_reg[277]  ( .D(nreg[277]), .CLK(clk), .RST(rst), .I(e_init[277]), 
        .Q(nreg[277]) );
  DFF \nreg_reg[276]  ( .D(nreg[276]), .CLK(clk), .RST(rst), .I(e_init[276]), 
        .Q(nreg[276]) );
  DFF \nreg_reg[275]  ( .D(nreg[275]), .CLK(clk), .RST(rst), .I(e_init[275]), 
        .Q(nreg[275]) );
  DFF \nreg_reg[274]  ( .D(nreg[274]), .CLK(clk), .RST(rst), .I(e_init[274]), 
        .Q(nreg[274]) );
  DFF \nreg_reg[273]  ( .D(nreg[273]), .CLK(clk), .RST(rst), .I(e_init[273]), 
        .Q(nreg[273]) );
  DFF \nreg_reg[272]  ( .D(nreg[272]), .CLK(clk), .RST(rst), .I(e_init[272]), 
        .Q(nreg[272]) );
  DFF \nreg_reg[271]  ( .D(nreg[271]), .CLK(clk), .RST(rst), .I(e_init[271]), 
        .Q(nreg[271]) );
  DFF \nreg_reg[270]  ( .D(nreg[270]), .CLK(clk), .RST(rst), .I(e_init[270]), 
        .Q(nreg[270]) );
  DFF \nreg_reg[269]  ( .D(nreg[269]), .CLK(clk), .RST(rst), .I(e_init[269]), 
        .Q(nreg[269]) );
  DFF \nreg_reg[268]  ( .D(nreg[268]), .CLK(clk), .RST(rst), .I(e_init[268]), 
        .Q(nreg[268]) );
  DFF \nreg_reg[267]  ( .D(nreg[267]), .CLK(clk), .RST(rst), .I(e_init[267]), 
        .Q(nreg[267]) );
  DFF \nreg_reg[266]  ( .D(nreg[266]), .CLK(clk), .RST(rst), .I(e_init[266]), 
        .Q(nreg[266]) );
  DFF \nreg_reg[265]  ( .D(nreg[265]), .CLK(clk), .RST(rst), .I(e_init[265]), 
        .Q(nreg[265]) );
  DFF \nreg_reg[264]  ( .D(nreg[264]), .CLK(clk), .RST(rst), .I(e_init[264]), 
        .Q(nreg[264]) );
  DFF \nreg_reg[263]  ( .D(nreg[263]), .CLK(clk), .RST(rst), .I(e_init[263]), 
        .Q(nreg[263]) );
  DFF \nreg_reg[262]  ( .D(nreg[262]), .CLK(clk), .RST(rst), .I(e_init[262]), 
        .Q(nreg[262]) );
  DFF \nreg_reg[261]  ( .D(nreg[261]), .CLK(clk), .RST(rst), .I(e_init[261]), 
        .Q(nreg[261]) );
  DFF \nreg_reg[260]  ( .D(nreg[260]), .CLK(clk), .RST(rst), .I(e_init[260]), 
        .Q(nreg[260]) );
  DFF \nreg_reg[259]  ( .D(nreg[259]), .CLK(clk), .RST(rst), .I(e_init[259]), 
        .Q(nreg[259]) );
  DFF \nreg_reg[258]  ( .D(nreg[258]), .CLK(clk), .RST(rst), .I(e_init[258]), 
        .Q(nreg[258]) );
  DFF \nreg_reg[257]  ( .D(nreg[257]), .CLK(clk), .RST(rst), .I(e_init[257]), 
        .Q(nreg[257]) );
  DFF \nreg_reg[256]  ( .D(nreg[256]), .CLK(clk), .RST(rst), .I(e_init[256]), 
        .Q(nreg[256]) );
  DFF \nreg_reg[255]  ( .D(nreg[255]), .CLK(clk), .RST(rst), .I(e_init[255]), 
        .Q(nreg[255]) );
  DFF \nreg_reg[254]  ( .D(nreg[254]), .CLK(clk), .RST(rst), .I(e_init[254]), 
        .Q(nreg[254]) );
  DFF \nreg_reg[253]  ( .D(nreg[253]), .CLK(clk), .RST(rst), .I(e_init[253]), 
        .Q(nreg[253]) );
  DFF \nreg_reg[252]  ( .D(nreg[252]), .CLK(clk), .RST(rst), .I(e_init[252]), 
        .Q(nreg[252]) );
  DFF \nreg_reg[251]  ( .D(nreg[251]), .CLK(clk), .RST(rst), .I(e_init[251]), 
        .Q(nreg[251]) );
  DFF \nreg_reg[250]  ( .D(nreg[250]), .CLK(clk), .RST(rst), .I(e_init[250]), 
        .Q(nreg[250]) );
  DFF \nreg_reg[249]  ( .D(nreg[249]), .CLK(clk), .RST(rst), .I(e_init[249]), 
        .Q(nreg[249]) );
  DFF \nreg_reg[248]  ( .D(nreg[248]), .CLK(clk), .RST(rst), .I(e_init[248]), 
        .Q(nreg[248]) );
  DFF \nreg_reg[247]  ( .D(nreg[247]), .CLK(clk), .RST(rst), .I(e_init[247]), 
        .Q(nreg[247]) );
  DFF \nreg_reg[246]  ( .D(nreg[246]), .CLK(clk), .RST(rst), .I(e_init[246]), 
        .Q(nreg[246]) );
  DFF \nreg_reg[245]  ( .D(nreg[245]), .CLK(clk), .RST(rst), .I(e_init[245]), 
        .Q(nreg[245]) );
  DFF \nreg_reg[244]  ( .D(nreg[244]), .CLK(clk), .RST(rst), .I(e_init[244]), 
        .Q(nreg[244]) );
  DFF \nreg_reg[243]  ( .D(nreg[243]), .CLK(clk), .RST(rst), .I(e_init[243]), 
        .Q(nreg[243]) );
  DFF \nreg_reg[242]  ( .D(nreg[242]), .CLK(clk), .RST(rst), .I(e_init[242]), 
        .Q(nreg[242]) );
  DFF \nreg_reg[241]  ( .D(nreg[241]), .CLK(clk), .RST(rst), .I(e_init[241]), 
        .Q(nreg[241]) );
  DFF \nreg_reg[240]  ( .D(nreg[240]), .CLK(clk), .RST(rst), .I(e_init[240]), 
        .Q(nreg[240]) );
  DFF \nreg_reg[239]  ( .D(nreg[239]), .CLK(clk), .RST(rst), .I(e_init[239]), 
        .Q(nreg[239]) );
  DFF \nreg_reg[238]  ( .D(nreg[238]), .CLK(clk), .RST(rst), .I(e_init[238]), 
        .Q(nreg[238]) );
  DFF \nreg_reg[237]  ( .D(nreg[237]), .CLK(clk), .RST(rst), .I(e_init[237]), 
        .Q(nreg[237]) );
  DFF \nreg_reg[236]  ( .D(nreg[236]), .CLK(clk), .RST(rst), .I(e_init[236]), 
        .Q(nreg[236]) );
  DFF \nreg_reg[235]  ( .D(nreg[235]), .CLK(clk), .RST(rst), .I(e_init[235]), 
        .Q(nreg[235]) );
  DFF \nreg_reg[234]  ( .D(nreg[234]), .CLK(clk), .RST(rst), .I(e_init[234]), 
        .Q(nreg[234]) );
  DFF \nreg_reg[233]  ( .D(nreg[233]), .CLK(clk), .RST(rst), .I(e_init[233]), 
        .Q(nreg[233]) );
  DFF \nreg_reg[232]  ( .D(nreg[232]), .CLK(clk), .RST(rst), .I(e_init[232]), 
        .Q(nreg[232]) );
  DFF \nreg_reg[231]  ( .D(nreg[231]), .CLK(clk), .RST(rst), .I(e_init[231]), 
        .Q(nreg[231]) );
  DFF \nreg_reg[230]  ( .D(nreg[230]), .CLK(clk), .RST(rst), .I(e_init[230]), 
        .Q(nreg[230]) );
  DFF \nreg_reg[229]  ( .D(nreg[229]), .CLK(clk), .RST(rst), .I(e_init[229]), 
        .Q(nreg[229]) );
  DFF \nreg_reg[228]  ( .D(nreg[228]), .CLK(clk), .RST(rst), .I(e_init[228]), 
        .Q(nreg[228]) );
  DFF \nreg_reg[227]  ( .D(nreg[227]), .CLK(clk), .RST(rst), .I(e_init[227]), 
        .Q(nreg[227]) );
  DFF \nreg_reg[226]  ( .D(nreg[226]), .CLK(clk), .RST(rst), .I(e_init[226]), 
        .Q(nreg[226]) );
  DFF \nreg_reg[225]  ( .D(nreg[225]), .CLK(clk), .RST(rst), .I(e_init[225]), 
        .Q(nreg[225]) );
  DFF \nreg_reg[224]  ( .D(nreg[224]), .CLK(clk), .RST(rst), .I(e_init[224]), 
        .Q(nreg[224]) );
  DFF \nreg_reg[223]  ( .D(nreg[223]), .CLK(clk), .RST(rst), .I(e_init[223]), 
        .Q(nreg[223]) );
  DFF \nreg_reg[222]  ( .D(nreg[222]), .CLK(clk), .RST(rst), .I(e_init[222]), 
        .Q(nreg[222]) );
  DFF \nreg_reg[221]  ( .D(nreg[221]), .CLK(clk), .RST(rst), .I(e_init[221]), 
        .Q(nreg[221]) );
  DFF \nreg_reg[220]  ( .D(nreg[220]), .CLK(clk), .RST(rst), .I(e_init[220]), 
        .Q(nreg[220]) );
  DFF \nreg_reg[219]  ( .D(nreg[219]), .CLK(clk), .RST(rst), .I(e_init[219]), 
        .Q(nreg[219]) );
  DFF \nreg_reg[218]  ( .D(nreg[218]), .CLK(clk), .RST(rst), .I(e_init[218]), 
        .Q(nreg[218]) );
  DFF \nreg_reg[217]  ( .D(nreg[217]), .CLK(clk), .RST(rst), .I(e_init[217]), 
        .Q(nreg[217]) );
  DFF \nreg_reg[216]  ( .D(nreg[216]), .CLK(clk), .RST(rst), .I(e_init[216]), 
        .Q(nreg[216]) );
  DFF \nreg_reg[215]  ( .D(nreg[215]), .CLK(clk), .RST(rst), .I(e_init[215]), 
        .Q(nreg[215]) );
  DFF \nreg_reg[214]  ( .D(nreg[214]), .CLK(clk), .RST(rst), .I(e_init[214]), 
        .Q(nreg[214]) );
  DFF \nreg_reg[213]  ( .D(nreg[213]), .CLK(clk), .RST(rst), .I(e_init[213]), 
        .Q(nreg[213]) );
  DFF \nreg_reg[212]  ( .D(nreg[212]), .CLK(clk), .RST(rst), .I(e_init[212]), 
        .Q(nreg[212]) );
  DFF \nreg_reg[211]  ( .D(nreg[211]), .CLK(clk), .RST(rst), .I(e_init[211]), 
        .Q(nreg[211]) );
  DFF \nreg_reg[210]  ( .D(nreg[210]), .CLK(clk), .RST(rst), .I(e_init[210]), 
        .Q(nreg[210]) );
  DFF \nreg_reg[209]  ( .D(nreg[209]), .CLK(clk), .RST(rst), .I(e_init[209]), 
        .Q(nreg[209]) );
  DFF \nreg_reg[208]  ( .D(nreg[208]), .CLK(clk), .RST(rst), .I(e_init[208]), 
        .Q(nreg[208]) );
  DFF \nreg_reg[207]  ( .D(nreg[207]), .CLK(clk), .RST(rst), .I(e_init[207]), 
        .Q(nreg[207]) );
  DFF \nreg_reg[206]  ( .D(nreg[206]), .CLK(clk), .RST(rst), .I(e_init[206]), 
        .Q(nreg[206]) );
  DFF \nreg_reg[205]  ( .D(nreg[205]), .CLK(clk), .RST(rst), .I(e_init[205]), 
        .Q(nreg[205]) );
  DFF \nreg_reg[204]  ( .D(nreg[204]), .CLK(clk), .RST(rst), .I(e_init[204]), 
        .Q(nreg[204]) );
  DFF \nreg_reg[203]  ( .D(nreg[203]), .CLK(clk), .RST(rst), .I(e_init[203]), 
        .Q(nreg[203]) );
  DFF \nreg_reg[202]  ( .D(nreg[202]), .CLK(clk), .RST(rst), .I(e_init[202]), 
        .Q(nreg[202]) );
  DFF \nreg_reg[201]  ( .D(nreg[201]), .CLK(clk), .RST(rst), .I(e_init[201]), 
        .Q(nreg[201]) );
  DFF \nreg_reg[200]  ( .D(nreg[200]), .CLK(clk), .RST(rst), .I(e_init[200]), 
        .Q(nreg[200]) );
  DFF \nreg_reg[199]  ( .D(nreg[199]), .CLK(clk), .RST(rst), .I(e_init[199]), 
        .Q(nreg[199]) );
  DFF \nreg_reg[198]  ( .D(nreg[198]), .CLK(clk), .RST(rst), .I(e_init[198]), 
        .Q(nreg[198]) );
  DFF \nreg_reg[197]  ( .D(nreg[197]), .CLK(clk), .RST(rst), .I(e_init[197]), 
        .Q(nreg[197]) );
  DFF \nreg_reg[196]  ( .D(nreg[196]), .CLK(clk), .RST(rst), .I(e_init[196]), 
        .Q(nreg[196]) );
  DFF \nreg_reg[195]  ( .D(nreg[195]), .CLK(clk), .RST(rst), .I(e_init[195]), 
        .Q(nreg[195]) );
  DFF \nreg_reg[194]  ( .D(nreg[194]), .CLK(clk), .RST(rst), .I(e_init[194]), 
        .Q(nreg[194]) );
  DFF \nreg_reg[193]  ( .D(nreg[193]), .CLK(clk), .RST(rst), .I(e_init[193]), 
        .Q(nreg[193]) );
  DFF \nreg_reg[192]  ( .D(nreg[192]), .CLK(clk), .RST(rst), .I(e_init[192]), 
        .Q(nreg[192]) );
  DFF \nreg_reg[191]  ( .D(nreg[191]), .CLK(clk), .RST(rst), .I(e_init[191]), 
        .Q(nreg[191]) );
  DFF \nreg_reg[190]  ( .D(nreg[190]), .CLK(clk), .RST(rst), .I(e_init[190]), 
        .Q(nreg[190]) );
  DFF \nreg_reg[189]  ( .D(nreg[189]), .CLK(clk), .RST(rst), .I(e_init[189]), 
        .Q(nreg[189]) );
  DFF \nreg_reg[188]  ( .D(nreg[188]), .CLK(clk), .RST(rst), .I(e_init[188]), 
        .Q(nreg[188]) );
  DFF \nreg_reg[187]  ( .D(nreg[187]), .CLK(clk), .RST(rst), .I(e_init[187]), 
        .Q(nreg[187]) );
  DFF \nreg_reg[186]  ( .D(nreg[186]), .CLK(clk), .RST(rst), .I(e_init[186]), 
        .Q(nreg[186]) );
  DFF \nreg_reg[185]  ( .D(nreg[185]), .CLK(clk), .RST(rst), .I(e_init[185]), 
        .Q(nreg[185]) );
  DFF \nreg_reg[184]  ( .D(nreg[184]), .CLK(clk), .RST(rst), .I(e_init[184]), 
        .Q(nreg[184]) );
  DFF \nreg_reg[183]  ( .D(nreg[183]), .CLK(clk), .RST(rst), .I(e_init[183]), 
        .Q(nreg[183]) );
  DFF \nreg_reg[182]  ( .D(nreg[182]), .CLK(clk), .RST(rst), .I(e_init[182]), 
        .Q(nreg[182]) );
  DFF \nreg_reg[181]  ( .D(nreg[181]), .CLK(clk), .RST(rst), .I(e_init[181]), 
        .Q(nreg[181]) );
  DFF \nreg_reg[180]  ( .D(nreg[180]), .CLK(clk), .RST(rst), .I(e_init[180]), 
        .Q(nreg[180]) );
  DFF \nreg_reg[179]  ( .D(nreg[179]), .CLK(clk), .RST(rst), .I(e_init[179]), 
        .Q(nreg[179]) );
  DFF \nreg_reg[178]  ( .D(nreg[178]), .CLK(clk), .RST(rst), .I(e_init[178]), 
        .Q(nreg[178]) );
  DFF \nreg_reg[177]  ( .D(nreg[177]), .CLK(clk), .RST(rst), .I(e_init[177]), 
        .Q(nreg[177]) );
  DFF \nreg_reg[176]  ( .D(nreg[176]), .CLK(clk), .RST(rst), .I(e_init[176]), 
        .Q(nreg[176]) );
  DFF \nreg_reg[175]  ( .D(nreg[175]), .CLK(clk), .RST(rst), .I(e_init[175]), 
        .Q(nreg[175]) );
  DFF \nreg_reg[174]  ( .D(nreg[174]), .CLK(clk), .RST(rst), .I(e_init[174]), 
        .Q(nreg[174]) );
  DFF \nreg_reg[173]  ( .D(nreg[173]), .CLK(clk), .RST(rst), .I(e_init[173]), 
        .Q(nreg[173]) );
  DFF \nreg_reg[172]  ( .D(nreg[172]), .CLK(clk), .RST(rst), .I(e_init[172]), 
        .Q(nreg[172]) );
  DFF \nreg_reg[171]  ( .D(nreg[171]), .CLK(clk), .RST(rst), .I(e_init[171]), 
        .Q(nreg[171]) );
  DFF \nreg_reg[170]  ( .D(nreg[170]), .CLK(clk), .RST(rst), .I(e_init[170]), 
        .Q(nreg[170]) );
  DFF \nreg_reg[169]  ( .D(nreg[169]), .CLK(clk), .RST(rst), .I(e_init[169]), 
        .Q(nreg[169]) );
  DFF \nreg_reg[168]  ( .D(nreg[168]), .CLK(clk), .RST(rst), .I(e_init[168]), 
        .Q(nreg[168]) );
  DFF \nreg_reg[167]  ( .D(nreg[167]), .CLK(clk), .RST(rst), .I(e_init[167]), 
        .Q(nreg[167]) );
  DFF \nreg_reg[166]  ( .D(nreg[166]), .CLK(clk), .RST(rst), .I(e_init[166]), 
        .Q(nreg[166]) );
  DFF \nreg_reg[165]  ( .D(nreg[165]), .CLK(clk), .RST(rst), .I(e_init[165]), 
        .Q(nreg[165]) );
  DFF \nreg_reg[164]  ( .D(nreg[164]), .CLK(clk), .RST(rst), .I(e_init[164]), 
        .Q(nreg[164]) );
  DFF \nreg_reg[163]  ( .D(nreg[163]), .CLK(clk), .RST(rst), .I(e_init[163]), 
        .Q(nreg[163]) );
  DFF \nreg_reg[162]  ( .D(nreg[162]), .CLK(clk), .RST(rst), .I(e_init[162]), 
        .Q(nreg[162]) );
  DFF \nreg_reg[161]  ( .D(nreg[161]), .CLK(clk), .RST(rst), .I(e_init[161]), 
        .Q(nreg[161]) );
  DFF \nreg_reg[160]  ( .D(nreg[160]), .CLK(clk), .RST(rst), .I(e_init[160]), 
        .Q(nreg[160]) );
  DFF \nreg_reg[159]  ( .D(nreg[159]), .CLK(clk), .RST(rst), .I(e_init[159]), 
        .Q(nreg[159]) );
  DFF \nreg_reg[158]  ( .D(nreg[158]), .CLK(clk), .RST(rst), .I(e_init[158]), 
        .Q(nreg[158]) );
  DFF \nreg_reg[157]  ( .D(nreg[157]), .CLK(clk), .RST(rst), .I(e_init[157]), 
        .Q(nreg[157]) );
  DFF \nreg_reg[156]  ( .D(nreg[156]), .CLK(clk), .RST(rst), .I(e_init[156]), 
        .Q(nreg[156]) );
  DFF \nreg_reg[155]  ( .D(nreg[155]), .CLK(clk), .RST(rst), .I(e_init[155]), 
        .Q(nreg[155]) );
  DFF \nreg_reg[154]  ( .D(nreg[154]), .CLK(clk), .RST(rst), .I(e_init[154]), 
        .Q(nreg[154]) );
  DFF \nreg_reg[153]  ( .D(nreg[153]), .CLK(clk), .RST(rst), .I(e_init[153]), 
        .Q(nreg[153]) );
  DFF \nreg_reg[152]  ( .D(nreg[152]), .CLK(clk), .RST(rst), .I(e_init[152]), 
        .Q(nreg[152]) );
  DFF \nreg_reg[151]  ( .D(nreg[151]), .CLK(clk), .RST(rst), .I(e_init[151]), 
        .Q(nreg[151]) );
  DFF \nreg_reg[150]  ( .D(nreg[150]), .CLK(clk), .RST(rst), .I(e_init[150]), 
        .Q(nreg[150]) );
  DFF \nreg_reg[149]  ( .D(nreg[149]), .CLK(clk), .RST(rst), .I(e_init[149]), 
        .Q(nreg[149]) );
  DFF \nreg_reg[148]  ( .D(nreg[148]), .CLK(clk), .RST(rst), .I(e_init[148]), 
        .Q(nreg[148]) );
  DFF \nreg_reg[147]  ( .D(nreg[147]), .CLK(clk), .RST(rst), .I(e_init[147]), 
        .Q(nreg[147]) );
  DFF \nreg_reg[146]  ( .D(nreg[146]), .CLK(clk), .RST(rst), .I(e_init[146]), 
        .Q(nreg[146]) );
  DFF \nreg_reg[145]  ( .D(nreg[145]), .CLK(clk), .RST(rst), .I(e_init[145]), 
        .Q(nreg[145]) );
  DFF \nreg_reg[144]  ( .D(nreg[144]), .CLK(clk), .RST(rst), .I(e_init[144]), 
        .Q(nreg[144]) );
  DFF \nreg_reg[143]  ( .D(nreg[143]), .CLK(clk), .RST(rst), .I(e_init[143]), 
        .Q(nreg[143]) );
  DFF \nreg_reg[142]  ( .D(nreg[142]), .CLK(clk), .RST(rst), .I(e_init[142]), 
        .Q(nreg[142]) );
  DFF \nreg_reg[141]  ( .D(nreg[141]), .CLK(clk), .RST(rst), .I(e_init[141]), 
        .Q(nreg[141]) );
  DFF \nreg_reg[140]  ( .D(nreg[140]), .CLK(clk), .RST(rst), .I(e_init[140]), 
        .Q(nreg[140]) );
  DFF \nreg_reg[139]  ( .D(nreg[139]), .CLK(clk), .RST(rst), .I(e_init[139]), 
        .Q(nreg[139]) );
  DFF \nreg_reg[138]  ( .D(nreg[138]), .CLK(clk), .RST(rst), .I(e_init[138]), 
        .Q(nreg[138]) );
  DFF \nreg_reg[137]  ( .D(nreg[137]), .CLK(clk), .RST(rst), .I(e_init[137]), 
        .Q(nreg[137]) );
  DFF \nreg_reg[136]  ( .D(nreg[136]), .CLK(clk), .RST(rst), .I(e_init[136]), 
        .Q(nreg[136]) );
  DFF \nreg_reg[135]  ( .D(nreg[135]), .CLK(clk), .RST(rst), .I(e_init[135]), 
        .Q(nreg[135]) );
  DFF \nreg_reg[134]  ( .D(nreg[134]), .CLK(clk), .RST(rst), .I(e_init[134]), 
        .Q(nreg[134]) );
  DFF \nreg_reg[133]  ( .D(nreg[133]), .CLK(clk), .RST(rst), .I(e_init[133]), 
        .Q(nreg[133]) );
  DFF \nreg_reg[132]  ( .D(nreg[132]), .CLK(clk), .RST(rst), .I(e_init[132]), 
        .Q(nreg[132]) );
  DFF \nreg_reg[131]  ( .D(nreg[131]), .CLK(clk), .RST(rst), .I(e_init[131]), 
        .Q(nreg[131]) );
  DFF \nreg_reg[130]  ( .D(nreg[130]), .CLK(clk), .RST(rst), .I(e_init[130]), 
        .Q(nreg[130]) );
  DFF \nreg_reg[129]  ( .D(nreg[129]), .CLK(clk), .RST(rst), .I(e_init[129]), 
        .Q(nreg[129]) );
  DFF \nreg_reg[128]  ( .D(nreg[128]), .CLK(clk), .RST(rst), .I(e_init[128]), 
        .Q(nreg[128]) );
  DFF \nreg_reg[127]  ( .D(nreg[127]), .CLK(clk), .RST(rst), .I(e_init[127]), 
        .Q(nreg[127]) );
  DFF \nreg_reg[126]  ( .D(nreg[126]), .CLK(clk), .RST(rst), .I(e_init[126]), 
        .Q(nreg[126]) );
  DFF \nreg_reg[125]  ( .D(nreg[125]), .CLK(clk), .RST(rst), .I(e_init[125]), 
        .Q(nreg[125]) );
  DFF \nreg_reg[124]  ( .D(nreg[124]), .CLK(clk), .RST(rst), .I(e_init[124]), 
        .Q(nreg[124]) );
  DFF \nreg_reg[123]  ( .D(nreg[123]), .CLK(clk), .RST(rst), .I(e_init[123]), 
        .Q(nreg[123]) );
  DFF \nreg_reg[122]  ( .D(nreg[122]), .CLK(clk), .RST(rst), .I(e_init[122]), 
        .Q(nreg[122]) );
  DFF \nreg_reg[121]  ( .D(nreg[121]), .CLK(clk), .RST(rst), .I(e_init[121]), 
        .Q(nreg[121]) );
  DFF \nreg_reg[120]  ( .D(nreg[120]), .CLK(clk), .RST(rst), .I(e_init[120]), 
        .Q(nreg[120]) );
  DFF \nreg_reg[119]  ( .D(nreg[119]), .CLK(clk), .RST(rst), .I(e_init[119]), 
        .Q(nreg[119]) );
  DFF \nreg_reg[118]  ( .D(nreg[118]), .CLK(clk), .RST(rst), .I(e_init[118]), 
        .Q(nreg[118]) );
  DFF \nreg_reg[117]  ( .D(nreg[117]), .CLK(clk), .RST(rst), .I(e_init[117]), 
        .Q(nreg[117]) );
  DFF \nreg_reg[116]  ( .D(nreg[116]), .CLK(clk), .RST(rst), .I(e_init[116]), 
        .Q(nreg[116]) );
  DFF \nreg_reg[115]  ( .D(nreg[115]), .CLK(clk), .RST(rst), .I(e_init[115]), 
        .Q(nreg[115]) );
  DFF \nreg_reg[114]  ( .D(nreg[114]), .CLK(clk), .RST(rst), .I(e_init[114]), 
        .Q(nreg[114]) );
  DFF \nreg_reg[113]  ( .D(nreg[113]), .CLK(clk), .RST(rst), .I(e_init[113]), 
        .Q(nreg[113]) );
  DFF \nreg_reg[112]  ( .D(nreg[112]), .CLK(clk), .RST(rst), .I(e_init[112]), 
        .Q(nreg[112]) );
  DFF \nreg_reg[111]  ( .D(nreg[111]), .CLK(clk), .RST(rst), .I(e_init[111]), 
        .Q(nreg[111]) );
  DFF \nreg_reg[110]  ( .D(nreg[110]), .CLK(clk), .RST(rst), .I(e_init[110]), 
        .Q(nreg[110]) );
  DFF \nreg_reg[109]  ( .D(nreg[109]), .CLK(clk), .RST(rst), .I(e_init[109]), 
        .Q(nreg[109]) );
  DFF \nreg_reg[108]  ( .D(nreg[108]), .CLK(clk), .RST(rst), .I(e_init[108]), 
        .Q(nreg[108]) );
  DFF \nreg_reg[107]  ( .D(nreg[107]), .CLK(clk), .RST(rst), .I(e_init[107]), 
        .Q(nreg[107]) );
  DFF \nreg_reg[106]  ( .D(nreg[106]), .CLK(clk), .RST(rst), .I(e_init[106]), 
        .Q(nreg[106]) );
  DFF \nreg_reg[105]  ( .D(nreg[105]), .CLK(clk), .RST(rst), .I(e_init[105]), 
        .Q(nreg[105]) );
  DFF \nreg_reg[104]  ( .D(nreg[104]), .CLK(clk), .RST(rst), .I(e_init[104]), 
        .Q(nreg[104]) );
  DFF \nreg_reg[103]  ( .D(nreg[103]), .CLK(clk), .RST(rst), .I(e_init[103]), 
        .Q(nreg[103]) );
  DFF \nreg_reg[102]  ( .D(nreg[102]), .CLK(clk), .RST(rst), .I(e_init[102]), 
        .Q(nreg[102]) );
  DFF \nreg_reg[101]  ( .D(nreg[101]), .CLK(clk), .RST(rst), .I(e_init[101]), 
        .Q(nreg[101]) );
  DFF \nreg_reg[100]  ( .D(nreg[100]), .CLK(clk), .RST(rst), .I(e_init[100]), 
        .Q(nreg[100]) );
  DFF \nreg_reg[99]  ( .D(nreg[99]), .CLK(clk), .RST(rst), .I(e_init[99]), .Q(
        nreg[99]) );
  DFF \nreg_reg[98]  ( .D(nreg[98]), .CLK(clk), .RST(rst), .I(e_init[98]), .Q(
        nreg[98]) );
  DFF \nreg_reg[97]  ( .D(nreg[97]), .CLK(clk), .RST(rst), .I(e_init[97]), .Q(
        nreg[97]) );
  DFF \nreg_reg[96]  ( .D(nreg[96]), .CLK(clk), .RST(rst), .I(e_init[96]), .Q(
        nreg[96]) );
  DFF \nreg_reg[95]  ( .D(nreg[95]), .CLK(clk), .RST(rst), .I(e_init[95]), .Q(
        nreg[95]) );
  DFF \nreg_reg[94]  ( .D(nreg[94]), .CLK(clk), .RST(rst), .I(e_init[94]), .Q(
        nreg[94]) );
  DFF \nreg_reg[93]  ( .D(nreg[93]), .CLK(clk), .RST(rst), .I(e_init[93]), .Q(
        nreg[93]) );
  DFF \nreg_reg[92]  ( .D(nreg[92]), .CLK(clk), .RST(rst), .I(e_init[92]), .Q(
        nreg[92]) );
  DFF \nreg_reg[91]  ( .D(nreg[91]), .CLK(clk), .RST(rst), .I(e_init[91]), .Q(
        nreg[91]) );
  DFF \nreg_reg[90]  ( .D(nreg[90]), .CLK(clk), .RST(rst), .I(e_init[90]), .Q(
        nreg[90]) );
  DFF \nreg_reg[89]  ( .D(nreg[89]), .CLK(clk), .RST(rst), .I(e_init[89]), .Q(
        nreg[89]) );
  DFF \nreg_reg[88]  ( .D(nreg[88]), .CLK(clk), .RST(rst), .I(e_init[88]), .Q(
        nreg[88]) );
  DFF \nreg_reg[87]  ( .D(nreg[87]), .CLK(clk), .RST(rst), .I(e_init[87]), .Q(
        nreg[87]) );
  DFF \nreg_reg[86]  ( .D(nreg[86]), .CLK(clk), .RST(rst), .I(e_init[86]), .Q(
        nreg[86]) );
  DFF \nreg_reg[85]  ( .D(nreg[85]), .CLK(clk), .RST(rst), .I(e_init[85]), .Q(
        nreg[85]) );
  DFF \nreg_reg[84]  ( .D(nreg[84]), .CLK(clk), .RST(rst), .I(e_init[84]), .Q(
        nreg[84]) );
  DFF \nreg_reg[83]  ( .D(nreg[83]), .CLK(clk), .RST(rst), .I(e_init[83]), .Q(
        nreg[83]) );
  DFF \nreg_reg[82]  ( .D(nreg[82]), .CLK(clk), .RST(rst), .I(e_init[82]), .Q(
        nreg[82]) );
  DFF \nreg_reg[81]  ( .D(nreg[81]), .CLK(clk), .RST(rst), .I(e_init[81]), .Q(
        nreg[81]) );
  DFF \nreg_reg[80]  ( .D(nreg[80]), .CLK(clk), .RST(rst), .I(e_init[80]), .Q(
        nreg[80]) );
  DFF \nreg_reg[79]  ( .D(nreg[79]), .CLK(clk), .RST(rst), .I(e_init[79]), .Q(
        nreg[79]) );
  DFF \nreg_reg[78]  ( .D(nreg[78]), .CLK(clk), .RST(rst), .I(e_init[78]), .Q(
        nreg[78]) );
  DFF \nreg_reg[77]  ( .D(nreg[77]), .CLK(clk), .RST(rst), .I(e_init[77]), .Q(
        nreg[77]) );
  DFF \nreg_reg[76]  ( .D(nreg[76]), .CLK(clk), .RST(rst), .I(e_init[76]), .Q(
        nreg[76]) );
  DFF \nreg_reg[75]  ( .D(nreg[75]), .CLK(clk), .RST(rst), .I(e_init[75]), .Q(
        nreg[75]) );
  DFF \nreg_reg[74]  ( .D(nreg[74]), .CLK(clk), .RST(rst), .I(e_init[74]), .Q(
        nreg[74]) );
  DFF \nreg_reg[73]  ( .D(nreg[73]), .CLK(clk), .RST(rst), .I(e_init[73]), .Q(
        nreg[73]) );
  DFF \nreg_reg[72]  ( .D(nreg[72]), .CLK(clk), .RST(rst), .I(e_init[72]), .Q(
        nreg[72]) );
  DFF \nreg_reg[71]  ( .D(nreg[71]), .CLK(clk), .RST(rst), .I(e_init[71]), .Q(
        nreg[71]) );
  DFF \nreg_reg[70]  ( .D(nreg[70]), .CLK(clk), .RST(rst), .I(e_init[70]), .Q(
        nreg[70]) );
  DFF \nreg_reg[69]  ( .D(nreg[69]), .CLK(clk), .RST(rst), .I(e_init[69]), .Q(
        nreg[69]) );
  DFF \nreg_reg[68]  ( .D(nreg[68]), .CLK(clk), .RST(rst), .I(e_init[68]), .Q(
        nreg[68]) );
  DFF \nreg_reg[67]  ( .D(nreg[67]), .CLK(clk), .RST(rst), .I(e_init[67]), .Q(
        nreg[67]) );
  DFF \nreg_reg[66]  ( .D(nreg[66]), .CLK(clk), .RST(rst), .I(e_init[66]), .Q(
        nreg[66]) );
  DFF \nreg_reg[65]  ( .D(nreg[65]), .CLK(clk), .RST(rst), .I(e_init[65]), .Q(
        nreg[65]) );
  DFF \nreg_reg[64]  ( .D(nreg[64]), .CLK(clk), .RST(rst), .I(e_init[64]), .Q(
        nreg[64]) );
  DFF \nreg_reg[63]  ( .D(nreg[63]), .CLK(clk), .RST(rst), .I(e_init[63]), .Q(
        nreg[63]) );
  DFF \nreg_reg[62]  ( .D(nreg[62]), .CLK(clk), .RST(rst), .I(e_init[62]), .Q(
        nreg[62]) );
  DFF \nreg_reg[61]  ( .D(nreg[61]), .CLK(clk), .RST(rst), .I(e_init[61]), .Q(
        nreg[61]) );
  DFF \nreg_reg[60]  ( .D(nreg[60]), .CLK(clk), .RST(rst), .I(e_init[60]), .Q(
        nreg[60]) );
  DFF \nreg_reg[59]  ( .D(nreg[59]), .CLK(clk), .RST(rst), .I(e_init[59]), .Q(
        nreg[59]) );
  DFF \nreg_reg[58]  ( .D(nreg[58]), .CLK(clk), .RST(rst), .I(e_init[58]), .Q(
        nreg[58]) );
  DFF \nreg_reg[57]  ( .D(nreg[57]), .CLK(clk), .RST(rst), .I(e_init[57]), .Q(
        nreg[57]) );
  DFF \nreg_reg[56]  ( .D(nreg[56]), .CLK(clk), .RST(rst), .I(e_init[56]), .Q(
        nreg[56]) );
  DFF \nreg_reg[55]  ( .D(nreg[55]), .CLK(clk), .RST(rst), .I(e_init[55]), .Q(
        nreg[55]) );
  DFF \nreg_reg[54]  ( .D(nreg[54]), .CLK(clk), .RST(rst), .I(e_init[54]), .Q(
        nreg[54]) );
  DFF \nreg_reg[53]  ( .D(nreg[53]), .CLK(clk), .RST(rst), .I(e_init[53]), .Q(
        nreg[53]) );
  DFF \nreg_reg[52]  ( .D(nreg[52]), .CLK(clk), .RST(rst), .I(e_init[52]), .Q(
        nreg[52]) );
  DFF \nreg_reg[51]  ( .D(nreg[51]), .CLK(clk), .RST(rst), .I(e_init[51]), .Q(
        nreg[51]) );
  DFF \nreg_reg[50]  ( .D(nreg[50]), .CLK(clk), .RST(rst), .I(e_init[50]), .Q(
        nreg[50]) );
  DFF \nreg_reg[49]  ( .D(nreg[49]), .CLK(clk), .RST(rst), .I(e_init[49]), .Q(
        nreg[49]) );
  DFF \nreg_reg[48]  ( .D(nreg[48]), .CLK(clk), .RST(rst), .I(e_init[48]), .Q(
        nreg[48]) );
  DFF \nreg_reg[47]  ( .D(nreg[47]), .CLK(clk), .RST(rst), .I(e_init[47]), .Q(
        nreg[47]) );
  DFF \nreg_reg[46]  ( .D(nreg[46]), .CLK(clk), .RST(rst), .I(e_init[46]), .Q(
        nreg[46]) );
  DFF \nreg_reg[45]  ( .D(nreg[45]), .CLK(clk), .RST(rst), .I(e_init[45]), .Q(
        nreg[45]) );
  DFF \nreg_reg[44]  ( .D(nreg[44]), .CLK(clk), .RST(rst), .I(e_init[44]), .Q(
        nreg[44]) );
  DFF \nreg_reg[43]  ( .D(nreg[43]), .CLK(clk), .RST(rst), .I(e_init[43]), .Q(
        nreg[43]) );
  DFF \nreg_reg[42]  ( .D(nreg[42]), .CLK(clk), .RST(rst), .I(e_init[42]), .Q(
        nreg[42]) );
  DFF \nreg_reg[41]  ( .D(nreg[41]), .CLK(clk), .RST(rst), .I(e_init[41]), .Q(
        nreg[41]) );
  DFF \nreg_reg[40]  ( .D(nreg[40]), .CLK(clk), .RST(rst), .I(e_init[40]), .Q(
        nreg[40]) );
  DFF \nreg_reg[39]  ( .D(nreg[39]), .CLK(clk), .RST(rst), .I(e_init[39]), .Q(
        nreg[39]) );
  DFF \nreg_reg[38]  ( .D(nreg[38]), .CLK(clk), .RST(rst), .I(e_init[38]), .Q(
        nreg[38]) );
  DFF \nreg_reg[37]  ( .D(nreg[37]), .CLK(clk), .RST(rst), .I(e_init[37]), .Q(
        nreg[37]) );
  DFF \nreg_reg[36]  ( .D(nreg[36]), .CLK(clk), .RST(rst), .I(e_init[36]), .Q(
        nreg[36]) );
  DFF \nreg_reg[35]  ( .D(nreg[35]), .CLK(clk), .RST(rst), .I(e_init[35]), .Q(
        nreg[35]) );
  DFF \nreg_reg[34]  ( .D(nreg[34]), .CLK(clk), .RST(rst), .I(e_init[34]), .Q(
        nreg[34]) );
  DFF \nreg_reg[33]  ( .D(nreg[33]), .CLK(clk), .RST(rst), .I(e_init[33]), .Q(
        nreg[33]) );
  DFF \nreg_reg[32]  ( .D(nreg[32]), .CLK(clk), .RST(rst), .I(e_init[32]), .Q(
        nreg[32]) );
  DFF \nreg_reg[31]  ( .D(nreg[31]), .CLK(clk), .RST(rst), .I(e_init[31]), .Q(
        nreg[31]) );
  DFF \nreg_reg[30]  ( .D(nreg[30]), .CLK(clk), .RST(rst), .I(e_init[30]), .Q(
        nreg[30]) );
  DFF \nreg_reg[29]  ( .D(nreg[29]), .CLK(clk), .RST(rst), .I(e_init[29]), .Q(
        nreg[29]) );
  DFF \nreg_reg[28]  ( .D(nreg[28]), .CLK(clk), .RST(rst), .I(e_init[28]), .Q(
        nreg[28]) );
  DFF \nreg_reg[27]  ( .D(nreg[27]), .CLK(clk), .RST(rst), .I(e_init[27]), .Q(
        nreg[27]) );
  DFF \nreg_reg[26]  ( .D(nreg[26]), .CLK(clk), .RST(rst), .I(e_init[26]), .Q(
        nreg[26]) );
  DFF \nreg_reg[25]  ( .D(nreg[25]), .CLK(clk), .RST(rst), .I(e_init[25]), .Q(
        nreg[25]) );
  DFF \nreg_reg[24]  ( .D(nreg[24]), .CLK(clk), .RST(rst), .I(e_init[24]), .Q(
        nreg[24]) );
  DFF \nreg_reg[23]  ( .D(nreg[23]), .CLK(clk), .RST(rst), .I(e_init[23]), .Q(
        nreg[23]) );
  DFF \nreg_reg[22]  ( .D(nreg[22]), .CLK(clk), .RST(rst), .I(e_init[22]), .Q(
        nreg[22]) );
  DFF \nreg_reg[21]  ( .D(nreg[21]), .CLK(clk), .RST(rst), .I(e_init[21]), .Q(
        nreg[21]) );
  DFF \nreg_reg[20]  ( .D(nreg[20]), .CLK(clk), .RST(rst), .I(e_init[20]), .Q(
        nreg[20]) );
  DFF \nreg_reg[19]  ( .D(nreg[19]), .CLK(clk), .RST(rst), .I(e_init[19]), .Q(
        nreg[19]) );
  DFF \nreg_reg[18]  ( .D(nreg[18]), .CLK(clk), .RST(rst), .I(e_init[18]), .Q(
        nreg[18]) );
  DFF \nreg_reg[17]  ( .D(nreg[17]), .CLK(clk), .RST(rst), .I(e_init[17]), .Q(
        nreg[17]) );
  DFF \nreg_reg[16]  ( .D(nreg[16]), .CLK(clk), .RST(rst), .I(e_init[16]), .Q(
        nreg[16]) );
  DFF \nreg_reg[15]  ( .D(nreg[15]), .CLK(clk), .RST(rst), .I(e_init[15]), .Q(
        nreg[15]) );
  DFF \nreg_reg[14]  ( .D(nreg[14]), .CLK(clk), .RST(rst), .I(e_init[14]), .Q(
        nreg[14]) );
  DFF \nreg_reg[13]  ( .D(nreg[13]), .CLK(clk), .RST(rst), .I(e_init[13]), .Q(
        nreg[13]) );
  DFF \nreg_reg[12]  ( .D(nreg[12]), .CLK(clk), .RST(rst), .I(e_init[12]), .Q(
        nreg[12]) );
  DFF \nreg_reg[11]  ( .D(nreg[11]), .CLK(clk), .RST(rst), .I(e_init[11]), .Q(
        nreg[11]) );
  DFF \nreg_reg[10]  ( .D(nreg[10]), .CLK(clk), .RST(rst), .I(e_init[10]), .Q(
        nreg[10]) );
  DFF \nreg_reg[9]  ( .D(nreg[9]), .CLK(clk), .RST(rst), .I(e_init[9]), .Q(
        nreg[9]) );
  DFF \nreg_reg[8]  ( .D(nreg[8]), .CLK(clk), .RST(rst), .I(e_init[8]), .Q(
        nreg[8]) );
  DFF \nreg_reg[7]  ( .D(nreg[7]), .CLK(clk), .RST(rst), .I(e_init[7]), .Q(
        nreg[7]) );
  DFF \nreg_reg[6]  ( .D(nreg[6]), .CLK(clk), .RST(rst), .I(e_init[6]), .Q(
        nreg[6]) );
  DFF \nreg_reg[5]  ( .D(nreg[5]), .CLK(clk), .RST(rst), .I(e_init[5]), .Q(
        nreg[5]) );
  DFF \nreg_reg[4]  ( .D(nreg[4]), .CLK(clk), .RST(rst), .I(e_init[4]), .Q(
        nreg[4]) );
  DFF \nreg_reg[3]  ( .D(nreg[3]), .CLK(clk), .RST(rst), .I(e_init[3]), .Q(
        nreg[3]) );
  DFF \nreg_reg[2]  ( .D(nreg[2]), .CLK(clk), .RST(rst), .I(e_init[2]), .Q(
        nreg[2]) );
  DFF \nreg_reg[1]  ( .D(nreg[1]), .CLK(clk), .RST(rst), .I(e_init[1]), .Q(
        nreg[1]) );
  DFF \nreg_reg[0]  ( .D(nreg[0]), .CLK(clk), .RST(rst), .I(e_init[0]), .Q(
        nreg[0]) );
  DFF mul_pow_reg ( .D(n8), .CLK(clk), .RST(rst), .I(1'b0), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(ereg_next[0]), .CLK(clk), .RST(rst), .I(e_init[1024]), 
        .Q(ein[0]) );
  DFF \ereg_reg[1]  ( .D(ereg_next[1]), .CLK(clk), .RST(rst), .I(e_init[1025]), 
        .Q(ein[1]) );
  DFF \ereg_reg[2]  ( .D(ereg_next[2]), .CLK(clk), .RST(rst), .I(e_init[1026]), 
        .Q(ein[2]) );
  DFF \ereg_reg[3]  ( .D(ereg_next[3]), .CLK(clk), .RST(rst), .I(e_init[1027]), 
        .Q(ein[3]) );
  DFF \ereg_reg[4]  ( .D(ereg_next[4]), .CLK(clk), .RST(rst), .I(e_init[1028]), 
        .Q(ein[4]) );
  DFF \ereg_reg[5]  ( .D(ereg_next[5]), .CLK(clk), .RST(rst), .I(e_init[1029]), 
        .Q(ein[5]) );
  DFF \ereg_reg[6]  ( .D(ereg_next[6]), .CLK(clk), .RST(rst), .I(e_init[1030]), 
        .Q(ein[6]) );
  DFF \ereg_reg[7]  ( .D(ereg_next[7]), .CLK(clk), .RST(rst), .I(e_init[1031]), 
        .Q(ein[7]) );
  DFF \ereg_reg[8]  ( .D(ereg_next[8]), .CLK(clk), .RST(rst), .I(e_init[1032]), 
        .Q(ein[8]) );
  DFF \ereg_reg[9]  ( .D(ereg_next[9]), .CLK(clk), .RST(rst), .I(e_init[1033]), 
        .Q(ein[9]) );
  DFF \ereg_reg[10]  ( .D(ereg_next[10]), .CLK(clk), .RST(rst), .I(
        e_init[1034]), .Q(ein[10]) );
  DFF \ereg_reg[11]  ( .D(ereg_next[11]), .CLK(clk), .RST(rst), .I(
        e_init[1035]), .Q(ein[11]) );
  DFF \ereg_reg[12]  ( .D(ereg_next[12]), .CLK(clk), .RST(rst), .I(
        e_init[1036]), .Q(ein[12]) );
  DFF \ereg_reg[13]  ( .D(ereg_next[13]), .CLK(clk), .RST(rst), .I(
        e_init[1037]), .Q(ein[13]) );
  DFF \ereg_reg[14]  ( .D(ereg_next[14]), .CLK(clk), .RST(rst), .I(
        e_init[1038]), .Q(ein[14]) );
  DFF \ereg_reg[15]  ( .D(ereg_next[15]), .CLK(clk), .RST(rst), .I(
        e_init[1039]), .Q(ein[15]) );
  DFF \ereg_reg[16]  ( .D(ereg_next[16]), .CLK(clk), .RST(rst), .I(
        e_init[1040]), .Q(ein[16]) );
  DFF \ereg_reg[17]  ( .D(ereg_next[17]), .CLK(clk), .RST(rst), .I(
        e_init[1041]), .Q(ein[17]) );
  DFF \ereg_reg[18]  ( .D(ereg_next[18]), .CLK(clk), .RST(rst), .I(
        e_init[1042]), .Q(ein[18]) );
  DFF \ereg_reg[19]  ( .D(ereg_next[19]), .CLK(clk), .RST(rst), .I(
        e_init[1043]), .Q(ein[19]) );
  DFF \ereg_reg[20]  ( .D(ereg_next[20]), .CLK(clk), .RST(rst), .I(
        e_init[1044]), .Q(ein[20]) );
  DFF \ereg_reg[21]  ( .D(ereg_next[21]), .CLK(clk), .RST(rst), .I(
        e_init[1045]), .Q(ein[21]) );
  DFF \ereg_reg[22]  ( .D(ereg_next[22]), .CLK(clk), .RST(rst), .I(
        e_init[1046]), .Q(ein[22]) );
  DFF \ereg_reg[23]  ( .D(ereg_next[23]), .CLK(clk), .RST(rst), .I(
        e_init[1047]), .Q(ein[23]) );
  DFF \ereg_reg[24]  ( .D(ereg_next[24]), .CLK(clk), .RST(rst), .I(
        e_init[1048]), .Q(ein[24]) );
  DFF \ereg_reg[25]  ( .D(ereg_next[25]), .CLK(clk), .RST(rst), .I(
        e_init[1049]), .Q(ein[25]) );
  DFF \ereg_reg[26]  ( .D(ereg_next[26]), .CLK(clk), .RST(rst), .I(
        e_init[1050]), .Q(ein[26]) );
  DFF \ereg_reg[27]  ( .D(ereg_next[27]), .CLK(clk), .RST(rst), .I(
        e_init[1051]), .Q(ein[27]) );
  DFF \ereg_reg[28]  ( .D(ereg_next[28]), .CLK(clk), .RST(rst), .I(
        e_init[1052]), .Q(ein[28]) );
  DFF \ereg_reg[29]  ( .D(ereg_next[29]), .CLK(clk), .RST(rst), .I(
        e_init[1053]), .Q(ein[29]) );
  DFF \ereg_reg[30]  ( .D(ereg_next[30]), .CLK(clk), .RST(rst), .I(
        e_init[1054]), .Q(ein[30]) );
  DFF \ereg_reg[31]  ( .D(ereg_next[31]), .CLK(clk), .RST(rst), .I(
        e_init[1055]), .Q(ein[31]) );
  DFF \ereg_reg[32]  ( .D(ereg_next[32]), .CLK(clk), .RST(rst), .I(
        e_init[1056]), .Q(ein[32]) );
  DFF \ereg_reg[33]  ( .D(ereg_next[33]), .CLK(clk), .RST(rst), .I(
        e_init[1057]), .Q(ein[33]) );
  DFF \ereg_reg[34]  ( .D(ereg_next[34]), .CLK(clk), .RST(rst), .I(
        e_init[1058]), .Q(ein[34]) );
  DFF \ereg_reg[35]  ( .D(ereg_next[35]), .CLK(clk), .RST(rst), .I(
        e_init[1059]), .Q(ein[35]) );
  DFF \ereg_reg[36]  ( .D(ereg_next[36]), .CLK(clk), .RST(rst), .I(
        e_init[1060]), .Q(ein[36]) );
  DFF \ereg_reg[37]  ( .D(ereg_next[37]), .CLK(clk), .RST(rst), .I(
        e_init[1061]), .Q(ein[37]) );
  DFF \ereg_reg[38]  ( .D(ereg_next[38]), .CLK(clk), .RST(rst), .I(
        e_init[1062]), .Q(ein[38]) );
  DFF \ereg_reg[39]  ( .D(ereg_next[39]), .CLK(clk), .RST(rst), .I(
        e_init[1063]), .Q(ein[39]) );
  DFF \ereg_reg[40]  ( .D(ereg_next[40]), .CLK(clk), .RST(rst), .I(
        e_init[1064]), .Q(ein[40]) );
  DFF \ereg_reg[41]  ( .D(ereg_next[41]), .CLK(clk), .RST(rst), .I(
        e_init[1065]), .Q(ein[41]) );
  DFF \ereg_reg[42]  ( .D(ereg_next[42]), .CLK(clk), .RST(rst), .I(
        e_init[1066]), .Q(ein[42]) );
  DFF \ereg_reg[43]  ( .D(ereg_next[43]), .CLK(clk), .RST(rst), .I(
        e_init[1067]), .Q(ein[43]) );
  DFF \ereg_reg[44]  ( .D(ereg_next[44]), .CLK(clk), .RST(rst), .I(
        e_init[1068]), .Q(ein[44]) );
  DFF \ereg_reg[45]  ( .D(ereg_next[45]), .CLK(clk), .RST(rst), .I(
        e_init[1069]), .Q(ein[45]) );
  DFF \ereg_reg[46]  ( .D(ereg_next[46]), .CLK(clk), .RST(rst), .I(
        e_init[1070]), .Q(ein[46]) );
  DFF \ereg_reg[47]  ( .D(ereg_next[47]), .CLK(clk), .RST(rst), .I(
        e_init[1071]), .Q(ein[47]) );
  DFF \ereg_reg[48]  ( .D(ereg_next[48]), .CLK(clk), .RST(rst), .I(
        e_init[1072]), .Q(ein[48]) );
  DFF \ereg_reg[49]  ( .D(ereg_next[49]), .CLK(clk), .RST(rst), .I(
        e_init[1073]), .Q(ein[49]) );
  DFF \ereg_reg[50]  ( .D(ereg_next[50]), .CLK(clk), .RST(rst), .I(
        e_init[1074]), .Q(ein[50]) );
  DFF \ereg_reg[51]  ( .D(ereg_next[51]), .CLK(clk), .RST(rst), .I(
        e_init[1075]), .Q(ein[51]) );
  DFF \ereg_reg[52]  ( .D(ereg_next[52]), .CLK(clk), .RST(rst), .I(
        e_init[1076]), .Q(ein[52]) );
  DFF \ereg_reg[53]  ( .D(ereg_next[53]), .CLK(clk), .RST(rst), .I(
        e_init[1077]), .Q(ein[53]) );
  DFF \ereg_reg[54]  ( .D(ereg_next[54]), .CLK(clk), .RST(rst), .I(
        e_init[1078]), .Q(ein[54]) );
  DFF \ereg_reg[55]  ( .D(ereg_next[55]), .CLK(clk), .RST(rst), .I(
        e_init[1079]), .Q(ein[55]) );
  DFF \ereg_reg[56]  ( .D(ereg_next[56]), .CLK(clk), .RST(rst), .I(
        e_init[1080]), .Q(ein[56]) );
  DFF \ereg_reg[57]  ( .D(ereg_next[57]), .CLK(clk), .RST(rst), .I(
        e_init[1081]), .Q(ein[57]) );
  DFF \ereg_reg[58]  ( .D(ereg_next[58]), .CLK(clk), .RST(rst), .I(
        e_init[1082]), .Q(ein[58]) );
  DFF \ereg_reg[59]  ( .D(ereg_next[59]), .CLK(clk), .RST(rst), .I(
        e_init[1083]), .Q(ein[59]) );
  DFF \ereg_reg[60]  ( .D(ereg_next[60]), .CLK(clk), .RST(rst), .I(
        e_init[1084]), .Q(ein[60]) );
  DFF \ereg_reg[61]  ( .D(ereg_next[61]), .CLK(clk), .RST(rst), .I(
        e_init[1085]), .Q(ein[61]) );
  DFF \ereg_reg[62]  ( .D(ereg_next[62]), .CLK(clk), .RST(rst), .I(
        e_init[1086]), .Q(ein[62]) );
  DFF \ereg_reg[63]  ( .D(ereg_next[63]), .CLK(clk), .RST(rst), .I(
        e_init[1087]), .Q(ein[63]) );
  DFF \ereg_reg[64]  ( .D(ereg_next[64]), .CLK(clk), .RST(rst), .I(
        e_init[1088]), .Q(ein[64]) );
  DFF \ereg_reg[65]  ( .D(ereg_next[65]), .CLK(clk), .RST(rst), .I(
        e_init[1089]), .Q(ein[65]) );
  DFF \ereg_reg[66]  ( .D(ereg_next[66]), .CLK(clk), .RST(rst), .I(
        e_init[1090]), .Q(ein[66]) );
  DFF \ereg_reg[67]  ( .D(ereg_next[67]), .CLK(clk), .RST(rst), .I(
        e_init[1091]), .Q(ein[67]) );
  DFF \ereg_reg[68]  ( .D(ereg_next[68]), .CLK(clk), .RST(rst), .I(
        e_init[1092]), .Q(ein[68]) );
  DFF \ereg_reg[69]  ( .D(ereg_next[69]), .CLK(clk), .RST(rst), .I(
        e_init[1093]), .Q(ein[69]) );
  DFF \ereg_reg[70]  ( .D(ereg_next[70]), .CLK(clk), .RST(rst), .I(
        e_init[1094]), .Q(ein[70]) );
  DFF \ereg_reg[71]  ( .D(ereg_next[71]), .CLK(clk), .RST(rst), .I(
        e_init[1095]), .Q(ein[71]) );
  DFF \ereg_reg[72]  ( .D(ereg_next[72]), .CLK(clk), .RST(rst), .I(
        e_init[1096]), .Q(ein[72]) );
  DFF \ereg_reg[73]  ( .D(ereg_next[73]), .CLK(clk), .RST(rst), .I(
        e_init[1097]), .Q(ein[73]) );
  DFF \ereg_reg[74]  ( .D(ereg_next[74]), .CLK(clk), .RST(rst), .I(
        e_init[1098]), .Q(ein[74]) );
  DFF \ereg_reg[75]  ( .D(ereg_next[75]), .CLK(clk), .RST(rst), .I(
        e_init[1099]), .Q(ein[75]) );
  DFF \ereg_reg[76]  ( .D(ereg_next[76]), .CLK(clk), .RST(rst), .I(
        e_init[1100]), .Q(ein[76]) );
  DFF \ereg_reg[77]  ( .D(ereg_next[77]), .CLK(clk), .RST(rst), .I(
        e_init[1101]), .Q(ein[77]) );
  DFF \ereg_reg[78]  ( .D(ereg_next[78]), .CLK(clk), .RST(rst), .I(
        e_init[1102]), .Q(ein[78]) );
  DFF \ereg_reg[79]  ( .D(ereg_next[79]), .CLK(clk), .RST(rst), .I(
        e_init[1103]), .Q(ein[79]) );
  DFF \ereg_reg[80]  ( .D(ereg_next[80]), .CLK(clk), .RST(rst), .I(
        e_init[1104]), .Q(ein[80]) );
  DFF \ereg_reg[81]  ( .D(ereg_next[81]), .CLK(clk), .RST(rst), .I(
        e_init[1105]), .Q(ein[81]) );
  DFF \ereg_reg[82]  ( .D(ereg_next[82]), .CLK(clk), .RST(rst), .I(
        e_init[1106]), .Q(ein[82]) );
  DFF \ereg_reg[83]  ( .D(ereg_next[83]), .CLK(clk), .RST(rst), .I(
        e_init[1107]), .Q(ein[83]) );
  DFF \ereg_reg[84]  ( .D(ereg_next[84]), .CLK(clk), .RST(rst), .I(
        e_init[1108]), .Q(ein[84]) );
  DFF \ereg_reg[85]  ( .D(ereg_next[85]), .CLK(clk), .RST(rst), .I(
        e_init[1109]), .Q(ein[85]) );
  DFF \ereg_reg[86]  ( .D(ereg_next[86]), .CLK(clk), .RST(rst), .I(
        e_init[1110]), .Q(ein[86]) );
  DFF \ereg_reg[87]  ( .D(ereg_next[87]), .CLK(clk), .RST(rst), .I(
        e_init[1111]), .Q(ein[87]) );
  DFF \ereg_reg[88]  ( .D(ereg_next[88]), .CLK(clk), .RST(rst), .I(
        e_init[1112]), .Q(ein[88]) );
  DFF \ereg_reg[89]  ( .D(ereg_next[89]), .CLK(clk), .RST(rst), .I(
        e_init[1113]), .Q(ein[89]) );
  DFF \ereg_reg[90]  ( .D(ereg_next[90]), .CLK(clk), .RST(rst), .I(
        e_init[1114]), .Q(ein[90]) );
  DFF \ereg_reg[91]  ( .D(ereg_next[91]), .CLK(clk), .RST(rst), .I(
        e_init[1115]), .Q(ein[91]) );
  DFF \ereg_reg[92]  ( .D(ereg_next[92]), .CLK(clk), .RST(rst), .I(
        e_init[1116]), .Q(ein[92]) );
  DFF \ereg_reg[93]  ( .D(ereg_next[93]), .CLK(clk), .RST(rst), .I(
        e_init[1117]), .Q(ein[93]) );
  DFF \ereg_reg[94]  ( .D(ereg_next[94]), .CLK(clk), .RST(rst), .I(
        e_init[1118]), .Q(ein[94]) );
  DFF \ereg_reg[95]  ( .D(ereg_next[95]), .CLK(clk), .RST(rst), .I(
        e_init[1119]), .Q(ein[95]) );
  DFF \ereg_reg[96]  ( .D(ereg_next[96]), .CLK(clk), .RST(rst), .I(
        e_init[1120]), .Q(ein[96]) );
  DFF \ereg_reg[97]  ( .D(ereg_next[97]), .CLK(clk), .RST(rst), .I(
        e_init[1121]), .Q(ein[97]) );
  DFF \ereg_reg[98]  ( .D(ereg_next[98]), .CLK(clk), .RST(rst), .I(
        e_init[1122]), .Q(ein[98]) );
  DFF \ereg_reg[99]  ( .D(ereg_next[99]), .CLK(clk), .RST(rst), .I(
        e_init[1123]), .Q(ein[99]) );
  DFF \ereg_reg[100]  ( .D(ereg_next[100]), .CLK(clk), .RST(rst), .I(
        e_init[1124]), .Q(ein[100]) );
  DFF \ereg_reg[101]  ( .D(ereg_next[101]), .CLK(clk), .RST(rst), .I(
        e_init[1125]), .Q(ein[101]) );
  DFF \ereg_reg[102]  ( .D(ereg_next[102]), .CLK(clk), .RST(rst), .I(
        e_init[1126]), .Q(ein[102]) );
  DFF \ereg_reg[103]  ( .D(ereg_next[103]), .CLK(clk), .RST(rst), .I(
        e_init[1127]), .Q(ein[103]) );
  DFF \ereg_reg[104]  ( .D(ereg_next[104]), .CLK(clk), .RST(rst), .I(
        e_init[1128]), .Q(ein[104]) );
  DFF \ereg_reg[105]  ( .D(ereg_next[105]), .CLK(clk), .RST(rst), .I(
        e_init[1129]), .Q(ein[105]) );
  DFF \ereg_reg[106]  ( .D(ereg_next[106]), .CLK(clk), .RST(rst), .I(
        e_init[1130]), .Q(ein[106]) );
  DFF \ereg_reg[107]  ( .D(ereg_next[107]), .CLK(clk), .RST(rst), .I(
        e_init[1131]), .Q(ein[107]) );
  DFF \ereg_reg[108]  ( .D(ereg_next[108]), .CLK(clk), .RST(rst), .I(
        e_init[1132]), .Q(ein[108]) );
  DFF \ereg_reg[109]  ( .D(ereg_next[109]), .CLK(clk), .RST(rst), .I(
        e_init[1133]), .Q(ein[109]) );
  DFF \ereg_reg[110]  ( .D(ereg_next[110]), .CLK(clk), .RST(rst), .I(
        e_init[1134]), .Q(ein[110]) );
  DFF \ereg_reg[111]  ( .D(ereg_next[111]), .CLK(clk), .RST(rst), .I(
        e_init[1135]), .Q(ein[111]) );
  DFF \ereg_reg[112]  ( .D(ereg_next[112]), .CLK(clk), .RST(rst), .I(
        e_init[1136]), .Q(ein[112]) );
  DFF \ereg_reg[113]  ( .D(ereg_next[113]), .CLK(clk), .RST(rst), .I(
        e_init[1137]), .Q(ein[113]) );
  DFF \ereg_reg[114]  ( .D(ereg_next[114]), .CLK(clk), .RST(rst), .I(
        e_init[1138]), .Q(ein[114]) );
  DFF \ereg_reg[115]  ( .D(ereg_next[115]), .CLK(clk), .RST(rst), .I(
        e_init[1139]), .Q(ein[115]) );
  DFF \ereg_reg[116]  ( .D(ereg_next[116]), .CLK(clk), .RST(rst), .I(
        e_init[1140]), .Q(ein[116]) );
  DFF \ereg_reg[117]  ( .D(ereg_next[117]), .CLK(clk), .RST(rst), .I(
        e_init[1141]), .Q(ein[117]) );
  DFF \ereg_reg[118]  ( .D(ereg_next[118]), .CLK(clk), .RST(rst), .I(
        e_init[1142]), .Q(ein[118]) );
  DFF \ereg_reg[119]  ( .D(ereg_next[119]), .CLK(clk), .RST(rst), .I(
        e_init[1143]), .Q(ein[119]) );
  DFF \ereg_reg[120]  ( .D(ereg_next[120]), .CLK(clk), .RST(rst), .I(
        e_init[1144]), .Q(ein[120]) );
  DFF \ereg_reg[121]  ( .D(ereg_next[121]), .CLK(clk), .RST(rst), .I(
        e_init[1145]), .Q(ein[121]) );
  DFF \ereg_reg[122]  ( .D(ereg_next[122]), .CLK(clk), .RST(rst), .I(
        e_init[1146]), .Q(ein[122]) );
  DFF \ereg_reg[123]  ( .D(ereg_next[123]), .CLK(clk), .RST(rst), .I(
        e_init[1147]), .Q(ein[123]) );
  DFF \ereg_reg[124]  ( .D(ereg_next[124]), .CLK(clk), .RST(rst), .I(
        e_init[1148]), .Q(ein[124]) );
  DFF \ereg_reg[125]  ( .D(ereg_next[125]), .CLK(clk), .RST(rst), .I(
        e_init[1149]), .Q(ein[125]) );
  DFF \ereg_reg[126]  ( .D(ereg_next[126]), .CLK(clk), .RST(rst), .I(
        e_init[1150]), .Q(ein[126]) );
  DFF \ereg_reg[127]  ( .D(ereg_next[127]), .CLK(clk), .RST(rst), .I(
        e_init[1151]), .Q(ein[127]) );
  DFF \ereg_reg[128]  ( .D(ereg_next[128]), .CLK(clk), .RST(rst), .I(
        e_init[1152]), .Q(ein[128]) );
  DFF \ereg_reg[129]  ( .D(ereg_next[129]), .CLK(clk), .RST(rst), .I(
        e_init[1153]), .Q(ein[129]) );
  DFF \ereg_reg[130]  ( .D(ereg_next[130]), .CLK(clk), .RST(rst), .I(
        e_init[1154]), .Q(ein[130]) );
  DFF \ereg_reg[131]  ( .D(ereg_next[131]), .CLK(clk), .RST(rst), .I(
        e_init[1155]), .Q(ein[131]) );
  DFF \ereg_reg[132]  ( .D(ereg_next[132]), .CLK(clk), .RST(rst), .I(
        e_init[1156]), .Q(ein[132]) );
  DFF \ereg_reg[133]  ( .D(ereg_next[133]), .CLK(clk), .RST(rst), .I(
        e_init[1157]), .Q(ein[133]) );
  DFF \ereg_reg[134]  ( .D(ereg_next[134]), .CLK(clk), .RST(rst), .I(
        e_init[1158]), .Q(ein[134]) );
  DFF \ereg_reg[135]  ( .D(ereg_next[135]), .CLK(clk), .RST(rst), .I(
        e_init[1159]), .Q(ein[135]) );
  DFF \ereg_reg[136]  ( .D(ereg_next[136]), .CLK(clk), .RST(rst), .I(
        e_init[1160]), .Q(ein[136]) );
  DFF \ereg_reg[137]  ( .D(ereg_next[137]), .CLK(clk), .RST(rst), .I(
        e_init[1161]), .Q(ein[137]) );
  DFF \ereg_reg[138]  ( .D(ereg_next[138]), .CLK(clk), .RST(rst), .I(
        e_init[1162]), .Q(ein[138]) );
  DFF \ereg_reg[139]  ( .D(ereg_next[139]), .CLK(clk), .RST(rst), .I(
        e_init[1163]), .Q(ein[139]) );
  DFF \ereg_reg[140]  ( .D(ereg_next[140]), .CLK(clk), .RST(rst), .I(
        e_init[1164]), .Q(ein[140]) );
  DFF \ereg_reg[141]  ( .D(ereg_next[141]), .CLK(clk), .RST(rst), .I(
        e_init[1165]), .Q(ein[141]) );
  DFF \ereg_reg[142]  ( .D(ereg_next[142]), .CLK(clk), .RST(rst), .I(
        e_init[1166]), .Q(ein[142]) );
  DFF \ereg_reg[143]  ( .D(ereg_next[143]), .CLK(clk), .RST(rst), .I(
        e_init[1167]), .Q(ein[143]) );
  DFF \ereg_reg[144]  ( .D(ereg_next[144]), .CLK(clk), .RST(rst), .I(
        e_init[1168]), .Q(ein[144]) );
  DFF \ereg_reg[145]  ( .D(ereg_next[145]), .CLK(clk), .RST(rst), .I(
        e_init[1169]), .Q(ein[145]) );
  DFF \ereg_reg[146]  ( .D(ereg_next[146]), .CLK(clk), .RST(rst), .I(
        e_init[1170]), .Q(ein[146]) );
  DFF \ereg_reg[147]  ( .D(ereg_next[147]), .CLK(clk), .RST(rst), .I(
        e_init[1171]), .Q(ein[147]) );
  DFF \ereg_reg[148]  ( .D(ereg_next[148]), .CLK(clk), .RST(rst), .I(
        e_init[1172]), .Q(ein[148]) );
  DFF \ereg_reg[149]  ( .D(ereg_next[149]), .CLK(clk), .RST(rst), .I(
        e_init[1173]), .Q(ein[149]) );
  DFF \ereg_reg[150]  ( .D(ereg_next[150]), .CLK(clk), .RST(rst), .I(
        e_init[1174]), .Q(ein[150]) );
  DFF \ereg_reg[151]  ( .D(ereg_next[151]), .CLK(clk), .RST(rst), .I(
        e_init[1175]), .Q(ein[151]) );
  DFF \ereg_reg[152]  ( .D(ereg_next[152]), .CLK(clk), .RST(rst), .I(
        e_init[1176]), .Q(ein[152]) );
  DFF \ereg_reg[153]  ( .D(ereg_next[153]), .CLK(clk), .RST(rst), .I(
        e_init[1177]), .Q(ein[153]) );
  DFF \ereg_reg[154]  ( .D(ereg_next[154]), .CLK(clk), .RST(rst), .I(
        e_init[1178]), .Q(ein[154]) );
  DFF \ereg_reg[155]  ( .D(ereg_next[155]), .CLK(clk), .RST(rst), .I(
        e_init[1179]), .Q(ein[155]) );
  DFF \ereg_reg[156]  ( .D(ereg_next[156]), .CLK(clk), .RST(rst), .I(
        e_init[1180]), .Q(ein[156]) );
  DFF \ereg_reg[157]  ( .D(ereg_next[157]), .CLK(clk), .RST(rst), .I(
        e_init[1181]), .Q(ein[157]) );
  DFF \ereg_reg[158]  ( .D(ereg_next[158]), .CLK(clk), .RST(rst), .I(
        e_init[1182]), .Q(ein[158]) );
  DFF \ereg_reg[159]  ( .D(ereg_next[159]), .CLK(clk), .RST(rst), .I(
        e_init[1183]), .Q(ein[159]) );
  DFF \ereg_reg[160]  ( .D(ereg_next[160]), .CLK(clk), .RST(rst), .I(
        e_init[1184]), .Q(ein[160]) );
  DFF \ereg_reg[161]  ( .D(ereg_next[161]), .CLK(clk), .RST(rst), .I(
        e_init[1185]), .Q(ein[161]) );
  DFF \ereg_reg[162]  ( .D(ereg_next[162]), .CLK(clk), .RST(rst), .I(
        e_init[1186]), .Q(ein[162]) );
  DFF \ereg_reg[163]  ( .D(ereg_next[163]), .CLK(clk), .RST(rst), .I(
        e_init[1187]), .Q(ein[163]) );
  DFF \ereg_reg[164]  ( .D(ereg_next[164]), .CLK(clk), .RST(rst), .I(
        e_init[1188]), .Q(ein[164]) );
  DFF \ereg_reg[165]  ( .D(ereg_next[165]), .CLK(clk), .RST(rst), .I(
        e_init[1189]), .Q(ein[165]) );
  DFF \ereg_reg[166]  ( .D(ereg_next[166]), .CLK(clk), .RST(rst), .I(
        e_init[1190]), .Q(ein[166]) );
  DFF \ereg_reg[167]  ( .D(ereg_next[167]), .CLK(clk), .RST(rst), .I(
        e_init[1191]), .Q(ein[167]) );
  DFF \ereg_reg[168]  ( .D(ereg_next[168]), .CLK(clk), .RST(rst), .I(
        e_init[1192]), .Q(ein[168]) );
  DFF \ereg_reg[169]  ( .D(ereg_next[169]), .CLK(clk), .RST(rst), .I(
        e_init[1193]), .Q(ein[169]) );
  DFF \ereg_reg[170]  ( .D(ereg_next[170]), .CLK(clk), .RST(rst), .I(
        e_init[1194]), .Q(ein[170]) );
  DFF \ereg_reg[171]  ( .D(ereg_next[171]), .CLK(clk), .RST(rst), .I(
        e_init[1195]), .Q(ein[171]) );
  DFF \ereg_reg[172]  ( .D(ereg_next[172]), .CLK(clk), .RST(rst), .I(
        e_init[1196]), .Q(ein[172]) );
  DFF \ereg_reg[173]  ( .D(ereg_next[173]), .CLK(clk), .RST(rst), .I(
        e_init[1197]), .Q(ein[173]) );
  DFF \ereg_reg[174]  ( .D(ereg_next[174]), .CLK(clk), .RST(rst), .I(
        e_init[1198]), .Q(ein[174]) );
  DFF \ereg_reg[175]  ( .D(ereg_next[175]), .CLK(clk), .RST(rst), .I(
        e_init[1199]), .Q(ein[175]) );
  DFF \ereg_reg[176]  ( .D(ereg_next[176]), .CLK(clk), .RST(rst), .I(
        e_init[1200]), .Q(ein[176]) );
  DFF \ereg_reg[177]  ( .D(ereg_next[177]), .CLK(clk), .RST(rst), .I(
        e_init[1201]), .Q(ein[177]) );
  DFF \ereg_reg[178]  ( .D(ereg_next[178]), .CLK(clk), .RST(rst), .I(
        e_init[1202]), .Q(ein[178]) );
  DFF \ereg_reg[179]  ( .D(ereg_next[179]), .CLK(clk), .RST(rst), .I(
        e_init[1203]), .Q(ein[179]) );
  DFF \ereg_reg[180]  ( .D(ereg_next[180]), .CLK(clk), .RST(rst), .I(
        e_init[1204]), .Q(ein[180]) );
  DFF \ereg_reg[181]  ( .D(ereg_next[181]), .CLK(clk), .RST(rst), .I(
        e_init[1205]), .Q(ein[181]) );
  DFF \ereg_reg[182]  ( .D(ereg_next[182]), .CLK(clk), .RST(rst), .I(
        e_init[1206]), .Q(ein[182]) );
  DFF \ereg_reg[183]  ( .D(ereg_next[183]), .CLK(clk), .RST(rst), .I(
        e_init[1207]), .Q(ein[183]) );
  DFF \ereg_reg[184]  ( .D(ereg_next[184]), .CLK(clk), .RST(rst), .I(
        e_init[1208]), .Q(ein[184]) );
  DFF \ereg_reg[185]  ( .D(ereg_next[185]), .CLK(clk), .RST(rst), .I(
        e_init[1209]), .Q(ein[185]) );
  DFF \ereg_reg[186]  ( .D(ereg_next[186]), .CLK(clk), .RST(rst), .I(
        e_init[1210]), .Q(ein[186]) );
  DFF \ereg_reg[187]  ( .D(ereg_next[187]), .CLK(clk), .RST(rst), .I(
        e_init[1211]), .Q(ein[187]) );
  DFF \ereg_reg[188]  ( .D(ereg_next[188]), .CLK(clk), .RST(rst), .I(
        e_init[1212]), .Q(ein[188]) );
  DFF \ereg_reg[189]  ( .D(ereg_next[189]), .CLK(clk), .RST(rst), .I(
        e_init[1213]), .Q(ein[189]) );
  DFF \ereg_reg[190]  ( .D(ereg_next[190]), .CLK(clk), .RST(rst), .I(
        e_init[1214]), .Q(ein[190]) );
  DFF \ereg_reg[191]  ( .D(ereg_next[191]), .CLK(clk), .RST(rst), .I(
        e_init[1215]), .Q(ein[191]) );
  DFF \ereg_reg[192]  ( .D(ereg_next[192]), .CLK(clk), .RST(rst), .I(
        e_init[1216]), .Q(ein[192]) );
  DFF \ereg_reg[193]  ( .D(ereg_next[193]), .CLK(clk), .RST(rst), .I(
        e_init[1217]), .Q(ein[193]) );
  DFF \ereg_reg[194]  ( .D(ereg_next[194]), .CLK(clk), .RST(rst), .I(
        e_init[1218]), .Q(ein[194]) );
  DFF \ereg_reg[195]  ( .D(ereg_next[195]), .CLK(clk), .RST(rst), .I(
        e_init[1219]), .Q(ein[195]) );
  DFF \ereg_reg[196]  ( .D(ereg_next[196]), .CLK(clk), .RST(rst), .I(
        e_init[1220]), .Q(ein[196]) );
  DFF \ereg_reg[197]  ( .D(ereg_next[197]), .CLK(clk), .RST(rst), .I(
        e_init[1221]), .Q(ein[197]) );
  DFF \ereg_reg[198]  ( .D(ereg_next[198]), .CLK(clk), .RST(rst), .I(
        e_init[1222]), .Q(ein[198]) );
  DFF \ereg_reg[199]  ( .D(ereg_next[199]), .CLK(clk), .RST(rst), .I(
        e_init[1223]), .Q(ein[199]) );
  DFF \ereg_reg[200]  ( .D(ereg_next[200]), .CLK(clk), .RST(rst), .I(
        e_init[1224]), .Q(ein[200]) );
  DFF \ereg_reg[201]  ( .D(ereg_next[201]), .CLK(clk), .RST(rst), .I(
        e_init[1225]), .Q(ein[201]) );
  DFF \ereg_reg[202]  ( .D(ereg_next[202]), .CLK(clk), .RST(rst), .I(
        e_init[1226]), .Q(ein[202]) );
  DFF \ereg_reg[203]  ( .D(ereg_next[203]), .CLK(clk), .RST(rst), .I(
        e_init[1227]), .Q(ein[203]) );
  DFF \ereg_reg[204]  ( .D(ereg_next[204]), .CLK(clk), .RST(rst), .I(
        e_init[1228]), .Q(ein[204]) );
  DFF \ereg_reg[205]  ( .D(ereg_next[205]), .CLK(clk), .RST(rst), .I(
        e_init[1229]), .Q(ein[205]) );
  DFF \ereg_reg[206]  ( .D(ereg_next[206]), .CLK(clk), .RST(rst), .I(
        e_init[1230]), .Q(ein[206]) );
  DFF \ereg_reg[207]  ( .D(ereg_next[207]), .CLK(clk), .RST(rst), .I(
        e_init[1231]), .Q(ein[207]) );
  DFF \ereg_reg[208]  ( .D(ereg_next[208]), .CLK(clk), .RST(rst), .I(
        e_init[1232]), .Q(ein[208]) );
  DFF \ereg_reg[209]  ( .D(ereg_next[209]), .CLK(clk), .RST(rst), .I(
        e_init[1233]), .Q(ein[209]) );
  DFF \ereg_reg[210]  ( .D(ereg_next[210]), .CLK(clk), .RST(rst), .I(
        e_init[1234]), .Q(ein[210]) );
  DFF \ereg_reg[211]  ( .D(ereg_next[211]), .CLK(clk), .RST(rst), .I(
        e_init[1235]), .Q(ein[211]) );
  DFF \ereg_reg[212]  ( .D(ereg_next[212]), .CLK(clk), .RST(rst), .I(
        e_init[1236]), .Q(ein[212]) );
  DFF \ereg_reg[213]  ( .D(ereg_next[213]), .CLK(clk), .RST(rst), .I(
        e_init[1237]), .Q(ein[213]) );
  DFF \ereg_reg[214]  ( .D(ereg_next[214]), .CLK(clk), .RST(rst), .I(
        e_init[1238]), .Q(ein[214]) );
  DFF \ereg_reg[215]  ( .D(ereg_next[215]), .CLK(clk), .RST(rst), .I(
        e_init[1239]), .Q(ein[215]) );
  DFF \ereg_reg[216]  ( .D(ereg_next[216]), .CLK(clk), .RST(rst), .I(
        e_init[1240]), .Q(ein[216]) );
  DFF \ereg_reg[217]  ( .D(ereg_next[217]), .CLK(clk), .RST(rst), .I(
        e_init[1241]), .Q(ein[217]) );
  DFF \ereg_reg[218]  ( .D(ereg_next[218]), .CLK(clk), .RST(rst), .I(
        e_init[1242]), .Q(ein[218]) );
  DFF \ereg_reg[219]  ( .D(ereg_next[219]), .CLK(clk), .RST(rst), .I(
        e_init[1243]), .Q(ein[219]) );
  DFF \ereg_reg[220]  ( .D(ereg_next[220]), .CLK(clk), .RST(rst), .I(
        e_init[1244]), .Q(ein[220]) );
  DFF \ereg_reg[221]  ( .D(ereg_next[221]), .CLK(clk), .RST(rst), .I(
        e_init[1245]), .Q(ein[221]) );
  DFF \ereg_reg[222]  ( .D(ereg_next[222]), .CLK(clk), .RST(rst), .I(
        e_init[1246]), .Q(ein[222]) );
  DFF \ereg_reg[223]  ( .D(ereg_next[223]), .CLK(clk), .RST(rst), .I(
        e_init[1247]), .Q(ein[223]) );
  DFF \ereg_reg[224]  ( .D(ereg_next[224]), .CLK(clk), .RST(rst), .I(
        e_init[1248]), .Q(ein[224]) );
  DFF \ereg_reg[225]  ( .D(ereg_next[225]), .CLK(clk), .RST(rst), .I(
        e_init[1249]), .Q(ein[225]) );
  DFF \ereg_reg[226]  ( .D(ereg_next[226]), .CLK(clk), .RST(rst), .I(
        e_init[1250]), .Q(ein[226]) );
  DFF \ereg_reg[227]  ( .D(ereg_next[227]), .CLK(clk), .RST(rst), .I(
        e_init[1251]), .Q(ein[227]) );
  DFF \ereg_reg[228]  ( .D(ereg_next[228]), .CLK(clk), .RST(rst), .I(
        e_init[1252]), .Q(ein[228]) );
  DFF \ereg_reg[229]  ( .D(ereg_next[229]), .CLK(clk), .RST(rst), .I(
        e_init[1253]), .Q(ein[229]) );
  DFF \ereg_reg[230]  ( .D(ereg_next[230]), .CLK(clk), .RST(rst), .I(
        e_init[1254]), .Q(ein[230]) );
  DFF \ereg_reg[231]  ( .D(ereg_next[231]), .CLK(clk), .RST(rst), .I(
        e_init[1255]), .Q(ein[231]) );
  DFF \ereg_reg[232]  ( .D(ereg_next[232]), .CLK(clk), .RST(rst), .I(
        e_init[1256]), .Q(ein[232]) );
  DFF \ereg_reg[233]  ( .D(ereg_next[233]), .CLK(clk), .RST(rst), .I(
        e_init[1257]), .Q(ein[233]) );
  DFF \ereg_reg[234]  ( .D(ereg_next[234]), .CLK(clk), .RST(rst), .I(
        e_init[1258]), .Q(ein[234]) );
  DFF \ereg_reg[235]  ( .D(ereg_next[235]), .CLK(clk), .RST(rst), .I(
        e_init[1259]), .Q(ein[235]) );
  DFF \ereg_reg[236]  ( .D(ereg_next[236]), .CLK(clk), .RST(rst), .I(
        e_init[1260]), .Q(ein[236]) );
  DFF \ereg_reg[237]  ( .D(ereg_next[237]), .CLK(clk), .RST(rst), .I(
        e_init[1261]), .Q(ein[237]) );
  DFF \ereg_reg[238]  ( .D(ereg_next[238]), .CLK(clk), .RST(rst), .I(
        e_init[1262]), .Q(ein[238]) );
  DFF \ereg_reg[239]  ( .D(ereg_next[239]), .CLK(clk), .RST(rst), .I(
        e_init[1263]), .Q(ein[239]) );
  DFF \ereg_reg[240]  ( .D(ereg_next[240]), .CLK(clk), .RST(rst), .I(
        e_init[1264]), .Q(ein[240]) );
  DFF \ereg_reg[241]  ( .D(ereg_next[241]), .CLK(clk), .RST(rst), .I(
        e_init[1265]), .Q(ein[241]) );
  DFF \ereg_reg[242]  ( .D(ereg_next[242]), .CLK(clk), .RST(rst), .I(
        e_init[1266]), .Q(ein[242]) );
  DFF \ereg_reg[243]  ( .D(ereg_next[243]), .CLK(clk), .RST(rst), .I(
        e_init[1267]), .Q(ein[243]) );
  DFF \ereg_reg[244]  ( .D(ereg_next[244]), .CLK(clk), .RST(rst), .I(
        e_init[1268]), .Q(ein[244]) );
  DFF \ereg_reg[245]  ( .D(ereg_next[245]), .CLK(clk), .RST(rst), .I(
        e_init[1269]), .Q(ein[245]) );
  DFF \ereg_reg[246]  ( .D(ereg_next[246]), .CLK(clk), .RST(rst), .I(
        e_init[1270]), .Q(ein[246]) );
  DFF \ereg_reg[247]  ( .D(ereg_next[247]), .CLK(clk), .RST(rst), .I(
        e_init[1271]), .Q(ein[247]) );
  DFF \ereg_reg[248]  ( .D(ereg_next[248]), .CLK(clk), .RST(rst), .I(
        e_init[1272]), .Q(ein[248]) );
  DFF \ereg_reg[249]  ( .D(ereg_next[249]), .CLK(clk), .RST(rst), .I(
        e_init[1273]), .Q(ein[249]) );
  DFF \ereg_reg[250]  ( .D(ereg_next[250]), .CLK(clk), .RST(rst), .I(
        e_init[1274]), .Q(ein[250]) );
  DFF \ereg_reg[251]  ( .D(ereg_next[251]), .CLK(clk), .RST(rst), .I(
        e_init[1275]), .Q(ein[251]) );
  DFF \ereg_reg[252]  ( .D(ereg_next[252]), .CLK(clk), .RST(rst), .I(
        e_init[1276]), .Q(ein[252]) );
  DFF \ereg_reg[253]  ( .D(ereg_next[253]), .CLK(clk), .RST(rst), .I(
        e_init[1277]), .Q(ein[253]) );
  DFF \ereg_reg[254]  ( .D(ereg_next[254]), .CLK(clk), .RST(rst), .I(
        e_init[1278]), .Q(ein[254]) );
  DFF \ereg_reg[255]  ( .D(ereg_next[255]), .CLK(clk), .RST(rst), .I(
        e_init[1279]), .Q(ein[255]) );
  DFF \ereg_reg[256]  ( .D(ereg_next[256]), .CLK(clk), .RST(rst), .I(
        e_init[1280]), .Q(ein[256]) );
  DFF \ereg_reg[257]  ( .D(ereg_next[257]), .CLK(clk), .RST(rst), .I(
        e_init[1281]), .Q(ein[257]) );
  DFF \ereg_reg[258]  ( .D(ereg_next[258]), .CLK(clk), .RST(rst), .I(
        e_init[1282]), .Q(ein[258]) );
  DFF \ereg_reg[259]  ( .D(ereg_next[259]), .CLK(clk), .RST(rst), .I(
        e_init[1283]), .Q(ein[259]) );
  DFF \ereg_reg[260]  ( .D(ereg_next[260]), .CLK(clk), .RST(rst), .I(
        e_init[1284]), .Q(ein[260]) );
  DFF \ereg_reg[261]  ( .D(ereg_next[261]), .CLK(clk), .RST(rst), .I(
        e_init[1285]), .Q(ein[261]) );
  DFF \ereg_reg[262]  ( .D(ereg_next[262]), .CLK(clk), .RST(rst), .I(
        e_init[1286]), .Q(ein[262]) );
  DFF \ereg_reg[263]  ( .D(ereg_next[263]), .CLK(clk), .RST(rst), .I(
        e_init[1287]), .Q(ein[263]) );
  DFF \ereg_reg[264]  ( .D(ereg_next[264]), .CLK(clk), .RST(rst), .I(
        e_init[1288]), .Q(ein[264]) );
  DFF \ereg_reg[265]  ( .D(ereg_next[265]), .CLK(clk), .RST(rst), .I(
        e_init[1289]), .Q(ein[265]) );
  DFF \ereg_reg[266]  ( .D(ereg_next[266]), .CLK(clk), .RST(rst), .I(
        e_init[1290]), .Q(ein[266]) );
  DFF \ereg_reg[267]  ( .D(ereg_next[267]), .CLK(clk), .RST(rst), .I(
        e_init[1291]), .Q(ein[267]) );
  DFF \ereg_reg[268]  ( .D(ereg_next[268]), .CLK(clk), .RST(rst), .I(
        e_init[1292]), .Q(ein[268]) );
  DFF \ereg_reg[269]  ( .D(ereg_next[269]), .CLK(clk), .RST(rst), .I(
        e_init[1293]), .Q(ein[269]) );
  DFF \ereg_reg[270]  ( .D(ereg_next[270]), .CLK(clk), .RST(rst), .I(
        e_init[1294]), .Q(ein[270]) );
  DFF \ereg_reg[271]  ( .D(ereg_next[271]), .CLK(clk), .RST(rst), .I(
        e_init[1295]), .Q(ein[271]) );
  DFF \ereg_reg[272]  ( .D(ereg_next[272]), .CLK(clk), .RST(rst), .I(
        e_init[1296]), .Q(ein[272]) );
  DFF \ereg_reg[273]  ( .D(ereg_next[273]), .CLK(clk), .RST(rst), .I(
        e_init[1297]), .Q(ein[273]) );
  DFF \ereg_reg[274]  ( .D(ereg_next[274]), .CLK(clk), .RST(rst), .I(
        e_init[1298]), .Q(ein[274]) );
  DFF \ereg_reg[275]  ( .D(ereg_next[275]), .CLK(clk), .RST(rst), .I(
        e_init[1299]), .Q(ein[275]) );
  DFF \ereg_reg[276]  ( .D(ereg_next[276]), .CLK(clk), .RST(rst), .I(
        e_init[1300]), .Q(ein[276]) );
  DFF \ereg_reg[277]  ( .D(ereg_next[277]), .CLK(clk), .RST(rst), .I(
        e_init[1301]), .Q(ein[277]) );
  DFF \ereg_reg[278]  ( .D(ereg_next[278]), .CLK(clk), .RST(rst), .I(
        e_init[1302]), .Q(ein[278]) );
  DFF \ereg_reg[279]  ( .D(ereg_next[279]), .CLK(clk), .RST(rst), .I(
        e_init[1303]), .Q(ein[279]) );
  DFF \ereg_reg[280]  ( .D(ereg_next[280]), .CLK(clk), .RST(rst), .I(
        e_init[1304]), .Q(ein[280]) );
  DFF \ereg_reg[281]  ( .D(ereg_next[281]), .CLK(clk), .RST(rst), .I(
        e_init[1305]), .Q(ein[281]) );
  DFF \ereg_reg[282]  ( .D(ereg_next[282]), .CLK(clk), .RST(rst), .I(
        e_init[1306]), .Q(ein[282]) );
  DFF \ereg_reg[283]  ( .D(ereg_next[283]), .CLK(clk), .RST(rst), .I(
        e_init[1307]), .Q(ein[283]) );
  DFF \ereg_reg[284]  ( .D(ereg_next[284]), .CLK(clk), .RST(rst), .I(
        e_init[1308]), .Q(ein[284]) );
  DFF \ereg_reg[285]  ( .D(ereg_next[285]), .CLK(clk), .RST(rst), .I(
        e_init[1309]), .Q(ein[285]) );
  DFF \ereg_reg[286]  ( .D(ereg_next[286]), .CLK(clk), .RST(rst), .I(
        e_init[1310]), .Q(ein[286]) );
  DFF \ereg_reg[287]  ( .D(ereg_next[287]), .CLK(clk), .RST(rst), .I(
        e_init[1311]), .Q(ein[287]) );
  DFF \ereg_reg[288]  ( .D(ereg_next[288]), .CLK(clk), .RST(rst), .I(
        e_init[1312]), .Q(ein[288]) );
  DFF \ereg_reg[289]  ( .D(ereg_next[289]), .CLK(clk), .RST(rst), .I(
        e_init[1313]), .Q(ein[289]) );
  DFF \ereg_reg[290]  ( .D(ereg_next[290]), .CLK(clk), .RST(rst), .I(
        e_init[1314]), .Q(ein[290]) );
  DFF \ereg_reg[291]  ( .D(ereg_next[291]), .CLK(clk), .RST(rst), .I(
        e_init[1315]), .Q(ein[291]) );
  DFF \ereg_reg[292]  ( .D(ereg_next[292]), .CLK(clk), .RST(rst), .I(
        e_init[1316]), .Q(ein[292]) );
  DFF \ereg_reg[293]  ( .D(ereg_next[293]), .CLK(clk), .RST(rst), .I(
        e_init[1317]), .Q(ein[293]) );
  DFF \ereg_reg[294]  ( .D(ereg_next[294]), .CLK(clk), .RST(rst), .I(
        e_init[1318]), .Q(ein[294]) );
  DFF \ereg_reg[295]  ( .D(ereg_next[295]), .CLK(clk), .RST(rst), .I(
        e_init[1319]), .Q(ein[295]) );
  DFF \ereg_reg[296]  ( .D(ereg_next[296]), .CLK(clk), .RST(rst), .I(
        e_init[1320]), .Q(ein[296]) );
  DFF \ereg_reg[297]  ( .D(ereg_next[297]), .CLK(clk), .RST(rst), .I(
        e_init[1321]), .Q(ein[297]) );
  DFF \ereg_reg[298]  ( .D(ereg_next[298]), .CLK(clk), .RST(rst), .I(
        e_init[1322]), .Q(ein[298]) );
  DFF \ereg_reg[299]  ( .D(ereg_next[299]), .CLK(clk), .RST(rst), .I(
        e_init[1323]), .Q(ein[299]) );
  DFF \ereg_reg[300]  ( .D(ereg_next[300]), .CLK(clk), .RST(rst), .I(
        e_init[1324]), .Q(ein[300]) );
  DFF \ereg_reg[301]  ( .D(ereg_next[301]), .CLK(clk), .RST(rst), .I(
        e_init[1325]), .Q(ein[301]) );
  DFF \ereg_reg[302]  ( .D(ereg_next[302]), .CLK(clk), .RST(rst), .I(
        e_init[1326]), .Q(ein[302]) );
  DFF \ereg_reg[303]  ( .D(ereg_next[303]), .CLK(clk), .RST(rst), .I(
        e_init[1327]), .Q(ein[303]) );
  DFF \ereg_reg[304]  ( .D(ereg_next[304]), .CLK(clk), .RST(rst), .I(
        e_init[1328]), .Q(ein[304]) );
  DFF \ereg_reg[305]  ( .D(ereg_next[305]), .CLK(clk), .RST(rst), .I(
        e_init[1329]), .Q(ein[305]) );
  DFF \ereg_reg[306]  ( .D(ereg_next[306]), .CLK(clk), .RST(rst), .I(
        e_init[1330]), .Q(ein[306]) );
  DFF \ereg_reg[307]  ( .D(ereg_next[307]), .CLK(clk), .RST(rst), .I(
        e_init[1331]), .Q(ein[307]) );
  DFF \ereg_reg[308]  ( .D(ereg_next[308]), .CLK(clk), .RST(rst), .I(
        e_init[1332]), .Q(ein[308]) );
  DFF \ereg_reg[309]  ( .D(ereg_next[309]), .CLK(clk), .RST(rst), .I(
        e_init[1333]), .Q(ein[309]) );
  DFF \ereg_reg[310]  ( .D(ereg_next[310]), .CLK(clk), .RST(rst), .I(
        e_init[1334]), .Q(ein[310]) );
  DFF \ereg_reg[311]  ( .D(ereg_next[311]), .CLK(clk), .RST(rst), .I(
        e_init[1335]), .Q(ein[311]) );
  DFF \ereg_reg[312]  ( .D(ereg_next[312]), .CLK(clk), .RST(rst), .I(
        e_init[1336]), .Q(ein[312]) );
  DFF \ereg_reg[313]  ( .D(ereg_next[313]), .CLK(clk), .RST(rst), .I(
        e_init[1337]), .Q(ein[313]) );
  DFF \ereg_reg[314]  ( .D(ereg_next[314]), .CLK(clk), .RST(rst), .I(
        e_init[1338]), .Q(ein[314]) );
  DFF \ereg_reg[315]  ( .D(ereg_next[315]), .CLK(clk), .RST(rst), .I(
        e_init[1339]), .Q(ein[315]) );
  DFF \ereg_reg[316]  ( .D(ereg_next[316]), .CLK(clk), .RST(rst), .I(
        e_init[1340]), .Q(ein[316]) );
  DFF \ereg_reg[317]  ( .D(ereg_next[317]), .CLK(clk), .RST(rst), .I(
        e_init[1341]), .Q(ein[317]) );
  DFF \ereg_reg[318]  ( .D(ereg_next[318]), .CLK(clk), .RST(rst), .I(
        e_init[1342]), .Q(ein[318]) );
  DFF \ereg_reg[319]  ( .D(ereg_next[319]), .CLK(clk), .RST(rst), .I(
        e_init[1343]), .Q(ein[319]) );
  DFF \ereg_reg[320]  ( .D(ereg_next[320]), .CLK(clk), .RST(rst), .I(
        e_init[1344]), .Q(ein[320]) );
  DFF \ereg_reg[321]  ( .D(ereg_next[321]), .CLK(clk), .RST(rst), .I(
        e_init[1345]), .Q(ein[321]) );
  DFF \ereg_reg[322]  ( .D(ereg_next[322]), .CLK(clk), .RST(rst), .I(
        e_init[1346]), .Q(ein[322]) );
  DFF \ereg_reg[323]  ( .D(ereg_next[323]), .CLK(clk), .RST(rst), .I(
        e_init[1347]), .Q(ein[323]) );
  DFF \ereg_reg[324]  ( .D(ereg_next[324]), .CLK(clk), .RST(rst), .I(
        e_init[1348]), .Q(ein[324]) );
  DFF \ereg_reg[325]  ( .D(ereg_next[325]), .CLK(clk), .RST(rst), .I(
        e_init[1349]), .Q(ein[325]) );
  DFF \ereg_reg[326]  ( .D(ereg_next[326]), .CLK(clk), .RST(rst), .I(
        e_init[1350]), .Q(ein[326]) );
  DFF \ereg_reg[327]  ( .D(ereg_next[327]), .CLK(clk), .RST(rst), .I(
        e_init[1351]), .Q(ein[327]) );
  DFF \ereg_reg[328]  ( .D(ereg_next[328]), .CLK(clk), .RST(rst), .I(
        e_init[1352]), .Q(ein[328]) );
  DFF \ereg_reg[329]  ( .D(ereg_next[329]), .CLK(clk), .RST(rst), .I(
        e_init[1353]), .Q(ein[329]) );
  DFF \ereg_reg[330]  ( .D(ereg_next[330]), .CLK(clk), .RST(rst), .I(
        e_init[1354]), .Q(ein[330]) );
  DFF \ereg_reg[331]  ( .D(ereg_next[331]), .CLK(clk), .RST(rst), .I(
        e_init[1355]), .Q(ein[331]) );
  DFF \ereg_reg[332]  ( .D(ereg_next[332]), .CLK(clk), .RST(rst), .I(
        e_init[1356]), .Q(ein[332]) );
  DFF \ereg_reg[333]  ( .D(ereg_next[333]), .CLK(clk), .RST(rst), .I(
        e_init[1357]), .Q(ein[333]) );
  DFF \ereg_reg[334]  ( .D(ereg_next[334]), .CLK(clk), .RST(rst), .I(
        e_init[1358]), .Q(ein[334]) );
  DFF \ereg_reg[335]  ( .D(ereg_next[335]), .CLK(clk), .RST(rst), .I(
        e_init[1359]), .Q(ein[335]) );
  DFF \ereg_reg[336]  ( .D(ereg_next[336]), .CLK(clk), .RST(rst), .I(
        e_init[1360]), .Q(ein[336]) );
  DFF \ereg_reg[337]  ( .D(ereg_next[337]), .CLK(clk), .RST(rst), .I(
        e_init[1361]), .Q(ein[337]) );
  DFF \ereg_reg[338]  ( .D(ereg_next[338]), .CLK(clk), .RST(rst), .I(
        e_init[1362]), .Q(ein[338]) );
  DFF \ereg_reg[339]  ( .D(ereg_next[339]), .CLK(clk), .RST(rst), .I(
        e_init[1363]), .Q(ein[339]) );
  DFF \ereg_reg[340]  ( .D(ereg_next[340]), .CLK(clk), .RST(rst), .I(
        e_init[1364]), .Q(ein[340]) );
  DFF \ereg_reg[341]  ( .D(ereg_next[341]), .CLK(clk), .RST(rst), .I(
        e_init[1365]), .Q(ein[341]) );
  DFF \ereg_reg[342]  ( .D(ereg_next[342]), .CLK(clk), .RST(rst), .I(
        e_init[1366]), .Q(ein[342]) );
  DFF \ereg_reg[343]  ( .D(ereg_next[343]), .CLK(clk), .RST(rst), .I(
        e_init[1367]), .Q(ein[343]) );
  DFF \ereg_reg[344]  ( .D(ereg_next[344]), .CLK(clk), .RST(rst), .I(
        e_init[1368]), .Q(ein[344]) );
  DFF \ereg_reg[345]  ( .D(ereg_next[345]), .CLK(clk), .RST(rst), .I(
        e_init[1369]), .Q(ein[345]) );
  DFF \ereg_reg[346]  ( .D(ereg_next[346]), .CLK(clk), .RST(rst), .I(
        e_init[1370]), .Q(ein[346]) );
  DFF \ereg_reg[347]  ( .D(ereg_next[347]), .CLK(clk), .RST(rst), .I(
        e_init[1371]), .Q(ein[347]) );
  DFF \ereg_reg[348]  ( .D(ereg_next[348]), .CLK(clk), .RST(rst), .I(
        e_init[1372]), .Q(ein[348]) );
  DFF \ereg_reg[349]  ( .D(ereg_next[349]), .CLK(clk), .RST(rst), .I(
        e_init[1373]), .Q(ein[349]) );
  DFF \ereg_reg[350]  ( .D(ereg_next[350]), .CLK(clk), .RST(rst), .I(
        e_init[1374]), .Q(ein[350]) );
  DFF \ereg_reg[351]  ( .D(ereg_next[351]), .CLK(clk), .RST(rst), .I(
        e_init[1375]), .Q(ein[351]) );
  DFF \ereg_reg[352]  ( .D(ereg_next[352]), .CLK(clk), .RST(rst), .I(
        e_init[1376]), .Q(ein[352]) );
  DFF \ereg_reg[353]  ( .D(ereg_next[353]), .CLK(clk), .RST(rst), .I(
        e_init[1377]), .Q(ein[353]) );
  DFF \ereg_reg[354]  ( .D(ereg_next[354]), .CLK(clk), .RST(rst), .I(
        e_init[1378]), .Q(ein[354]) );
  DFF \ereg_reg[355]  ( .D(ereg_next[355]), .CLK(clk), .RST(rst), .I(
        e_init[1379]), .Q(ein[355]) );
  DFF \ereg_reg[356]  ( .D(ereg_next[356]), .CLK(clk), .RST(rst), .I(
        e_init[1380]), .Q(ein[356]) );
  DFF \ereg_reg[357]  ( .D(ereg_next[357]), .CLK(clk), .RST(rst), .I(
        e_init[1381]), .Q(ein[357]) );
  DFF \ereg_reg[358]  ( .D(ereg_next[358]), .CLK(clk), .RST(rst), .I(
        e_init[1382]), .Q(ein[358]) );
  DFF \ereg_reg[359]  ( .D(ereg_next[359]), .CLK(clk), .RST(rst), .I(
        e_init[1383]), .Q(ein[359]) );
  DFF \ereg_reg[360]  ( .D(ereg_next[360]), .CLK(clk), .RST(rst), .I(
        e_init[1384]), .Q(ein[360]) );
  DFF \ereg_reg[361]  ( .D(ereg_next[361]), .CLK(clk), .RST(rst), .I(
        e_init[1385]), .Q(ein[361]) );
  DFF \ereg_reg[362]  ( .D(ereg_next[362]), .CLK(clk), .RST(rst), .I(
        e_init[1386]), .Q(ein[362]) );
  DFF \ereg_reg[363]  ( .D(ereg_next[363]), .CLK(clk), .RST(rst), .I(
        e_init[1387]), .Q(ein[363]) );
  DFF \ereg_reg[364]  ( .D(ereg_next[364]), .CLK(clk), .RST(rst), .I(
        e_init[1388]), .Q(ein[364]) );
  DFF \ereg_reg[365]  ( .D(ereg_next[365]), .CLK(clk), .RST(rst), .I(
        e_init[1389]), .Q(ein[365]) );
  DFF \ereg_reg[366]  ( .D(ereg_next[366]), .CLK(clk), .RST(rst), .I(
        e_init[1390]), .Q(ein[366]) );
  DFF \ereg_reg[367]  ( .D(ereg_next[367]), .CLK(clk), .RST(rst), .I(
        e_init[1391]), .Q(ein[367]) );
  DFF \ereg_reg[368]  ( .D(ereg_next[368]), .CLK(clk), .RST(rst), .I(
        e_init[1392]), .Q(ein[368]) );
  DFF \ereg_reg[369]  ( .D(ereg_next[369]), .CLK(clk), .RST(rst), .I(
        e_init[1393]), .Q(ein[369]) );
  DFF \ereg_reg[370]  ( .D(ereg_next[370]), .CLK(clk), .RST(rst), .I(
        e_init[1394]), .Q(ein[370]) );
  DFF \ereg_reg[371]  ( .D(ereg_next[371]), .CLK(clk), .RST(rst), .I(
        e_init[1395]), .Q(ein[371]) );
  DFF \ereg_reg[372]  ( .D(ereg_next[372]), .CLK(clk), .RST(rst), .I(
        e_init[1396]), .Q(ein[372]) );
  DFF \ereg_reg[373]  ( .D(ereg_next[373]), .CLK(clk), .RST(rst), .I(
        e_init[1397]), .Q(ein[373]) );
  DFF \ereg_reg[374]  ( .D(ereg_next[374]), .CLK(clk), .RST(rst), .I(
        e_init[1398]), .Q(ein[374]) );
  DFF \ereg_reg[375]  ( .D(ereg_next[375]), .CLK(clk), .RST(rst), .I(
        e_init[1399]), .Q(ein[375]) );
  DFF \ereg_reg[376]  ( .D(ereg_next[376]), .CLK(clk), .RST(rst), .I(
        e_init[1400]), .Q(ein[376]) );
  DFF \ereg_reg[377]  ( .D(ereg_next[377]), .CLK(clk), .RST(rst), .I(
        e_init[1401]), .Q(ein[377]) );
  DFF \ereg_reg[378]  ( .D(ereg_next[378]), .CLK(clk), .RST(rst), .I(
        e_init[1402]), .Q(ein[378]) );
  DFF \ereg_reg[379]  ( .D(ereg_next[379]), .CLK(clk), .RST(rst), .I(
        e_init[1403]), .Q(ein[379]) );
  DFF \ereg_reg[380]  ( .D(ereg_next[380]), .CLK(clk), .RST(rst), .I(
        e_init[1404]), .Q(ein[380]) );
  DFF \ereg_reg[381]  ( .D(ereg_next[381]), .CLK(clk), .RST(rst), .I(
        e_init[1405]), .Q(ein[381]) );
  DFF \ereg_reg[382]  ( .D(ereg_next[382]), .CLK(clk), .RST(rst), .I(
        e_init[1406]), .Q(ein[382]) );
  DFF \ereg_reg[383]  ( .D(ereg_next[383]), .CLK(clk), .RST(rst), .I(
        e_init[1407]), .Q(ein[383]) );
  DFF \ereg_reg[384]  ( .D(ereg_next[384]), .CLK(clk), .RST(rst), .I(
        e_init[1408]), .Q(ein[384]) );
  DFF \ereg_reg[385]  ( .D(ereg_next[385]), .CLK(clk), .RST(rst), .I(
        e_init[1409]), .Q(ein[385]) );
  DFF \ereg_reg[386]  ( .D(ereg_next[386]), .CLK(clk), .RST(rst), .I(
        e_init[1410]), .Q(ein[386]) );
  DFF \ereg_reg[387]  ( .D(ereg_next[387]), .CLK(clk), .RST(rst), .I(
        e_init[1411]), .Q(ein[387]) );
  DFF \ereg_reg[388]  ( .D(ereg_next[388]), .CLK(clk), .RST(rst), .I(
        e_init[1412]), .Q(ein[388]) );
  DFF \ereg_reg[389]  ( .D(ereg_next[389]), .CLK(clk), .RST(rst), .I(
        e_init[1413]), .Q(ein[389]) );
  DFF \ereg_reg[390]  ( .D(ereg_next[390]), .CLK(clk), .RST(rst), .I(
        e_init[1414]), .Q(ein[390]) );
  DFF \ereg_reg[391]  ( .D(ereg_next[391]), .CLK(clk), .RST(rst), .I(
        e_init[1415]), .Q(ein[391]) );
  DFF \ereg_reg[392]  ( .D(ereg_next[392]), .CLK(clk), .RST(rst), .I(
        e_init[1416]), .Q(ein[392]) );
  DFF \ereg_reg[393]  ( .D(ereg_next[393]), .CLK(clk), .RST(rst), .I(
        e_init[1417]), .Q(ein[393]) );
  DFF \ereg_reg[394]  ( .D(ereg_next[394]), .CLK(clk), .RST(rst), .I(
        e_init[1418]), .Q(ein[394]) );
  DFF \ereg_reg[395]  ( .D(ereg_next[395]), .CLK(clk), .RST(rst), .I(
        e_init[1419]), .Q(ein[395]) );
  DFF \ereg_reg[396]  ( .D(ereg_next[396]), .CLK(clk), .RST(rst), .I(
        e_init[1420]), .Q(ein[396]) );
  DFF \ereg_reg[397]  ( .D(ereg_next[397]), .CLK(clk), .RST(rst), .I(
        e_init[1421]), .Q(ein[397]) );
  DFF \ereg_reg[398]  ( .D(ereg_next[398]), .CLK(clk), .RST(rst), .I(
        e_init[1422]), .Q(ein[398]) );
  DFF \ereg_reg[399]  ( .D(ereg_next[399]), .CLK(clk), .RST(rst), .I(
        e_init[1423]), .Q(ein[399]) );
  DFF \ereg_reg[400]  ( .D(ereg_next[400]), .CLK(clk), .RST(rst), .I(
        e_init[1424]), .Q(ein[400]) );
  DFF \ereg_reg[401]  ( .D(ereg_next[401]), .CLK(clk), .RST(rst), .I(
        e_init[1425]), .Q(ein[401]) );
  DFF \ereg_reg[402]  ( .D(ereg_next[402]), .CLK(clk), .RST(rst), .I(
        e_init[1426]), .Q(ein[402]) );
  DFF \ereg_reg[403]  ( .D(ereg_next[403]), .CLK(clk), .RST(rst), .I(
        e_init[1427]), .Q(ein[403]) );
  DFF \ereg_reg[404]  ( .D(ereg_next[404]), .CLK(clk), .RST(rst), .I(
        e_init[1428]), .Q(ein[404]) );
  DFF \ereg_reg[405]  ( .D(ereg_next[405]), .CLK(clk), .RST(rst), .I(
        e_init[1429]), .Q(ein[405]) );
  DFF \ereg_reg[406]  ( .D(ereg_next[406]), .CLK(clk), .RST(rst), .I(
        e_init[1430]), .Q(ein[406]) );
  DFF \ereg_reg[407]  ( .D(ereg_next[407]), .CLK(clk), .RST(rst), .I(
        e_init[1431]), .Q(ein[407]) );
  DFF \ereg_reg[408]  ( .D(ereg_next[408]), .CLK(clk), .RST(rst), .I(
        e_init[1432]), .Q(ein[408]) );
  DFF \ereg_reg[409]  ( .D(ereg_next[409]), .CLK(clk), .RST(rst), .I(
        e_init[1433]), .Q(ein[409]) );
  DFF \ereg_reg[410]  ( .D(ereg_next[410]), .CLK(clk), .RST(rst), .I(
        e_init[1434]), .Q(ein[410]) );
  DFF \ereg_reg[411]  ( .D(ereg_next[411]), .CLK(clk), .RST(rst), .I(
        e_init[1435]), .Q(ein[411]) );
  DFF \ereg_reg[412]  ( .D(ereg_next[412]), .CLK(clk), .RST(rst), .I(
        e_init[1436]), .Q(ein[412]) );
  DFF \ereg_reg[413]  ( .D(ereg_next[413]), .CLK(clk), .RST(rst), .I(
        e_init[1437]), .Q(ein[413]) );
  DFF \ereg_reg[414]  ( .D(ereg_next[414]), .CLK(clk), .RST(rst), .I(
        e_init[1438]), .Q(ein[414]) );
  DFF \ereg_reg[415]  ( .D(ereg_next[415]), .CLK(clk), .RST(rst), .I(
        e_init[1439]), .Q(ein[415]) );
  DFF \ereg_reg[416]  ( .D(ereg_next[416]), .CLK(clk), .RST(rst), .I(
        e_init[1440]), .Q(ein[416]) );
  DFF \ereg_reg[417]  ( .D(ereg_next[417]), .CLK(clk), .RST(rst), .I(
        e_init[1441]), .Q(ein[417]) );
  DFF \ereg_reg[418]  ( .D(ereg_next[418]), .CLK(clk), .RST(rst), .I(
        e_init[1442]), .Q(ein[418]) );
  DFF \ereg_reg[419]  ( .D(ereg_next[419]), .CLK(clk), .RST(rst), .I(
        e_init[1443]), .Q(ein[419]) );
  DFF \ereg_reg[420]  ( .D(ereg_next[420]), .CLK(clk), .RST(rst), .I(
        e_init[1444]), .Q(ein[420]) );
  DFF \ereg_reg[421]  ( .D(ereg_next[421]), .CLK(clk), .RST(rst), .I(
        e_init[1445]), .Q(ein[421]) );
  DFF \ereg_reg[422]  ( .D(ereg_next[422]), .CLK(clk), .RST(rst), .I(
        e_init[1446]), .Q(ein[422]) );
  DFF \ereg_reg[423]  ( .D(ereg_next[423]), .CLK(clk), .RST(rst), .I(
        e_init[1447]), .Q(ein[423]) );
  DFF \ereg_reg[424]  ( .D(ereg_next[424]), .CLK(clk), .RST(rst), .I(
        e_init[1448]), .Q(ein[424]) );
  DFF \ereg_reg[425]  ( .D(ereg_next[425]), .CLK(clk), .RST(rst), .I(
        e_init[1449]), .Q(ein[425]) );
  DFF \ereg_reg[426]  ( .D(ereg_next[426]), .CLK(clk), .RST(rst), .I(
        e_init[1450]), .Q(ein[426]) );
  DFF \ereg_reg[427]  ( .D(ereg_next[427]), .CLK(clk), .RST(rst), .I(
        e_init[1451]), .Q(ein[427]) );
  DFF \ereg_reg[428]  ( .D(ereg_next[428]), .CLK(clk), .RST(rst), .I(
        e_init[1452]), .Q(ein[428]) );
  DFF \ereg_reg[429]  ( .D(ereg_next[429]), .CLK(clk), .RST(rst), .I(
        e_init[1453]), .Q(ein[429]) );
  DFF \ereg_reg[430]  ( .D(ereg_next[430]), .CLK(clk), .RST(rst), .I(
        e_init[1454]), .Q(ein[430]) );
  DFF \ereg_reg[431]  ( .D(ereg_next[431]), .CLK(clk), .RST(rst), .I(
        e_init[1455]), .Q(ein[431]) );
  DFF \ereg_reg[432]  ( .D(ereg_next[432]), .CLK(clk), .RST(rst), .I(
        e_init[1456]), .Q(ein[432]) );
  DFF \ereg_reg[433]  ( .D(ereg_next[433]), .CLK(clk), .RST(rst), .I(
        e_init[1457]), .Q(ein[433]) );
  DFF \ereg_reg[434]  ( .D(ereg_next[434]), .CLK(clk), .RST(rst), .I(
        e_init[1458]), .Q(ein[434]) );
  DFF \ereg_reg[435]  ( .D(ereg_next[435]), .CLK(clk), .RST(rst), .I(
        e_init[1459]), .Q(ein[435]) );
  DFF \ereg_reg[436]  ( .D(ereg_next[436]), .CLK(clk), .RST(rst), .I(
        e_init[1460]), .Q(ein[436]) );
  DFF \ereg_reg[437]  ( .D(ereg_next[437]), .CLK(clk), .RST(rst), .I(
        e_init[1461]), .Q(ein[437]) );
  DFF \ereg_reg[438]  ( .D(ereg_next[438]), .CLK(clk), .RST(rst), .I(
        e_init[1462]), .Q(ein[438]) );
  DFF \ereg_reg[439]  ( .D(ereg_next[439]), .CLK(clk), .RST(rst), .I(
        e_init[1463]), .Q(ein[439]) );
  DFF \ereg_reg[440]  ( .D(ereg_next[440]), .CLK(clk), .RST(rst), .I(
        e_init[1464]), .Q(ein[440]) );
  DFF \ereg_reg[441]  ( .D(ereg_next[441]), .CLK(clk), .RST(rst), .I(
        e_init[1465]), .Q(ein[441]) );
  DFF \ereg_reg[442]  ( .D(ereg_next[442]), .CLK(clk), .RST(rst), .I(
        e_init[1466]), .Q(ein[442]) );
  DFF \ereg_reg[443]  ( .D(ereg_next[443]), .CLK(clk), .RST(rst), .I(
        e_init[1467]), .Q(ein[443]) );
  DFF \ereg_reg[444]  ( .D(ereg_next[444]), .CLK(clk), .RST(rst), .I(
        e_init[1468]), .Q(ein[444]) );
  DFF \ereg_reg[445]  ( .D(ereg_next[445]), .CLK(clk), .RST(rst), .I(
        e_init[1469]), .Q(ein[445]) );
  DFF \ereg_reg[446]  ( .D(ereg_next[446]), .CLK(clk), .RST(rst), .I(
        e_init[1470]), .Q(ein[446]) );
  DFF \ereg_reg[447]  ( .D(ereg_next[447]), .CLK(clk), .RST(rst), .I(
        e_init[1471]), .Q(ein[447]) );
  DFF \ereg_reg[448]  ( .D(ereg_next[448]), .CLK(clk), .RST(rst), .I(
        e_init[1472]), .Q(ein[448]) );
  DFF \ereg_reg[449]  ( .D(ereg_next[449]), .CLK(clk), .RST(rst), .I(
        e_init[1473]), .Q(ein[449]) );
  DFF \ereg_reg[450]  ( .D(ereg_next[450]), .CLK(clk), .RST(rst), .I(
        e_init[1474]), .Q(ein[450]) );
  DFF \ereg_reg[451]  ( .D(ereg_next[451]), .CLK(clk), .RST(rst), .I(
        e_init[1475]), .Q(ein[451]) );
  DFF \ereg_reg[452]  ( .D(ereg_next[452]), .CLK(clk), .RST(rst), .I(
        e_init[1476]), .Q(ein[452]) );
  DFF \ereg_reg[453]  ( .D(ereg_next[453]), .CLK(clk), .RST(rst), .I(
        e_init[1477]), .Q(ein[453]) );
  DFF \ereg_reg[454]  ( .D(ereg_next[454]), .CLK(clk), .RST(rst), .I(
        e_init[1478]), .Q(ein[454]) );
  DFF \ereg_reg[455]  ( .D(ereg_next[455]), .CLK(clk), .RST(rst), .I(
        e_init[1479]), .Q(ein[455]) );
  DFF \ereg_reg[456]  ( .D(ereg_next[456]), .CLK(clk), .RST(rst), .I(
        e_init[1480]), .Q(ein[456]) );
  DFF \ereg_reg[457]  ( .D(ereg_next[457]), .CLK(clk), .RST(rst), .I(
        e_init[1481]), .Q(ein[457]) );
  DFF \ereg_reg[458]  ( .D(ereg_next[458]), .CLK(clk), .RST(rst), .I(
        e_init[1482]), .Q(ein[458]) );
  DFF \ereg_reg[459]  ( .D(ereg_next[459]), .CLK(clk), .RST(rst), .I(
        e_init[1483]), .Q(ein[459]) );
  DFF \ereg_reg[460]  ( .D(ereg_next[460]), .CLK(clk), .RST(rst), .I(
        e_init[1484]), .Q(ein[460]) );
  DFF \ereg_reg[461]  ( .D(ereg_next[461]), .CLK(clk), .RST(rst), .I(
        e_init[1485]), .Q(ein[461]) );
  DFF \ereg_reg[462]  ( .D(ereg_next[462]), .CLK(clk), .RST(rst), .I(
        e_init[1486]), .Q(ein[462]) );
  DFF \ereg_reg[463]  ( .D(ereg_next[463]), .CLK(clk), .RST(rst), .I(
        e_init[1487]), .Q(ein[463]) );
  DFF \ereg_reg[464]  ( .D(ereg_next[464]), .CLK(clk), .RST(rst), .I(
        e_init[1488]), .Q(ein[464]) );
  DFF \ereg_reg[465]  ( .D(ereg_next[465]), .CLK(clk), .RST(rst), .I(
        e_init[1489]), .Q(ein[465]) );
  DFF \ereg_reg[466]  ( .D(ereg_next[466]), .CLK(clk), .RST(rst), .I(
        e_init[1490]), .Q(ein[466]) );
  DFF \ereg_reg[467]  ( .D(ereg_next[467]), .CLK(clk), .RST(rst), .I(
        e_init[1491]), .Q(ein[467]) );
  DFF \ereg_reg[468]  ( .D(ereg_next[468]), .CLK(clk), .RST(rst), .I(
        e_init[1492]), .Q(ein[468]) );
  DFF \ereg_reg[469]  ( .D(ereg_next[469]), .CLK(clk), .RST(rst), .I(
        e_init[1493]), .Q(ein[469]) );
  DFF \ereg_reg[470]  ( .D(ereg_next[470]), .CLK(clk), .RST(rst), .I(
        e_init[1494]), .Q(ein[470]) );
  DFF \ereg_reg[471]  ( .D(ereg_next[471]), .CLK(clk), .RST(rst), .I(
        e_init[1495]), .Q(ein[471]) );
  DFF \ereg_reg[472]  ( .D(ereg_next[472]), .CLK(clk), .RST(rst), .I(
        e_init[1496]), .Q(ein[472]) );
  DFF \ereg_reg[473]  ( .D(ereg_next[473]), .CLK(clk), .RST(rst), .I(
        e_init[1497]), .Q(ein[473]) );
  DFF \ereg_reg[474]  ( .D(ereg_next[474]), .CLK(clk), .RST(rst), .I(
        e_init[1498]), .Q(ein[474]) );
  DFF \ereg_reg[475]  ( .D(ereg_next[475]), .CLK(clk), .RST(rst), .I(
        e_init[1499]), .Q(ein[475]) );
  DFF \ereg_reg[476]  ( .D(ereg_next[476]), .CLK(clk), .RST(rst), .I(
        e_init[1500]), .Q(ein[476]) );
  DFF \ereg_reg[477]  ( .D(ereg_next[477]), .CLK(clk), .RST(rst), .I(
        e_init[1501]), .Q(ein[477]) );
  DFF \ereg_reg[478]  ( .D(ereg_next[478]), .CLK(clk), .RST(rst), .I(
        e_init[1502]), .Q(ein[478]) );
  DFF \ereg_reg[479]  ( .D(ereg_next[479]), .CLK(clk), .RST(rst), .I(
        e_init[1503]), .Q(ein[479]) );
  DFF \ereg_reg[480]  ( .D(ereg_next[480]), .CLK(clk), .RST(rst), .I(
        e_init[1504]), .Q(ein[480]) );
  DFF \ereg_reg[481]  ( .D(ereg_next[481]), .CLK(clk), .RST(rst), .I(
        e_init[1505]), .Q(ein[481]) );
  DFF \ereg_reg[482]  ( .D(ereg_next[482]), .CLK(clk), .RST(rst), .I(
        e_init[1506]), .Q(ein[482]) );
  DFF \ereg_reg[483]  ( .D(ereg_next[483]), .CLK(clk), .RST(rst), .I(
        e_init[1507]), .Q(ein[483]) );
  DFF \ereg_reg[484]  ( .D(ereg_next[484]), .CLK(clk), .RST(rst), .I(
        e_init[1508]), .Q(ein[484]) );
  DFF \ereg_reg[485]  ( .D(ereg_next[485]), .CLK(clk), .RST(rst), .I(
        e_init[1509]), .Q(ein[485]) );
  DFF \ereg_reg[486]  ( .D(ereg_next[486]), .CLK(clk), .RST(rst), .I(
        e_init[1510]), .Q(ein[486]) );
  DFF \ereg_reg[487]  ( .D(ereg_next[487]), .CLK(clk), .RST(rst), .I(
        e_init[1511]), .Q(ein[487]) );
  DFF \ereg_reg[488]  ( .D(ereg_next[488]), .CLK(clk), .RST(rst), .I(
        e_init[1512]), .Q(ein[488]) );
  DFF \ereg_reg[489]  ( .D(ereg_next[489]), .CLK(clk), .RST(rst), .I(
        e_init[1513]), .Q(ein[489]) );
  DFF \ereg_reg[490]  ( .D(ereg_next[490]), .CLK(clk), .RST(rst), .I(
        e_init[1514]), .Q(ein[490]) );
  DFF \ereg_reg[491]  ( .D(ereg_next[491]), .CLK(clk), .RST(rst), .I(
        e_init[1515]), .Q(ein[491]) );
  DFF \ereg_reg[492]  ( .D(ereg_next[492]), .CLK(clk), .RST(rst), .I(
        e_init[1516]), .Q(ein[492]) );
  DFF \ereg_reg[493]  ( .D(ereg_next[493]), .CLK(clk), .RST(rst), .I(
        e_init[1517]), .Q(ein[493]) );
  DFF \ereg_reg[494]  ( .D(ereg_next[494]), .CLK(clk), .RST(rst), .I(
        e_init[1518]), .Q(ein[494]) );
  DFF \ereg_reg[495]  ( .D(ereg_next[495]), .CLK(clk), .RST(rst), .I(
        e_init[1519]), .Q(ein[495]) );
  DFF \ereg_reg[496]  ( .D(ereg_next[496]), .CLK(clk), .RST(rst), .I(
        e_init[1520]), .Q(ein[496]) );
  DFF \ereg_reg[497]  ( .D(ereg_next[497]), .CLK(clk), .RST(rst), .I(
        e_init[1521]), .Q(ein[497]) );
  DFF \ereg_reg[498]  ( .D(ereg_next[498]), .CLK(clk), .RST(rst), .I(
        e_init[1522]), .Q(ein[498]) );
  DFF \ereg_reg[499]  ( .D(ereg_next[499]), .CLK(clk), .RST(rst), .I(
        e_init[1523]), .Q(ein[499]) );
  DFF \ereg_reg[500]  ( .D(ereg_next[500]), .CLK(clk), .RST(rst), .I(
        e_init[1524]), .Q(ein[500]) );
  DFF \ereg_reg[501]  ( .D(ereg_next[501]), .CLK(clk), .RST(rst), .I(
        e_init[1525]), .Q(ein[501]) );
  DFF \ereg_reg[502]  ( .D(ereg_next[502]), .CLK(clk), .RST(rst), .I(
        e_init[1526]), .Q(ein[502]) );
  DFF \ereg_reg[503]  ( .D(ereg_next[503]), .CLK(clk), .RST(rst), .I(
        e_init[1527]), .Q(ein[503]) );
  DFF \ereg_reg[504]  ( .D(ereg_next[504]), .CLK(clk), .RST(rst), .I(
        e_init[1528]), .Q(ein[504]) );
  DFF \ereg_reg[505]  ( .D(ereg_next[505]), .CLK(clk), .RST(rst), .I(
        e_init[1529]), .Q(ein[505]) );
  DFF \ereg_reg[506]  ( .D(ereg_next[506]), .CLK(clk), .RST(rst), .I(
        e_init[1530]), .Q(ein[506]) );
  DFF \ereg_reg[507]  ( .D(ereg_next[507]), .CLK(clk), .RST(rst), .I(
        e_init[1531]), .Q(ein[507]) );
  DFF \ereg_reg[508]  ( .D(ereg_next[508]), .CLK(clk), .RST(rst), .I(
        e_init[1532]), .Q(ein[508]) );
  DFF \ereg_reg[509]  ( .D(ereg_next[509]), .CLK(clk), .RST(rst), .I(
        e_init[1533]), .Q(ein[509]) );
  DFF \ereg_reg[510]  ( .D(ereg_next[510]), .CLK(clk), .RST(rst), .I(
        e_init[1534]), .Q(ein[510]) );
  DFF \ereg_reg[511]  ( .D(ereg_next[511]), .CLK(clk), .RST(rst), .I(
        e_init[1535]), .Q(ein[511]) );
  DFF \ereg_reg[512]  ( .D(ereg_next[512]), .CLK(clk), .RST(rst), .I(
        e_init[1536]), .Q(ein[512]) );
  DFF \ereg_reg[513]  ( .D(ereg_next[513]), .CLK(clk), .RST(rst), .I(
        e_init[1537]), .Q(ein[513]) );
  DFF \ereg_reg[514]  ( .D(ereg_next[514]), .CLK(clk), .RST(rst), .I(
        e_init[1538]), .Q(ein[514]) );
  DFF \ereg_reg[515]  ( .D(ereg_next[515]), .CLK(clk), .RST(rst), .I(
        e_init[1539]), .Q(ein[515]) );
  DFF \ereg_reg[516]  ( .D(ereg_next[516]), .CLK(clk), .RST(rst), .I(
        e_init[1540]), .Q(ein[516]) );
  DFF \ereg_reg[517]  ( .D(ereg_next[517]), .CLK(clk), .RST(rst), .I(
        e_init[1541]), .Q(ein[517]) );
  DFF \ereg_reg[518]  ( .D(ereg_next[518]), .CLK(clk), .RST(rst), .I(
        e_init[1542]), .Q(ein[518]) );
  DFF \ereg_reg[519]  ( .D(ereg_next[519]), .CLK(clk), .RST(rst), .I(
        e_init[1543]), .Q(ein[519]) );
  DFF \ereg_reg[520]  ( .D(ereg_next[520]), .CLK(clk), .RST(rst), .I(
        e_init[1544]), .Q(ein[520]) );
  DFF \ereg_reg[521]  ( .D(ereg_next[521]), .CLK(clk), .RST(rst), .I(
        e_init[1545]), .Q(ein[521]) );
  DFF \ereg_reg[522]  ( .D(ereg_next[522]), .CLK(clk), .RST(rst), .I(
        e_init[1546]), .Q(ein[522]) );
  DFF \ereg_reg[523]  ( .D(ereg_next[523]), .CLK(clk), .RST(rst), .I(
        e_init[1547]), .Q(ein[523]) );
  DFF \ereg_reg[524]  ( .D(ereg_next[524]), .CLK(clk), .RST(rst), .I(
        e_init[1548]), .Q(ein[524]) );
  DFF \ereg_reg[525]  ( .D(ereg_next[525]), .CLK(clk), .RST(rst), .I(
        e_init[1549]), .Q(ein[525]) );
  DFF \ereg_reg[526]  ( .D(ereg_next[526]), .CLK(clk), .RST(rst), .I(
        e_init[1550]), .Q(ein[526]) );
  DFF \ereg_reg[527]  ( .D(ereg_next[527]), .CLK(clk), .RST(rst), .I(
        e_init[1551]), .Q(ein[527]) );
  DFF \ereg_reg[528]  ( .D(ereg_next[528]), .CLK(clk), .RST(rst), .I(
        e_init[1552]), .Q(ein[528]) );
  DFF \ereg_reg[529]  ( .D(ereg_next[529]), .CLK(clk), .RST(rst), .I(
        e_init[1553]), .Q(ein[529]) );
  DFF \ereg_reg[530]  ( .D(ereg_next[530]), .CLK(clk), .RST(rst), .I(
        e_init[1554]), .Q(ein[530]) );
  DFF \ereg_reg[531]  ( .D(ereg_next[531]), .CLK(clk), .RST(rst), .I(
        e_init[1555]), .Q(ein[531]) );
  DFF \ereg_reg[532]  ( .D(ereg_next[532]), .CLK(clk), .RST(rst), .I(
        e_init[1556]), .Q(ein[532]) );
  DFF \ereg_reg[533]  ( .D(ereg_next[533]), .CLK(clk), .RST(rst), .I(
        e_init[1557]), .Q(ein[533]) );
  DFF \ereg_reg[534]  ( .D(ereg_next[534]), .CLK(clk), .RST(rst), .I(
        e_init[1558]), .Q(ein[534]) );
  DFF \ereg_reg[535]  ( .D(ereg_next[535]), .CLK(clk), .RST(rst), .I(
        e_init[1559]), .Q(ein[535]) );
  DFF \ereg_reg[536]  ( .D(ereg_next[536]), .CLK(clk), .RST(rst), .I(
        e_init[1560]), .Q(ein[536]) );
  DFF \ereg_reg[537]  ( .D(ereg_next[537]), .CLK(clk), .RST(rst), .I(
        e_init[1561]), .Q(ein[537]) );
  DFF \ereg_reg[538]  ( .D(ereg_next[538]), .CLK(clk), .RST(rst), .I(
        e_init[1562]), .Q(ein[538]) );
  DFF \ereg_reg[539]  ( .D(ereg_next[539]), .CLK(clk), .RST(rst), .I(
        e_init[1563]), .Q(ein[539]) );
  DFF \ereg_reg[540]  ( .D(ereg_next[540]), .CLK(clk), .RST(rst), .I(
        e_init[1564]), .Q(ein[540]) );
  DFF \ereg_reg[541]  ( .D(ereg_next[541]), .CLK(clk), .RST(rst), .I(
        e_init[1565]), .Q(ein[541]) );
  DFF \ereg_reg[542]  ( .D(ereg_next[542]), .CLK(clk), .RST(rst), .I(
        e_init[1566]), .Q(ein[542]) );
  DFF \ereg_reg[543]  ( .D(ereg_next[543]), .CLK(clk), .RST(rst), .I(
        e_init[1567]), .Q(ein[543]) );
  DFF \ereg_reg[544]  ( .D(ereg_next[544]), .CLK(clk), .RST(rst), .I(
        e_init[1568]), .Q(ein[544]) );
  DFF \ereg_reg[545]  ( .D(ereg_next[545]), .CLK(clk), .RST(rst), .I(
        e_init[1569]), .Q(ein[545]) );
  DFF \ereg_reg[546]  ( .D(ereg_next[546]), .CLK(clk), .RST(rst), .I(
        e_init[1570]), .Q(ein[546]) );
  DFF \ereg_reg[547]  ( .D(ereg_next[547]), .CLK(clk), .RST(rst), .I(
        e_init[1571]), .Q(ein[547]) );
  DFF \ereg_reg[548]  ( .D(ereg_next[548]), .CLK(clk), .RST(rst), .I(
        e_init[1572]), .Q(ein[548]) );
  DFF \ereg_reg[549]  ( .D(ereg_next[549]), .CLK(clk), .RST(rst), .I(
        e_init[1573]), .Q(ein[549]) );
  DFF \ereg_reg[550]  ( .D(ereg_next[550]), .CLK(clk), .RST(rst), .I(
        e_init[1574]), .Q(ein[550]) );
  DFF \ereg_reg[551]  ( .D(ereg_next[551]), .CLK(clk), .RST(rst), .I(
        e_init[1575]), .Q(ein[551]) );
  DFF \ereg_reg[552]  ( .D(ereg_next[552]), .CLK(clk), .RST(rst), .I(
        e_init[1576]), .Q(ein[552]) );
  DFF \ereg_reg[553]  ( .D(ereg_next[553]), .CLK(clk), .RST(rst), .I(
        e_init[1577]), .Q(ein[553]) );
  DFF \ereg_reg[554]  ( .D(ereg_next[554]), .CLK(clk), .RST(rst), .I(
        e_init[1578]), .Q(ein[554]) );
  DFF \ereg_reg[555]  ( .D(ereg_next[555]), .CLK(clk), .RST(rst), .I(
        e_init[1579]), .Q(ein[555]) );
  DFF \ereg_reg[556]  ( .D(ereg_next[556]), .CLK(clk), .RST(rst), .I(
        e_init[1580]), .Q(ein[556]) );
  DFF \ereg_reg[557]  ( .D(ereg_next[557]), .CLK(clk), .RST(rst), .I(
        e_init[1581]), .Q(ein[557]) );
  DFF \ereg_reg[558]  ( .D(ereg_next[558]), .CLK(clk), .RST(rst), .I(
        e_init[1582]), .Q(ein[558]) );
  DFF \ereg_reg[559]  ( .D(ereg_next[559]), .CLK(clk), .RST(rst), .I(
        e_init[1583]), .Q(ein[559]) );
  DFF \ereg_reg[560]  ( .D(ereg_next[560]), .CLK(clk), .RST(rst), .I(
        e_init[1584]), .Q(ein[560]) );
  DFF \ereg_reg[561]  ( .D(ereg_next[561]), .CLK(clk), .RST(rst), .I(
        e_init[1585]), .Q(ein[561]) );
  DFF \ereg_reg[562]  ( .D(ereg_next[562]), .CLK(clk), .RST(rst), .I(
        e_init[1586]), .Q(ein[562]) );
  DFF \ereg_reg[563]  ( .D(ereg_next[563]), .CLK(clk), .RST(rst), .I(
        e_init[1587]), .Q(ein[563]) );
  DFF \ereg_reg[564]  ( .D(ereg_next[564]), .CLK(clk), .RST(rst), .I(
        e_init[1588]), .Q(ein[564]) );
  DFF \ereg_reg[565]  ( .D(ereg_next[565]), .CLK(clk), .RST(rst), .I(
        e_init[1589]), .Q(ein[565]) );
  DFF \ereg_reg[566]  ( .D(ereg_next[566]), .CLK(clk), .RST(rst), .I(
        e_init[1590]), .Q(ein[566]) );
  DFF \ereg_reg[567]  ( .D(ereg_next[567]), .CLK(clk), .RST(rst), .I(
        e_init[1591]), .Q(ein[567]) );
  DFF \ereg_reg[568]  ( .D(ereg_next[568]), .CLK(clk), .RST(rst), .I(
        e_init[1592]), .Q(ein[568]) );
  DFF \ereg_reg[569]  ( .D(ereg_next[569]), .CLK(clk), .RST(rst), .I(
        e_init[1593]), .Q(ein[569]) );
  DFF \ereg_reg[570]  ( .D(ereg_next[570]), .CLK(clk), .RST(rst), .I(
        e_init[1594]), .Q(ein[570]) );
  DFF \ereg_reg[571]  ( .D(ereg_next[571]), .CLK(clk), .RST(rst), .I(
        e_init[1595]), .Q(ein[571]) );
  DFF \ereg_reg[572]  ( .D(ereg_next[572]), .CLK(clk), .RST(rst), .I(
        e_init[1596]), .Q(ein[572]) );
  DFF \ereg_reg[573]  ( .D(ereg_next[573]), .CLK(clk), .RST(rst), .I(
        e_init[1597]), .Q(ein[573]) );
  DFF \ereg_reg[574]  ( .D(ereg_next[574]), .CLK(clk), .RST(rst), .I(
        e_init[1598]), .Q(ein[574]) );
  DFF \ereg_reg[575]  ( .D(ereg_next[575]), .CLK(clk), .RST(rst), .I(
        e_init[1599]), .Q(ein[575]) );
  DFF \ereg_reg[576]  ( .D(ereg_next[576]), .CLK(clk), .RST(rst), .I(
        e_init[1600]), .Q(ein[576]) );
  DFF \ereg_reg[577]  ( .D(ereg_next[577]), .CLK(clk), .RST(rst), .I(
        e_init[1601]), .Q(ein[577]) );
  DFF \ereg_reg[578]  ( .D(ereg_next[578]), .CLK(clk), .RST(rst), .I(
        e_init[1602]), .Q(ein[578]) );
  DFF \ereg_reg[579]  ( .D(ereg_next[579]), .CLK(clk), .RST(rst), .I(
        e_init[1603]), .Q(ein[579]) );
  DFF \ereg_reg[580]  ( .D(ereg_next[580]), .CLK(clk), .RST(rst), .I(
        e_init[1604]), .Q(ein[580]) );
  DFF \ereg_reg[581]  ( .D(ereg_next[581]), .CLK(clk), .RST(rst), .I(
        e_init[1605]), .Q(ein[581]) );
  DFF \ereg_reg[582]  ( .D(ereg_next[582]), .CLK(clk), .RST(rst), .I(
        e_init[1606]), .Q(ein[582]) );
  DFF \ereg_reg[583]  ( .D(ereg_next[583]), .CLK(clk), .RST(rst), .I(
        e_init[1607]), .Q(ein[583]) );
  DFF \ereg_reg[584]  ( .D(ereg_next[584]), .CLK(clk), .RST(rst), .I(
        e_init[1608]), .Q(ein[584]) );
  DFF \ereg_reg[585]  ( .D(ereg_next[585]), .CLK(clk), .RST(rst), .I(
        e_init[1609]), .Q(ein[585]) );
  DFF \ereg_reg[586]  ( .D(ereg_next[586]), .CLK(clk), .RST(rst), .I(
        e_init[1610]), .Q(ein[586]) );
  DFF \ereg_reg[587]  ( .D(ereg_next[587]), .CLK(clk), .RST(rst), .I(
        e_init[1611]), .Q(ein[587]) );
  DFF \ereg_reg[588]  ( .D(ereg_next[588]), .CLK(clk), .RST(rst), .I(
        e_init[1612]), .Q(ein[588]) );
  DFF \ereg_reg[589]  ( .D(ereg_next[589]), .CLK(clk), .RST(rst), .I(
        e_init[1613]), .Q(ein[589]) );
  DFF \ereg_reg[590]  ( .D(ereg_next[590]), .CLK(clk), .RST(rst), .I(
        e_init[1614]), .Q(ein[590]) );
  DFF \ereg_reg[591]  ( .D(ereg_next[591]), .CLK(clk), .RST(rst), .I(
        e_init[1615]), .Q(ein[591]) );
  DFF \ereg_reg[592]  ( .D(ereg_next[592]), .CLK(clk), .RST(rst), .I(
        e_init[1616]), .Q(ein[592]) );
  DFF \ereg_reg[593]  ( .D(ereg_next[593]), .CLK(clk), .RST(rst), .I(
        e_init[1617]), .Q(ein[593]) );
  DFF \ereg_reg[594]  ( .D(ereg_next[594]), .CLK(clk), .RST(rst), .I(
        e_init[1618]), .Q(ein[594]) );
  DFF \ereg_reg[595]  ( .D(ereg_next[595]), .CLK(clk), .RST(rst), .I(
        e_init[1619]), .Q(ein[595]) );
  DFF \ereg_reg[596]  ( .D(ereg_next[596]), .CLK(clk), .RST(rst), .I(
        e_init[1620]), .Q(ein[596]) );
  DFF \ereg_reg[597]  ( .D(ereg_next[597]), .CLK(clk), .RST(rst), .I(
        e_init[1621]), .Q(ein[597]) );
  DFF \ereg_reg[598]  ( .D(ereg_next[598]), .CLK(clk), .RST(rst), .I(
        e_init[1622]), .Q(ein[598]) );
  DFF \ereg_reg[599]  ( .D(ereg_next[599]), .CLK(clk), .RST(rst), .I(
        e_init[1623]), .Q(ein[599]) );
  DFF \ereg_reg[600]  ( .D(ereg_next[600]), .CLK(clk), .RST(rst), .I(
        e_init[1624]), .Q(ein[600]) );
  DFF \ereg_reg[601]  ( .D(ereg_next[601]), .CLK(clk), .RST(rst), .I(
        e_init[1625]), .Q(ein[601]) );
  DFF \ereg_reg[602]  ( .D(ereg_next[602]), .CLK(clk), .RST(rst), .I(
        e_init[1626]), .Q(ein[602]) );
  DFF \ereg_reg[603]  ( .D(ereg_next[603]), .CLK(clk), .RST(rst), .I(
        e_init[1627]), .Q(ein[603]) );
  DFF \ereg_reg[604]  ( .D(ereg_next[604]), .CLK(clk), .RST(rst), .I(
        e_init[1628]), .Q(ein[604]) );
  DFF \ereg_reg[605]  ( .D(ereg_next[605]), .CLK(clk), .RST(rst), .I(
        e_init[1629]), .Q(ein[605]) );
  DFF \ereg_reg[606]  ( .D(ereg_next[606]), .CLK(clk), .RST(rst), .I(
        e_init[1630]), .Q(ein[606]) );
  DFF \ereg_reg[607]  ( .D(ereg_next[607]), .CLK(clk), .RST(rst), .I(
        e_init[1631]), .Q(ein[607]) );
  DFF \ereg_reg[608]  ( .D(ereg_next[608]), .CLK(clk), .RST(rst), .I(
        e_init[1632]), .Q(ein[608]) );
  DFF \ereg_reg[609]  ( .D(ereg_next[609]), .CLK(clk), .RST(rst), .I(
        e_init[1633]), .Q(ein[609]) );
  DFF \ereg_reg[610]  ( .D(ereg_next[610]), .CLK(clk), .RST(rst), .I(
        e_init[1634]), .Q(ein[610]) );
  DFF \ereg_reg[611]  ( .D(ereg_next[611]), .CLK(clk), .RST(rst), .I(
        e_init[1635]), .Q(ein[611]) );
  DFF \ereg_reg[612]  ( .D(ereg_next[612]), .CLK(clk), .RST(rst), .I(
        e_init[1636]), .Q(ein[612]) );
  DFF \ereg_reg[613]  ( .D(ereg_next[613]), .CLK(clk), .RST(rst), .I(
        e_init[1637]), .Q(ein[613]) );
  DFF \ereg_reg[614]  ( .D(ereg_next[614]), .CLK(clk), .RST(rst), .I(
        e_init[1638]), .Q(ein[614]) );
  DFF \ereg_reg[615]  ( .D(ereg_next[615]), .CLK(clk), .RST(rst), .I(
        e_init[1639]), .Q(ein[615]) );
  DFF \ereg_reg[616]  ( .D(ereg_next[616]), .CLK(clk), .RST(rst), .I(
        e_init[1640]), .Q(ein[616]) );
  DFF \ereg_reg[617]  ( .D(ereg_next[617]), .CLK(clk), .RST(rst), .I(
        e_init[1641]), .Q(ein[617]) );
  DFF \ereg_reg[618]  ( .D(ereg_next[618]), .CLK(clk), .RST(rst), .I(
        e_init[1642]), .Q(ein[618]) );
  DFF \ereg_reg[619]  ( .D(ereg_next[619]), .CLK(clk), .RST(rst), .I(
        e_init[1643]), .Q(ein[619]) );
  DFF \ereg_reg[620]  ( .D(ereg_next[620]), .CLK(clk), .RST(rst), .I(
        e_init[1644]), .Q(ein[620]) );
  DFF \ereg_reg[621]  ( .D(ereg_next[621]), .CLK(clk), .RST(rst), .I(
        e_init[1645]), .Q(ein[621]) );
  DFF \ereg_reg[622]  ( .D(ereg_next[622]), .CLK(clk), .RST(rst), .I(
        e_init[1646]), .Q(ein[622]) );
  DFF \ereg_reg[623]  ( .D(ereg_next[623]), .CLK(clk), .RST(rst), .I(
        e_init[1647]), .Q(ein[623]) );
  DFF \ereg_reg[624]  ( .D(ereg_next[624]), .CLK(clk), .RST(rst), .I(
        e_init[1648]), .Q(ein[624]) );
  DFF \ereg_reg[625]  ( .D(ereg_next[625]), .CLK(clk), .RST(rst), .I(
        e_init[1649]), .Q(ein[625]) );
  DFF \ereg_reg[626]  ( .D(ereg_next[626]), .CLK(clk), .RST(rst), .I(
        e_init[1650]), .Q(ein[626]) );
  DFF \ereg_reg[627]  ( .D(ereg_next[627]), .CLK(clk), .RST(rst), .I(
        e_init[1651]), .Q(ein[627]) );
  DFF \ereg_reg[628]  ( .D(ereg_next[628]), .CLK(clk), .RST(rst), .I(
        e_init[1652]), .Q(ein[628]) );
  DFF \ereg_reg[629]  ( .D(ereg_next[629]), .CLK(clk), .RST(rst), .I(
        e_init[1653]), .Q(ein[629]) );
  DFF \ereg_reg[630]  ( .D(ereg_next[630]), .CLK(clk), .RST(rst), .I(
        e_init[1654]), .Q(ein[630]) );
  DFF \ereg_reg[631]  ( .D(ereg_next[631]), .CLK(clk), .RST(rst), .I(
        e_init[1655]), .Q(ein[631]) );
  DFF \ereg_reg[632]  ( .D(ereg_next[632]), .CLK(clk), .RST(rst), .I(
        e_init[1656]), .Q(ein[632]) );
  DFF \ereg_reg[633]  ( .D(ereg_next[633]), .CLK(clk), .RST(rst), .I(
        e_init[1657]), .Q(ein[633]) );
  DFF \ereg_reg[634]  ( .D(ereg_next[634]), .CLK(clk), .RST(rst), .I(
        e_init[1658]), .Q(ein[634]) );
  DFF \ereg_reg[635]  ( .D(ereg_next[635]), .CLK(clk), .RST(rst), .I(
        e_init[1659]), .Q(ein[635]) );
  DFF \ereg_reg[636]  ( .D(ereg_next[636]), .CLK(clk), .RST(rst), .I(
        e_init[1660]), .Q(ein[636]) );
  DFF \ereg_reg[637]  ( .D(ereg_next[637]), .CLK(clk), .RST(rst), .I(
        e_init[1661]), .Q(ein[637]) );
  DFF \ereg_reg[638]  ( .D(ereg_next[638]), .CLK(clk), .RST(rst), .I(
        e_init[1662]), .Q(ein[638]) );
  DFF \ereg_reg[639]  ( .D(ereg_next[639]), .CLK(clk), .RST(rst), .I(
        e_init[1663]), .Q(ein[639]) );
  DFF \ereg_reg[640]  ( .D(ereg_next[640]), .CLK(clk), .RST(rst), .I(
        e_init[1664]), .Q(ein[640]) );
  DFF \ereg_reg[641]  ( .D(ereg_next[641]), .CLK(clk), .RST(rst), .I(
        e_init[1665]), .Q(ein[641]) );
  DFF \ereg_reg[642]  ( .D(ereg_next[642]), .CLK(clk), .RST(rst), .I(
        e_init[1666]), .Q(ein[642]) );
  DFF \ereg_reg[643]  ( .D(ereg_next[643]), .CLK(clk), .RST(rst), .I(
        e_init[1667]), .Q(ein[643]) );
  DFF \ereg_reg[644]  ( .D(ereg_next[644]), .CLK(clk), .RST(rst), .I(
        e_init[1668]), .Q(ein[644]) );
  DFF \ereg_reg[645]  ( .D(ereg_next[645]), .CLK(clk), .RST(rst), .I(
        e_init[1669]), .Q(ein[645]) );
  DFF \ereg_reg[646]  ( .D(ereg_next[646]), .CLK(clk), .RST(rst), .I(
        e_init[1670]), .Q(ein[646]) );
  DFF \ereg_reg[647]  ( .D(ereg_next[647]), .CLK(clk), .RST(rst), .I(
        e_init[1671]), .Q(ein[647]) );
  DFF \ereg_reg[648]  ( .D(ereg_next[648]), .CLK(clk), .RST(rst), .I(
        e_init[1672]), .Q(ein[648]) );
  DFF \ereg_reg[649]  ( .D(ereg_next[649]), .CLK(clk), .RST(rst), .I(
        e_init[1673]), .Q(ein[649]) );
  DFF \ereg_reg[650]  ( .D(ereg_next[650]), .CLK(clk), .RST(rst), .I(
        e_init[1674]), .Q(ein[650]) );
  DFF \ereg_reg[651]  ( .D(ereg_next[651]), .CLK(clk), .RST(rst), .I(
        e_init[1675]), .Q(ein[651]) );
  DFF \ereg_reg[652]  ( .D(ereg_next[652]), .CLK(clk), .RST(rst), .I(
        e_init[1676]), .Q(ein[652]) );
  DFF \ereg_reg[653]  ( .D(ereg_next[653]), .CLK(clk), .RST(rst), .I(
        e_init[1677]), .Q(ein[653]) );
  DFF \ereg_reg[654]  ( .D(ereg_next[654]), .CLK(clk), .RST(rst), .I(
        e_init[1678]), .Q(ein[654]) );
  DFF \ereg_reg[655]  ( .D(ereg_next[655]), .CLK(clk), .RST(rst), .I(
        e_init[1679]), .Q(ein[655]) );
  DFF \ereg_reg[656]  ( .D(ereg_next[656]), .CLK(clk), .RST(rst), .I(
        e_init[1680]), .Q(ein[656]) );
  DFF \ereg_reg[657]  ( .D(ereg_next[657]), .CLK(clk), .RST(rst), .I(
        e_init[1681]), .Q(ein[657]) );
  DFF \ereg_reg[658]  ( .D(ereg_next[658]), .CLK(clk), .RST(rst), .I(
        e_init[1682]), .Q(ein[658]) );
  DFF \ereg_reg[659]  ( .D(ereg_next[659]), .CLK(clk), .RST(rst), .I(
        e_init[1683]), .Q(ein[659]) );
  DFF \ereg_reg[660]  ( .D(ereg_next[660]), .CLK(clk), .RST(rst), .I(
        e_init[1684]), .Q(ein[660]) );
  DFF \ereg_reg[661]  ( .D(ereg_next[661]), .CLK(clk), .RST(rst), .I(
        e_init[1685]), .Q(ein[661]) );
  DFF \ereg_reg[662]  ( .D(ereg_next[662]), .CLK(clk), .RST(rst), .I(
        e_init[1686]), .Q(ein[662]) );
  DFF \ereg_reg[663]  ( .D(ereg_next[663]), .CLK(clk), .RST(rst), .I(
        e_init[1687]), .Q(ein[663]) );
  DFF \ereg_reg[664]  ( .D(ereg_next[664]), .CLK(clk), .RST(rst), .I(
        e_init[1688]), .Q(ein[664]) );
  DFF \ereg_reg[665]  ( .D(ereg_next[665]), .CLK(clk), .RST(rst), .I(
        e_init[1689]), .Q(ein[665]) );
  DFF \ereg_reg[666]  ( .D(ereg_next[666]), .CLK(clk), .RST(rst), .I(
        e_init[1690]), .Q(ein[666]) );
  DFF \ereg_reg[667]  ( .D(ereg_next[667]), .CLK(clk), .RST(rst), .I(
        e_init[1691]), .Q(ein[667]) );
  DFF \ereg_reg[668]  ( .D(ereg_next[668]), .CLK(clk), .RST(rst), .I(
        e_init[1692]), .Q(ein[668]) );
  DFF \ereg_reg[669]  ( .D(ereg_next[669]), .CLK(clk), .RST(rst), .I(
        e_init[1693]), .Q(ein[669]) );
  DFF \ereg_reg[670]  ( .D(ereg_next[670]), .CLK(clk), .RST(rst), .I(
        e_init[1694]), .Q(ein[670]) );
  DFF \ereg_reg[671]  ( .D(ereg_next[671]), .CLK(clk), .RST(rst), .I(
        e_init[1695]), .Q(ein[671]) );
  DFF \ereg_reg[672]  ( .D(ereg_next[672]), .CLK(clk), .RST(rst), .I(
        e_init[1696]), .Q(ein[672]) );
  DFF \ereg_reg[673]  ( .D(ereg_next[673]), .CLK(clk), .RST(rst), .I(
        e_init[1697]), .Q(ein[673]) );
  DFF \ereg_reg[674]  ( .D(ereg_next[674]), .CLK(clk), .RST(rst), .I(
        e_init[1698]), .Q(ein[674]) );
  DFF \ereg_reg[675]  ( .D(ereg_next[675]), .CLK(clk), .RST(rst), .I(
        e_init[1699]), .Q(ein[675]) );
  DFF \ereg_reg[676]  ( .D(ereg_next[676]), .CLK(clk), .RST(rst), .I(
        e_init[1700]), .Q(ein[676]) );
  DFF \ereg_reg[677]  ( .D(ereg_next[677]), .CLK(clk), .RST(rst), .I(
        e_init[1701]), .Q(ein[677]) );
  DFF \ereg_reg[678]  ( .D(ereg_next[678]), .CLK(clk), .RST(rst), .I(
        e_init[1702]), .Q(ein[678]) );
  DFF \ereg_reg[679]  ( .D(ereg_next[679]), .CLK(clk), .RST(rst), .I(
        e_init[1703]), .Q(ein[679]) );
  DFF \ereg_reg[680]  ( .D(ereg_next[680]), .CLK(clk), .RST(rst), .I(
        e_init[1704]), .Q(ein[680]) );
  DFF \ereg_reg[681]  ( .D(ereg_next[681]), .CLK(clk), .RST(rst), .I(
        e_init[1705]), .Q(ein[681]) );
  DFF \ereg_reg[682]  ( .D(ereg_next[682]), .CLK(clk), .RST(rst), .I(
        e_init[1706]), .Q(ein[682]) );
  DFF \ereg_reg[683]  ( .D(ereg_next[683]), .CLK(clk), .RST(rst), .I(
        e_init[1707]), .Q(ein[683]) );
  DFF \ereg_reg[684]  ( .D(ereg_next[684]), .CLK(clk), .RST(rst), .I(
        e_init[1708]), .Q(ein[684]) );
  DFF \ereg_reg[685]  ( .D(ereg_next[685]), .CLK(clk), .RST(rst), .I(
        e_init[1709]), .Q(ein[685]) );
  DFF \ereg_reg[686]  ( .D(ereg_next[686]), .CLK(clk), .RST(rst), .I(
        e_init[1710]), .Q(ein[686]) );
  DFF \ereg_reg[687]  ( .D(ereg_next[687]), .CLK(clk), .RST(rst), .I(
        e_init[1711]), .Q(ein[687]) );
  DFF \ereg_reg[688]  ( .D(ereg_next[688]), .CLK(clk), .RST(rst), .I(
        e_init[1712]), .Q(ein[688]) );
  DFF \ereg_reg[689]  ( .D(ereg_next[689]), .CLK(clk), .RST(rst), .I(
        e_init[1713]), .Q(ein[689]) );
  DFF \ereg_reg[690]  ( .D(ereg_next[690]), .CLK(clk), .RST(rst), .I(
        e_init[1714]), .Q(ein[690]) );
  DFF \ereg_reg[691]  ( .D(ereg_next[691]), .CLK(clk), .RST(rst), .I(
        e_init[1715]), .Q(ein[691]) );
  DFF \ereg_reg[692]  ( .D(ereg_next[692]), .CLK(clk), .RST(rst), .I(
        e_init[1716]), .Q(ein[692]) );
  DFF \ereg_reg[693]  ( .D(ereg_next[693]), .CLK(clk), .RST(rst), .I(
        e_init[1717]), .Q(ein[693]) );
  DFF \ereg_reg[694]  ( .D(ereg_next[694]), .CLK(clk), .RST(rst), .I(
        e_init[1718]), .Q(ein[694]) );
  DFF \ereg_reg[695]  ( .D(ereg_next[695]), .CLK(clk), .RST(rst), .I(
        e_init[1719]), .Q(ein[695]) );
  DFF \ereg_reg[696]  ( .D(ereg_next[696]), .CLK(clk), .RST(rst), .I(
        e_init[1720]), .Q(ein[696]) );
  DFF \ereg_reg[697]  ( .D(ereg_next[697]), .CLK(clk), .RST(rst), .I(
        e_init[1721]), .Q(ein[697]) );
  DFF \ereg_reg[698]  ( .D(ereg_next[698]), .CLK(clk), .RST(rst), .I(
        e_init[1722]), .Q(ein[698]) );
  DFF \ereg_reg[699]  ( .D(ereg_next[699]), .CLK(clk), .RST(rst), .I(
        e_init[1723]), .Q(ein[699]) );
  DFF \ereg_reg[700]  ( .D(ereg_next[700]), .CLK(clk), .RST(rst), .I(
        e_init[1724]), .Q(ein[700]) );
  DFF \ereg_reg[701]  ( .D(ereg_next[701]), .CLK(clk), .RST(rst), .I(
        e_init[1725]), .Q(ein[701]) );
  DFF \ereg_reg[702]  ( .D(ereg_next[702]), .CLK(clk), .RST(rst), .I(
        e_init[1726]), .Q(ein[702]) );
  DFF \ereg_reg[703]  ( .D(ereg_next[703]), .CLK(clk), .RST(rst), .I(
        e_init[1727]), .Q(ein[703]) );
  DFF \ereg_reg[704]  ( .D(ereg_next[704]), .CLK(clk), .RST(rst), .I(
        e_init[1728]), .Q(ein[704]) );
  DFF \ereg_reg[705]  ( .D(ereg_next[705]), .CLK(clk), .RST(rst), .I(
        e_init[1729]), .Q(ein[705]) );
  DFF \ereg_reg[706]  ( .D(ereg_next[706]), .CLK(clk), .RST(rst), .I(
        e_init[1730]), .Q(ein[706]) );
  DFF \ereg_reg[707]  ( .D(ereg_next[707]), .CLK(clk), .RST(rst), .I(
        e_init[1731]), .Q(ein[707]) );
  DFF \ereg_reg[708]  ( .D(ereg_next[708]), .CLK(clk), .RST(rst), .I(
        e_init[1732]), .Q(ein[708]) );
  DFF \ereg_reg[709]  ( .D(ereg_next[709]), .CLK(clk), .RST(rst), .I(
        e_init[1733]), .Q(ein[709]) );
  DFF \ereg_reg[710]  ( .D(ereg_next[710]), .CLK(clk), .RST(rst), .I(
        e_init[1734]), .Q(ein[710]) );
  DFF \ereg_reg[711]  ( .D(ereg_next[711]), .CLK(clk), .RST(rst), .I(
        e_init[1735]), .Q(ein[711]) );
  DFF \ereg_reg[712]  ( .D(ereg_next[712]), .CLK(clk), .RST(rst), .I(
        e_init[1736]), .Q(ein[712]) );
  DFF \ereg_reg[713]  ( .D(ereg_next[713]), .CLK(clk), .RST(rst), .I(
        e_init[1737]), .Q(ein[713]) );
  DFF \ereg_reg[714]  ( .D(ereg_next[714]), .CLK(clk), .RST(rst), .I(
        e_init[1738]), .Q(ein[714]) );
  DFF \ereg_reg[715]  ( .D(ereg_next[715]), .CLK(clk), .RST(rst), .I(
        e_init[1739]), .Q(ein[715]) );
  DFF \ereg_reg[716]  ( .D(ereg_next[716]), .CLK(clk), .RST(rst), .I(
        e_init[1740]), .Q(ein[716]) );
  DFF \ereg_reg[717]  ( .D(ereg_next[717]), .CLK(clk), .RST(rst), .I(
        e_init[1741]), .Q(ein[717]) );
  DFF \ereg_reg[718]  ( .D(ereg_next[718]), .CLK(clk), .RST(rst), .I(
        e_init[1742]), .Q(ein[718]) );
  DFF \ereg_reg[719]  ( .D(ereg_next[719]), .CLK(clk), .RST(rst), .I(
        e_init[1743]), .Q(ein[719]) );
  DFF \ereg_reg[720]  ( .D(ereg_next[720]), .CLK(clk), .RST(rst), .I(
        e_init[1744]), .Q(ein[720]) );
  DFF \ereg_reg[721]  ( .D(ereg_next[721]), .CLK(clk), .RST(rst), .I(
        e_init[1745]), .Q(ein[721]) );
  DFF \ereg_reg[722]  ( .D(ereg_next[722]), .CLK(clk), .RST(rst), .I(
        e_init[1746]), .Q(ein[722]) );
  DFF \ereg_reg[723]  ( .D(ereg_next[723]), .CLK(clk), .RST(rst), .I(
        e_init[1747]), .Q(ein[723]) );
  DFF \ereg_reg[724]  ( .D(ereg_next[724]), .CLK(clk), .RST(rst), .I(
        e_init[1748]), .Q(ein[724]) );
  DFF \ereg_reg[725]  ( .D(ereg_next[725]), .CLK(clk), .RST(rst), .I(
        e_init[1749]), .Q(ein[725]) );
  DFF \ereg_reg[726]  ( .D(ereg_next[726]), .CLK(clk), .RST(rst), .I(
        e_init[1750]), .Q(ein[726]) );
  DFF \ereg_reg[727]  ( .D(ereg_next[727]), .CLK(clk), .RST(rst), .I(
        e_init[1751]), .Q(ein[727]) );
  DFF \ereg_reg[728]  ( .D(ereg_next[728]), .CLK(clk), .RST(rst), .I(
        e_init[1752]), .Q(ein[728]) );
  DFF \ereg_reg[729]  ( .D(ereg_next[729]), .CLK(clk), .RST(rst), .I(
        e_init[1753]), .Q(ein[729]) );
  DFF \ereg_reg[730]  ( .D(ereg_next[730]), .CLK(clk), .RST(rst), .I(
        e_init[1754]), .Q(ein[730]) );
  DFF \ereg_reg[731]  ( .D(ereg_next[731]), .CLK(clk), .RST(rst), .I(
        e_init[1755]), .Q(ein[731]) );
  DFF \ereg_reg[732]  ( .D(ereg_next[732]), .CLK(clk), .RST(rst), .I(
        e_init[1756]), .Q(ein[732]) );
  DFF \ereg_reg[733]  ( .D(ereg_next[733]), .CLK(clk), .RST(rst), .I(
        e_init[1757]), .Q(ein[733]) );
  DFF \ereg_reg[734]  ( .D(ereg_next[734]), .CLK(clk), .RST(rst), .I(
        e_init[1758]), .Q(ein[734]) );
  DFF \ereg_reg[735]  ( .D(ereg_next[735]), .CLK(clk), .RST(rst), .I(
        e_init[1759]), .Q(ein[735]) );
  DFF \ereg_reg[736]  ( .D(ereg_next[736]), .CLK(clk), .RST(rst), .I(
        e_init[1760]), .Q(ein[736]) );
  DFF \ereg_reg[737]  ( .D(ereg_next[737]), .CLK(clk), .RST(rst), .I(
        e_init[1761]), .Q(ein[737]) );
  DFF \ereg_reg[738]  ( .D(ereg_next[738]), .CLK(clk), .RST(rst), .I(
        e_init[1762]), .Q(ein[738]) );
  DFF \ereg_reg[739]  ( .D(ereg_next[739]), .CLK(clk), .RST(rst), .I(
        e_init[1763]), .Q(ein[739]) );
  DFF \ereg_reg[740]  ( .D(ereg_next[740]), .CLK(clk), .RST(rst), .I(
        e_init[1764]), .Q(ein[740]) );
  DFF \ereg_reg[741]  ( .D(ereg_next[741]), .CLK(clk), .RST(rst), .I(
        e_init[1765]), .Q(ein[741]) );
  DFF \ereg_reg[742]  ( .D(ereg_next[742]), .CLK(clk), .RST(rst), .I(
        e_init[1766]), .Q(ein[742]) );
  DFF \ereg_reg[743]  ( .D(ereg_next[743]), .CLK(clk), .RST(rst), .I(
        e_init[1767]), .Q(ein[743]) );
  DFF \ereg_reg[744]  ( .D(ereg_next[744]), .CLK(clk), .RST(rst), .I(
        e_init[1768]), .Q(ein[744]) );
  DFF \ereg_reg[745]  ( .D(ereg_next[745]), .CLK(clk), .RST(rst), .I(
        e_init[1769]), .Q(ein[745]) );
  DFF \ereg_reg[746]  ( .D(ereg_next[746]), .CLK(clk), .RST(rst), .I(
        e_init[1770]), .Q(ein[746]) );
  DFF \ereg_reg[747]  ( .D(ereg_next[747]), .CLK(clk), .RST(rst), .I(
        e_init[1771]), .Q(ein[747]) );
  DFF \ereg_reg[748]  ( .D(ereg_next[748]), .CLK(clk), .RST(rst), .I(
        e_init[1772]), .Q(ein[748]) );
  DFF \ereg_reg[749]  ( .D(ereg_next[749]), .CLK(clk), .RST(rst), .I(
        e_init[1773]), .Q(ein[749]) );
  DFF \ereg_reg[750]  ( .D(ereg_next[750]), .CLK(clk), .RST(rst), .I(
        e_init[1774]), .Q(ein[750]) );
  DFF \ereg_reg[751]  ( .D(ereg_next[751]), .CLK(clk), .RST(rst), .I(
        e_init[1775]), .Q(ein[751]) );
  DFF \ereg_reg[752]  ( .D(ereg_next[752]), .CLK(clk), .RST(rst), .I(
        e_init[1776]), .Q(ein[752]) );
  DFF \ereg_reg[753]  ( .D(ereg_next[753]), .CLK(clk), .RST(rst), .I(
        e_init[1777]), .Q(ein[753]) );
  DFF \ereg_reg[754]  ( .D(ereg_next[754]), .CLK(clk), .RST(rst), .I(
        e_init[1778]), .Q(ein[754]) );
  DFF \ereg_reg[755]  ( .D(ereg_next[755]), .CLK(clk), .RST(rst), .I(
        e_init[1779]), .Q(ein[755]) );
  DFF \ereg_reg[756]  ( .D(ereg_next[756]), .CLK(clk), .RST(rst), .I(
        e_init[1780]), .Q(ein[756]) );
  DFF \ereg_reg[757]  ( .D(ereg_next[757]), .CLK(clk), .RST(rst), .I(
        e_init[1781]), .Q(ein[757]) );
  DFF \ereg_reg[758]  ( .D(ereg_next[758]), .CLK(clk), .RST(rst), .I(
        e_init[1782]), .Q(ein[758]) );
  DFF \ereg_reg[759]  ( .D(ereg_next[759]), .CLK(clk), .RST(rst), .I(
        e_init[1783]), .Q(ein[759]) );
  DFF \ereg_reg[760]  ( .D(ereg_next[760]), .CLK(clk), .RST(rst), .I(
        e_init[1784]), .Q(ein[760]) );
  DFF \ereg_reg[761]  ( .D(ereg_next[761]), .CLK(clk), .RST(rst), .I(
        e_init[1785]), .Q(ein[761]) );
  DFF \ereg_reg[762]  ( .D(ereg_next[762]), .CLK(clk), .RST(rst), .I(
        e_init[1786]), .Q(ein[762]) );
  DFF \ereg_reg[763]  ( .D(ereg_next[763]), .CLK(clk), .RST(rst), .I(
        e_init[1787]), .Q(ein[763]) );
  DFF \ereg_reg[764]  ( .D(ereg_next[764]), .CLK(clk), .RST(rst), .I(
        e_init[1788]), .Q(ein[764]) );
  DFF \ereg_reg[765]  ( .D(ereg_next[765]), .CLK(clk), .RST(rst), .I(
        e_init[1789]), .Q(ein[765]) );
  DFF \ereg_reg[766]  ( .D(ereg_next[766]), .CLK(clk), .RST(rst), .I(
        e_init[1790]), .Q(ein[766]) );
  DFF \ereg_reg[767]  ( .D(ereg_next[767]), .CLK(clk), .RST(rst), .I(
        e_init[1791]), .Q(ein[767]) );
  DFF \ereg_reg[768]  ( .D(ereg_next[768]), .CLK(clk), .RST(rst), .I(
        e_init[1792]), .Q(ein[768]) );
  DFF \ereg_reg[769]  ( .D(ereg_next[769]), .CLK(clk), .RST(rst), .I(
        e_init[1793]), .Q(ein[769]) );
  DFF \ereg_reg[770]  ( .D(ereg_next[770]), .CLK(clk), .RST(rst), .I(
        e_init[1794]), .Q(ein[770]) );
  DFF \ereg_reg[771]  ( .D(ereg_next[771]), .CLK(clk), .RST(rst), .I(
        e_init[1795]), .Q(ein[771]) );
  DFF \ereg_reg[772]  ( .D(ereg_next[772]), .CLK(clk), .RST(rst), .I(
        e_init[1796]), .Q(ein[772]) );
  DFF \ereg_reg[773]  ( .D(ereg_next[773]), .CLK(clk), .RST(rst), .I(
        e_init[1797]), .Q(ein[773]) );
  DFF \ereg_reg[774]  ( .D(ereg_next[774]), .CLK(clk), .RST(rst), .I(
        e_init[1798]), .Q(ein[774]) );
  DFF \ereg_reg[775]  ( .D(ereg_next[775]), .CLK(clk), .RST(rst), .I(
        e_init[1799]), .Q(ein[775]) );
  DFF \ereg_reg[776]  ( .D(ereg_next[776]), .CLK(clk), .RST(rst), .I(
        e_init[1800]), .Q(ein[776]) );
  DFF \ereg_reg[777]  ( .D(ereg_next[777]), .CLK(clk), .RST(rst), .I(
        e_init[1801]), .Q(ein[777]) );
  DFF \ereg_reg[778]  ( .D(ereg_next[778]), .CLK(clk), .RST(rst), .I(
        e_init[1802]), .Q(ein[778]) );
  DFF \ereg_reg[779]  ( .D(ereg_next[779]), .CLK(clk), .RST(rst), .I(
        e_init[1803]), .Q(ein[779]) );
  DFF \ereg_reg[780]  ( .D(ereg_next[780]), .CLK(clk), .RST(rst), .I(
        e_init[1804]), .Q(ein[780]) );
  DFF \ereg_reg[781]  ( .D(ereg_next[781]), .CLK(clk), .RST(rst), .I(
        e_init[1805]), .Q(ein[781]) );
  DFF \ereg_reg[782]  ( .D(ereg_next[782]), .CLK(clk), .RST(rst), .I(
        e_init[1806]), .Q(ein[782]) );
  DFF \ereg_reg[783]  ( .D(ereg_next[783]), .CLK(clk), .RST(rst), .I(
        e_init[1807]), .Q(ein[783]) );
  DFF \ereg_reg[784]  ( .D(ereg_next[784]), .CLK(clk), .RST(rst), .I(
        e_init[1808]), .Q(ein[784]) );
  DFF \ereg_reg[785]  ( .D(ereg_next[785]), .CLK(clk), .RST(rst), .I(
        e_init[1809]), .Q(ein[785]) );
  DFF \ereg_reg[786]  ( .D(ereg_next[786]), .CLK(clk), .RST(rst), .I(
        e_init[1810]), .Q(ein[786]) );
  DFF \ereg_reg[787]  ( .D(ereg_next[787]), .CLK(clk), .RST(rst), .I(
        e_init[1811]), .Q(ein[787]) );
  DFF \ereg_reg[788]  ( .D(ereg_next[788]), .CLK(clk), .RST(rst), .I(
        e_init[1812]), .Q(ein[788]) );
  DFF \ereg_reg[789]  ( .D(ereg_next[789]), .CLK(clk), .RST(rst), .I(
        e_init[1813]), .Q(ein[789]) );
  DFF \ereg_reg[790]  ( .D(ereg_next[790]), .CLK(clk), .RST(rst), .I(
        e_init[1814]), .Q(ein[790]) );
  DFF \ereg_reg[791]  ( .D(ereg_next[791]), .CLK(clk), .RST(rst), .I(
        e_init[1815]), .Q(ein[791]) );
  DFF \ereg_reg[792]  ( .D(ereg_next[792]), .CLK(clk), .RST(rst), .I(
        e_init[1816]), .Q(ein[792]) );
  DFF \ereg_reg[793]  ( .D(ereg_next[793]), .CLK(clk), .RST(rst), .I(
        e_init[1817]), .Q(ein[793]) );
  DFF \ereg_reg[794]  ( .D(ereg_next[794]), .CLK(clk), .RST(rst), .I(
        e_init[1818]), .Q(ein[794]) );
  DFF \ereg_reg[795]  ( .D(ereg_next[795]), .CLK(clk), .RST(rst), .I(
        e_init[1819]), .Q(ein[795]) );
  DFF \ereg_reg[796]  ( .D(ereg_next[796]), .CLK(clk), .RST(rst), .I(
        e_init[1820]), .Q(ein[796]) );
  DFF \ereg_reg[797]  ( .D(ereg_next[797]), .CLK(clk), .RST(rst), .I(
        e_init[1821]), .Q(ein[797]) );
  DFF \ereg_reg[798]  ( .D(ereg_next[798]), .CLK(clk), .RST(rst), .I(
        e_init[1822]), .Q(ein[798]) );
  DFF \ereg_reg[799]  ( .D(ereg_next[799]), .CLK(clk), .RST(rst), .I(
        e_init[1823]), .Q(ein[799]) );
  DFF \ereg_reg[800]  ( .D(ereg_next[800]), .CLK(clk), .RST(rst), .I(
        e_init[1824]), .Q(ein[800]) );
  DFF \ereg_reg[801]  ( .D(ereg_next[801]), .CLK(clk), .RST(rst), .I(
        e_init[1825]), .Q(ein[801]) );
  DFF \ereg_reg[802]  ( .D(ereg_next[802]), .CLK(clk), .RST(rst), .I(
        e_init[1826]), .Q(ein[802]) );
  DFF \ereg_reg[803]  ( .D(ereg_next[803]), .CLK(clk), .RST(rst), .I(
        e_init[1827]), .Q(ein[803]) );
  DFF \ereg_reg[804]  ( .D(ereg_next[804]), .CLK(clk), .RST(rst), .I(
        e_init[1828]), .Q(ein[804]) );
  DFF \ereg_reg[805]  ( .D(ereg_next[805]), .CLK(clk), .RST(rst), .I(
        e_init[1829]), .Q(ein[805]) );
  DFF \ereg_reg[806]  ( .D(ereg_next[806]), .CLK(clk), .RST(rst), .I(
        e_init[1830]), .Q(ein[806]) );
  DFF \ereg_reg[807]  ( .D(ereg_next[807]), .CLK(clk), .RST(rst), .I(
        e_init[1831]), .Q(ein[807]) );
  DFF \ereg_reg[808]  ( .D(ereg_next[808]), .CLK(clk), .RST(rst), .I(
        e_init[1832]), .Q(ein[808]) );
  DFF \ereg_reg[809]  ( .D(ereg_next[809]), .CLK(clk), .RST(rst), .I(
        e_init[1833]), .Q(ein[809]) );
  DFF \ereg_reg[810]  ( .D(ereg_next[810]), .CLK(clk), .RST(rst), .I(
        e_init[1834]), .Q(ein[810]) );
  DFF \ereg_reg[811]  ( .D(ereg_next[811]), .CLK(clk), .RST(rst), .I(
        e_init[1835]), .Q(ein[811]) );
  DFF \ereg_reg[812]  ( .D(ereg_next[812]), .CLK(clk), .RST(rst), .I(
        e_init[1836]), .Q(ein[812]) );
  DFF \ereg_reg[813]  ( .D(ereg_next[813]), .CLK(clk), .RST(rst), .I(
        e_init[1837]), .Q(ein[813]) );
  DFF \ereg_reg[814]  ( .D(ereg_next[814]), .CLK(clk), .RST(rst), .I(
        e_init[1838]), .Q(ein[814]) );
  DFF \ereg_reg[815]  ( .D(ereg_next[815]), .CLK(clk), .RST(rst), .I(
        e_init[1839]), .Q(ein[815]) );
  DFF \ereg_reg[816]  ( .D(ereg_next[816]), .CLK(clk), .RST(rst), .I(
        e_init[1840]), .Q(ein[816]) );
  DFF \ereg_reg[817]  ( .D(ereg_next[817]), .CLK(clk), .RST(rst), .I(
        e_init[1841]), .Q(ein[817]) );
  DFF \ereg_reg[818]  ( .D(ereg_next[818]), .CLK(clk), .RST(rst), .I(
        e_init[1842]), .Q(ein[818]) );
  DFF \ereg_reg[819]  ( .D(ereg_next[819]), .CLK(clk), .RST(rst), .I(
        e_init[1843]), .Q(ein[819]) );
  DFF \ereg_reg[820]  ( .D(ereg_next[820]), .CLK(clk), .RST(rst), .I(
        e_init[1844]), .Q(ein[820]) );
  DFF \ereg_reg[821]  ( .D(ereg_next[821]), .CLK(clk), .RST(rst), .I(
        e_init[1845]), .Q(ein[821]) );
  DFF \ereg_reg[822]  ( .D(ereg_next[822]), .CLK(clk), .RST(rst), .I(
        e_init[1846]), .Q(ein[822]) );
  DFF \ereg_reg[823]  ( .D(ereg_next[823]), .CLK(clk), .RST(rst), .I(
        e_init[1847]), .Q(ein[823]) );
  DFF \ereg_reg[824]  ( .D(ereg_next[824]), .CLK(clk), .RST(rst), .I(
        e_init[1848]), .Q(ein[824]) );
  DFF \ereg_reg[825]  ( .D(ereg_next[825]), .CLK(clk), .RST(rst), .I(
        e_init[1849]), .Q(ein[825]) );
  DFF \ereg_reg[826]  ( .D(ereg_next[826]), .CLK(clk), .RST(rst), .I(
        e_init[1850]), .Q(ein[826]) );
  DFF \ereg_reg[827]  ( .D(ereg_next[827]), .CLK(clk), .RST(rst), .I(
        e_init[1851]), .Q(ein[827]) );
  DFF \ereg_reg[828]  ( .D(ereg_next[828]), .CLK(clk), .RST(rst), .I(
        e_init[1852]), .Q(ein[828]) );
  DFF \ereg_reg[829]  ( .D(ereg_next[829]), .CLK(clk), .RST(rst), .I(
        e_init[1853]), .Q(ein[829]) );
  DFF \ereg_reg[830]  ( .D(ereg_next[830]), .CLK(clk), .RST(rst), .I(
        e_init[1854]), .Q(ein[830]) );
  DFF \ereg_reg[831]  ( .D(ereg_next[831]), .CLK(clk), .RST(rst), .I(
        e_init[1855]), .Q(ein[831]) );
  DFF \ereg_reg[832]  ( .D(ereg_next[832]), .CLK(clk), .RST(rst), .I(
        e_init[1856]), .Q(ein[832]) );
  DFF \ereg_reg[833]  ( .D(ereg_next[833]), .CLK(clk), .RST(rst), .I(
        e_init[1857]), .Q(ein[833]) );
  DFF \ereg_reg[834]  ( .D(ereg_next[834]), .CLK(clk), .RST(rst), .I(
        e_init[1858]), .Q(ein[834]) );
  DFF \ereg_reg[835]  ( .D(ereg_next[835]), .CLK(clk), .RST(rst), .I(
        e_init[1859]), .Q(ein[835]) );
  DFF \ereg_reg[836]  ( .D(ereg_next[836]), .CLK(clk), .RST(rst), .I(
        e_init[1860]), .Q(ein[836]) );
  DFF \ereg_reg[837]  ( .D(ereg_next[837]), .CLK(clk), .RST(rst), .I(
        e_init[1861]), .Q(ein[837]) );
  DFF \ereg_reg[838]  ( .D(ereg_next[838]), .CLK(clk), .RST(rst), .I(
        e_init[1862]), .Q(ein[838]) );
  DFF \ereg_reg[839]  ( .D(ereg_next[839]), .CLK(clk), .RST(rst), .I(
        e_init[1863]), .Q(ein[839]) );
  DFF \ereg_reg[840]  ( .D(ereg_next[840]), .CLK(clk), .RST(rst), .I(
        e_init[1864]), .Q(ein[840]) );
  DFF \ereg_reg[841]  ( .D(ereg_next[841]), .CLK(clk), .RST(rst), .I(
        e_init[1865]), .Q(ein[841]) );
  DFF \ereg_reg[842]  ( .D(ereg_next[842]), .CLK(clk), .RST(rst), .I(
        e_init[1866]), .Q(ein[842]) );
  DFF \ereg_reg[843]  ( .D(ereg_next[843]), .CLK(clk), .RST(rst), .I(
        e_init[1867]), .Q(ein[843]) );
  DFF \ereg_reg[844]  ( .D(ereg_next[844]), .CLK(clk), .RST(rst), .I(
        e_init[1868]), .Q(ein[844]) );
  DFF \ereg_reg[845]  ( .D(ereg_next[845]), .CLK(clk), .RST(rst), .I(
        e_init[1869]), .Q(ein[845]) );
  DFF \ereg_reg[846]  ( .D(ereg_next[846]), .CLK(clk), .RST(rst), .I(
        e_init[1870]), .Q(ein[846]) );
  DFF \ereg_reg[847]  ( .D(ereg_next[847]), .CLK(clk), .RST(rst), .I(
        e_init[1871]), .Q(ein[847]) );
  DFF \ereg_reg[848]  ( .D(ereg_next[848]), .CLK(clk), .RST(rst), .I(
        e_init[1872]), .Q(ein[848]) );
  DFF \ereg_reg[849]  ( .D(ereg_next[849]), .CLK(clk), .RST(rst), .I(
        e_init[1873]), .Q(ein[849]) );
  DFF \ereg_reg[850]  ( .D(ereg_next[850]), .CLK(clk), .RST(rst), .I(
        e_init[1874]), .Q(ein[850]) );
  DFF \ereg_reg[851]  ( .D(ereg_next[851]), .CLK(clk), .RST(rst), .I(
        e_init[1875]), .Q(ein[851]) );
  DFF \ereg_reg[852]  ( .D(ereg_next[852]), .CLK(clk), .RST(rst), .I(
        e_init[1876]), .Q(ein[852]) );
  DFF \ereg_reg[853]  ( .D(ereg_next[853]), .CLK(clk), .RST(rst), .I(
        e_init[1877]), .Q(ein[853]) );
  DFF \ereg_reg[854]  ( .D(ereg_next[854]), .CLK(clk), .RST(rst), .I(
        e_init[1878]), .Q(ein[854]) );
  DFF \ereg_reg[855]  ( .D(ereg_next[855]), .CLK(clk), .RST(rst), .I(
        e_init[1879]), .Q(ein[855]) );
  DFF \ereg_reg[856]  ( .D(ereg_next[856]), .CLK(clk), .RST(rst), .I(
        e_init[1880]), .Q(ein[856]) );
  DFF \ereg_reg[857]  ( .D(ereg_next[857]), .CLK(clk), .RST(rst), .I(
        e_init[1881]), .Q(ein[857]) );
  DFF \ereg_reg[858]  ( .D(ereg_next[858]), .CLK(clk), .RST(rst), .I(
        e_init[1882]), .Q(ein[858]) );
  DFF \ereg_reg[859]  ( .D(ereg_next[859]), .CLK(clk), .RST(rst), .I(
        e_init[1883]), .Q(ein[859]) );
  DFF \ereg_reg[860]  ( .D(ereg_next[860]), .CLK(clk), .RST(rst), .I(
        e_init[1884]), .Q(ein[860]) );
  DFF \ereg_reg[861]  ( .D(ereg_next[861]), .CLK(clk), .RST(rst), .I(
        e_init[1885]), .Q(ein[861]) );
  DFF \ereg_reg[862]  ( .D(ereg_next[862]), .CLK(clk), .RST(rst), .I(
        e_init[1886]), .Q(ein[862]) );
  DFF \ereg_reg[863]  ( .D(ereg_next[863]), .CLK(clk), .RST(rst), .I(
        e_init[1887]), .Q(ein[863]) );
  DFF \ereg_reg[864]  ( .D(ereg_next[864]), .CLK(clk), .RST(rst), .I(
        e_init[1888]), .Q(ein[864]) );
  DFF \ereg_reg[865]  ( .D(ereg_next[865]), .CLK(clk), .RST(rst), .I(
        e_init[1889]), .Q(ein[865]) );
  DFF \ereg_reg[866]  ( .D(ereg_next[866]), .CLK(clk), .RST(rst), .I(
        e_init[1890]), .Q(ein[866]) );
  DFF \ereg_reg[867]  ( .D(ereg_next[867]), .CLK(clk), .RST(rst), .I(
        e_init[1891]), .Q(ein[867]) );
  DFF \ereg_reg[868]  ( .D(ereg_next[868]), .CLK(clk), .RST(rst), .I(
        e_init[1892]), .Q(ein[868]) );
  DFF \ereg_reg[869]  ( .D(ereg_next[869]), .CLK(clk), .RST(rst), .I(
        e_init[1893]), .Q(ein[869]) );
  DFF \ereg_reg[870]  ( .D(ereg_next[870]), .CLK(clk), .RST(rst), .I(
        e_init[1894]), .Q(ein[870]) );
  DFF \ereg_reg[871]  ( .D(ereg_next[871]), .CLK(clk), .RST(rst), .I(
        e_init[1895]), .Q(ein[871]) );
  DFF \ereg_reg[872]  ( .D(ereg_next[872]), .CLK(clk), .RST(rst), .I(
        e_init[1896]), .Q(ein[872]) );
  DFF \ereg_reg[873]  ( .D(ereg_next[873]), .CLK(clk), .RST(rst), .I(
        e_init[1897]), .Q(ein[873]) );
  DFF \ereg_reg[874]  ( .D(ereg_next[874]), .CLK(clk), .RST(rst), .I(
        e_init[1898]), .Q(ein[874]) );
  DFF \ereg_reg[875]  ( .D(ereg_next[875]), .CLK(clk), .RST(rst), .I(
        e_init[1899]), .Q(ein[875]) );
  DFF \ereg_reg[876]  ( .D(ereg_next[876]), .CLK(clk), .RST(rst), .I(
        e_init[1900]), .Q(ein[876]) );
  DFF \ereg_reg[877]  ( .D(ereg_next[877]), .CLK(clk), .RST(rst), .I(
        e_init[1901]), .Q(ein[877]) );
  DFF \ereg_reg[878]  ( .D(ereg_next[878]), .CLK(clk), .RST(rst), .I(
        e_init[1902]), .Q(ein[878]) );
  DFF \ereg_reg[879]  ( .D(ereg_next[879]), .CLK(clk), .RST(rst), .I(
        e_init[1903]), .Q(ein[879]) );
  DFF \ereg_reg[880]  ( .D(ereg_next[880]), .CLK(clk), .RST(rst), .I(
        e_init[1904]), .Q(ein[880]) );
  DFF \ereg_reg[881]  ( .D(ereg_next[881]), .CLK(clk), .RST(rst), .I(
        e_init[1905]), .Q(ein[881]) );
  DFF \ereg_reg[882]  ( .D(ereg_next[882]), .CLK(clk), .RST(rst), .I(
        e_init[1906]), .Q(ein[882]) );
  DFF \ereg_reg[883]  ( .D(ereg_next[883]), .CLK(clk), .RST(rst), .I(
        e_init[1907]), .Q(ein[883]) );
  DFF \ereg_reg[884]  ( .D(ereg_next[884]), .CLK(clk), .RST(rst), .I(
        e_init[1908]), .Q(ein[884]) );
  DFF \ereg_reg[885]  ( .D(ereg_next[885]), .CLK(clk), .RST(rst), .I(
        e_init[1909]), .Q(ein[885]) );
  DFF \ereg_reg[886]  ( .D(ereg_next[886]), .CLK(clk), .RST(rst), .I(
        e_init[1910]), .Q(ein[886]) );
  DFF \ereg_reg[887]  ( .D(ereg_next[887]), .CLK(clk), .RST(rst), .I(
        e_init[1911]), .Q(ein[887]) );
  DFF \ereg_reg[888]  ( .D(ereg_next[888]), .CLK(clk), .RST(rst), .I(
        e_init[1912]), .Q(ein[888]) );
  DFF \ereg_reg[889]  ( .D(ereg_next[889]), .CLK(clk), .RST(rst), .I(
        e_init[1913]), .Q(ein[889]) );
  DFF \ereg_reg[890]  ( .D(ereg_next[890]), .CLK(clk), .RST(rst), .I(
        e_init[1914]), .Q(ein[890]) );
  DFF \ereg_reg[891]  ( .D(ereg_next[891]), .CLK(clk), .RST(rst), .I(
        e_init[1915]), .Q(ein[891]) );
  DFF \ereg_reg[892]  ( .D(ereg_next[892]), .CLK(clk), .RST(rst), .I(
        e_init[1916]), .Q(ein[892]) );
  DFF \ereg_reg[893]  ( .D(ereg_next[893]), .CLK(clk), .RST(rst), .I(
        e_init[1917]), .Q(ein[893]) );
  DFF \ereg_reg[894]  ( .D(ereg_next[894]), .CLK(clk), .RST(rst), .I(
        e_init[1918]), .Q(ein[894]) );
  DFF \ereg_reg[895]  ( .D(ereg_next[895]), .CLK(clk), .RST(rst), .I(
        e_init[1919]), .Q(ein[895]) );
  DFF \ereg_reg[896]  ( .D(ereg_next[896]), .CLK(clk), .RST(rst), .I(
        e_init[1920]), .Q(ein[896]) );
  DFF \ereg_reg[897]  ( .D(ereg_next[897]), .CLK(clk), .RST(rst), .I(
        e_init[1921]), .Q(ein[897]) );
  DFF \ereg_reg[898]  ( .D(ereg_next[898]), .CLK(clk), .RST(rst), .I(
        e_init[1922]), .Q(ein[898]) );
  DFF \ereg_reg[899]  ( .D(ereg_next[899]), .CLK(clk), .RST(rst), .I(
        e_init[1923]), .Q(ein[899]) );
  DFF \ereg_reg[900]  ( .D(ereg_next[900]), .CLK(clk), .RST(rst), .I(
        e_init[1924]), .Q(ein[900]) );
  DFF \ereg_reg[901]  ( .D(ereg_next[901]), .CLK(clk), .RST(rst), .I(
        e_init[1925]), .Q(ein[901]) );
  DFF \ereg_reg[902]  ( .D(ereg_next[902]), .CLK(clk), .RST(rst), .I(
        e_init[1926]), .Q(ein[902]) );
  DFF \ereg_reg[903]  ( .D(ereg_next[903]), .CLK(clk), .RST(rst), .I(
        e_init[1927]), .Q(ein[903]) );
  DFF \ereg_reg[904]  ( .D(ereg_next[904]), .CLK(clk), .RST(rst), .I(
        e_init[1928]), .Q(ein[904]) );
  DFF \ereg_reg[905]  ( .D(ereg_next[905]), .CLK(clk), .RST(rst), .I(
        e_init[1929]), .Q(ein[905]) );
  DFF \ereg_reg[906]  ( .D(ereg_next[906]), .CLK(clk), .RST(rst), .I(
        e_init[1930]), .Q(ein[906]) );
  DFF \ereg_reg[907]  ( .D(ereg_next[907]), .CLK(clk), .RST(rst), .I(
        e_init[1931]), .Q(ein[907]) );
  DFF \ereg_reg[908]  ( .D(ereg_next[908]), .CLK(clk), .RST(rst), .I(
        e_init[1932]), .Q(ein[908]) );
  DFF \ereg_reg[909]  ( .D(ereg_next[909]), .CLK(clk), .RST(rst), .I(
        e_init[1933]), .Q(ein[909]) );
  DFF \ereg_reg[910]  ( .D(ereg_next[910]), .CLK(clk), .RST(rst), .I(
        e_init[1934]), .Q(ein[910]) );
  DFF \ereg_reg[911]  ( .D(ereg_next[911]), .CLK(clk), .RST(rst), .I(
        e_init[1935]), .Q(ein[911]) );
  DFF \ereg_reg[912]  ( .D(ereg_next[912]), .CLK(clk), .RST(rst), .I(
        e_init[1936]), .Q(ein[912]) );
  DFF \ereg_reg[913]  ( .D(ereg_next[913]), .CLK(clk), .RST(rst), .I(
        e_init[1937]), .Q(ein[913]) );
  DFF \ereg_reg[914]  ( .D(ereg_next[914]), .CLK(clk), .RST(rst), .I(
        e_init[1938]), .Q(ein[914]) );
  DFF \ereg_reg[915]  ( .D(ereg_next[915]), .CLK(clk), .RST(rst), .I(
        e_init[1939]), .Q(ein[915]) );
  DFF \ereg_reg[916]  ( .D(ereg_next[916]), .CLK(clk), .RST(rst), .I(
        e_init[1940]), .Q(ein[916]) );
  DFF \ereg_reg[917]  ( .D(ereg_next[917]), .CLK(clk), .RST(rst), .I(
        e_init[1941]), .Q(ein[917]) );
  DFF \ereg_reg[918]  ( .D(ereg_next[918]), .CLK(clk), .RST(rst), .I(
        e_init[1942]), .Q(ein[918]) );
  DFF \ereg_reg[919]  ( .D(ereg_next[919]), .CLK(clk), .RST(rst), .I(
        e_init[1943]), .Q(ein[919]) );
  DFF \ereg_reg[920]  ( .D(ereg_next[920]), .CLK(clk), .RST(rst), .I(
        e_init[1944]), .Q(ein[920]) );
  DFF \ereg_reg[921]  ( .D(ereg_next[921]), .CLK(clk), .RST(rst), .I(
        e_init[1945]), .Q(ein[921]) );
  DFF \ereg_reg[922]  ( .D(ereg_next[922]), .CLK(clk), .RST(rst), .I(
        e_init[1946]), .Q(ein[922]) );
  DFF \ereg_reg[923]  ( .D(ereg_next[923]), .CLK(clk), .RST(rst), .I(
        e_init[1947]), .Q(ein[923]) );
  DFF \ereg_reg[924]  ( .D(ereg_next[924]), .CLK(clk), .RST(rst), .I(
        e_init[1948]), .Q(ein[924]) );
  DFF \ereg_reg[925]  ( .D(ereg_next[925]), .CLK(clk), .RST(rst), .I(
        e_init[1949]), .Q(ein[925]) );
  DFF \ereg_reg[926]  ( .D(ereg_next[926]), .CLK(clk), .RST(rst), .I(
        e_init[1950]), .Q(ein[926]) );
  DFF \ereg_reg[927]  ( .D(ereg_next[927]), .CLK(clk), .RST(rst), .I(
        e_init[1951]), .Q(ein[927]) );
  DFF \ereg_reg[928]  ( .D(ereg_next[928]), .CLK(clk), .RST(rst), .I(
        e_init[1952]), .Q(ein[928]) );
  DFF \ereg_reg[929]  ( .D(ereg_next[929]), .CLK(clk), .RST(rst), .I(
        e_init[1953]), .Q(ein[929]) );
  DFF \ereg_reg[930]  ( .D(ereg_next[930]), .CLK(clk), .RST(rst), .I(
        e_init[1954]), .Q(ein[930]) );
  DFF \ereg_reg[931]  ( .D(ereg_next[931]), .CLK(clk), .RST(rst), .I(
        e_init[1955]), .Q(ein[931]) );
  DFF \ereg_reg[932]  ( .D(ereg_next[932]), .CLK(clk), .RST(rst), .I(
        e_init[1956]), .Q(ein[932]) );
  DFF \ereg_reg[933]  ( .D(ereg_next[933]), .CLK(clk), .RST(rst), .I(
        e_init[1957]), .Q(ein[933]) );
  DFF \ereg_reg[934]  ( .D(ereg_next[934]), .CLK(clk), .RST(rst), .I(
        e_init[1958]), .Q(ein[934]) );
  DFF \ereg_reg[935]  ( .D(ereg_next[935]), .CLK(clk), .RST(rst), .I(
        e_init[1959]), .Q(ein[935]) );
  DFF \ereg_reg[936]  ( .D(ereg_next[936]), .CLK(clk), .RST(rst), .I(
        e_init[1960]), .Q(ein[936]) );
  DFF \ereg_reg[937]  ( .D(ereg_next[937]), .CLK(clk), .RST(rst), .I(
        e_init[1961]), .Q(ein[937]) );
  DFF \ereg_reg[938]  ( .D(ereg_next[938]), .CLK(clk), .RST(rst), .I(
        e_init[1962]), .Q(ein[938]) );
  DFF \ereg_reg[939]  ( .D(ereg_next[939]), .CLK(clk), .RST(rst), .I(
        e_init[1963]), .Q(ein[939]) );
  DFF \ereg_reg[940]  ( .D(ereg_next[940]), .CLK(clk), .RST(rst), .I(
        e_init[1964]), .Q(ein[940]) );
  DFF \ereg_reg[941]  ( .D(ereg_next[941]), .CLK(clk), .RST(rst), .I(
        e_init[1965]), .Q(ein[941]) );
  DFF \ereg_reg[942]  ( .D(ereg_next[942]), .CLK(clk), .RST(rst), .I(
        e_init[1966]), .Q(ein[942]) );
  DFF \ereg_reg[943]  ( .D(ereg_next[943]), .CLK(clk), .RST(rst), .I(
        e_init[1967]), .Q(ein[943]) );
  DFF \ereg_reg[944]  ( .D(ereg_next[944]), .CLK(clk), .RST(rst), .I(
        e_init[1968]), .Q(ein[944]) );
  DFF \ereg_reg[945]  ( .D(ereg_next[945]), .CLK(clk), .RST(rst), .I(
        e_init[1969]), .Q(ein[945]) );
  DFF \ereg_reg[946]  ( .D(ereg_next[946]), .CLK(clk), .RST(rst), .I(
        e_init[1970]), .Q(ein[946]) );
  DFF \ereg_reg[947]  ( .D(ereg_next[947]), .CLK(clk), .RST(rst), .I(
        e_init[1971]), .Q(ein[947]) );
  DFF \ereg_reg[948]  ( .D(ereg_next[948]), .CLK(clk), .RST(rst), .I(
        e_init[1972]), .Q(ein[948]) );
  DFF \ereg_reg[949]  ( .D(ereg_next[949]), .CLK(clk), .RST(rst), .I(
        e_init[1973]), .Q(ein[949]) );
  DFF \ereg_reg[950]  ( .D(ereg_next[950]), .CLK(clk), .RST(rst), .I(
        e_init[1974]), .Q(ein[950]) );
  DFF \ereg_reg[951]  ( .D(ereg_next[951]), .CLK(clk), .RST(rst), .I(
        e_init[1975]), .Q(ein[951]) );
  DFF \ereg_reg[952]  ( .D(ereg_next[952]), .CLK(clk), .RST(rst), .I(
        e_init[1976]), .Q(ein[952]) );
  DFF \ereg_reg[953]  ( .D(ereg_next[953]), .CLK(clk), .RST(rst), .I(
        e_init[1977]), .Q(ein[953]) );
  DFF \ereg_reg[954]  ( .D(ereg_next[954]), .CLK(clk), .RST(rst), .I(
        e_init[1978]), .Q(ein[954]) );
  DFF \ereg_reg[955]  ( .D(ereg_next[955]), .CLK(clk), .RST(rst), .I(
        e_init[1979]), .Q(ein[955]) );
  DFF \ereg_reg[956]  ( .D(ereg_next[956]), .CLK(clk), .RST(rst), .I(
        e_init[1980]), .Q(ein[956]) );
  DFF \ereg_reg[957]  ( .D(ereg_next[957]), .CLK(clk), .RST(rst), .I(
        e_init[1981]), .Q(ein[957]) );
  DFF \ereg_reg[958]  ( .D(ereg_next[958]), .CLK(clk), .RST(rst), .I(
        e_init[1982]), .Q(ein[958]) );
  DFF \ereg_reg[959]  ( .D(ereg_next[959]), .CLK(clk), .RST(rst), .I(
        e_init[1983]), .Q(ein[959]) );
  DFF \ereg_reg[960]  ( .D(ereg_next[960]), .CLK(clk), .RST(rst), .I(
        e_init[1984]), .Q(ein[960]) );
  DFF \ereg_reg[961]  ( .D(ereg_next[961]), .CLK(clk), .RST(rst), .I(
        e_init[1985]), .Q(ein[961]) );
  DFF \ereg_reg[962]  ( .D(ereg_next[962]), .CLK(clk), .RST(rst), .I(
        e_init[1986]), .Q(ein[962]) );
  DFF \ereg_reg[963]  ( .D(ereg_next[963]), .CLK(clk), .RST(rst), .I(
        e_init[1987]), .Q(ein[963]) );
  DFF \ereg_reg[964]  ( .D(ereg_next[964]), .CLK(clk), .RST(rst), .I(
        e_init[1988]), .Q(ein[964]) );
  DFF \ereg_reg[965]  ( .D(ereg_next[965]), .CLK(clk), .RST(rst), .I(
        e_init[1989]), .Q(ein[965]) );
  DFF \ereg_reg[966]  ( .D(ereg_next[966]), .CLK(clk), .RST(rst), .I(
        e_init[1990]), .Q(ein[966]) );
  DFF \ereg_reg[967]  ( .D(ereg_next[967]), .CLK(clk), .RST(rst), .I(
        e_init[1991]), .Q(ein[967]) );
  DFF \ereg_reg[968]  ( .D(ereg_next[968]), .CLK(clk), .RST(rst), .I(
        e_init[1992]), .Q(ein[968]) );
  DFF \ereg_reg[969]  ( .D(ereg_next[969]), .CLK(clk), .RST(rst), .I(
        e_init[1993]), .Q(ein[969]) );
  DFF \ereg_reg[970]  ( .D(ereg_next[970]), .CLK(clk), .RST(rst), .I(
        e_init[1994]), .Q(ein[970]) );
  DFF \ereg_reg[971]  ( .D(ereg_next[971]), .CLK(clk), .RST(rst), .I(
        e_init[1995]), .Q(ein[971]) );
  DFF \ereg_reg[972]  ( .D(ereg_next[972]), .CLK(clk), .RST(rst), .I(
        e_init[1996]), .Q(ein[972]) );
  DFF \ereg_reg[973]  ( .D(ereg_next[973]), .CLK(clk), .RST(rst), .I(
        e_init[1997]), .Q(ein[973]) );
  DFF \ereg_reg[974]  ( .D(ereg_next[974]), .CLK(clk), .RST(rst), .I(
        e_init[1998]), .Q(ein[974]) );
  DFF \ereg_reg[975]  ( .D(ereg_next[975]), .CLK(clk), .RST(rst), .I(
        e_init[1999]), .Q(ein[975]) );
  DFF \ereg_reg[976]  ( .D(ereg_next[976]), .CLK(clk), .RST(rst), .I(
        e_init[2000]), .Q(ein[976]) );
  DFF \ereg_reg[977]  ( .D(ereg_next[977]), .CLK(clk), .RST(rst), .I(
        e_init[2001]), .Q(ein[977]) );
  DFF \ereg_reg[978]  ( .D(ereg_next[978]), .CLK(clk), .RST(rst), .I(
        e_init[2002]), .Q(ein[978]) );
  DFF \ereg_reg[979]  ( .D(ereg_next[979]), .CLK(clk), .RST(rst), .I(
        e_init[2003]), .Q(ein[979]) );
  DFF \ereg_reg[980]  ( .D(ereg_next[980]), .CLK(clk), .RST(rst), .I(
        e_init[2004]), .Q(ein[980]) );
  DFF \ereg_reg[981]  ( .D(ereg_next[981]), .CLK(clk), .RST(rst), .I(
        e_init[2005]), .Q(ein[981]) );
  DFF \ereg_reg[982]  ( .D(ereg_next[982]), .CLK(clk), .RST(rst), .I(
        e_init[2006]), .Q(ein[982]) );
  DFF \ereg_reg[983]  ( .D(ereg_next[983]), .CLK(clk), .RST(rst), .I(
        e_init[2007]), .Q(ein[983]) );
  DFF \ereg_reg[984]  ( .D(ereg_next[984]), .CLK(clk), .RST(rst), .I(
        e_init[2008]), .Q(ein[984]) );
  DFF \ereg_reg[985]  ( .D(ereg_next[985]), .CLK(clk), .RST(rst), .I(
        e_init[2009]), .Q(ein[985]) );
  DFF \ereg_reg[986]  ( .D(ereg_next[986]), .CLK(clk), .RST(rst), .I(
        e_init[2010]), .Q(ein[986]) );
  DFF \ereg_reg[987]  ( .D(ereg_next[987]), .CLK(clk), .RST(rst), .I(
        e_init[2011]), .Q(ein[987]) );
  DFF \ereg_reg[988]  ( .D(ereg_next[988]), .CLK(clk), .RST(rst), .I(
        e_init[2012]), .Q(ein[988]) );
  DFF \ereg_reg[989]  ( .D(ereg_next[989]), .CLK(clk), .RST(rst), .I(
        e_init[2013]), .Q(ein[989]) );
  DFF \ereg_reg[990]  ( .D(ereg_next[990]), .CLK(clk), .RST(rst), .I(
        e_init[2014]), .Q(ein[990]) );
  DFF \ereg_reg[991]  ( .D(ereg_next[991]), .CLK(clk), .RST(rst), .I(
        e_init[2015]), .Q(ein[991]) );
  DFF \ereg_reg[992]  ( .D(ereg_next[992]), .CLK(clk), .RST(rst), .I(
        e_init[2016]), .Q(ein[992]) );
  DFF \ereg_reg[993]  ( .D(ereg_next[993]), .CLK(clk), .RST(rst), .I(
        e_init[2017]), .Q(ein[993]) );
  DFF \ereg_reg[994]  ( .D(ereg_next[994]), .CLK(clk), .RST(rst), .I(
        e_init[2018]), .Q(ein[994]) );
  DFF \ereg_reg[995]  ( .D(ereg_next[995]), .CLK(clk), .RST(rst), .I(
        e_init[2019]), .Q(ein[995]) );
  DFF \ereg_reg[996]  ( .D(ereg_next[996]), .CLK(clk), .RST(rst), .I(
        e_init[2020]), .Q(ein[996]) );
  DFF \ereg_reg[997]  ( .D(ereg_next[997]), .CLK(clk), .RST(rst), .I(
        e_init[2021]), .Q(ein[997]) );
  DFF \ereg_reg[998]  ( .D(ereg_next[998]), .CLK(clk), .RST(rst), .I(
        e_init[2022]), .Q(ein[998]) );
  DFF \ereg_reg[999]  ( .D(ereg_next[999]), .CLK(clk), .RST(rst), .I(
        e_init[2023]), .Q(ein[999]) );
  DFF \ereg_reg[1000]  ( .D(ereg_next[1000]), .CLK(clk), .RST(rst), .I(
        e_init[2024]), .Q(ein[1000]) );
  DFF \ereg_reg[1001]  ( .D(ereg_next[1001]), .CLK(clk), .RST(rst), .I(
        e_init[2025]), .Q(ein[1001]) );
  DFF \ereg_reg[1002]  ( .D(ereg_next[1002]), .CLK(clk), .RST(rst), .I(
        e_init[2026]), .Q(ein[1002]) );
  DFF \ereg_reg[1003]  ( .D(ereg_next[1003]), .CLK(clk), .RST(rst), .I(
        e_init[2027]), .Q(ein[1003]) );
  DFF \ereg_reg[1004]  ( .D(ereg_next[1004]), .CLK(clk), .RST(rst), .I(
        e_init[2028]), .Q(ein[1004]) );
  DFF \ereg_reg[1005]  ( .D(ereg_next[1005]), .CLK(clk), .RST(rst), .I(
        e_init[2029]), .Q(ein[1005]) );
  DFF \ereg_reg[1006]  ( .D(ereg_next[1006]), .CLK(clk), .RST(rst), .I(
        e_init[2030]), .Q(ein[1006]) );
  DFF \ereg_reg[1007]  ( .D(ereg_next[1007]), .CLK(clk), .RST(rst), .I(
        e_init[2031]), .Q(ein[1007]) );
  DFF \ereg_reg[1008]  ( .D(ereg_next[1008]), .CLK(clk), .RST(rst), .I(
        e_init[2032]), .Q(ein[1008]) );
  DFF \ereg_reg[1009]  ( .D(ereg_next[1009]), .CLK(clk), .RST(rst), .I(
        e_init[2033]), .Q(ein[1009]) );
  DFF \ereg_reg[1010]  ( .D(ereg_next[1010]), .CLK(clk), .RST(rst), .I(
        e_init[2034]), .Q(ein[1010]) );
  DFF \ereg_reg[1011]  ( .D(ereg_next[1011]), .CLK(clk), .RST(rst), .I(
        e_init[2035]), .Q(ein[1011]) );
  DFF \ereg_reg[1012]  ( .D(ereg_next[1012]), .CLK(clk), .RST(rst), .I(
        e_init[2036]), .Q(ein[1012]) );
  DFF \ereg_reg[1013]  ( .D(ereg_next[1013]), .CLK(clk), .RST(rst), .I(
        e_init[2037]), .Q(ein[1013]) );
  DFF \ereg_reg[1014]  ( .D(ereg_next[1014]), .CLK(clk), .RST(rst), .I(
        e_init[2038]), .Q(ein[1014]) );
  DFF \ereg_reg[1015]  ( .D(ereg_next[1015]), .CLK(clk), .RST(rst), .I(
        e_init[2039]), .Q(ein[1015]) );
  DFF \ereg_reg[1016]  ( .D(ereg_next[1016]), .CLK(clk), .RST(rst), .I(
        e_init[2040]), .Q(ein[1016]) );
  DFF \ereg_reg[1017]  ( .D(ereg_next[1017]), .CLK(clk), .RST(rst), .I(
        e_init[2041]), .Q(ein[1017]) );
  DFF \ereg_reg[1018]  ( .D(ereg_next[1018]), .CLK(clk), .RST(rst), .I(
        e_init[2042]), .Q(ein[1018]) );
  DFF \ereg_reg[1019]  ( .D(ereg_next[1019]), .CLK(clk), .RST(rst), .I(
        e_init[2043]), .Q(ein[1019]) );
  DFF \ereg_reg[1020]  ( .D(ereg_next[1020]), .CLK(clk), .RST(rst), .I(
        e_init[2044]), .Q(ein[1020]) );
  DFF \ereg_reg[1021]  ( .D(ereg_next[1021]), .CLK(clk), .RST(rst), .I(
        e_init[2045]), .Q(ein[1021]) );
  DFF \ereg_reg[1022]  ( .D(ereg_next[1022]), .CLK(clk), .RST(rst), .I(
        e_init[2046]), .Q(ein[1022]) );
  DFF \ereg_reg[1023]  ( .D(ereg_next[1023]), .CLK(clk), .RST(rst), .I(
        e_init[2047]), .Q(ein[1023]) );
  DFF first_one_reg ( .D(n6), .CLK(clk), .RST(rst), .I(1'b0), .Q(first_one) );
  DFF \mreg_reg[1023]  ( .D(mreg[1023]), .CLK(clk), .RST(rst), .I(g_init[1023]), .Q(mreg[1023]) );
  DFF \mreg_reg[1022]  ( .D(mreg[1022]), .CLK(clk), .RST(rst), .I(g_init[1022]), .Q(mreg[1022]) );
  DFF \mreg_reg[1021]  ( .D(mreg[1021]), .CLK(clk), .RST(rst), .I(g_init[1021]), .Q(mreg[1021]) );
  DFF \mreg_reg[1020]  ( .D(mreg[1020]), .CLK(clk), .RST(rst), .I(g_init[1020]), .Q(mreg[1020]) );
  DFF \mreg_reg[1019]  ( .D(mreg[1019]), .CLK(clk), .RST(rst), .I(g_init[1019]), .Q(mreg[1019]) );
  DFF \mreg_reg[1018]  ( .D(mreg[1018]), .CLK(clk), .RST(rst), .I(g_init[1018]), .Q(mreg[1018]) );
  DFF \mreg_reg[1017]  ( .D(mreg[1017]), .CLK(clk), .RST(rst), .I(g_init[1017]), .Q(mreg[1017]) );
  DFF \mreg_reg[1016]  ( .D(mreg[1016]), .CLK(clk), .RST(rst), .I(g_init[1016]), .Q(mreg[1016]) );
  DFF \mreg_reg[1015]  ( .D(mreg[1015]), .CLK(clk), .RST(rst), .I(g_init[1015]), .Q(mreg[1015]) );
  DFF \mreg_reg[1014]  ( .D(mreg[1014]), .CLK(clk), .RST(rst), .I(g_init[1014]), .Q(mreg[1014]) );
  DFF \mreg_reg[1013]  ( .D(mreg[1013]), .CLK(clk), .RST(rst), .I(g_init[1013]), .Q(mreg[1013]) );
  DFF \mreg_reg[1012]  ( .D(mreg[1012]), .CLK(clk), .RST(rst), .I(g_init[1012]), .Q(mreg[1012]) );
  DFF \mreg_reg[1011]  ( .D(mreg[1011]), .CLK(clk), .RST(rst), .I(g_init[1011]), .Q(mreg[1011]) );
  DFF \mreg_reg[1010]  ( .D(mreg[1010]), .CLK(clk), .RST(rst), .I(g_init[1010]), .Q(mreg[1010]) );
  DFF \mreg_reg[1009]  ( .D(mreg[1009]), .CLK(clk), .RST(rst), .I(g_init[1009]), .Q(mreg[1009]) );
  DFF \mreg_reg[1008]  ( .D(mreg[1008]), .CLK(clk), .RST(rst), .I(g_init[1008]), .Q(mreg[1008]) );
  DFF \mreg_reg[1007]  ( .D(mreg[1007]), .CLK(clk), .RST(rst), .I(g_init[1007]), .Q(mreg[1007]) );
  DFF \mreg_reg[1006]  ( .D(mreg[1006]), .CLK(clk), .RST(rst), .I(g_init[1006]), .Q(mreg[1006]) );
  DFF \mreg_reg[1005]  ( .D(mreg[1005]), .CLK(clk), .RST(rst), .I(g_init[1005]), .Q(mreg[1005]) );
  DFF \mreg_reg[1004]  ( .D(mreg[1004]), .CLK(clk), .RST(rst), .I(g_init[1004]), .Q(mreg[1004]) );
  DFF \mreg_reg[1003]  ( .D(mreg[1003]), .CLK(clk), .RST(rst), .I(g_init[1003]), .Q(mreg[1003]) );
  DFF \mreg_reg[1002]  ( .D(mreg[1002]), .CLK(clk), .RST(rst), .I(g_init[1002]), .Q(mreg[1002]) );
  DFF \mreg_reg[1001]  ( .D(mreg[1001]), .CLK(clk), .RST(rst), .I(g_init[1001]), .Q(mreg[1001]) );
  DFF \mreg_reg[1000]  ( .D(mreg[1000]), .CLK(clk), .RST(rst), .I(g_init[1000]), .Q(mreg[1000]) );
  DFF \mreg_reg[999]  ( .D(mreg[999]), .CLK(clk), .RST(rst), .I(g_init[999]), 
        .Q(mreg[999]) );
  DFF \mreg_reg[998]  ( .D(mreg[998]), .CLK(clk), .RST(rst), .I(g_init[998]), 
        .Q(mreg[998]) );
  DFF \mreg_reg[997]  ( .D(mreg[997]), .CLK(clk), .RST(rst), .I(g_init[997]), 
        .Q(mreg[997]) );
  DFF \mreg_reg[996]  ( .D(mreg[996]), .CLK(clk), .RST(rst), .I(g_init[996]), 
        .Q(mreg[996]) );
  DFF \mreg_reg[995]  ( .D(mreg[995]), .CLK(clk), .RST(rst), .I(g_init[995]), 
        .Q(mreg[995]) );
  DFF \mreg_reg[994]  ( .D(mreg[994]), .CLK(clk), .RST(rst), .I(g_init[994]), 
        .Q(mreg[994]) );
  DFF \mreg_reg[993]  ( .D(mreg[993]), .CLK(clk), .RST(rst), .I(g_init[993]), 
        .Q(mreg[993]) );
  DFF \mreg_reg[992]  ( .D(mreg[992]), .CLK(clk), .RST(rst), .I(g_init[992]), 
        .Q(mreg[992]) );
  DFF \mreg_reg[991]  ( .D(mreg[991]), .CLK(clk), .RST(rst), .I(g_init[991]), 
        .Q(mreg[991]) );
  DFF \mreg_reg[990]  ( .D(mreg[990]), .CLK(clk), .RST(rst), .I(g_init[990]), 
        .Q(mreg[990]) );
  DFF \mreg_reg[989]  ( .D(mreg[989]), .CLK(clk), .RST(rst), .I(g_init[989]), 
        .Q(mreg[989]) );
  DFF \mreg_reg[988]  ( .D(mreg[988]), .CLK(clk), .RST(rst), .I(g_init[988]), 
        .Q(mreg[988]) );
  DFF \mreg_reg[987]  ( .D(mreg[987]), .CLK(clk), .RST(rst), .I(g_init[987]), 
        .Q(mreg[987]) );
  DFF \mreg_reg[986]  ( .D(mreg[986]), .CLK(clk), .RST(rst), .I(g_init[986]), 
        .Q(mreg[986]) );
  DFF \mreg_reg[985]  ( .D(mreg[985]), .CLK(clk), .RST(rst), .I(g_init[985]), 
        .Q(mreg[985]) );
  DFF \mreg_reg[984]  ( .D(mreg[984]), .CLK(clk), .RST(rst), .I(g_init[984]), 
        .Q(mreg[984]) );
  DFF \mreg_reg[983]  ( .D(mreg[983]), .CLK(clk), .RST(rst), .I(g_init[983]), 
        .Q(mreg[983]) );
  DFF \mreg_reg[982]  ( .D(mreg[982]), .CLK(clk), .RST(rst), .I(g_init[982]), 
        .Q(mreg[982]) );
  DFF \mreg_reg[981]  ( .D(mreg[981]), .CLK(clk), .RST(rst), .I(g_init[981]), 
        .Q(mreg[981]) );
  DFF \mreg_reg[980]  ( .D(mreg[980]), .CLK(clk), .RST(rst), .I(g_init[980]), 
        .Q(mreg[980]) );
  DFF \mreg_reg[979]  ( .D(mreg[979]), .CLK(clk), .RST(rst), .I(g_init[979]), 
        .Q(mreg[979]) );
  DFF \mreg_reg[978]  ( .D(mreg[978]), .CLK(clk), .RST(rst), .I(g_init[978]), 
        .Q(mreg[978]) );
  DFF \mreg_reg[977]  ( .D(mreg[977]), .CLK(clk), .RST(rst), .I(g_init[977]), 
        .Q(mreg[977]) );
  DFF \mreg_reg[976]  ( .D(mreg[976]), .CLK(clk), .RST(rst), .I(g_init[976]), 
        .Q(mreg[976]) );
  DFF \mreg_reg[975]  ( .D(mreg[975]), .CLK(clk), .RST(rst), .I(g_init[975]), 
        .Q(mreg[975]) );
  DFF \mreg_reg[974]  ( .D(mreg[974]), .CLK(clk), .RST(rst), .I(g_init[974]), 
        .Q(mreg[974]) );
  DFF \mreg_reg[973]  ( .D(mreg[973]), .CLK(clk), .RST(rst), .I(g_init[973]), 
        .Q(mreg[973]) );
  DFF \mreg_reg[972]  ( .D(mreg[972]), .CLK(clk), .RST(rst), .I(g_init[972]), 
        .Q(mreg[972]) );
  DFF \mreg_reg[971]  ( .D(mreg[971]), .CLK(clk), .RST(rst), .I(g_init[971]), 
        .Q(mreg[971]) );
  DFF \mreg_reg[970]  ( .D(mreg[970]), .CLK(clk), .RST(rst), .I(g_init[970]), 
        .Q(mreg[970]) );
  DFF \mreg_reg[969]  ( .D(mreg[969]), .CLK(clk), .RST(rst), .I(g_init[969]), 
        .Q(mreg[969]) );
  DFF \mreg_reg[968]  ( .D(mreg[968]), .CLK(clk), .RST(rst), .I(g_init[968]), 
        .Q(mreg[968]) );
  DFF \mreg_reg[967]  ( .D(mreg[967]), .CLK(clk), .RST(rst), .I(g_init[967]), 
        .Q(mreg[967]) );
  DFF \mreg_reg[966]  ( .D(mreg[966]), .CLK(clk), .RST(rst), .I(g_init[966]), 
        .Q(mreg[966]) );
  DFF \mreg_reg[965]  ( .D(mreg[965]), .CLK(clk), .RST(rst), .I(g_init[965]), 
        .Q(mreg[965]) );
  DFF \mreg_reg[964]  ( .D(mreg[964]), .CLK(clk), .RST(rst), .I(g_init[964]), 
        .Q(mreg[964]) );
  DFF \mreg_reg[963]  ( .D(mreg[963]), .CLK(clk), .RST(rst), .I(g_init[963]), 
        .Q(mreg[963]) );
  DFF \mreg_reg[962]  ( .D(mreg[962]), .CLK(clk), .RST(rst), .I(g_init[962]), 
        .Q(mreg[962]) );
  DFF \mreg_reg[961]  ( .D(mreg[961]), .CLK(clk), .RST(rst), .I(g_init[961]), 
        .Q(mreg[961]) );
  DFF \mreg_reg[960]  ( .D(mreg[960]), .CLK(clk), .RST(rst), .I(g_init[960]), 
        .Q(mreg[960]) );
  DFF \mreg_reg[959]  ( .D(mreg[959]), .CLK(clk), .RST(rst), .I(g_init[959]), 
        .Q(mreg[959]) );
  DFF \mreg_reg[958]  ( .D(mreg[958]), .CLK(clk), .RST(rst), .I(g_init[958]), 
        .Q(mreg[958]) );
  DFF \mreg_reg[957]  ( .D(mreg[957]), .CLK(clk), .RST(rst), .I(g_init[957]), 
        .Q(mreg[957]) );
  DFF \mreg_reg[956]  ( .D(mreg[956]), .CLK(clk), .RST(rst), .I(g_init[956]), 
        .Q(mreg[956]) );
  DFF \mreg_reg[955]  ( .D(mreg[955]), .CLK(clk), .RST(rst), .I(g_init[955]), 
        .Q(mreg[955]) );
  DFF \mreg_reg[954]  ( .D(mreg[954]), .CLK(clk), .RST(rst), .I(g_init[954]), 
        .Q(mreg[954]) );
  DFF \mreg_reg[953]  ( .D(mreg[953]), .CLK(clk), .RST(rst), .I(g_init[953]), 
        .Q(mreg[953]) );
  DFF \mreg_reg[952]  ( .D(mreg[952]), .CLK(clk), .RST(rst), .I(g_init[952]), 
        .Q(mreg[952]) );
  DFF \mreg_reg[951]  ( .D(mreg[951]), .CLK(clk), .RST(rst), .I(g_init[951]), 
        .Q(mreg[951]) );
  DFF \mreg_reg[950]  ( .D(mreg[950]), .CLK(clk), .RST(rst), .I(g_init[950]), 
        .Q(mreg[950]) );
  DFF \mreg_reg[949]  ( .D(mreg[949]), .CLK(clk), .RST(rst), .I(g_init[949]), 
        .Q(mreg[949]) );
  DFF \mreg_reg[948]  ( .D(mreg[948]), .CLK(clk), .RST(rst), .I(g_init[948]), 
        .Q(mreg[948]) );
  DFF \mreg_reg[947]  ( .D(mreg[947]), .CLK(clk), .RST(rst), .I(g_init[947]), 
        .Q(mreg[947]) );
  DFF \mreg_reg[946]  ( .D(mreg[946]), .CLK(clk), .RST(rst), .I(g_init[946]), 
        .Q(mreg[946]) );
  DFF \mreg_reg[945]  ( .D(mreg[945]), .CLK(clk), .RST(rst), .I(g_init[945]), 
        .Q(mreg[945]) );
  DFF \mreg_reg[944]  ( .D(mreg[944]), .CLK(clk), .RST(rst), .I(g_init[944]), 
        .Q(mreg[944]) );
  DFF \mreg_reg[943]  ( .D(mreg[943]), .CLK(clk), .RST(rst), .I(g_init[943]), 
        .Q(mreg[943]) );
  DFF \mreg_reg[942]  ( .D(mreg[942]), .CLK(clk), .RST(rst), .I(g_init[942]), 
        .Q(mreg[942]) );
  DFF \mreg_reg[941]  ( .D(mreg[941]), .CLK(clk), .RST(rst), .I(g_init[941]), 
        .Q(mreg[941]) );
  DFF \mreg_reg[940]  ( .D(mreg[940]), .CLK(clk), .RST(rst), .I(g_init[940]), 
        .Q(mreg[940]) );
  DFF \mreg_reg[939]  ( .D(mreg[939]), .CLK(clk), .RST(rst), .I(g_init[939]), 
        .Q(mreg[939]) );
  DFF \mreg_reg[938]  ( .D(mreg[938]), .CLK(clk), .RST(rst), .I(g_init[938]), 
        .Q(mreg[938]) );
  DFF \mreg_reg[937]  ( .D(mreg[937]), .CLK(clk), .RST(rst), .I(g_init[937]), 
        .Q(mreg[937]) );
  DFF \mreg_reg[936]  ( .D(mreg[936]), .CLK(clk), .RST(rst), .I(g_init[936]), 
        .Q(mreg[936]) );
  DFF \mreg_reg[935]  ( .D(mreg[935]), .CLK(clk), .RST(rst), .I(g_init[935]), 
        .Q(mreg[935]) );
  DFF \mreg_reg[934]  ( .D(mreg[934]), .CLK(clk), .RST(rst), .I(g_init[934]), 
        .Q(mreg[934]) );
  DFF \mreg_reg[933]  ( .D(mreg[933]), .CLK(clk), .RST(rst), .I(g_init[933]), 
        .Q(mreg[933]) );
  DFF \mreg_reg[932]  ( .D(mreg[932]), .CLK(clk), .RST(rst), .I(g_init[932]), 
        .Q(mreg[932]) );
  DFF \mreg_reg[931]  ( .D(mreg[931]), .CLK(clk), .RST(rst), .I(g_init[931]), 
        .Q(mreg[931]) );
  DFF \mreg_reg[930]  ( .D(mreg[930]), .CLK(clk), .RST(rst), .I(g_init[930]), 
        .Q(mreg[930]) );
  DFF \mreg_reg[929]  ( .D(mreg[929]), .CLK(clk), .RST(rst), .I(g_init[929]), 
        .Q(mreg[929]) );
  DFF \mreg_reg[928]  ( .D(mreg[928]), .CLK(clk), .RST(rst), .I(g_init[928]), 
        .Q(mreg[928]) );
  DFF \mreg_reg[927]  ( .D(mreg[927]), .CLK(clk), .RST(rst), .I(g_init[927]), 
        .Q(mreg[927]) );
  DFF \mreg_reg[926]  ( .D(mreg[926]), .CLK(clk), .RST(rst), .I(g_init[926]), 
        .Q(mreg[926]) );
  DFF \mreg_reg[925]  ( .D(mreg[925]), .CLK(clk), .RST(rst), .I(g_init[925]), 
        .Q(mreg[925]) );
  DFF \mreg_reg[924]  ( .D(mreg[924]), .CLK(clk), .RST(rst), .I(g_init[924]), 
        .Q(mreg[924]) );
  DFF \mreg_reg[923]  ( .D(mreg[923]), .CLK(clk), .RST(rst), .I(g_init[923]), 
        .Q(mreg[923]) );
  DFF \mreg_reg[922]  ( .D(mreg[922]), .CLK(clk), .RST(rst), .I(g_init[922]), 
        .Q(mreg[922]) );
  DFF \mreg_reg[921]  ( .D(mreg[921]), .CLK(clk), .RST(rst), .I(g_init[921]), 
        .Q(mreg[921]) );
  DFF \mreg_reg[920]  ( .D(mreg[920]), .CLK(clk), .RST(rst), .I(g_init[920]), 
        .Q(mreg[920]) );
  DFF \mreg_reg[919]  ( .D(mreg[919]), .CLK(clk), .RST(rst), .I(g_init[919]), 
        .Q(mreg[919]) );
  DFF \mreg_reg[918]  ( .D(mreg[918]), .CLK(clk), .RST(rst), .I(g_init[918]), 
        .Q(mreg[918]) );
  DFF \mreg_reg[917]  ( .D(mreg[917]), .CLK(clk), .RST(rst), .I(g_init[917]), 
        .Q(mreg[917]) );
  DFF \mreg_reg[916]  ( .D(mreg[916]), .CLK(clk), .RST(rst), .I(g_init[916]), 
        .Q(mreg[916]) );
  DFF \mreg_reg[915]  ( .D(mreg[915]), .CLK(clk), .RST(rst), .I(g_init[915]), 
        .Q(mreg[915]) );
  DFF \mreg_reg[914]  ( .D(mreg[914]), .CLK(clk), .RST(rst), .I(g_init[914]), 
        .Q(mreg[914]) );
  DFF \mreg_reg[913]  ( .D(mreg[913]), .CLK(clk), .RST(rst), .I(g_init[913]), 
        .Q(mreg[913]) );
  DFF \mreg_reg[912]  ( .D(mreg[912]), .CLK(clk), .RST(rst), .I(g_init[912]), 
        .Q(mreg[912]) );
  DFF \mreg_reg[911]  ( .D(mreg[911]), .CLK(clk), .RST(rst), .I(g_init[911]), 
        .Q(mreg[911]) );
  DFF \mreg_reg[910]  ( .D(mreg[910]), .CLK(clk), .RST(rst), .I(g_init[910]), 
        .Q(mreg[910]) );
  DFF \mreg_reg[909]  ( .D(mreg[909]), .CLK(clk), .RST(rst), .I(g_init[909]), 
        .Q(mreg[909]) );
  DFF \mreg_reg[908]  ( .D(mreg[908]), .CLK(clk), .RST(rst), .I(g_init[908]), 
        .Q(mreg[908]) );
  DFF \mreg_reg[907]  ( .D(mreg[907]), .CLK(clk), .RST(rst), .I(g_init[907]), 
        .Q(mreg[907]) );
  DFF \mreg_reg[906]  ( .D(mreg[906]), .CLK(clk), .RST(rst), .I(g_init[906]), 
        .Q(mreg[906]) );
  DFF \mreg_reg[905]  ( .D(mreg[905]), .CLK(clk), .RST(rst), .I(g_init[905]), 
        .Q(mreg[905]) );
  DFF \mreg_reg[904]  ( .D(mreg[904]), .CLK(clk), .RST(rst), .I(g_init[904]), 
        .Q(mreg[904]) );
  DFF \mreg_reg[903]  ( .D(mreg[903]), .CLK(clk), .RST(rst), .I(g_init[903]), 
        .Q(mreg[903]) );
  DFF \mreg_reg[902]  ( .D(mreg[902]), .CLK(clk), .RST(rst), .I(g_init[902]), 
        .Q(mreg[902]) );
  DFF \mreg_reg[901]  ( .D(mreg[901]), .CLK(clk), .RST(rst), .I(g_init[901]), 
        .Q(mreg[901]) );
  DFF \mreg_reg[900]  ( .D(mreg[900]), .CLK(clk), .RST(rst), .I(g_init[900]), 
        .Q(mreg[900]) );
  DFF \mreg_reg[899]  ( .D(mreg[899]), .CLK(clk), .RST(rst), .I(g_init[899]), 
        .Q(mreg[899]) );
  DFF \mreg_reg[898]  ( .D(mreg[898]), .CLK(clk), .RST(rst), .I(g_init[898]), 
        .Q(mreg[898]) );
  DFF \mreg_reg[897]  ( .D(mreg[897]), .CLK(clk), .RST(rst), .I(g_init[897]), 
        .Q(mreg[897]) );
  DFF \mreg_reg[896]  ( .D(mreg[896]), .CLK(clk), .RST(rst), .I(g_init[896]), 
        .Q(mreg[896]) );
  DFF \mreg_reg[895]  ( .D(mreg[895]), .CLK(clk), .RST(rst), .I(g_init[895]), 
        .Q(mreg[895]) );
  DFF \mreg_reg[894]  ( .D(mreg[894]), .CLK(clk), .RST(rst), .I(g_init[894]), 
        .Q(mreg[894]) );
  DFF \mreg_reg[893]  ( .D(mreg[893]), .CLK(clk), .RST(rst), .I(g_init[893]), 
        .Q(mreg[893]) );
  DFF \mreg_reg[892]  ( .D(mreg[892]), .CLK(clk), .RST(rst), .I(g_init[892]), 
        .Q(mreg[892]) );
  DFF \mreg_reg[891]  ( .D(mreg[891]), .CLK(clk), .RST(rst), .I(g_init[891]), 
        .Q(mreg[891]) );
  DFF \mreg_reg[890]  ( .D(mreg[890]), .CLK(clk), .RST(rst), .I(g_init[890]), 
        .Q(mreg[890]) );
  DFF \mreg_reg[889]  ( .D(mreg[889]), .CLK(clk), .RST(rst), .I(g_init[889]), 
        .Q(mreg[889]) );
  DFF \mreg_reg[888]  ( .D(mreg[888]), .CLK(clk), .RST(rst), .I(g_init[888]), 
        .Q(mreg[888]) );
  DFF \mreg_reg[887]  ( .D(mreg[887]), .CLK(clk), .RST(rst), .I(g_init[887]), 
        .Q(mreg[887]) );
  DFF \mreg_reg[886]  ( .D(mreg[886]), .CLK(clk), .RST(rst), .I(g_init[886]), 
        .Q(mreg[886]) );
  DFF \mreg_reg[885]  ( .D(mreg[885]), .CLK(clk), .RST(rst), .I(g_init[885]), 
        .Q(mreg[885]) );
  DFF \mreg_reg[884]  ( .D(mreg[884]), .CLK(clk), .RST(rst), .I(g_init[884]), 
        .Q(mreg[884]) );
  DFF \mreg_reg[883]  ( .D(mreg[883]), .CLK(clk), .RST(rst), .I(g_init[883]), 
        .Q(mreg[883]) );
  DFF \mreg_reg[882]  ( .D(mreg[882]), .CLK(clk), .RST(rst), .I(g_init[882]), 
        .Q(mreg[882]) );
  DFF \mreg_reg[881]  ( .D(mreg[881]), .CLK(clk), .RST(rst), .I(g_init[881]), 
        .Q(mreg[881]) );
  DFF \mreg_reg[880]  ( .D(mreg[880]), .CLK(clk), .RST(rst), .I(g_init[880]), 
        .Q(mreg[880]) );
  DFF \mreg_reg[879]  ( .D(mreg[879]), .CLK(clk), .RST(rst), .I(g_init[879]), 
        .Q(mreg[879]) );
  DFF \mreg_reg[878]  ( .D(mreg[878]), .CLK(clk), .RST(rst), .I(g_init[878]), 
        .Q(mreg[878]) );
  DFF \mreg_reg[877]  ( .D(mreg[877]), .CLK(clk), .RST(rst), .I(g_init[877]), 
        .Q(mreg[877]) );
  DFF \mreg_reg[876]  ( .D(mreg[876]), .CLK(clk), .RST(rst), .I(g_init[876]), 
        .Q(mreg[876]) );
  DFF \mreg_reg[875]  ( .D(mreg[875]), .CLK(clk), .RST(rst), .I(g_init[875]), 
        .Q(mreg[875]) );
  DFF \mreg_reg[874]  ( .D(mreg[874]), .CLK(clk), .RST(rst), .I(g_init[874]), 
        .Q(mreg[874]) );
  DFF \mreg_reg[873]  ( .D(mreg[873]), .CLK(clk), .RST(rst), .I(g_init[873]), 
        .Q(mreg[873]) );
  DFF \mreg_reg[872]  ( .D(mreg[872]), .CLK(clk), .RST(rst), .I(g_init[872]), 
        .Q(mreg[872]) );
  DFF \mreg_reg[871]  ( .D(mreg[871]), .CLK(clk), .RST(rst), .I(g_init[871]), 
        .Q(mreg[871]) );
  DFF \mreg_reg[870]  ( .D(mreg[870]), .CLK(clk), .RST(rst), .I(g_init[870]), 
        .Q(mreg[870]) );
  DFF \mreg_reg[869]  ( .D(mreg[869]), .CLK(clk), .RST(rst), .I(g_init[869]), 
        .Q(mreg[869]) );
  DFF \mreg_reg[868]  ( .D(mreg[868]), .CLK(clk), .RST(rst), .I(g_init[868]), 
        .Q(mreg[868]) );
  DFF \mreg_reg[867]  ( .D(mreg[867]), .CLK(clk), .RST(rst), .I(g_init[867]), 
        .Q(mreg[867]) );
  DFF \mreg_reg[866]  ( .D(mreg[866]), .CLK(clk), .RST(rst), .I(g_init[866]), 
        .Q(mreg[866]) );
  DFF \mreg_reg[865]  ( .D(mreg[865]), .CLK(clk), .RST(rst), .I(g_init[865]), 
        .Q(mreg[865]) );
  DFF \mreg_reg[864]  ( .D(mreg[864]), .CLK(clk), .RST(rst), .I(g_init[864]), 
        .Q(mreg[864]) );
  DFF \mreg_reg[863]  ( .D(mreg[863]), .CLK(clk), .RST(rst), .I(g_init[863]), 
        .Q(mreg[863]) );
  DFF \mreg_reg[862]  ( .D(mreg[862]), .CLK(clk), .RST(rst), .I(g_init[862]), 
        .Q(mreg[862]) );
  DFF \mreg_reg[861]  ( .D(mreg[861]), .CLK(clk), .RST(rst), .I(g_init[861]), 
        .Q(mreg[861]) );
  DFF \mreg_reg[860]  ( .D(mreg[860]), .CLK(clk), .RST(rst), .I(g_init[860]), 
        .Q(mreg[860]) );
  DFF \mreg_reg[859]  ( .D(mreg[859]), .CLK(clk), .RST(rst), .I(g_init[859]), 
        .Q(mreg[859]) );
  DFF \mreg_reg[858]  ( .D(mreg[858]), .CLK(clk), .RST(rst), .I(g_init[858]), 
        .Q(mreg[858]) );
  DFF \mreg_reg[857]  ( .D(mreg[857]), .CLK(clk), .RST(rst), .I(g_init[857]), 
        .Q(mreg[857]) );
  DFF \mreg_reg[856]  ( .D(mreg[856]), .CLK(clk), .RST(rst), .I(g_init[856]), 
        .Q(mreg[856]) );
  DFF \mreg_reg[855]  ( .D(mreg[855]), .CLK(clk), .RST(rst), .I(g_init[855]), 
        .Q(mreg[855]) );
  DFF \mreg_reg[854]  ( .D(mreg[854]), .CLK(clk), .RST(rst), .I(g_init[854]), 
        .Q(mreg[854]) );
  DFF \mreg_reg[853]  ( .D(mreg[853]), .CLK(clk), .RST(rst), .I(g_init[853]), 
        .Q(mreg[853]) );
  DFF \mreg_reg[852]  ( .D(mreg[852]), .CLK(clk), .RST(rst), .I(g_init[852]), 
        .Q(mreg[852]) );
  DFF \mreg_reg[851]  ( .D(mreg[851]), .CLK(clk), .RST(rst), .I(g_init[851]), 
        .Q(mreg[851]) );
  DFF \mreg_reg[850]  ( .D(mreg[850]), .CLK(clk), .RST(rst), .I(g_init[850]), 
        .Q(mreg[850]) );
  DFF \mreg_reg[849]  ( .D(mreg[849]), .CLK(clk), .RST(rst), .I(g_init[849]), 
        .Q(mreg[849]) );
  DFF \mreg_reg[848]  ( .D(mreg[848]), .CLK(clk), .RST(rst), .I(g_init[848]), 
        .Q(mreg[848]) );
  DFF \mreg_reg[847]  ( .D(mreg[847]), .CLK(clk), .RST(rst), .I(g_init[847]), 
        .Q(mreg[847]) );
  DFF \mreg_reg[846]  ( .D(mreg[846]), .CLK(clk), .RST(rst), .I(g_init[846]), 
        .Q(mreg[846]) );
  DFF \mreg_reg[845]  ( .D(mreg[845]), .CLK(clk), .RST(rst), .I(g_init[845]), 
        .Q(mreg[845]) );
  DFF \mreg_reg[844]  ( .D(mreg[844]), .CLK(clk), .RST(rst), .I(g_init[844]), 
        .Q(mreg[844]) );
  DFF \mreg_reg[843]  ( .D(mreg[843]), .CLK(clk), .RST(rst), .I(g_init[843]), 
        .Q(mreg[843]) );
  DFF \mreg_reg[842]  ( .D(mreg[842]), .CLK(clk), .RST(rst), .I(g_init[842]), 
        .Q(mreg[842]) );
  DFF \mreg_reg[841]  ( .D(mreg[841]), .CLK(clk), .RST(rst), .I(g_init[841]), 
        .Q(mreg[841]) );
  DFF \mreg_reg[840]  ( .D(mreg[840]), .CLK(clk), .RST(rst), .I(g_init[840]), 
        .Q(mreg[840]) );
  DFF \mreg_reg[839]  ( .D(mreg[839]), .CLK(clk), .RST(rst), .I(g_init[839]), 
        .Q(mreg[839]) );
  DFF \mreg_reg[838]  ( .D(mreg[838]), .CLK(clk), .RST(rst), .I(g_init[838]), 
        .Q(mreg[838]) );
  DFF \mreg_reg[837]  ( .D(mreg[837]), .CLK(clk), .RST(rst), .I(g_init[837]), 
        .Q(mreg[837]) );
  DFF \mreg_reg[836]  ( .D(mreg[836]), .CLK(clk), .RST(rst), .I(g_init[836]), 
        .Q(mreg[836]) );
  DFF \mreg_reg[835]  ( .D(mreg[835]), .CLK(clk), .RST(rst), .I(g_init[835]), 
        .Q(mreg[835]) );
  DFF \mreg_reg[834]  ( .D(mreg[834]), .CLK(clk), .RST(rst), .I(g_init[834]), 
        .Q(mreg[834]) );
  DFF \mreg_reg[833]  ( .D(mreg[833]), .CLK(clk), .RST(rst), .I(g_init[833]), 
        .Q(mreg[833]) );
  DFF \mreg_reg[832]  ( .D(mreg[832]), .CLK(clk), .RST(rst), .I(g_init[832]), 
        .Q(mreg[832]) );
  DFF \mreg_reg[831]  ( .D(mreg[831]), .CLK(clk), .RST(rst), .I(g_init[831]), 
        .Q(mreg[831]) );
  DFF \mreg_reg[830]  ( .D(mreg[830]), .CLK(clk), .RST(rst), .I(g_init[830]), 
        .Q(mreg[830]) );
  DFF \mreg_reg[829]  ( .D(mreg[829]), .CLK(clk), .RST(rst), .I(g_init[829]), 
        .Q(mreg[829]) );
  DFF \mreg_reg[828]  ( .D(mreg[828]), .CLK(clk), .RST(rst), .I(g_init[828]), 
        .Q(mreg[828]) );
  DFF \mreg_reg[827]  ( .D(mreg[827]), .CLK(clk), .RST(rst), .I(g_init[827]), 
        .Q(mreg[827]) );
  DFF \mreg_reg[826]  ( .D(mreg[826]), .CLK(clk), .RST(rst), .I(g_init[826]), 
        .Q(mreg[826]) );
  DFF \mreg_reg[825]  ( .D(mreg[825]), .CLK(clk), .RST(rst), .I(g_init[825]), 
        .Q(mreg[825]) );
  DFF \mreg_reg[824]  ( .D(mreg[824]), .CLK(clk), .RST(rst), .I(g_init[824]), 
        .Q(mreg[824]) );
  DFF \mreg_reg[823]  ( .D(mreg[823]), .CLK(clk), .RST(rst), .I(g_init[823]), 
        .Q(mreg[823]) );
  DFF \mreg_reg[822]  ( .D(mreg[822]), .CLK(clk), .RST(rst), .I(g_init[822]), 
        .Q(mreg[822]) );
  DFF \mreg_reg[821]  ( .D(mreg[821]), .CLK(clk), .RST(rst), .I(g_init[821]), 
        .Q(mreg[821]) );
  DFF \mreg_reg[820]  ( .D(mreg[820]), .CLK(clk), .RST(rst), .I(g_init[820]), 
        .Q(mreg[820]) );
  DFF \mreg_reg[819]  ( .D(mreg[819]), .CLK(clk), .RST(rst), .I(g_init[819]), 
        .Q(mreg[819]) );
  DFF \mreg_reg[818]  ( .D(mreg[818]), .CLK(clk), .RST(rst), .I(g_init[818]), 
        .Q(mreg[818]) );
  DFF \mreg_reg[817]  ( .D(mreg[817]), .CLK(clk), .RST(rst), .I(g_init[817]), 
        .Q(mreg[817]) );
  DFF \mreg_reg[816]  ( .D(mreg[816]), .CLK(clk), .RST(rst), .I(g_init[816]), 
        .Q(mreg[816]) );
  DFF \mreg_reg[815]  ( .D(mreg[815]), .CLK(clk), .RST(rst), .I(g_init[815]), 
        .Q(mreg[815]) );
  DFF \mreg_reg[814]  ( .D(mreg[814]), .CLK(clk), .RST(rst), .I(g_init[814]), 
        .Q(mreg[814]) );
  DFF \mreg_reg[813]  ( .D(mreg[813]), .CLK(clk), .RST(rst), .I(g_init[813]), 
        .Q(mreg[813]) );
  DFF \mreg_reg[812]  ( .D(mreg[812]), .CLK(clk), .RST(rst), .I(g_init[812]), 
        .Q(mreg[812]) );
  DFF \mreg_reg[811]  ( .D(mreg[811]), .CLK(clk), .RST(rst), .I(g_init[811]), 
        .Q(mreg[811]) );
  DFF \mreg_reg[810]  ( .D(mreg[810]), .CLK(clk), .RST(rst), .I(g_init[810]), 
        .Q(mreg[810]) );
  DFF \mreg_reg[809]  ( .D(mreg[809]), .CLK(clk), .RST(rst), .I(g_init[809]), 
        .Q(mreg[809]) );
  DFF \mreg_reg[808]  ( .D(mreg[808]), .CLK(clk), .RST(rst), .I(g_init[808]), 
        .Q(mreg[808]) );
  DFF \mreg_reg[807]  ( .D(mreg[807]), .CLK(clk), .RST(rst), .I(g_init[807]), 
        .Q(mreg[807]) );
  DFF \mreg_reg[806]  ( .D(mreg[806]), .CLK(clk), .RST(rst), .I(g_init[806]), 
        .Q(mreg[806]) );
  DFF \mreg_reg[805]  ( .D(mreg[805]), .CLK(clk), .RST(rst), .I(g_init[805]), 
        .Q(mreg[805]) );
  DFF \mreg_reg[804]  ( .D(mreg[804]), .CLK(clk), .RST(rst), .I(g_init[804]), 
        .Q(mreg[804]) );
  DFF \mreg_reg[803]  ( .D(mreg[803]), .CLK(clk), .RST(rst), .I(g_init[803]), 
        .Q(mreg[803]) );
  DFF \mreg_reg[802]  ( .D(mreg[802]), .CLK(clk), .RST(rst), .I(g_init[802]), 
        .Q(mreg[802]) );
  DFF \mreg_reg[801]  ( .D(mreg[801]), .CLK(clk), .RST(rst), .I(g_init[801]), 
        .Q(mreg[801]) );
  DFF \mreg_reg[800]  ( .D(mreg[800]), .CLK(clk), .RST(rst), .I(g_init[800]), 
        .Q(mreg[800]) );
  DFF \mreg_reg[799]  ( .D(mreg[799]), .CLK(clk), .RST(rst), .I(g_init[799]), 
        .Q(mreg[799]) );
  DFF \mreg_reg[798]  ( .D(mreg[798]), .CLK(clk), .RST(rst), .I(g_init[798]), 
        .Q(mreg[798]) );
  DFF \mreg_reg[797]  ( .D(mreg[797]), .CLK(clk), .RST(rst), .I(g_init[797]), 
        .Q(mreg[797]) );
  DFF \mreg_reg[796]  ( .D(mreg[796]), .CLK(clk), .RST(rst), .I(g_init[796]), 
        .Q(mreg[796]) );
  DFF \mreg_reg[795]  ( .D(mreg[795]), .CLK(clk), .RST(rst), .I(g_init[795]), 
        .Q(mreg[795]) );
  DFF \mreg_reg[794]  ( .D(mreg[794]), .CLK(clk), .RST(rst), .I(g_init[794]), 
        .Q(mreg[794]) );
  DFF \mreg_reg[793]  ( .D(mreg[793]), .CLK(clk), .RST(rst), .I(g_init[793]), 
        .Q(mreg[793]) );
  DFF \mreg_reg[792]  ( .D(mreg[792]), .CLK(clk), .RST(rst), .I(g_init[792]), 
        .Q(mreg[792]) );
  DFF \mreg_reg[791]  ( .D(mreg[791]), .CLK(clk), .RST(rst), .I(g_init[791]), 
        .Q(mreg[791]) );
  DFF \mreg_reg[790]  ( .D(mreg[790]), .CLK(clk), .RST(rst), .I(g_init[790]), 
        .Q(mreg[790]) );
  DFF \mreg_reg[789]  ( .D(mreg[789]), .CLK(clk), .RST(rst), .I(g_init[789]), 
        .Q(mreg[789]) );
  DFF \mreg_reg[788]  ( .D(mreg[788]), .CLK(clk), .RST(rst), .I(g_init[788]), 
        .Q(mreg[788]) );
  DFF \mreg_reg[787]  ( .D(mreg[787]), .CLK(clk), .RST(rst), .I(g_init[787]), 
        .Q(mreg[787]) );
  DFF \mreg_reg[786]  ( .D(mreg[786]), .CLK(clk), .RST(rst), .I(g_init[786]), 
        .Q(mreg[786]) );
  DFF \mreg_reg[785]  ( .D(mreg[785]), .CLK(clk), .RST(rst), .I(g_init[785]), 
        .Q(mreg[785]) );
  DFF \mreg_reg[784]  ( .D(mreg[784]), .CLK(clk), .RST(rst), .I(g_init[784]), 
        .Q(mreg[784]) );
  DFF \mreg_reg[783]  ( .D(mreg[783]), .CLK(clk), .RST(rst), .I(g_init[783]), 
        .Q(mreg[783]) );
  DFF \mreg_reg[782]  ( .D(mreg[782]), .CLK(clk), .RST(rst), .I(g_init[782]), 
        .Q(mreg[782]) );
  DFF \mreg_reg[781]  ( .D(mreg[781]), .CLK(clk), .RST(rst), .I(g_init[781]), 
        .Q(mreg[781]) );
  DFF \mreg_reg[780]  ( .D(mreg[780]), .CLK(clk), .RST(rst), .I(g_init[780]), 
        .Q(mreg[780]) );
  DFF \mreg_reg[779]  ( .D(mreg[779]), .CLK(clk), .RST(rst), .I(g_init[779]), 
        .Q(mreg[779]) );
  DFF \mreg_reg[778]  ( .D(mreg[778]), .CLK(clk), .RST(rst), .I(g_init[778]), 
        .Q(mreg[778]) );
  DFF \mreg_reg[777]  ( .D(mreg[777]), .CLK(clk), .RST(rst), .I(g_init[777]), 
        .Q(mreg[777]) );
  DFF \mreg_reg[776]  ( .D(mreg[776]), .CLK(clk), .RST(rst), .I(g_init[776]), 
        .Q(mreg[776]) );
  DFF \mreg_reg[775]  ( .D(mreg[775]), .CLK(clk), .RST(rst), .I(g_init[775]), 
        .Q(mreg[775]) );
  DFF \mreg_reg[774]  ( .D(mreg[774]), .CLK(clk), .RST(rst), .I(g_init[774]), 
        .Q(mreg[774]) );
  DFF \mreg_reg[773]  ( .D(mreg[773]), .CLK(clk), .RST(rst), .I(g_init[773]), 
        .Q(mreg[773]) );
  DFF \mreg_reg[772]  ( .D(mreg[772]), .CLK(clk), .RST(rst), .I(g_init[772]), 
        .Q(mreg[772]) );
  DFF \mreg_reg[771]  ( .D(mreg[771]), .CLK(clk), .RST(rst), .I(g_init[771]), 
        .Q(mreg[771]) );
  DFF \mreg_reg[770]  ( .D(mreg[770]), .CLK(clk), .RST(rst), .I(g_init[770]), 
        .Q(mreg[770]) );
  DFF \mreg_reg[769]  ( .D(mreg[769]), .CLK(clk), .RST(rst), .I(g_init[769]), 
        .Q(mreg[769]) );
  DFF \mreg_reg[768]  ( .D(mreg[768]), .CLK(clk), .RST(rst), .I(g_init[768]), 
        .Q(mreg[768]) );
  DFF \mreg_reg[767]  ( .D(mreg[767]), .CLK(clk), .RST(rst), .I(g_init[767]), 
        .Q(mreg[767]) );
  DFF \mreg_reg[766]  ( .D(mreg[766]), .CLK(clk), .RST(rst), .I(g_init[766]), 
        .Q(mreg[766]) );
  DFF \mreg_reg[765]  ( .D(mreg[765]), .CLK(clk), .RST(rst), .I(g_init[765]), 
        .Q(mreg[765]) );
  DFF \mreg_reg[764]  ( .D(mreg[764]), .CLK(clk), .RST(rst), .I(g_init[764]), 
        .Q(mreg[764]) );
  DFF \mreg_reg[763]  ( .D(mreg[763]), .CLK(clk), .RST(rst), .I(g_init[763]), 
        .Q(mreg[763]) );
  DFF \mreg_reg[762]  ( .D(mreg[762]), .CLK(clk), .RST(rst), .I(g_init[762]), 
        .Q(mreg[762]) );
  DFF \mreg_reg[761]  ( .D(mreg[761]), .CLK(clk), .RST(rst), .I(g_init[761]), 
        .Q(mreg[761]) );
  DFF \mreg_reg[760]  ( .D(mreg[760]), .CLK(clk), .RST(rst), .I(g_init[760]), 
        .Q(mreg[760]) );
  DFF \mreg_reg[759]  ( .D(mreg[759]), .CLK(clk), .RST(rst), .I(g_init[759]), 
        .Q(mreg[759]) );
  DFF \mreg_reg[758]  ( .D(mreg[758]), .CLK(clk), .RST(rst), .I(g_init[758]), 
        .Q(mreg[758]) );
  DFF \mreg_reg[757]  ( .D(mreg[757]), .CLK(clk), .RST(rst), .I(g_init[757]), 
        .Q(mreg[757]) );
  DFF \mreg_reg[756]  ( .D(mreg[756]), .CLK(clk), .RST(rst), .I(g_init[756]), 
        .Q(mreg[756]) );
  DFF \mreg_reg[755]  ( .D(mreg[755]), .CLK(clk), .RST(rst), .I(g_init[755]), 
        .Q(mreg[755]) );
  DFF \mreg_reg[754]  ( .D(mreg[754]), .CLK(clk), .RST(rst), .I(g_init[754]), 
        .Q(mreg[754]) );
  DFF \mreg_reg[753]  ( .D(mreg[753]), .CLK(clk), .RST(rst), .I(g_init[753]), 
        .Q(mreg[753]) );
  DFF \mreg_reg[752]  ( .D(mreg[752]), .CLK(clk), .RST(rst), .I(g_init[752]), 
        .Q(mreg[752]) );
  DFF \mreg_reg[751]  ( .D(mreg[751]), .CLK(clk), .RST(rst), .I(g_init[751]), 
        .Q(mreg[751]) );
  DFF \mreg_reg[750]  ( .D(mreg[750]), .CLK(clk), .RST(rst), .I(g_init[750]), 
        .Q(mreg[750]) );
  DFF \mreg_reg[749]  ( .D(mreg[749]), .CLK(clk), .RST(rst), .I(g_init[749]), 
        .Q(mreg[749]) );
  DFF \mreg_reg[748]  ( .D(mreg[748]), .CLK(clk), .RST(rst), .I(g_init[748]), 
        .Q(mreg[748]) );
  DFF \mreg_reg[747]  ( .D(mreg[747]), .CLK(clk), .RST(rst), .I(g_init[747]), 
        .Q(mreg[747]) );
  DFF \mreg_reg[746]  ( .D(mreg[746]), .CLK(clk), .RST(rst), .I(g_init[746]), 
        .Q(mreg[746]) );
  DFF \mreg_reg[745]  ( .D(mreg[745]), .CLK(clk), .RST(rst), .I(g_init[745]), 
        .Q(mreg[745]) );
  DFF \mreg_reg[744]  ( .D(mreg[744]), .CLK(clk), .RST(rst), .I(g_init[744]), 
        .Q(mreg[744]) );
  DFF \mreg_reg[743]  ( .D(mreg[743]), .CLK(clk), .RST(rst), .I(g_init[743]), 
        .Q(mreg[743]) );
  DFF \mreg_reg[742]  ( .D(mreg[742]), .CLK(clk), .RST(rst), .I(g_init[742]), 
        .Q(mreg[742]) );
  DFF \mreg_reg[741]  ( .D(mreg[741]), .CLK(clk), .RST(rst), .I(g_init[741]), 
        .Q(mreg[741]) );
  DFF \mreg_reg[740]  ( .D(mreg[740]), .CLK(clk), .RST(rst), .I(g_init[740]), 
        .Q(mreg[740]) );
  DFF \mreg_reg[739]  ( .D(mreg[739]), .CLK(clk), .RST(rst), .I(g_init[739]), 
        .Q(mreg[739]) );
  DFF \mreg_reg[738]  ( .D(mreg[738]), .CLK(clk), .RST(rst), .I(g_init[738]), 
        .Q(mreg[738]) );
  DFF \mreg_reg[737]  ( .D(mreg[737]), .CLK(clk), .RST(rst), .I(g_init[737]), 
        .Q(mreg[737]) );
  DFF \mreg_reg[736]  ( .D(mreg[736]), .CLK(clk), .RST(rst), .I(g_init[736]), 
        .Q(mreg[736]) );
  DFF \mreg_reg[735]  ( .D(mreg[735]), .CLK(clk), .RST(rst), .I(g_init[735]), 
        .Q(mreg[735]) );
  DFF \mreg_reg[734]  ( .D(mreg[734]), .CLK(clk), .RST(rst), .I(g_init[734]), 
        .Q(mreg[734]) );
  DFF \mreg_reg[733]  ( .D(mreg[733]), .CLK(clk), .RST(rst), .I(g_init[733]), 
        .Q(mreg[733]) );
  DFF \mreg_reg[732]  ( .D(mreg[732]), .CLK(clk), .RST(rst), .I(g_init[732]), 
        .Q(mreg[732]) );
  DFF \mreg_reg[731]  ( .D(mreg[731]), .CLK(clk), .RST(rst), .I(g_init[731]), 
        .Q(mreg[731]) );
  DFF \mreg_reg[730]  ( .D(mreg[730]), .CLK(clk), .RST(rst), .I(g_init[730]), 
        .Q(mreg[730]) );
  DFF \mreg_reg[729]  ( .D(mreg[729]), .CLK(clk), .RST(rst), .I(g_init[729]), 
        .Q(mreg[729]) );
  DFF \mreg_reg[728]  ( .D(mreg[728]), .CLK(clk), .RST(rst), .I(g_init[728]), 
        .Q(mreg[728]) );
  DFF \mreg_reg[727]  ( .D(mreg[727]), .CLK(clk), .RST(rst), .I(g_init[727]), 
        .Q(mreg[727]) );
  DFF \mreg_reg[726]  ( .D(mreg[726]), .CLK(clk), .RST(rst), .I(g_init[726]), 
        .Q(mreg[726]) );
  DFF \mreg_reg[725]  ( .D(mreg[725]), .CLK(clk), .RST(rst), .I(g_init[725]), 
        .Q(mreg[725]) );
  DFF \mreg_reg[724]  ( .D(mreg[724]), .CLK(clk), .RST(rst), .I(g_init[724]), 
        .Q(mreg[724]) );
  DFF \mreg_reg[723]  ( .D(mreg[723]), .CLK(clk), .RST(rst), .I(g_init[723]), 
        .Q(mreg[723]) );
  DFF \mreg_reg[722]  ( .D(mreg[722]), .CLK(clk), .RST(rst), .I(g_init[722]), 
        .Q(mreg[722]) );
  DFF \mreg_reg[721]  ( .D(mreg[721]), .CLK(clk), .RST(rst), .I(g_init[721]), 
        .Q(mreg[721]) );
  DFF \mreg_reg[720]  ( .D(mreg[720]), .CLK(clk), .RST(rst), .I(g_init[720]), 
        .Q(mreg[720]) );
  DFF \mreg_reg[719]  ( .D(mreg[719]), .CLK(clk), .RST(rst), .I(g_init[719]), 
        .Q(mreg[719]) );
  DFF \mreg_reg[718]  ( .D(mreg[718]), .CLK(clk), .RST(rst), .I(g_init[718]), 
        .Q(mreg[718]) );
  DFF \mreg_reg[717]  ( .D(mreg[717]), .CLK(clk), .RST(rst), .I(g_init[717]), 
        .Q(mreg[717]) );
  DFF \mreg_reg[716]  ( .D(mreg[716]), .CLK(clk), .RST(rst), .I(g_init[716]), 
        .Q(mreg[716]) );
  DFF \mreg_reg[715]  ( .D(mreg[715]), .CLK(clk), .RST(rst), .I(g_init[715]), 
        .Q(mreg[715]) );
  DFF \mreg_reg[714]  ( .D(mreg[714]), .CLK(clk), .RST(rst), .I(g_init[714]), 
        .Q(mreg[714]) );
  DFF \mreg_reg[713]  ( .D(mreg[713]), .CLK(clk), .RST(rst), .I(g_init[713]), 
        .Q(mreg[713]) );
  DFF \mreg_reg[712]  ( .D(mreg[712]), .CLK(clk), .RST(rst), .I(g_init[712]), 
        .Q(mreg[712]) );
  DFF \mreg_reg[711]  ( .D(mreg[711]), .CLK(clk), .RST(rst), .I(g_init[711]), 
        .Q(mreg[711]) );
  DFF \mreg_reg[710]  ( .D(mreg[710]), .CLK(clk), .RST(rst), .I(g_init[710]), 
        .Q(mreg[710]) );
  DFF \mreg_reg[709]  ( .D(mreg[709]), .CLK(clk), .RST(rst), .I(g_init[709]), 
        .Q(mreg[709]) );
  DFF \mreg_reg[708]  ( .D(mreg[708]), .CLK(clk), .RST(rst), .I(g_init[708]), 
        .Q(mreg[708]) );
  DFF \mreg_reg[707]  ( .D(mreg[707]), .CLK(clk), .RST(rst), .I(g_init[707]), 
        .Q(mreg[707]) );
  DFF \mreg_reg[706]  ( .D(mreg[706]), .CLK(clk), .RST(rst), .I(g_init[706]), 
        .Q(mreg[706]) );
  DFF \mreg_reg[705]  ( .D(mreg[705]), .CLK(clk), .RST(rst), .I(g_init[705]), 
        .Q(mreg[705]) );
  DFF \mreg_reg[704]  ( .D(mreg[704]), .CLK(clk), .RST(rst), .I(g_init[704]), 
        .Q(mreg[704]) );
  DFF \mreg_reg[703]  ( .D(mreg[703]), .CLK(clk), .RST(rst), .I(g_init[703]), 
        .Q(mreg[703]) );
  DFF \mreg_reg[702]  ( .D(mreg[702]), .CLK(clk), .RST(rst), .I(g_init[702]), 
        .Q(mreg[702]) );
  DFF \mreg_reg[701]  ( .D(mreg[701]), .CLK(clk), .RST(rst), .I(g_init[701]), 
        .Q(mreg[701]) );
  DFF \mreg_reg[700]  ( .D(mreg[700]), .CLK(clk), .RST(rst), .I(g_init[700]), 
        .Q(mreg[700]) );
  DFF \mreg_reg[699]  ( .D(mreg[699]), .CLK(clk), .RST(rst), .I(g_init[699]), 
        .Q(mreg[699]) );
  DFF \mreg_reg[698]  ( .D(mreg[698]), .CLK(clk), .RST(rst), .I(g_init[698]), 
        .Q(mreg[698]) );
  DFF \mreg_reg[697]  ( .D(mreg[697]), .CLK(clk), .RST(rst), .I(g_init[697]), 
        .Q(mreg[697]) );
  DFF \mreg_reg[696]  ( .D(mreg[696]), .CLK(clk), .RST(rst), .I(g_init[696]), 
        .Q(mreg[696]) );
  DFF \mreg_reg[695]  ( .D(mreg[695]), .CLK(clk), .RST(rst), .I(g_init[695]), 
        .Q(mreg[695]) );
  DFF \mreg_reg[694]  ( .D(mreg[694]), .CLK(clk), .RST(rst), .I(g_init[694]), 
        .Q(mreg[694]) );
  DFF \mreg_reg[693]  ( .D(mreg[693]), .CLK(clk), .RST(rst), .I(g_init[693]), 
        .Q(mreg[693]) );
  DFF \mreg_reg[692]  ( .D(mreg[692]), .CLK(clk), .RST(rst), .I(g_init[692]), 
        .Q(mreg[692]) );
  DFF \mreg_reg[691]  ( .D(mreg[691]), .CLK(clk), .RST(rst), .I(g_init[691]), 
        .Q(mreg[691]) );
  DFF \mreg_reg[690]  ( .D(mreg[690]), .CLK(clk), .RST(rst), .I(g_init[690]), 
        .Q(mreg[690]) );
  DFF \mreg_reg[689]  ( .D(mreg[689]), .CLK(clk), .RST(rst), .I(g_init[689]), 
        .Q(mreg[689]) );
  DFF \mreg_reg[688]  ( .D(mreg[688]), .CLK(clk), .RST(rst), .I(g_init[688]), 
        .Q(mreg[688]) );
  DFF \mreg_reg[687]  ( .D(mreg[687]), .CLK(clk), .RST(rst), .I(g_init[687]), 
        .Q(mreg[687]) );
  DFF \mreg_reg[686]  ( .D(mreg[686]), .CLK(clk), .RST(rst), .I(g_init[686]), 
        .Q(mreg[686]) );
  DFF \mreg_reg[685]  ( .D(mreg[685]), .CLK(clk), .RST(rst), .I(g_init[685]), 
        .Q(mreg[685]) );
  DFF \mreg_reg[684]  ( .D(mreg[684]), .CLK(clk), .RST(rst), .I(g_init[684]), 
        .Q(mreg[684]) );
  DFF \mreg_reg[683]  ( .D(mreg[683]), .CLK(clk), .RST(rst), .I(g_init[683]), 
        .Q(mreg[683]) );
  DFF \mreg_reg[682]  ( .D(mreg[682]), .CLK(clk), .RST(rst), .I(g_init[682]), 
        .Q(mreg[682]) );
  DFF \mreg_reg[681]  ( .D(mreg[681]), .CLK(clk), .RST(rst), .I(g_init[681]), 
        .Q(mreg[681]) );
  DFF \mreg_reg[680]  ( .D(mreg[680]), .CLK(clk), .RST(rst), .I(g_init[680]), 
        .Q(mreg[680]) );
  DFF \mreg_reg[679]  ( .D(mreg[679]), .CLK(clk), .RST(rst), .I(g_init[679]), 
        .Q(mreg[679]) );
  DFF \mreg_reg[678]  ( .D(mreg[678]), .CLK(clk), .RST(rst), .I(g_init[678]), 
        .Q(mreg[678]) );
  DFF \mreg_reg[677]  ( .D(mreg[677]), .CLK(clk), .RST(rst), .I(g_init[677]), 
        .Q(mreg[677]) );
  DFF \mreg_reg[676]  ( .D(mreg[676]), .CLK(clk), .RST(rst), .I(g_init[676]), 
        .Q(mreg[676]) );
  DFF \mreg_reg[675]  ( .D(mreg[675]), .CLK(clk), .RST(rst), .I(g_init[675]), 
        .Q(mreg[675]) );
  DFF \mreg_reg[674]  ( .D(mreg[674]), .CLK(clk), .RST(rst), .I(g_init[674]), 
        .Q(mreg[674]) );
  DFF \mreg_reg[673]  ( .D(mreg[673]), .CLK(clk), .RST(rst), .I(g_init[673]), 
        .Q(mreg[673]) );
  DFF \mreg_reg[672]  ( .D(mreg[672]), .CLK(clk), .RST(rst), .I(g_init[672]), 
        .Q(mreg[672]) );
  DFF \mreg_reg[671]  ( .D(mreg[671]), .CLK(clk), .RST(rst), .I(g_init[671]), 
        .Q(mreg[671]) );
  DFF \mreg_reg[670]  ( .D(mreg[670]), .CLK(clk), .RST(rst), .I(g_init[670]), 
        .Q(mreg[670]) );
  DFF \mreg_reg[669]  ( .D(mreg[669]), .CLK(clk), .RST(rst), .I(g_init[669]), 
        .Q(mreg[669]) );
  DFF \mreg_reg[668]  ( .D(mreg[668]), .CLK(clk), .RST(rst), .I(g_init[668]), 
        .Q(mreg[668]) );
  DFF \mreg_reg[667]  ( .D(mreg[667]), .CLK(clk), .RST(rst), .I(g_init[667]), 
        .Q(mreg[667]) );
  DFF \mreg_reg[666]  ( .D(mreg[666]), .CLK(clk), .RST(rst), .I(g_init[666]), 
        .Q(mreg[666]) );
  DFF \mreg_reg[665]  ( .D(mreg[665]), .CLK(clk), .RST(rst), .I(g_init[665]), 
        .Q(mreg[665]) );
  DFF \mreg_reg[664]  ( .D(mreg[664]), .CLK(clk), .RST(rst), .I(g_init[664]), 
        .Q(mreg[664]) );
  DFF \mreg_reg[663]  ( .D(mreg[663]), .CLK(clk), .RST(rst), .I(g_init[663]), 
        .Q(mreg[663]) );
  DFF \mreg_reg[662]  ( .D(mreg[662]), .CLK(clk), .RST(rst), .I(g_init[662]), 
        .Q(mreg[662]) );
  DFF \mreg_reg[661]  ( .D(mreg[661]), .CLK(clk), .RST(rst), .I(g_init[661]), 
        .Q(mreg[661]) );
  DFF \mreg_reg[660]  ( .D(mreg[660]), .CLK(clk), .RST(rst), .I(g_init[660]), 
        .Q(mreg[660]) );
  DFF \mreg_reg[659]  ( .D(mreg[659]), .CLK(clk), .RST(rst), .I(g_init[659]), 
        .Q(mreg[659]) );
  DFF \mreg_reg[658]  ( .D(mreg[658]), .CLK(clk), .RST(rst), .I(g_init[658]), 
        .Q(mreg[658]) );
  DFF \mreg_reg[657]  ( .D(mreg[657]), .CLK(clk), .RST(rst), .I(g_init[657]), 
        .Q(mreg[657]) );
  DFF \mreg_reg[656]  ( .D(mreg[656]), .CLK(clk), .RST(rst), .I(g_init[656]), 
        .Q(mreg[656]) );
  DFF \mreg_reg[655]  ( .D(mreg[655]), .CLK(clk), .RST(rst), .I(g_init[655]), 
        .Q(mreg[655]) );
  DFF \mreg_reg[654]  ( .D(mreg[654]), .CLK(clk), .RST(rst), .I(g_init[654]), 
        .Q(mreg[654]) );
  DFF \mreg_reg[653]  ( .D(mreg[653]), .CLK(clk), .RST(rst), .I(g_init[653]), 
        .Q(mreg[653]) );
  DFF \mreg_reg[652]  ( .D(mreg[652]), .CLK(clk), .RST(rst), .I(g_init[652]), 
        .Q(mreg[652]) );
  DFF \mreg_reg[651]  ( .D(mreg[651]), .CLK(clk), .RST(rst), .I(g_init[651]), 
        .Q(mreg[651]) );
  DFF \mreg_reg[650]  ( .D(mreg[650]), .CLK(clk), .RST(rst), .I(g_init[650]), 
        .Q(mreg[650]) );
  DFF \mreg_reg[649]  ( .D(mreg[649]), .CLK(clk), .RST(rst), .I(g_init[649]), 
        .Q(mreg[649]) );
  DFF \mreg_reg[648]  ( .D(mreg[648]), .CLK(clk), .RST(rst), .I(g_init[648]), 
        .Q(mreg[648]) );
  DFF \mreg_reg[647]  ( .D(mreg[647]), .CLK(clk), .RST(rst), .I(g_init[647]), 
        .Q(mreg[647]) );
  DFF \mreg_reg[646]  ( .D(mreg[646]), .CLK(clk), .RST(rst), .I(g_init[646]), 
        .Q(mreg[646]) );
  DFF \mreg_reg[645]  ( .D(mreg[645]), .CLK(clk), .RST(rst), .I(g_init[645]), 
        .Q(mreg[645]) );
  DFF \mreg_reg[644]  ( .D(mreg[644]), .CLK(clk), .RST(rst), .I(g_init[644]), 
        .Q(mreg[644]) );
  DFF \mreg_reg[643]  ( .D(mreg[643]), .CLK(clk), .RST(rst), .I(g_init[643]), 
        .Q(mreg[643]) );
  DFF \mreg_reg[642]  ( .D(mreg[642]), .CLK(clk), .RST(rst), .I(g_init[642]), 
        .Q(mreg[642]) );
  DFF \mreg_reg[641]  ( .D(mreg[641]), .CLK(clk), .RST(rst), .I(g_init[641]), 
        .Q(mreg[641]) );
  DFF \mreg_reg[640]  ( .D(mreg[640]), .CLK(clk), .RST(rst), .I(g_init[640]), 
        .Q(mreg[640]) );
  DFF \mreg_reg[639]  ( .D(mreg[639]), .CLK(clk), .RST(rst), .I(g_init[639]), 
        .Q(mreg[639]) );
  DFF \mreg_reg[638]  ( .D(mreg[638]), .CLK(clk), .RST(rst), .I(g_init[638]), 
        .Q(mreg[638]) );
  DFF \mreg_reg[637]  ( .D(mreg[637]), .CLK(clk), .RST(rst), .I(g_init[637]), 
        .Q(mreg[637]) );
  DFF \mreg_reg[636]  ( .D(mreg[636]), .CLK(clk), .RST(rst), .I(g_init[636]), 
        .Q(mreg[636]) );
  DFF \mreg_reg[635]  ( .D(mreg[635]), .CLK(clk), .RST(rst), .I(g_init[635]), 
        .Q(mreg[635]) );
  DFF \mreg_reg[634]  ( .D(mreg[634]), .CLK(clk), .RST(rst), .I(g_init[634]), 
        .Q(mreg[634]) );
  DFF \mreg_reg[633]  ( .D(mreg[633]), .CLK(clk), .RST(rst), .I(g_init[633]), 
        .Q(mreg[633]) );
  DFF \mreg_reg[632]  ( .D(mreg[632]), .CLK(clk), .RST(rst), .I(g_init[632]), 
        .Q(mreg[632]) );
  DFF \mreg_reg[631]  ( .D(mreg[631]), .CLK(clk), .RST(rst), .I(g_init[631]), 
        .Q(mreg[631]) );
  DFF \mreg_reg[630]  ( .D(mreg[630]), .CLK(clk), .RST(rst), .I(g_init[630]), 
        .Q(mreg[630]) );
  DFF \mreg_reg[629]  ( .D(mreg[629]), .CLK(clk), .RST(rst), .I(g_init[629]), 
        .Q(mreg[629]) );
  DFF \mreg_reg[628]  ( .D(mreg[628]), .CLK(clk), .RST(rst), .I(g_init[628]), 
        .Q(mreg[628]) );
  DFF \mreg_reg[627]  ( .D(mreg[627]), .CLK(clk), .RST(rst), .I(g_init[627]), 
        .Q(mreg[627]) );
  DFF \mreg_reg[626]  ( .D(mreg[626]), .CLK(clk), .RST(rst), .I(g_init[626]), 
        .Q(mreg[626]) );
  DFF \mreg_reg[625]  ( .D(mreg[625]), .CLK(clk), .RST(rst), .I(g_init[625]), 
        .Q(mreg[625]) );
  DFF \mreg_reg[624]  ( .D(mreg[624]), .CLK(clk), .RST(rst), .I(g_init[624]), 
        .Q(mreg[624]) );
  DFF \mreg_reg[623]  ( .D(mreg[623]), .CLK(clk), .RST(rst), .I(g_init[623]), 
        .Q(mreg[623]) );
  DFF \mreg_reg[622]  ( .D(mreg[622]), .CLK(clk), .RST(rst), .I(g_init[622]), 
        .Q(mreg[622]) );
  DFF \mreg_reg[621]  ( .D(mreg[621]), .CLK(clk), .RST(rst), .I(g_init[621]), 
        .Q(mreg[621]) );
  DFF \mreg_reg[620]  ( .D(mreg[620]), .CLK(clk), .RST(rst), .I(g_init[620]), 
        .Q(mreg[620]) );
  DFF \mreg_reg[619]  ( .D(mreg[619]), .CLK(clk), .RST(rst), .I(g_init[619]), 
        .Q(mreg[619]) );
  DFF \mreg_reg[618]  ( .D(mreg[618]), .CLK(clk), .RST(rst), .I(g_init[618]), 
        .Q(mreg[618]) );
  DFF \mreg_reg[617]  ( .D(mreg[617]), .CLK(clk), .RST(rst), .I(g_init[617]), 
        .Q(mreg[617]) );
  DFF \mreg_reg[616]  ( .D(mreg[616]), .CLK(clk), .RST(rst), .I(g_init[616]), 
        .Q(mreg[616]) );
  DFF \mreg_reg[615]  ( .D(mreg[615]), .CLK(clk), .RST(rst), .I(g_init[615]), 
        .Q(mreg[615]) );
  DFF \mreg_reg[614]  ( .D(mreg[614]), .CLK(clk), .RST(rst), .I(g_init[614]), 
        .Q(mreg[614]) );
  DFF \mreg_reg[613]  ( .D(mreg[613]), .CLK(clk), .RST(rst), .I(g_init[613]), 
        .Q(mreg[613]) );
  DFF \mreg_reg[612]  ( .D(mreg[612]), .CLK(clk), .RST(rst), .I(g_init[612]), 
        .Q(mreg[612]) );
  DFF \mreg_reg[611]  ( .D(mreg[611]), .CLK(clk), .RST(rst), .I(g_init[611]), 
        .Q(mreg[611]) );
  DFF \mreg_reg[610]  ( .D(mreg[610]), .CLK(clk), .RST(rst), .I(g_init[610]), 
        .Q(mreg[610]) );
  DFF \mreg_reg[609]  ( .D(mreg[609]), .CLK(clk), .RST(rst), .I(g_init[609]), 
        .Q(mreg[609]) );
  DFF \mreg_reg[608]  ( .D(mreg[608]), .CLK(clk), .RST(rst), .I(g_init[608]), 
        .Q(mreg[608]) );
  DFF \mreg_reg[607]  ( .D(mreg[607]), .CLK(clk), .RST(rst), .I(g_init[607]), 
        .Q(mreg[607]) );
  DFF \mreg_reg[606]  ( .D(mreg[606]), .CLK(clk), .RST(rst), .I(g_init[606]), 
        .Q(mreg[606]) );
  DFF \mreg_reg[605]  ( .D(mreg[605]), .CLK(clk), .RST(rst), .I(g_init[605]), 
        .Q(mreg[605]) );
  DFF \mreg_reg[604]  ( .D(mreg[604]), .CLK(clk), .RST(rst), .I(g_init[604]), 
        .Q(mreg[604]) );
  DFF \mreg_reg[603]  ( .D(mreg[603]), .CLK(clk), .RST(rst), .I(g_init[603]), 
        .Q(mreg[603]) );
  DFF \mreg_reg[602]  ( .D(mreg[602]), .CLK(clk), .RST(rst), .I(g_init[602]), 
        .Q(mreg[602]) );
  DFF \mreg_reg[601]  ( .D(mreg[601]), .CLK(clk), .RST(rst), .I(g_init[601]), 
        .Q(mreg[601]) );
  DFF \mreg_reg[600]  ( .D(mreg[600]), .CLK(clk), .RST(rst), .I(g_init[600]), 
        .Q(mreg[600]) );
  DFF \mreg_reg[599]  ( .D(mreg[599]), .CLK(clk), .RST(rst), .I(g_init[599]), 
        .Q(mreg[599]) );
  DFF \mreg_reg[598]  ( .D(mreg[598]), .CLK(clk), .RST(rst), .I(g_init[598]), 
        .Q(mreg[598]) );
  DFF \mreg_reg[597]  ( .D(mreg[597]), .CLK(clk), .RST(rst), .I(g_init[597]), 
        .Q(mreg[597]) );
  DFF \mreg_reg[596]  ( .D(mreg[596]), .CLK(clk), .RST(rst), .I(g_init[596]), 
        .Q(mreg[596]) );
  DFF \mreg_reg[595]  ( .D(mreg[595]), .CLK(clk), .RST(rst), .I(g_init[595]), 
        .Q(mreg[595]) );
  DFF \mreg_reg[594]  ( .D(mreg[594]), .CLK(clk), .RST(rst), .I(g_init[594]), 
        .Q(mreg[594]) );
  DFF \mreg_reg[593]  ( .D(mreg[593]), .CLK(clk), .RST(rst), .I(g_init[593]), 
        .Q(mreg[593]) );
  DFF \mreg_reg[592]  ( .D(mreg[592]), .CLK(clk), .RST(rst), .I(g_init[592]), 
        .Q(mreg[592]) );
  DFF \mreg_reg[591]  ( .D(mreg[591]), .CLK(clk), .RST(rst), .I(g_init[591]), 
        .Q(mreg[591]) );
  DFF \mreg_reg[590]  ( .D(mreg[590]), .CLK(clk), .RST(rst), .I(g_init[590]), 
        .Q(mreg[590]) );
  DFF \mreg_reg[589]  ( .D(mreg[589]), .CLK(clk), .RST(rst), .I(g_init[589]), 
        .Q(mreg[589]) );
  DFF \mreg_reg[588]  ( .D(mreg[588]), .CLK(clk), .RST(rst), .I(g_init[588]), 
        .Q(mreg[588]) );
  DFF \mreg_reg[587]  ( .D(mreg[587]), .CLK(clk), .RST(rst), .I(g_init[587]), 
        .Q(mreg[587]) );
  DFF \mreg_reg[586]  ( .D(mreg[586]), .CLK(clk), .RST(rst), .I(g_init[586]), 
        .Q(mreg[586]) );
  DFF \mreg_reg[585]  ( .D(mreg[585]), .CLK(clk), .RST(rst), .I(g_init[585]), 
        .Q(mreg[585]) );
  DFF \mreg_reg[584]  ( .D(mreg[584]), .CLK(clk), .RST(rst), .I(g_init[584]), 
        .Q(mreg[584]) );
  DFF \mreg_reg[583]  ( .D(mreg[583]), .CLK(clk), .RST(rst), .I(g_init[583]), 
        .Q(mreg[583]) );
  DFF \mreg_reg[582]  ( .D(mreg[582]), .CLK(clk), .RST(rst), .I(g_init[582]), 
        .Q(mreg[582]) );
  DFF \mreg_reg[581]  ( .D(mreg[581]), .CLK(clk), .RST(rst), .I(g_init[581]), 
        .Q(mreg[581]) );
  DFF \mreg_reg[580]  ( .D(mreg[580]), .CLK(clk), .RST(rst), .I(g_init[580]), 
        .Q(mreg[580]) );
  DFF \mreg_reg[579]  ( .D(mreg[579]), .CLK(clk), .RST(rst), .I(g_init[579]), 
        .Q(mreg[579]) );
  DFF \mreg_reg[578]  ( .D(mreg[578]), .CLK(clk), .RST(rst), .I(g_init[578]), 
        .Q(mreg[578]) );
  DFF \mreg_reg[577]  ( .D(mreg[577]), .CLK(clk), .RST(rst), .I(g_init[577]), 
        .Q(mreg[577]) );
  DFF \mreg_reg[576]  ( .D(mreg[576]), .CLK(clk), .RST(rst), .I(g_init[576]), 
        .Q(mreg[576]) );
  DFF \mreg_reg[575]  ( .D(mreg[575]), .CLK(clk), .RST(rst), .I(g_init[575]), 
        .Q(mreg[575]) );
  DFF \mreg_reg[574]  ( .D(mreg[574]), .CLK(clk), .RST(rst), .I(g_init[574]), 
        .Q(mreg[574]) );
  DFF \mreg_reg[573]  ( .D(mreg[573]), .CLK(clk), .RST(rst), .I(g_init[573]), 
        .Q(mreg[573]) );
  DFF \mreg_reg[572]  ( .D(mreg[572]), .CLK(clk), .RST(rst), .I(g_init[572]), 
        .Q(mreg[572]) );
  DFF \mreg_reg[571]  ( .D(mreg[571]), .CLK(clk), .RST(rst), .I(g_init[571]), 
        .Q(mreg[571]) );
  DFF \mreg_reg[570]  ( .D(mreg[570]), .CLK(clk), .RST(rst), .I(g_init[570]), 
        .Q(mreg[570]) );
  DFF \mreg_reg[569]  ( .D(mreg[569]), .CLK(clk), .RST(rst), .I(g_init[569]), 
        .Q(mreg[569]) );
  DFF \mreg_reg[568]  ( .D(mreg[568]), .CLK(clk), .RST(rst), .I(g_init[568]), 
        .Q(mreg[568]) );
  DFF \mreg_reg[567]  ( .D(mreg[567]), .CLK(clk), .RST(rst), .I(g_init[567]), 
        .Q(mreg[567]) );
  DFF \mreg_reg[566]  ( .D(mreg[566]), .CLK(clk), .RST(rst), .I(g_init[566]), 
        .Q(mreg[566]) );
  DFF \mreg_reg[565]  ( .D(mreg[565]), .CLK(clk), .RST(rst), .I(g_init[565]), 
        .Q(mreg[565]) );
  DFF \mreg_reg[564]  ( .D(mreg[564]), .CLK(clk), .RST(rst), .I(g_init[564]), 
        .Q(mreg[564]) );
  DFF \mreg_reg[563]  ( .D(mreg[563]), .CLK(clk), .RST(rst), .I(g_init[563]), 
        .Q(mreg[563]) );
  DFF \mreg_reg[562]  ( .D(mreg[562]), .CLK(clk), .RST(rst), .I(g_init[562]), 
        .Q(mreg[562]) );
  DFF \mreg_reg[561]  ( .D(mreg[561]), .CLK(clk), .RST(rst), .I(g_init[561]), 
        .Q(mreg[561]) );
  DFF \mreg_reg[560]  ( .D(mreg[560]), .CLK(clk), .RST(rst), .I(g_init[560]), 
        .Q(mreg[560]) );
  DFF \mreg_reg[559]  ( .D(mreg[559]), .CLK(clk), .RST(rst), .I(g_init[559]), 
        .Q(mreg[559]) );
  DFF \mreg_reg[558]  ( .D(mreg[558]), .CLK(clk), .RST(rst), .I(g_init[558]), 
        .Q(mreg[558]) );
  DFF \mreg_reg[557]  ( .D(mreg[557]), .CLK(clk), .RST(rst), .I(g_init[557]), 
        .Q(mreg[557]) );
  DFF \mreg_reg[556]  ( .D(mreg[556]), .CLK(clk), .RST(rst), .I(g_init[556]), 
        .Q(mreg[556]) );
  DFF \mreg_reg[555]  ( .D(mreg[555]), .CLK(clk), .RST(rst), .I(g_init[555]), 
        .Q(mreg[555]) );
  DFF \mreg_reg[554]  ( .D(mreg[554]), .CLK(clk), .RST(rst), .I(g_init[554]), 
        .Q(mreg[554]) );
  DFF \mreg_reg[553]  ( .D(mreg[553]), .CLK(clk), .RST(rst), .I(g_init[553]), 
        .Q(mreg[553]) );
  DFF \mreg_reg[552]  ( .D(mreg[552]), .CLK(clk), .RST(rst), .I(g_init[552]), 
        .Q(mreg[552]) );
  DFF \mreg_reg[551]  ( .D(mreg[551]), .CLK(clk), .RST(rst), .I(g_init[551]), 
        .Q(mreg[551]) );
  DFF \mreg_reg[550]  ( .D(mreg[550]), .CLK(clk), .RST(rst), .I(g_init[550]), 
        .Q(mreg[550]) );
  DFF \mreg_reg[549]  ( .D(mreg[549]), .CLK(clk), .RST(rst), .I(g_init[549]), 
        .Q(mreg[549]) );
  DFF \mreg_reg[548]  ( .D(mreg[548]), .CLK(clk), .RST(rst), .I(g_init[548]), 
        .Q(mreg[548]) );
  DFF \mreg_reg[547]  ( .D(mreg[547]), .CLK(clk), .RST(rst), .I(g_init[547]), 
        .Q(mreg[547]) );
  DFF \mreg_reg[546]  ( .D(mreg[546]), .CLK(clk), .RST(rst), .I(g_init[546]), 
        .Q(mreg[546]) );
  DFF \mreg_reg[545]  ( .D(mreg[545]), .CLK(clk), .RST(rst), .I(g_init[545]), 
        .Q(mreg[545]) );
  DFF \mreg_reg[544]  ( .D(mreg[544]), .CLK(clk), .RST(rst), .I(g_init[544]), 
        .Q(mreg[544]) );
  DFF \mreg_reg[543]  ( .D(mreg[543]), .CLK(clk), .RST(rst), .I(g_init[543]), 
        .Q(mreg[543]) );
  DFF \mreg_reg[542]  ( .D(mreg[542]), .CLK(clk), .RST(rst), .I(g_init[542]), 
        .Q(mreg[542]) );
  DFF \mreg_reg[541]  ( .D(mreg[541]), .CLK(clk), .RST(rst), .I(g_init[541]), 
        .Q(mreg[541]) );
  DFF \mreg_reg[540]  ( .D(mreg[540]), .CLK(clk), .RST(rst), .I(g_init[540]), 
        .Q(mreg[540]) );
  DFF \mreg_reg[539]  ( .D(mreg[539]), .CLK(clk), .RST(rst), .I(g_init[539]), 
        .Q(mreg[539]) );
  DFF \mreg_reg[538]  ( .D(mreg[538]), .CLK(clk), .RST(rst), .I(g_init[538]), 
        .Q(mreg[538]) );
  DFF \mreg_reg[537]  ( .D(mreg[537]), .CLK(clk), .RST(rst), .I(g_init[537]), 
        .Q(mreg[537]) );
  DFF \mreg_reg[536]  ( .D(mreg[536]), .CLK(clk), .RST(rst), .I(g_init[536]), 
        .Q(mreg[536]) );
  DFF \mreg_reg[535]  ( .D(mreg[535]), .CLK(clk), .RST(rst), .I(g_init[535]), 
        .Q(mreg[535]) );
  DFF \mreg_reg[534]  ( .D(mreg[534]), .CLK(clk), .RST(rst), .I(g_init[534]), 
        .Q(mreg[534]) );
  DFF \mreg_reg[533]  ( .D(mreg[533]), .CLK(clk), .RST(rst), .I(g_init[533]), 
        .Q(mreg[533]) );
  DFF \mreg_reg[532]  ( .D(mreg[532]), .CLK(clk), .RST(rst), .I(g_init[532]), 
        .Q(mreg[532]) );
  DFF \mreg_reg[531]  ( .D(mreg[531]), .CLK(clk), .RST(rst), .I(g_init[531]), 
        .Q(mreg[531]) );
  DFF \mreg_reg[530]  ( .D(mreg[530]), .CLK(clk), .RST(rst), .I(g_init[530]), 
        .Q(mreg[530]) );
  DFF \mreg_reg[529]  ( .D(mreg[529]), .CLK(clk), .RST(rst), .I(g_init[529]), 
        .Q(mreg[529]) );
  DFF \mreg_reg[528]  ( .D(mreg[528]), .CLK(clk), .RST(rst), .I(g_init[528]), 
        .Q(mreg[528]) );
  DFF \mreg_reg[527]  ( .D(mreg[527]), .CLK(clk), .RST(rst), .I(g_init[527]), 
        .Q(mreg[527]) );
  DFF \mreg_reg[526]  ( .D(mreg[526]), .CLK(clk), .RST(rst), .I(g_init[526]), 
        .Q(mreg[526]) );
  DFF \mreg_reg[525]  ( .D(mreg[525]), .CLK(clk), .RST(rst), .I(g_init[525]), 
        .Q(mreg[525]) );
  DFF \mreg_reg[524]  ( .D(mreg[524]), .CLK(clk), .RST(rst), .I(g_init[524]), 
        .Q(mreg[524]) );
  DFF \mreg_reg[523]  ( .D(mreg[523]), .CLK(clk), .RST(rst), .I(g_init[523]), 
        .Q(mreg[523]) );
  DFF \mreg_reg[522]  ( .D(mreg[522]), .CLK(clk), .RST(rst), .I(g_init[522]), 
        .Q(mreg[522]) );
  DFF \mreg_reg[521]  ( .D(mreg[521]), .CLK(clk), .RST(rst), .I(g_init[521]), 
        .Q(mreg[521]) );
  DFF \mreg_reg[520]  ( .D(mreg[520]), .CLK(clk), .RST(rst), .I(g_init[520]), 
        .Q(mreg[520]) );
  DFF \mreg_reg[519]  ( .D(mreg[519]), .CLK(clk), .RST(rst), .I(g_init[519]), 
        .Q(mreg[519]) );
  DFF \mreg_reg[518]  ( .D(mreg[518]), .CLK(clk), .RST(rst), .I(g_init[518]), 
        .Q(mreg[518]) );
  DFF \mreg_reg[517]  ( .D(mreg[517]), .CLK(clk), .RST(rst), .I(g_init[517]), 
        .Q(mreg[517]) );
  DFF \mreg_reg[516]  ( .D(mreg[516]), .CLK(clk), .RST(rst), .I(g_init[516]), 
        .Q(mreg[516]) );
  DFF \mreg_reg[515]  ( .D(mreg[515]), .CLK(clk), .RST(rst), .I(g_init[515]), 
        .Q(mreg[515]) );
  DFF \mreg_reg[514]  ( .D(mreg[514]), .CLK(clk), .RST(rst), .I(g_init[514]), 
        .Q(mreg[514]) );
  DFF \mreg_reg[513]  ( .D(mreg[513]), .CLK(clk), .RST(rst), .I(g_init[513]), 
        .Q(mreg[513]) );
  DFF \mreg_reg[512]  ( .D(mreg[512]), .CLK(clk), .RST(rst), .I(g_init[512]), 
        .Q(mreg[512]) );
  DFF \mreg_reg[511]  ( .D(mreg[511]), .CLK(clk), .RST(rst), .I(g_init[511]), 
        .Q(mreg[511]) );
  DFF \mreg_reg[510]  ( .D(mreg[510]), .CLK(clk), .RST(rst), .I(g_init[510]), 
        .Q(mreg[510]) );
  DFF \mreg_reg[509]  ( .D(mreg[509]), .CLK(clk), .RST(rst), .I(g_init[509]), 
        .Q(mreg[509]) );
  DFF \mreg_reg[508]  ( .D(mreg[508]), .CLK(clk), .RST(rst), .I(g_init[508]), 
        .Q(mreg[508]) );
  DFF \mreg_reg[507]  ( .D(mreg[507]), .CLK(clk), .RST(rst), .I(g_init[507]), 
        .Q(mreg[507]) );
  DFF \mreg_reg[506]  ( .D(mreg[506]), .CLK(clk), .RST(rst), .I(g_init[506]), 
        .Q(mreg[506]) );
  DFF \mreg_reg[505]  ( .D(mreg[505]), .CLK(clk), .RST(rst), .I(g_init[505]), 
        .Q(mreg[505]) );
  DFF \mreg_reg[504]  ( .D(mreg[504]), .CLK(clk), .RST(rst), .I(g_init[504]), 
        .Q(mreg[504]) );
  DFF \mreg_reg[503]  ( .D(mreg[503]), .CLK(clk), .RST(rst), .I(g_init[503]), 
        .Q(mreg[503]) );
  DFF \mreg_reg[502]  ( .D(mreg[502]), .CLK(clk), .RST(rst), .I(g_init[502]), 
        .Q(mreg[502]) );
  DFF \mreg_reg[501]  ( .D(mreg[501]), .CLK(clk), .RST(rst), .I(g_init[501]), 
        .Q(mreg[501]) );
  DFF \mreg_reg[500]  ( .D(mreg[500]), .CLK(clk), .RST(rst), .I(g_init[500]), 
        .Q(mreg[500]) );
  DFF \mreg_reg[499]  ( .D(mreg[499]), .CLK(clk), .RST(rst), .I(g_init[499]), 
        .Q(mreg[499]) );
  DFF \mreg_reg[498]  ( .D(mreg[498]), .CLK(clk), .RST(rst), .I(g_init[498]), 
        .Q(mreg[498]) );
  DFF \mreg_reg[497]  ( .D(mreg[497]), .CLK(clk), .RST(rst), .I(g_init[497]), 
        .Q(mreg[497]) );
  DFF \mreg_reg[496]  ( .D(mreg[496]), .CLK(clk), .RST(rst), .I(g_init[496]), 
        .Q(mreg[496]) );
  DFF \mreg_reg[495]  ( .D(mreg[495]), .CLK(clk), .RST(rst), .I(g_init[495]), 
        .Q(mreg[495]) );
  DFF \mreg_reg[494]  ( .D(mreg[494]), .CLK(clk), .RST(rst), .I(g_init[494]), 
        .Q(mreg[494]) );
  DFF \mreg_reg[493]  ( .D(mreg[493]), .CLK(clk), .RST(rst), .I(g_init[493]), 
        .Q(mreg[493]) );
  DFF \mreg_reg[492]  ( .D(mreg[492]), .CLK(clk), .RST(rst), .I(g_init[492]), 
        .Q(mreg[492]) );
  DFF \mreg_reg[491]  ( .D(mreg[491]), .CLK(clk), .RST(rst), .I(g_init[491]), 
        .Q(mreg[491]) );
  DFF \mreg_reg[490]  ( .D(mreg[490]), .CLK(clk), .RST(rst), .I(g_init[490]), 
        .Q(mreg[490]) );
  DFF \mreg_reg[489]  ( .D(mreg[489]), .CLK(clk), .RST(rst), .I(g_init[489]), 
        .Q(mreg[489]) );
  DFF \mreg_reg[488]  ( .D(mreg[488]), .CLK(clk), .RST(rst), .I(g_init[488]), 
        .Q(mreg[488]) );
  DFF \mreg_reg[487]  ( .D(mreg[487]), .CLK(clk), .RST(rst), .I(g_init[487]), 
        .Q(mreg[487]) );
  DFF \mreg_reg[486]  ( .D(mreg[486]), .CLK(clk), .RST(rst), .I(g_init[486]), 
        .Q(mreg[486]) );
  DFF \mreg_reg[485]  ( .D(mreg[485]), .CLK(clk), .RST(rst), .I(g_init[485]), 
        .Q(mreg[485]) );
  DFF \mreg_reg[484]  ( .D(mreg[484]), .CLK(clk), .RST(rst), .I(g_init[484]), 
        .Q(mreg[484]) );
  DFF \mreg_reg[483]  ( .D(mreg[483]), .CLK(clk), .RST(rst), .I(g_init[483]), 
        .Q(mreg[483]) );
  DFF \mreg_reg[482]  ( .D(mreg[482]), .CLK(clk), .RST(rst), .I(g_init[482]), 
        .Q(mreg[482]) );
  DFF \mreg_reg[481]  ( .D(mreg[481]), .CLK(clk), .RST(rst), .I(g_init[481]), 
        .Q(mreg[481]) );
  DFF \mreg_reg[480]  ( .D(mreg[480]), .CLK(clk), .RST(rst), .I(g_init[480]), 
        .Q(mreg[480]) );
  DFF \mreg_reg[479]  ( .D(mreg[479]), .CLK(clk), .RST(rst), .I(g_init[479]), 
        .Q(mreg[479]) );
  DFF \mreg_reg[478]  ( .D(mreg[478]), .CLK(clk), .RST(rst), .I(g_init[478]), 
        .Q(mreg[478]) );
  DFF \mreg_reg[477]  ( .D(mreg[477]), .CLK(clk), .RST(rst), .I(g_init[477]), 
        .Q(mreg[477]) );
  DFF \mreg_reg[476]  ( .D(mreg[476]), .CLK(clk), .RST(rst), .I(g_init[476]), 
        .Q(mreg[476]) );
  DFF \mreg_reg[475]  ( .D(mreg[475]), .CLK(clk), .RST(rst), .I(g_init[475]), 
        .Q(mreg[475]) );
  DFF \mreg_reg[474]  ( .D(mreg[474]), .CLK(clk), .RST(rst), .I(g_init[474]), 
        .Q(mreg[474]) );
  DFF \mreg_reg[473]  ( .D(mreg[473]), .CLK(clk), .RST(rst), .I(g_init[473]), 
        .Q(mreg[473]) );
  DFF \mreg_reg[472]  ( .D(mreg[472]), .CLK(clk), .RST(rst), .I(g_init[472]), 
        .Q(mreg[472]) );
  DFF \mreg_reg[471]  ( .D(mreg[471]), .CLK(clk), .RST(rst), .I(g_init[471]), 
        .Q(mreg[471]) );
  DFF \mreg_reg[470]  ( .D(mreg[470]), .CLK(clk), .RST(rst), .I(g_init[470]), 
        .Q(mreg[470]) );
  DFF \mreg_reg[469]  ( .D(mreg[469]), .CLK(clk), .RST(rst), .I(g_init[469]), 
        .Q(mreg[469]) );
  DFF \mreg_reg[468]  ( .D(mreg[468]), .CLK(clk), .RST(rst), .I(g_init[468]), 
        .Q(mreg[468]) );
  DFF \mreg_reg[467]  ( .D(mreg[467]), .CLK(clk), .RST(rst), .I(g_init[467]), 
        .Q(mreg[467]) );
  DFF \mreg_reg[466]  ( .D(mreg[466]), .CLK(clk), .RST(rst), .I(g_init[466]), 
        .Q(mreg[466]) );
  DFF \mreg_reg[465]  ( .D(mreg[465]), .CLK(clk), .RST(rst), .I(g_init[465]), 
        .Q(mreg[465]) );
  DFF \mreg_reg[464]  ( .D(mreg[464]), .CLK(clk), .RST(rst), .I(g_init[464]), 
        .Q(mreg[464]) );
  DFF \mreg_reg[463]  ( .D(mreg[463]), .CLK(clk), .RST(rst), .I(g_init[463]), 
        .Q(mreg[463]) );
  DFF \mreg_reg[462]  ( .D(mreg[462]), .CLK(clk), .RST(rst), .I(g_init[462]), 
        .Q(mreg[462]) );
  DFF \mreg_reg[461]  ( .D(mreg[461]), .CLK(clk), .RST(rst), .I(g_init[461]), 
        .Q(mreg[461]) );
  DFF \mreg_reg[460]  ( .D(mreg[460]), .CLK(clk), .RST(rst), .I(g_init[460]), 
        .Q(mreg[460]) );
  DFF \mreg_reg[459]  ( .D(mreg[459]), .CLK(clk), .RST(rst), .I(g_init[459]), 
        .Q(mreg[459]) );
  DFF \mreg_reg[458]  ( .D(mreg[458]), .CLK(clk), .RST(rst), .I(g_init[458]), 
        .Q(mreg[458]) );
  DFF \mreg_reg[457]  ( .D(mreg[457]), .CLK(clk), .RST(rst), .I(g_init[457]), 
        .Q(mreg[457]) );
  DFF \mreg_reg[456]  ( .D(mreg[456]), .CLK(clk), .RST(rst), .I(g_init[456]), 
        .Q(mreg[456]) );
  DFF \mreg_reg[455]  ( .D(mreg[455]), .CLK(clk), .RST(rst), .I(g_init[455]), 
        .Q(mreg[455]) );
  DFF \mreg_reg[454]  ( .D(mreg[454]), .CLK(clk), .RST(rst), .I(g_init[454]), 
        .Q(mreg[454]) );
  DFF \mreg_reg[453]  ( .D(mreg[453]), .CLK(clk), .RST(rst), .I(g_init[453]), 
        .Q(mreg[453]) );
  DFF \mreg_reg[452]  ( .D(mreg[452]), .CLK(clk), .RST(rst), .I(g_init[452]), 
        .Q(mreg[452]) );
  DFF \mreg_reg[451]  ( .D(mreg[451]), .CLK(clk), .RST(rst), .I(g_init[451]), 
        .Q(mreg[451]) );
  DFF \mreg_reg[450]  ( .D(mreg[450]), .CLK(clk), .RST(rst), .I(g_init[450]), 
        .Q(mreg[450]) );
  DFF \mreg_reg[449]  ( .D(mreg[449]), .CLK(clk), .RST(rst), .I(g_init[449]), 
        .Q(mreg[449]) );
  DFF \mreg_reg[448]  ( .D(mreg[448]), .CLK(clk), .RST(rst), .I(g_init[448]), 
        .Q(mreg[448]) );
  DFF \mreg_reg[447]  ( .D(mreg[447]), .CLK(clk), .RST(rst), .I(g_init[447]), 
        .Q(mreg[447]) );
  DFF \mreg_reg[446]  ( .D(mreg[446]), .CLK(clk), .RST(rst), .I(g_init[446]), 
        .Q(mreg[446]) );
  DFF \mreg_reg[445]  ( .D(mreg[445]), .CLK(clk), .RST(rst), .I(g_init[445]), 
        .Q(mreg[445]) );
  DFF \mreg_reg[444]  ( .D(mreg[444]), .CLK(clk), .RST(rst), .I(g_init[444]), 
        .Q(mreg[444]) );
  DFF \mreg_reg[443]  ( .D(mreg[443]), .CLK(clk), .RST(rst), .I(g_init[443]), 
        .Q(mreg[443]) );
  DFF \mreg_reg[442]  ( .D(mreg[442]), .CLK(clk), .RST(rst), .I(g_init[442]), 
        .Q(mreg[442]) );
  DFF \mreg_reg[441]  ( .D(mreg[441]), .CLK(clk), .RST(rst), .I(g_init[441]), 
        .Q(mreg[441]) );
  DFF \mreg_reg[440]  ( .D(mreg[440]), .CLK(clk), .RST(rst), .I(g_init[440]), 
        .Q(mreg[440]) );
  DFF \mreg_reg[439]  ( .D(mreg[439]), .CLK(clk), .RST(rst), .I(g_init[439]), 
        .Q(mreg[439]) );
  DFF \mreg_reg[438]  ( .D(mreg[438]), .CLK(clk), .RST(rst), .I(g_init[438]), 
        .Q(mreg[438]) );
  DFF \mreg_reg[437]  ( .D(mreg[437]), .CLK(clk), .RST(rst), .I(g_init[437]), 
        .Q(mreg[437]) );
  DFF \mreg_reg[436]  ( .D(mreg[436]), .CLK(clk), .RST(rst), .I(g_init[436]), 
        .Q(mreg[436]) );
  DFF \mreg_reg[435]  ( .D(mreg[435]), .CLK(clk), .RST(rst), .I(g_init[435]), 
        .Q(mreg[435]) );
  DFF \mreg_reg[434]  ( .D(mreg[434]), .CLK(clk), .RST(rst), .I(g_init[434]), 
        .Q(mreg[434]) );
  DFF \mreg_reg[433]  ( .D(mreg[433]), .CLK(clk), .RST(rst), .I(g_init[433]), 
        .Q(mreg[433]) );
  DFF \mreg_reg[432]  ( .D(mreg[432]), .CLK(clk), .RST(rst), .I(g_init[432]), 
        .Q(mreg[432]) );
  DFF \mreg_reg[431]  ( .D(mreg[431]), .CLK(clk), .RST(rst), .I(g_init[431]), 
        .Q(mreg[431]) );
  DFF \mreg_reg[430]  ( .D(mreg[430]), .CLK(clk), .RST(rst), .I(g_init[430]), 
        .Q(mreg[430]) );
  DFF \mreg_reg[429]  ( .D(mreg[429]), .CLK(clk), .RST(rst), .I(g_init[429]), 
        .Q(mreg[429]) );
  DFF \mreg_reg[428]  ( .D(mreg[428]), .CLK(clk), .RST(rst), .I(g_init[428]), 
        .Q(mreg[428]) );
  DFF \mreg_reg[427]  ( .D(mreg[427]), .CLK(clk), .RST(rst), .I(g_init[427]), 
        .Q(mreg[427]) );
  DFF \mreg_reg[426]  ( .D(mreg[426]), .CLK(clk), .RST(rst), .I(g_init[426]), 
        .Q(mreg[426]) );
  DFF \mreg_reg[425]  ( .D(mreg[425]), .CLK(clk), .RST(rst), .I(g_init[425]), 
        .Q(mreg[425]) );
  DFF \mreg_reg[424]  ( .D(mreg[424]), .CLK(clk), .RST(rst), .I(g_init[424]), 
        .Q(mreg[424]) );
  DFF \mreg_reg[423]  ( .D(mreg[423]), .CLK(clk), .RST(rst), .I(g_init[423]), 
        .Q(mreg[423]) );
  DFF \mreg_reg[422]  ( .D(mreg[422]), .CLK(clk), .RST(rst), .I(g_init[422]), 
        .Q(mreg[422]) );
  DFF \mreg_reg[421]  ( .D(mreg[421]), .CLK(clk), .RST(rst), .I(g_init[421]), 
        .Q(mreg[421]) );
  DFF \mreg_reg[420]  ( .D(mreg[420]), .CLK(clk), .RST(rst), .I(g_init[420]), 
        .Q(mreg[420]) );
  DFF \mreg_reg[419]  ( .D(mreg[419]), .CLK(clk), .RST(rst), .I(g_init[419]), 
        .Q(mreg[419]) );
  DFF \mreg_reg[418]  ( .D(mreg[418]), .CLK(clk), .RST(rst), .I(g_init[418]), 
        .Q(mreg[418]) );
  DFF \mreg_reg[417]  ( .D(mreg[417]), .CLK(clk), .RST(rst), .I(g_init[417]), 
        .Q(mreg[417]) );
  DFF \mreg_reg[416]  ( .D(mreg[416]), .CLK(clk), .RST(rst), .I(g_init[416]), 
        .Q(mreg[416]) );
  DFF \mreg_reg[415]  ( .D(mreg[415]), .CLK(clk), .RST(rst), .I(g_init[415]), 
        .Q(mreg[415]) );
  DFF \mreg_reg[414]  ( .D(mreg[414]), .CLK(clk), .RST(rst), .I(g_init[414]), 
        .Q(mreg[414]) );
  DFF \mreg_reg[413]  ( .D(mreg[413]), .CLK(clk), .RST(rst), .I(g_init[413]), 
        .Q(mreg[413]) );
  DFF \mreg_reg[412]  ( .D(mreg[412]), .CLK(clk), .RST(rst), .I(g_init[412]), 
        .Q(mreg[412]) );
  DFF \mreg_reg[411]  ( .D(mreg[411]), .CLK(clk), .RST(rst), .I(g_init[411]), 
        .Q(mreg[411]) );
  DFF \mreg_reg[410]  ( .D(mreg[410]), .CLK(clk), .RST(rst), .I(g_init[410]), 
        .Q(mreg[410]) );
  DFF \mreg_reg[409]  ( .D(mreg[409]), .CLK(clk), .RST(rst), .I(g_init[409]), 
        .Q(mreg[409]) );
  DFF \mreg_reg[408]  ( .D(mreg[408]), .CLK(clk), .RST(rst), .I(g_init[408]), 
        .Q(mreg[408]) );
  DFF \mreg_reg[407]  ( .D(mreg[407]), .CLK(clk), .RST(rst), .I(g_init[407]), 
        .Q(mreg[407]) );
  DFF \mreg_reg[406]  ( .D(mreg[406]), .CLK(clk), .RST(rst), .I(g_init[406]), 
        .Q(mreg[406]) );
  DFF \mreg_reg[405]  ( .D(mreg[405]), .CLK(clk), .RST(rst), .I(g_init[405]), 
        .Q(mreg[405]) );
  DFF \mreg_reg[404]  ( .D(mreg[404]), .CLK(clk), .RST(rst), .I(g_init[404]), 
        .Q(mreg[404]) );
  DFF \mreg_reg[403]  ( .D(mreg[403]), .CLK(clk), .RST(rst), .I(g_init[403]), 
        .Q(mreg[403]) );
  DFF \mreg_reg[402]  ( .D(mreg[402]), .CLK(clk), .RST(rst), .I(g_init[402]), 
        .Q(mreg[402]) );
  DFF \mreg_reg[401]  ( .D(mreg[401]), .CLK(clk), .RST(rst), .I(g_init[401]), 
        .Q(mreg[401]) );
  DFF \mreg_reg[400]  ( .D(mreg[400]), .CLK(clk), .RST(rst), .I(g_init[400]), 
        .Q(mreg[400]) );
  DFF \mreg_reg[399]  ( .D(mreg[399]), .CLK(clk), .RST(rst), .I(g_init[399]), 
        .Q(mreg[399]) );
  DFF \mreg_reg[398]  ( .D(mreg[398]), .CLK(clk), .RST(rst), .I(g_init[398]), 
        .Q(mreg[398]) );
  DFF \mreg_reg[397]  ( .D(mreg[397]), .CLK(clk), .RST(rst), .I(g_init[397]), 
        .Q(mreg[397]) );
  DFF \mreg_reg[396]  ( .D(mreg[396]), .CLK(clk), .RST(rst), .I(g_init[396]), 
        .Q(mreg[396]) );
  DFF \mreg_reg[395]  ( .D(mreg[395]), .CLK(clk), .RST(rst), .I(g_init[395]), 
        .Q(mreg[395]) );
  DFF \mreg_reg[394]  ( .D(mreg[394]), .CLK(clk), .RST(rst), .I(g_init[394]), 
        .Q(mreg[394]) );
  DFF \mreg_reg[393]  ( .D(mreg[393]), .CLK(clk), .RST(rst), .I(g_init[393]), 
        .Q(mreg[393]) );
  DFF \mreg_reg[392]  ( .D(mreg[392]), .CLK(clk), .RST(rst), .I(g_init[392]), 
        .Q(mreg[392]) );
  DFF \mreg_reg[391]  ( .D(mreg[391]), .CLK(clk), .RST(rst), .I(g_init[391]), 
        .Q(mreg[391]) );
  DFF \mreg_reg[390]  ( .D(mreg[390]), .CLK(clk), .RST(rst), .I(g_init[390]), 
        .Q(mreg[390]) );
  DFF \mreg_reg[389]  ( .D(mreg[389]), .CLK(clk), .RST(rst), .I(g_init[389]), 
        .Q(mreg[389]) );
  DFF \mreg_reg[388]  ( .D(mreg[388]), .CLK(clk), .RST(rst), .I(g_init[388]), 
        .Q(mreg[388]) );
  DFF \mreg_reg[387]  ( .D(mreg[387]), .CLK(clk), .RST(rst), .I(g_init[387]), 
        .Q(mreg[387]) );
  DFF \mreg_reg[386]  ( .D(mreg[386]), .CLK(clk), .RST(rst), .I(g_init[386]), 
        .Q(mreg[386]) );
  DFF \mreg_reg[385]  ( .D(mreg[385]), .CLK(clk), .RST(rst), .I(g_init[385]), 
        .Q(mreg[385]) );
  DFF \mreg_reg[384]  ( .D(mreg[384]), .CLK(clk), .RST(rst), .I(g_init[384]), 
        .Q(mreg[384]) );
  DFF \mreg_reg[383]  ( .D(mreg[383]), .CLK(clk), .RST(rst), .I(g_init[383]), 
        .Q(mreg[383]) );
  DFF \mreg_reg[382]  ( .D(mreg[382]), .CLK(clk), .RST(rst), .I(g_init[382]), 
        .Q(mreg[382]) );
  DFF \mreg_reg[381]  ( .D(mreg[381]), .CLK(clk), .RST(rst), .I(g_init[381]), 
        .Q(mreg[381]) );
  DFF \mreg_reg[380]  ( .D(mreg[380]), .CLK(clk), .RST(rst), .I(g_init[380]), 
        .Q(mreg[380]) );
  DFF \mreg_reg[379]  ( .D(mreg[379]), .CLK(clk), .RST(rst), .I(g_init[379]), 
        .Q(mreg[379]) );
  DFF \mreg_reg[378]  ( .D(mreg[378]), .CLK(clk), .RST(rst), .I(g_init[378]), 
        .Q(mreg[378]) );
  DFF \mreg_reg[377]  ( .D(mreg[377]), .CLK(clk), .RST(rst), .I(g_init[377]), 
        .Q(mreg[377]) );
  DFF \mreg_reg[376]  ( .D(mreg[376]), .CLK(clk), .RST(rst), .I(g_init[376]), 
        .Q(mreg[376]) );
  DFF \mreg_reg[375]  ( .D(mreg[375]), .CLK(clk), .RST(rst), .I(g_init[375]), 
        .Q(mreg[375]) );
  DFF \mreg_reg[374]  ( .D(mreg[374]), .CLK(clk), .RST(rst), .I(g_init[374]), 
        .Q(mreg[374]) );
  DFF \mreg_reg[373]  ( .D(mreg[373]), .CLK(clk), .RST(rst), .I(g_init[373]), 
        .Q(mreg[373]) );
  DFF \mreg_reg[372]  ( .D(mreg[372]), .CLK(clk), .RST(rst), .I(g_init[372]), 
        .Q(mreg[372]) );
  DFF \mreg_reg[371]  ( .D(mreg[371]), .CLK(clk), .RST(rst), .I(g_init[371]), 
        .Q(mreg[371]) );
  DFF \mreg_reg[370]  ( .D(mreg[370]), .CLK(clk), .RST(rst), .I(g_init[370]), 
        .Q(mreg[370]) );
  DFF \mreg_reg[369]  ( .D(mreg[369]), .CLK(clk), .RST(rst), .I(g_init[369]), 
        .Q(mreg[369]) );
  DFF \mreg_reg[368]  ( .D(mreg[368]), .CLK(clk), .RST(rst), .I(g_init[368]), 
        .Q(mreg[368]) );
  DFF \mreg_reg[367]  ( .D(mreg[367]), .CLK(clk), .RST(rst), .I(g_init[367]), 
        .Q(mreg[367]) );
  DFF \mreg_reg[366]  ( .D(mreg[366]), .CLK(clk), .RST(rst), .I(g_init[366]), 
        .Q(mreg[366]) );
  DFF \mreg_reg[365]  ( .D(mreg[365]), .CLK(clk), .RST(rst), .I(g_init[365]), 
        .Q(mreg[365]) );
  DFF \mreg_reg[364]  ( .D(mreg[364]), .CLK(clk), .RST(rst), .I(g_init[364]), 
        .Q(mreg[364]) );
  DFF \mreg_reg[363]  ( .D(mreg[363]), .CLK(clk), .RST(rst), .I(g_init[363]), 
        .Q(mreg[363]) );
  DFF \mreg_reg[362]  ( .D(mreg[362]), .CLK(clk), .RST(rst), .I(g_init[362]), 
        .Q(mreg[362]) );
  DFF \mreg_reg[361]  ( .D(mreg[361]), .CLK(clk), .RST(rst), .I(g_init[361]), 
        .Q(mreg[361]) );
  DFF \mreg_reg[360]  ( .D(mreg[360]), .CLK(clk), .RST(rst), .I(g_init[360]), 
        .Q(mreg[360]) );
  DFF \mreg_reg[359]  ( .D(mreg[359]), .CLK(clk), .RST(rst), .I(g_init[359]), 
        .Q(mreg[359]) );
  DFF \mreg_reg[358]  ( .D(mreg[358]), .CLK(clk), .RST(rst), .I(g_init[358]), 
        .Q(mreg[358]) );
  DFF \mreg_reg[357]  ( .D(mreg[357]), .CLK(clk), .RST(rst), .I(g_init[357]), 
        .Q(mreg[357]) );
  DFF \mreg_reg[356]  ( .D(mreg[356]), .CLK(clk), .RST(rst), .I(g_init[356]), 
        .Q(mreg[356]) );
  DFF \mreg_reg[355]  ( .D(mreg[355]), .CLK(clk), .RST(rst), .I(g_init[355]), 
        .Q(mreg[355]) );
  DFF \mreg_reg[354]  ( .D(mreg[354]), .CLK(clk), .RST(rst), .I(g_init[354]), 
        .Q(mreg[354]) );
  DFF \mreg_reg[353]  ( .D(mreg[353]), .CLK(clk), .RST(rst), .I(g_init[353]), 
        .Q(mreg[353]) );
  DFF \mreg_reg[352]  ( .D(mreg[352]), .CLK(clk), .RST(rst), .I(g_init[352]), 
        .Q(mreg[352]) );
  DFF \mreg_reg[351]  ( .D(mreg[351]), .CLK(clk), .RST(rst), .I(g_init[351]), 
        .Q(mreg[351]) );
  DFF \mreg_reg[350]  ( .D(mreg[350]), .CLK(clk), .RST(rst), .I(g_init[350]), 
        .Q(mreg[350]) );
  DFF \mreg_reg[349]  ( .D(mreg[349]), .CLK(clk), .RST(rst), .I(g_init[349]), 
        .Q(mreg[349]) );
  DFF \mreg_reg[348]  ( .D(mreg[348]), .CLK(clk), .RST(rst), .I(g_init[348]), 
        .Q(mreg[348]) );
  DFF \mreg_reg[347]  ( .D(mreg[347]), .CLK(clk), .RST(rst), .I(g_init[347]), 
        .Q(mreg[347]) );
  DFF \mreg_reg[346]  ( .D(mreg[346]), .CLK(clk), .RST(rst), .I(g_init[346]), 
        .Q(mreg[346]) );
  DFF \mreg_reg[345]  ( .D(mreg[345]), .CLK(clk), .RST(rst), .I(g_init[345]), 
        .Q(mreg[345]) );
  DFF \mreg_reg[344]  ( .D(mreg[344]), .CLK(clk), .RST(rst), .I(g_init[344]), 
        .Q(mreg[344]) );
  DFF \mreg_reg[343]  ( .D(mreg[343]), .CLK(clk), .RST(rst), .I(g_init[343]), 
        .Q(mreg[343]) );
  DFF \mreg_reg[342]  ( .D(mreg[342]), .CLK(clk), .RST(rst), .I(g_init[342]), 
        .Q(mreg[342]) );
  DFF \mreg_reg[341]  ( .D(mreg[341]), .CLK(clk), .RST(rst), .I(g_init[341]), 
        .Q(mreg[341]) );
  DFF \mreg_reg[340]  ( .D(mreg[340]), .CLK(clk), .RST(rst), .I(g_init[340]), 
        .Q(mreg[340]) );
  DFF \mreg_reg[339]  ( .D(mreg[339]), .CLK(clk), .RST(rst), .I(g_init[339]), 
        .Q(mreg[339]) );
  DFF \mreg_reg[338]  ( .D(mreg[338]), .CLK(clk), .RST(rst), .I(g_init[338]), 
        .Q(mreg[338]) );
  DFF \mreg_reg[337]  ( .D(mreg[337]), .CLK(clk), .RST(rst), .I(g_init[337]), 
        .Q(mreg[337]) );
  DFF \mreg_reg[336]  ( .D(mreg[336]), .CLK(clk), .RST(rst), .I(g_init[336]), 
        .Q(mreg[336]) );
  DFF \mreg_reg[335]  ( .D(mreg[335]), .CLK(clk), .RST(rst), .I(g_init[335]), 
        .Q(mreg[335]) );
  DFF \mreg_reg[334]  ( .D(mreg[334]), .CLK(clk), .RST(rst), .I(g_init[334]), 
        .Q(mreg[334]) );
  DFF \mreg_reg[333]  ( .D(mreg[333]), .CLK(clk), .RST(rst), .I(g_init[333]), 
        .Q(mreg[333]) );
  DFF \mreg_reg[332]  ( .D(mreg[332]), .CLK(clk), .RST(rst), .I(g_init[332]), 
        .Q(mreg[332]) );
  DFF \mreg_reg[331]  ( .D(mreg[331]), .CLK(clk), .RST(rst), .I(g_init[331]), 
        .Q(mreg[331]) );
  DFF \mreg_reg[330]  ( .D(mreg[330]), .CLK(clk), .RST(rst), .I(g_init[330]), 
        .Q(mreg[330]) );
  DFF \mreg_reg[329]  ( .D(mreg[329]), .CLK(clk), .RST(rst), .I(g_init[329]), 
        .Q(mreg[329]) );
  DFF \mreg_reg[328]  ( .D(mreg[328]), .CLK(clk), .RST(rst), .I(g_init[328]), 
        .Q(mreg[328]) );
  DFF \mreg_reg[327]  ( .D(mreg[327]), .CLK(clk), .RST(rst), .I(g_init[327]), 
        .Q(mreg[327]) );
  DFF \mreg_reg[326]  ( .D(mreg[326]), .CLK(clk), .RST(rst), .I(g_init[326]), 
        .Q(mreg[326]) );
  DFF \mreg_reg[325]  ( .D(mreg[325]), .CLK(clk), .RST(rst), .I(g_init[325]), 
        .Q(mreg[325]) );
  DFF \mreg_reg[324]  ( .D(mreg[324]), .CLK(clk), .RST(rst), .I(g_init[324]), 
        .Q(mreg[324]) );
  DFF \mreg_reg[323]  ( .D(mreg[323]), .CLK(clk), .RST(rst), .I(g_init[323]), 
        .Q(mreg[323]) );
  DFF \mreg_reg[322]  ( .D(mreg[322]), .CLK(clk), .RST(rst), .I(g_init[322]), 
        .Q(mreg[322]) );
  DFF \mreg_reg[321]  ( .D(mreg[321]), .CLK(clk), .RST(rst), .I(g_init[321]), 
        .Q(mreg[321]) );
  DFF \mreg_reg[320]  ( .D(mreg[320]), .CLK(clk), .RST(rst), .I(g_init[320]), 
        .Q(mreg[320]) );
  DFF \mreg_reg[319]  ( .D(mreg[319]), .CLK(clk), .RST(rst), .I(g_init[319]), 
        .Q(mreg[319]) );
  DFF \mreg_reg[318]  ( .D(mreg[318]), .CLK(clk), .RST(rst), .I(g_init[318]), 
        .Q(mreg[318]) );
  DFF \mreg_reg[317]  ( .D(mreg[317]), .CLK(clk), .RST(rst), .I(g_init[317]), 
        .Q(mreg[317]) );
  DFF \mreg_reg[316]  ( .D(mreg[316]), .CLK(clk), .RST(rst), .I(g_init[316]), 
        .Q(mreg[316]) );
  DFF \mreg_reg[315]  ( .D(mreg[315]), .CLK(clk), .RST(rst), .I(g_init[315]), 
        .Q(mreg[315]) );
  DFF \mreg_reg[314]  ( .D(mreg[314]), .CLK(clk), .RST(rst), .I(g_init[314]), 
        .Q(mreg[314]) );
  DFF \mreg_reg[313]  ( .D(mreg[313]), .CLK(clk), .RST(rst), .I(g_init[313]), 
        .Q(mreg[313]) );
  DFF \mreg_reg[312]  ( .D(mreg[312]), .CLK(clk), .RST(rst), .I(g_init[312]), 
        .Q(mreg[312]) );
  DFF \mreg_reg[311]  ( .D(mreg[311]), .CLK(clk), .RST(rst), .I(g_init[311]), 
        .Q(mreg[311]) );
  DFF \mreg_reg[310]  ( .D(mreg[310]), .CLK(clk), .RST(rst), .I(g_init[310]), 
        .Q(mreg[310]) );
  DFF \mreg_reg[309]  ( .D(mreg[309]), .CLK(clk), .RST(rst), .I(g_init[309]), 
        .Q(mreg[309]) );
  DFF \mreg_reg[308]  ( .D(mreg[308]), .CLK(clk), .RST(rst), .I(g_init[308]), 
        .Q(mreg[308]) );
  DFF \mreg_reg[307]  ( .D(mreg[307]), .CLK(clk), .RST(rst), .I(g_init[307]), 
        .Q(mreg[307]) );
  DFF \mreg_reg[306]  ( .D(mreg[306]), .CLK(clk), .RST(rst), .I(g_init[306]), 
        .Q(mreg[306]) );
  DFF \mreg_reg[305]  ( .D(mreg[305]), .CLK(clk), .RST(rst), .I(g_init[305]), 
        .Q(mreg[305]) );
  DFF \mreg_reg[304]  ( .D(mreg[304]), .CLK(clk), .RST(rst), .I(g_init[304]), 
        .Q(mreg[304]) );
  DFF \mreg_reg[303]  ( .D(mreg[303]), .CLK(clk), .RST(rst), .I(g_init[303]), 
        .Q(mreg[303]) );
  DFF \mreg_reg[302]  ( .D(mreg[302]), .CLK(clk), .RST(rst), .I(g_init[302]), 
        .Q(mreg[302]) );
  DFF \mreg_reg[301]  ( .D(mreg[301]), .CLK(clk), .RST(rst), .I(g_init[301]), 
        .Q(mreg[301]) );
  DFF \mreg_reg[300]  ( .D(mreg[300]), .CLK(clk), .RST(rst), .I(g_init[300]), 
        .Q(mreg[300]) );
  DFF \mreg_reg[299]  ( .D(mreg[299]), .CLK(clk), .RST(rst), .I(g_init[299]), 
        .Q(mreg[299]) );
  DFF \mreg_reg[298]  ( .D(mreg[298]), .CLK(clk), .RST(rst), .I(g_init[298]), 
        .Q(mreg[298]) );
  DFF \mreg_reg[297]  ( .D(mreg[297]), .CLK(clk), .RST(rst), .I(g_init[297]), 
        .Q(mreg[297]) );
  DFF \mreg_reg[296]  ( .D(mreg[296]), .CLK(clk), .RST(rst), .I(g_init[296]), 
        .Q(mreg[296]) );
  DFF \mreg_reg[295]  ( .D(mreg[295]), .CLK(clk), .RST(rst), .I(g_init[295]), 
        .Q(mreg[295]) );
  DFF \mreg_reg[294]  ( .D(mreg[294]), .CLK(clk), .RST(rst), .I(g_init[294]), 
        .Q(mreg[294]) );
  DFF \mreg_reg[293]  ( .D(mreg[293]), .CLK(clk), .RST(rst), .I(g_init[293]), 
        .Q(mreg[293]) );
  DFF \mreg_reg[292]  ( .D(mreg[292]), .CLK(clk), .RST(rst), .I(g_init[292]), 
        .Q(mreg[292]) );
  DFF \mreg_reg[291]  ( .D(mreg[291]), .CLK(clk), .RST(rst), .I(g_init[291]), 
        .Q(mreg[291]) );
  DFF \mreg_reg[290]  ( .D(mreg[290]), .CLK(clk), .RST(rst), .I(g_init[290]), 
        .Q(mreg[290]) );
  DFF \mreg_reg[289]  ( .D(mreg[289]), .CLK(clk), .RST(rst), .I(g_init[289]), 
        .Q(mreg[289]) );
  DFF \mreg_reg[288]  ( .D(mreg[288]), .CLK(clk), .RST(rst), .I(g_init[288]), 
        .Q(mreg[288]) );
  DFF \mreg_reg[287]  ( .D(mreg[287]), .CLK(clk), .RST(rst), .I(g_init[287]), 
        .Q(mreg[287]) );
  DFF \mreg_reg[286]  ( .D(mreg[286]), .CLK(clk), .RST(rst), .I(g_init[286]), 
        .Q(mreg[286]) );
  DFF \mreg_reg[285]  ( .D(mreg[285]), .CLK(clk), .RST(rst), .I(g_init[285]), 
        .Q(mreg[285]) );
  DFF \mreg_reg[284]  ( .D(mreg[284]), .CLK(clk), .RST(rst), .I(g_init[284]), 
        .Q(mreg[284]) );
  DFF \mreg_reg[283]  ( .D(mreg[283]), .CLK(clk), .RST(rst), .I(g_init[283]), 
        .Q(mreg[283]) );
  DFF \mreg_reg[282]  ( .D(mreg[282]), .CLK(clk), .RST(rst), .I(g_init[282]), 
        .Q(mreg[282]) );
  DFF \mreg_reg[281]  ( .D(mreg[281]), .CLK(clk), .RST(rst), .I(g_init[281]), 
        .Q(mreg[281]) );
  DFF \mreg_reg[280]  ( .D(mreg[280]), .CLK(clk), .RST(rst), .I(g_init[280]), 
        .Q(mreg[280]) );
  DFF \mreg_reg[279]  ( .D(mreg[279]), .CLK(clk), .RST(rst), .I(g_init[279]), 
        .Q(mreg[279]) );
  DFF \mreg_reg[278]  ( .D(mreg[278]), .CLK(clk), .RST(rst), .I(g_init[278]), 
        .Q(mreg[278]) );
  DFF \mreg_reg[277]  ( .D(mreg[277]), .CLK(clk), .RST(rst), .I(g_init[277]), 
        .Q(mreg[277]) );
  DFF \mreg_reg[276]  ( .D(mreg[276]), .CLK(clk), .RST(rst), .I(g_init[276]), 
        .Q(mreg[276]) );
  DFF \mreg_reg[275]  ( .D(mreg[275]), .CLK(clk), .RST(rst), .I(g_init[275]), 
        .Q(mreg[275]) );
  DFF \mreg_reg[274]  ( .D(mreg[274]), .CLK(clk), .RST(rst), .I(g_init[274]), 
        .Q(mreg[274]) );
  DFF \mreg_reg[273]  ( .D(mreg[273]), .CLK(clk), .RST(rst), .I(g_init[273]), 
        .Q(mreg[273]) );
  DFF \mreg_reg[272]  ( .D(mreg[272]), .CLK(clk), .RST(rst), .I(g_init[272]), 
        .Q(mreg[272]) );
  DFF \mreg_reg[271]  ( .D(mreg[271]), .CLK(clk), .RST(rst), .I(g_init[271]), 
        .Q(mreg[271]) );
  DFF \mreg_reg[270]  ( .D(mreg[270]), .CLK(clk), .RST(rst), .I(g_init[270]), 
        .Q(mreg[270]) );
  DFF \mreg_reg[269]  ( .D(mreg[269]), .CLK(clk), .RST(rst), .I(g_init[269]), 
        .Q(mreg[269]) );
  DFF \mreg_reg[268]  ( .D(mreg[268]), .CLK(clk), .RST(rst), .I(g_init[268]), 
        .Q(mreg[268]) );
  DFF \mreg_reg[267]  ( .D(mreg[267]), .CLK(clk), .RST(rst), .I(g_init[267]), 
        .Q(mreg[267]) );
  DFF \mreg_reg[266]  ( .D(mreg[266]), .CLK(clk), .RST(rst), .I(g_init[266]), 
        .Q(mreg[266]) );
  DFF \mreg_reg[265]  ( .D(mreg[265]), .CLK(clk), .RST(rst), .I(g_init[265]), 
        .Q(mreg[265]) );
  DFF \mreg_reg[264]  ( .D(mreg[264]), .CLK(clk), .RST(rst), .I(g_init[264]), 
        .Q(mreg[264]) );
  DFF \mreg_reg[263]  ( .D(mreg[263]), .CLK(clk), .RST(rst), .I(g_init[263]), 
        .Q(mreg[263]) );
  DFF \mreg_reg[262]  ( .D(mreg[262]), .CLK(clk), .RST(rst), .I(g_init[262]), 
        .Q(mreg[262]) );
  DFF \mreg_reg[261]  ( .D(mreg[261]), .CLK(clk), .RST(rst), .I(g_init[261]), 
        .Q(mreg[261]) );
  DFF \mreg_reg[260]  ( .D(mreg[260]), .CLK(clk), .RST(rst), .I(g_init[260]), 
        .Q(mreg[260]) );
  DFF \mreg_reg[259]  ( .D(mreg[259]), .CLK(clk), .RST(rst), .I(g_init[259]), 
        .Q(mreg[259]) );
  DFF \mreg_reg[258]  ( .D(mreg[258]), .CLK(clk), .RST(rst), .I(g_init[258]), 
        .Q(mreg[258]) );
  DFF \mreg_reg[257]  ( .D(mreg[257]), .CLK(clk), .RST(rst), .I(g_init[257]), 
        .Q(mreg[257]) );
  DFF \mreg_reg[256]  ( .D(mreg[256]), .CLK(clk), .RST(rst), .I(g_init[256]), 
        .Q(mreg[256]) );
  DFF \mreg_reg[255]  ( .D(mreg[255]), .CLK(clk), .RST(rst), .I(g_init[255]), 
        .Q(mreg[255]) );
  DFF \mreg_reg[254]  ( .D(mreg[254]), .CLK(clk), .RST(rst), .I(g_init[254]), 
        .Q(mreg[254]) );
  DFF \mreg_reg[253]  ( .D(mreg[253]), .CLK(clk), .RST(rst), .I(g_init[253]), 
        .Q(mreg[253]) );
  DFF \mreg_reg[252]  ( .D(mreg[252]), .CLK(clk), .RST(rst), .I(g_init[252]), 
        .Q(mreg[252]) );
  DFF \mreg_reg[251]  ( .D(mreg[251]), .CLK(clk), .RST(rst), .I(g_init[251]), 
        .Q(mreg[251]) );
  DFF \mreg_reg[250]  ( .D(mreg[250]), .CLK(clk), .RST(rst), .I(g_init[250]), 
        .Q(mreg[250]) );
  DFF \mreg_reg[249]  ( .D(mreg[249]), .CLK(clk), .RST(rst), .I(g_init[249]), 
        .Q(mreg[249]) );
  DFF \mreg_reg[248]  ( .D(mreg[248]), .CLK(clk), .RST(rst), .I(g_init[248]), 
        .Q(mreg[248]) );
  DFF \mreg_reg[247]  ( .D(mreg[247]), .CLK(clk), .RST(rst), .I(g_init[247]), 
        .Q(mreg[247]) );
  DFF \mreg_reg[246]  ( .D(mreg[246]), .CLK(clk), .RST(rst), .I(g_init[246]), 
        .Q(mreg[246]) );
  DFF \mreg_reg[245]  ( .D(mreg[245]), .CLK(clk), .RST(rst), .I(g_init[245]), 
        .Q(mreg[245]) );
  DFF \mreg_reg[244]  ( .D(mreg[244]), .CLK(clk), .RST(rst), .I(g_init[244]), 
        .Q(mreg[244]) );
  DFF \mreg_reg[243]  ( .D(mreg[243]), .CLK(clk), .RST(rst), .I(g_init[243]), 
        .Q(mreg[243]) );
  DFF \mreg_reg[242]  ( .D(mreg[242]), .CLK(clk), .RST(rst), .I(g_init[242]), 
        .Q(mreg[242]) );
  DFF \mreg_reg[241]  ( .D(mreg[241]), .CLK(clk), .RST(rst), .I(g_init[241]), 
        .Q(mreg[241]) );
  DFF \mreg_reg[240]  ( .D(mreg[240]), .CLK(clk), .RST(rst), .I(g_init[240]), 
        .Q(mreg[240]) );
  DFF \mreg_reg[239]  ( .D(mreg[239]), .CLK(clk), .RST(rst), .I(g_init[239]), 
        .Q(mreg[239]) );
  DFF \mreg_reg[238]  ( .D(mreg[238]), .CLK(clk), .RST(rst), .I(g_init[238]), 
        .Q(mreg[238]) );
  DFF \mreg_reg[237]  ( .D(mreg[237]), .CLK(clk), .RST(rst), .I(g_init[237]), 
        .Q(mreg[237]) );
  DFF \mreg_reg[236]  ( .D(mreg[236]), .CLK(clk), .RST(rst), .I(g_init[236]), 
        .Q(mreg[236]) );
  DFF \mreg_reg[235]  ( .D(mreg[235]), .CLK(clk), .RST(rst), .I(g_init[235]), 
        .Q(mreg[235]) );
  DFF \mreg_reg[234]  ( .D(mreg[234]), .CLK(clk), .RST(rst), .I(g_init[234]), 
        .Q(mreg[234]) );
  DFF \mreg_reg[233]  ( .D(mreg[233]), .CLK(clk), .RST(rst), .I(g_init[233]), 
        .Q(mreg[233]) );
  DFF \mreg_reg[232]  ( .D(mreg[232]), .CLK(clk), .RST(rst), .I(g_init[232]), 
        .Q(mreg[232]) );
  DFF \mreg_reg[231]  ( .D(mreg[231]), .CLK(clk), .RST(rst), .I(g_init[231]), 
        .Q(mreg[231]) );
  DFF \mreg_reg[230]  ( .D(mreg[230]), .CLK(clk), .RST(rst), .I(g_init[230]), 
        .Q(mreg[230]) );
  DFF \mreg_reg[229]  ( .D(mreg[229]), .CLK(clk), .RST(rst), .I(g_init[229]), 
        .Q(mreg[229]) );
  DFF \mreg_reg[228]  ( .D(mreg[228]), .CLK(clk), .RST(rst), .I(g_init[228]), 
        .Q(mreg[228]) );
  DFF \mreg_reg[227]  ( .D(mreg[227]), .CLK(clk), .RST(rst), .I(g_init[227]), 
        .Q(mreg[227]) );
  DFF \mreg_reg[226]  ( .D(mreg[226]), .CLK(clk), .RST(rst), .I(g_init[226]), 
        .Q(mreg[226]) );
  DFF \mreg_reg[225]  ( .D(mreg[225]), .CLK(clk), .RST(rst), .I(g_init[225]), 
        .Q(mreg[225]) );
  DFF \mreg_reg[224]  ( .D(mreg[224]), .CLK(clk), .RST(rst), .I(g_init[224]), 
        .Q(mreg[224]) );
  DFF \mreg_reg[223]  ( .D(mreg[223]), .CLK(clk), .RST(rst), .I(g_init[223]), 
        .Q(mreg[223]) );
  DFF \mreg_reg[222]  ( .D(mreg[222]), .CLK(clk), .RST(rst), .I(g_init[222]), 
        .Q(mreg[222]) );
  DFF \mreg_reg[221]  ( .D(mreg[221]), .CLK(clk), .RST(rst), .I(g_init[221]), 
        .Q(mreg[221]) );
  DFF \mreg_reg[220]  ( .D(mreg[220]), .CLK(clk), .RST(rst), .I(g_init[220]), 
        .Q(mreg[220]) );
  DFF \mreg_reg[219]  ( .D(mreg[219]), .CLK(clk), .RST(rst), .I(g_init[219]), 
        .Q(mreg[219]) );
  DFF \mreg_reg[218]  ( .D(mreg[218]), .CLK(clk), .RST(rst), .I(g_init[218]), 
        .Q(mreg[218]) );
  DFF \mreg_reg[217]  ( .D(mreg[217]), .CLK(clk), .RST(rst), .I(g_init[217]), 
        .Q(mreg[217]) );
  DFF \mreg_reg[216]  ( .D(mreg[216]), .CLK(clk), .RST(rst), .I(g_init[216]), 
        .Q(mreg[216]) );
  DFF \mreg_reg[215]  ( .D(mreg[215]), .CLK(clk), .RST(rst), .I(g_init[215]), 
        .Q(mreg[215]) );
  DFF \mreg_reg[214]  ( .D(mreg[214]), .CLK(clk), .RST(rst), .I(g_init[214]), 
        .Q(mreg[214]) );
  DFF \mreg_reg[213]  ( .D(mreg[213]), .CLK(clk), .RST(rst), .I(g_init[213]), 
        .Q(mreg[213]) );
  DFF \mreg_reg[212]  ( .D(mreg[212]), .CLK(clk), .RST(rst), .I(g_init[212]), 
        .Q(mreg[212]) );
  DFF \mreg_reg[211]  ( .D(mreg[211]), .CLK(clk), .RST(rst), .I(g_init[211]), 
        .Q(mreg[211]) );
  DFF \mreg_reg[210]  ( .D(mreg[210]), .CLK(clk), .RST(rst), .I(g_init[210]), 
        .Q(mreg[210]) );
  DFF \mreg_reg[209]  ( .D(mreg[209]), .CLK(clk), .RST(rst), .I(g_init[209]), 
        .Q(mreg[209]) );
  DFF \mreg_reg[208]  ( .D(mreg[208]), .CLK(clk), .RST(rst), .I(g_init[208]), 
        .Q(mreg[208]) );
  DFF \mreg_reg[207]  ( .D(mreg[207]), .CLK(clk), .RST(rst), .I(g_init[207]), 
        .Q(mreg[207]) );
  DFF \mreg_reg[206]  ( .D(mreg[206]), .CLK(clk), .RST(rst), .I(g_init[206]), 
        .Q(mreg[206]) );
  DFF \mreg_reg[205]  ( .D(mreg[205]), .CLK(clk), .RST(rst), .I(g_init[205]), 
        .Q(mreg[205]) );
  DFF \mreg_reg[204]  ( .D(mreg[204]), .CLK(clk), .RST(rst), .I(g_init[204]), 
        .Q(mreg[204]) );
  DFF \mreg_reg[203]  ( .D(mreg[203]), .CLK(clk), .RST(rst), .I(g_init[203]), 
        .Q(mreg[203]) );
  DFF \mreg_reg[202]  ( .D(mreg[202]), .CLK(clk), .RST(rst), .I(g_init[202]), 
        .Q(mreg[202]) );
  DFF \mreg_reg[201]  ( .D(mreg[201]), .CLK(clk), .RST(rst), .I(g_init[201]), 
        .Q(mreg[201]) );
  DFF \mreg_reg[200]  ( .D(mreg[200]), .CLK(clk), .RST(rst), .I(g_init[200]), 
        .Q(mreg[200]) );
  DFF \mreg_reg[199]  ( .D(mreg[199]), .CLK(clk), .RST(rst), .I(g_init[199]), 
        .Q(mreg[199]) );
  DFF \mreg_reg[198]  ( .D(mreg[198]), .CLK(clk), .RST(rst), .I(g_init[198]), 
        .Q(mreg[198]) );
  DFF \mreg_reg[197]  ( .D(mreg[197]), .CLK(clk), .RST(rst), .I(g_init[197]), 
        .Q(mreg[197]) );
  DFF \mreg_reg[196]  ( .D(mreg[196]), .CLK(clk), .RST(rst), .I(g_init[196]), 
        .Q(mreg[196]) );
  DFF \mreg_reg[195]  ( .D(mreg[195]), .CLK(clk), .RST(rst), .I(g_init[195]), 
        .Q(mreg[195]) );
  DFF \mreg_reg[194]  ( .D(mreg[194]), .CLK(clk), .RST(rst), .I(g_init[194]), 
        .Q(mreg[194]) );
  DFF \mreg_reg[193]  ( .D(mreg[193]), .CLK(clk), .RST(rst), .I(g_init[193]), 
        .Q(mreg[193]) );
  DFF \mreg_reg[192]  ( .D(mreg[192]), .CLK(clk), .RST(rst), .I(g_init[192]), 
        .Q(mreg[192]) );
  DFF \mreg_reg[191]  ( .D(mreg[191]), .CLK(clk), .RST(rst), .I(g_init[191]), 
        .Q(mreg[191]) );
  DFF \mreg_reg[190]  ( .D(mreg[190]), .CLK(clk), .RST(rst), .I(g_init[190]), 
        .Q(mreg[190]) );
  DFF \mreg_reg[189]  ( .D(mreg[189]), .CLK(clk), .RST(rst), .I(g_init[189]), 
        .Q(mreg[189]) );
  DFF \mreg_reg[188]  ( .D(mreg[188]), .CLK(clk), .RST(rst), .I(g_init[188]), 
        .Q(mreg[188]) );
  DFF \mreg_reg[187]  ( .D(mreg[187]), .CLK(clk), .RST(rst), .I(g_init[187]), 
        .Q(mreg[187]) );
  DFF \mreg_reg[186]  ( .D(mreg[186]), .CLK(clk), .RST(rst), .I(g_init[186]), 
        .Q(mreg[186]) );
  DFF \mreg_reg[185]  ( .D(mreg[185]), .CLK(clk), .RST(rst), .I(g_init[185]), 
        .Q(mreg[185]) );
  DFF \mreg_reg[184]  ( .D(mreg[184]), .CLK(clk), .RST(rst), .I(g_init[184]), 
        .Q(mreg[184]) );
  DFF \mreg_reg[183]  ( .D(mreg[183]), .CLK(clk), .RST(rst), .I(g_init[183]), 
        .Q(mreg[183]) );
  DFF \mreg_reg[182]  ( .D(mreg[182]), .CLK(clk), .RST(rst), .I(g_init[182]), 
        .Q(mreg[182]) );
  DFF \mreg_reg[181]  ( .D(mreg[181]), .CLK(clk), .RST(rst), .I(g_init[181]), 
        .Q(mreg[181]) );
  DFF \mreg_reg[180]  ( .D(mreg[180]), .CLK(clk), .RST(rst), .I(g_init[180]), 
        .Q(mreg[180]) );
  DFF \mreg_reg[179]  ( .D(mreg[179]), .CLK(clk), .RST(rst), .I(g_init[179]), 
        .Q(mreg[179]) );
  DFF \mreg_reg[178]  ( .D(mreg[178]), .CLK(clk), .RST(rst), .I(g_init[178]), 
        .Q(mreg[178]) );
  DFF \mreg_reg[177]  ( .D(mreg[177]), .CLK(clk), .RST(rst), .I(g_init[177]), 
        .Q(mreg[177]) );
  DFF \mreg_reg[176]  ( .D(mreg[176]), .CLK(clk), .RST(rst), .I(g_init[176]), 
        .Q(mreg[176]) );
  DFF \mreg_reg[175]  ( .D(mreg[175]), .CLK(clk), .RST(rst), .I(g_init[175]), 
        .Q(mreg[175]) );
  DFF \mreg_reg[174]  ( .D(mreg[174]), .CLK(clk), .RST(rst), .I(g_init[174]), 
        .Q(mreg[174]) );
  DFF \mreg_reg[173]  ( .D(mreg[173]), .CLK(clk), .RST(rst), .I(g_init[173]), 
        .Q(mreg[173]) );
  DFF \mreg_reg[172]  ( .D(mreg[172]), .CLK(clk), .RST(rst), .I(g_init[172]), 
        .Q(mreg[172]) );
  DFF \mreg_reg[171]  ( .D(mreg[171]), .CLK(clk), .RST(rst), .I(g_init[171]), 
        .Q(mreg[171]) );
  DFF \mreg_reg[170]  ( .D(mreg[170]), .CLK(clk), .RST(rst), .I(g_init[170]), 
        .Q(mreg[170]) );
  DFF \mreg_reg[169]  ( .D(mreg[169]), .CLK(clk), .RST(rst), .I(g_init[169]), 
        .Q(mreg[169]) );
  DFF \mreg_reg[168]  ( .D(mreg[168]), .CLK(clk), .RST(rst), .I(g_init[168]), 
        .Q(mreg[168]) );
  DFF \mreg_reg[167]  ( .D(mreg[167]), .CLK(clk), .RST(rst), .I(g_init[167]), 
        .Q(mreg[167]) );
  DFF \mreg_reg[166]  ( .D(mreg[166]), .CLK(clk), .RST(rst), .I(g_init[166]), 
        .Q(mreg[166]) );
  DFF \mreg_reg[165]  ( .D(mreg[165]), .CLK(clk), .RST(rst), .I(g_init[165]), 
        .Q(mreg[165]) );
  DFF \mreg_reg[164]  ( .D(mreg[164]), .CLK(clk), .RST(rst), .I(g_init[164]), 
        .Q(mreg[164]) );
  DFF \mreg_reg[163]  ( .D(mreg[163]), .CLK(clk), .RST(rst), .I(g_init[163]), 
        .Q(mreg[163]) );
  DFF \mreg_reg[162]  ( .D(mreg[162]), .CLK(clk), .RST(rst), .I(g_init[162]), 
        .Q(mreg[162]) );
  DFF \mreg_reg[161]  ( .D(mreg[161]), .CLK(clk), .RST(rst), .I(g_init[161]), 
        .Q(mreg[161]) );
  DFF \mreg_reg[160]  ( .D(mreg[160]), .CLK(clk), .RST(rst), .I(g_init[160]), 
        .Q(mreg[160]) );
  DFF \mreg_reg[159]  ( .D(mreg[159]), .CLK(clk), .RST(rst), .I(g_init[159]), 
        .Q(mreg[159]) );
  DFF \mreg_reg[158]  ( .D(mreg[158]), .CLK(clk), .RST(rst), .I(g_init[158]), 
        .Q(mreg[158]) );
  DFF \mreg_reg[157]  ( .D(mreg[157]), .CLK(clk), .RST(rst), .I(g_init[157]), 
        .Q(mreg[157]) );
  DFF \mreg_reg[156]  ( .D(mreg[156]), .CLK(clk), .RST(rst), .I(g_init[156]), 
        .Q(mreg[156]) );
  DFF \mreg_reg[155]  ( .D(mreg[155]), .CLK(clk), .RST(rst), .I(g_init[155]), 
        .Q(mreg[155]) );
  DFF \mreg_reg[154]  ( .D(mreg[154]), .CLK(clk), .RST(rst), .I(g_init[154]), 
        .Q(mreg[154]) );
  DFF \mreg_reg[153]  ( .D(mreg[153]), .CLK(clk), .RST(rst), .I(g_init[153]), 
        .Q(mreg[153]) );
  DFF \mreg_reg[152]  ( .D(mreg[152]), .CLK(clk), .RST(rst), .I(g_init[152]), 
        .Q(mreg[152]) );
  DFF \mreg_reg[151]  ( .D(mreg[151]), .CLK(clk), .RST(rst), .I(g_init[151]), 
        .Q(mreg[151]) );
  DFF \mreg_reg[150]  ( .D(mreg[150]), .CLK(clk), .RST(rst), .I(g_init[150]), 
        .Q(mreg[150]) );
  DFF \mreg_reg[149]  ( .D(mreg[149]), .CLK(clk), .RST(rst), .I(g_init[149]), 
        .Q(mreg[149]) );
  DFF \mreg_reg[148]  ( .D(mreg[148]), .CLK(clk), .RST(rst), .I(g_init[148]), 
        .Q(mreg[148]) );
  DFF \mreg_reg[147]  ( .D(mreg[147]), .CLK(clk), .RST(rst), .I(g_init[147]), 
        .Q(mreg[147]) );
  DFF \mreg_reg[146]  ( .D(mreg[146]), .CLK(clk), .RST(rst), .I(g_init[146]), 
        .Q(mreg[146]) );
  DFF \mreg_reg[145]  ( .D(mreg[145]), .CLK(clk), .RST(rst), .I(g_init[145]), 
        .Q(mreg[145]) );
  DFF \mreg_reg[144]  ( .D(mreg[144]), .CLK(clk), .RST(rst), .I(g_init[144]), 
        .Q(mreg[144]) );
  DFF \mreg_reg[143]  ( .D(mreg[143]), .CLK(clk), .RST(rst), .I(g_init[143]), 
        .Q(mreg[143]) );
  DFF \mreg_reg[142]  ( .D(mreg[142]), .CLK(clk), .RST(rst), .I(g_init[142]), 
        .Q(mreg[142]) );
  DFF \mreg_reg[141]  ( .D(mreg[141]), .CLK(clk), .RST(rst), .I(g_init[141]), 
        .Q(mreg[141]) );
  DFF \mreg_reg[140]  ( .D(mreg[140]), .CLK(clk), .RST(rst), .I(g_init[140]), 
        .Q(mreg[140]) );
  DFF \mreg_reg[139]  ( .D(mreg[139]), .CLK(clk), .RST(rst), .I(g_init[139]), 
        .Q(mreg[139]) );
  DFF \mreg_reg[138]  ( .D(mreg[138]), .CLK(clk), .RST(rst), .I(g_init[138]), 
        .Q(mreg[138]) );
  DFF \mreg_reg[137]  ( .D(mreg[137]), .CLK(clk), .RST(rst), .I(g_init[137]), 
        .Q(mreg[137]) );
  DFF \mreg_reg[136]  ( .D(mreg[136]), .CLK(clk), .RST(rst), .I(g_init[136]), 
        .Q(mreg[136]) );
  DFF \mreg_reg[135]  ( .D(mreg[135]), .CLK(clk), .RST(rst), .I(g_init[135]), 
        .Q(mreg[135]) );
  DFF \mreg_reg[134]  ( .D(mreg[134]), .CLK(clk), .RST(rst), .I(g_init[134]), 
        .Q(mreg[134]) );
  DFF \mreg_reg[133]  ( .D(mreg[133]), .CLK(clk), .RST(rst), .I(g_init[133]), 
        .Q(mreg[133]) );
  DFF \mreg_reg[132]  ( .D(mreg[132]), .CLK(clk), .RST(rst), .I(g_init[132]), 
        .Q(mreg[132]) );
  DFF \mreg_reg[131]  ( .D(mreg[131]), .CLK(clk), .RST(rst), .I(g_init[131]), 
        .Q(mreg[131]) );
  DFF \mreg_reg[130]  ( .D(mreg[130]), .CLK(clk), .RST(rst), .I(g_init[130]), 
        .Q(mreg[130]) );
  DFF \mreg_reg[129]  ( .D(mreg[129]), .CLK(clk), .RST(rst), .I(g_init[129]), 
        .Q(mreg[129]) );
  DFF \mreg_reg[128]  ( .D(mreg[128]), .CLK(clk), .RST(rst), .I(g_init[128]), 
        .Q(mreg[128]) );
  DFF \mreg_reg[127]  ( .D(mreg[127]), .CLK(clk), .RST(rst), .I(g_init[127]), 
        .Q(mreg[127]) );
  DFF \mreg_reg[126]  ( .D(mreg[126]), .CLK(clk), .RST(rst), .I(g_init[126]), 
        .Q(mreg[126]) );
  DFF \mreg_reg[125]  ( .D(mreg[125]), .CLK(clk), .RST(rst), .I(g_init[125]), 
        .Q(mreg[125]) );
  DFF \mreg_reg[124]  ( .D(mreg[124]), .CLK(clk), .RST(rst), .I(g_init[124]), 
        .Q(mreg[124]) );
  DFF \mreg_reg[123]  ( .D(mreg[123]), .CLK(clk), .RST(rst), .I(g_init[123]), 
        .Q(mreg[123]) );
  DFF \mreg_reg[122]  ( .D(mreg[122]), .CLK(clk), .RST(rst), .I(g_init[122]), 
        .Q(mreg[122]) );
  DFF \mreg_reg[121]  ( .D(mreg[121]), .CLK(clk), .RST(rst), .I(g_init[121]), 
        .Q(mreg[121]) );
  DFF \mreg_reg[120]  ( .D(mreg[120]), .CLK(clk), .RST(rst), .I(g_init[120]), 
        .Q(mreg[120]) );
  DFF \mreg_reg[119]  ( .D(mreg[119]), .CLK(clk), .RST(rst), .I(g_init[119]), 
        .Q(mreg[119]) );
  DFF \mreg_reg[118]  ( .D(mreg[118]), .CLK(clk), .RST(rst), .I(g_init[118]), 
        .Q(mreg[118]) );
  DFF \mreg_reg[117]  ( .D(mreg[117]), .CLK(clk), .RST(rst), .I(g_init[117]), 
        .Q(mreg[117]) );
  DFF \mreg_reg[116]  ( .D(mreg[116]), .CLK(clk), .RST(rst), .I(g_init[116]), 
        .Q(mreg[116]) );
  DFF \mreg_reg[115]  ( .D(mreg[115]), .CLK(clk), .RST(rst), .I(g_init[115]), 
        .Q(mreg[115]) );
  DFF \mreg_reg[114]  ( .D(mreg[114]), .CLK(clk), .RST(rst), .I(g_init[114]), 
        .Q(mreg[114]) );
  DFF \mreg_reg[113]  ( .D(mreg[113]), .CLK(clk), .RST(rst), .I(g_init[113]), 
        .Q(mreg[113]) );
  DFF \mreg_reg[112]  ( .D(mreg[112]), .CLK(clk), .RST(rst), .I(g_init[112]), 
        .Q(mreg[112]) );
  DFF \mreg_reg[111]  ( .D(mreg[111]), .CLK(clk), .RST(rst), .I(g_init[111]), 
        .Q(mreg[111]) );
  DFF \mreg_reg[110]  ( .D(mreg[110]), .CLK(clk), .RST(rst), .I(g_init[110]), 
        .Q(mreg[110]) );
  DFF \mreg_reg[109]  ( .D(mreg[109]), .CLK(clk), .RST(rst), .I(g_init[109]), 
        .Q(mreg[109]) );
  DFF \mreg_reg[108]  ( .D(mreg[108]), .CLK(clk), .RST(rst), .I(g_init[108]), 
        .Q(mreg[108]) );
  DFF \mreg_reg[107]  ( .D(mreg[107]), .CLK(clk), .RST(rst), .I(g_init[107]), 
        .Q(mreg[107]) );
  DFF \mreg_reg[106]  ( .D(mreg[106]), .CLK(clk), .RST(rst), .I(g_init[106]), 
        .Q(mreg[106]) );
  DFF \mreg_reg[105]  ( .D(mreg[105]), .CLK(clk), .RST(rst), .I(g_init[105]), 
        .Q(mreg[105]) );
  DFF \mreg_reg[104]  ( .D(mreg[104]), .CLK(clk), .RST(rst), .I(g_init[104]), 
        .Q(mreg[104]) );
  DFF \mreg_reg[103]  ( .D(mreg[103]), .CLK(clk), .RST(rst), .I(g_init[103]), 
        .Q(mreg[103]) );
  DFF \mreg_reg[102]  ( .D(mreg[102]), .CLK(clk), .RST(rst), .I(g_init[102]), 
        .Q(mreg[102]) );
  DFF \mreg_reg[101]  ( .D(mreg[101]), .CLK(clk), .RST(rst), .I(g_init[101]), 
        .Q(mreg[101]) );
  DFF \mreg_reg[100]  ( .D(mreg[100]), .CLK(clk), .RST(rst), .I(g_init[100]), 
        .Q(mreg[100]) );
  DFF \mreg_reg[99]  ( .D(mreg[99]), .CLK(clk), .RST(rst), .I(g_init[99]), .Q(
        mreg[99]) );
  DFF \mreg_reg[98]  ( .D(mreg[98]), .CLK(clk), .RST(rst), .I(g_init[98]), .Q(
        mreg[98]) );
  DFF \mreg_reg[97]  ( .D(mreg[97]), .CLK(clk), .RST(rst), .I(g_init[97]), .Q(
        mreg[97]) );
  DFF \mreg_reg[96]  ( .D(mreg[96]), .CLK(clk), .RST(rst), .I(g_init[96]), .Q(
        mreg[96]) );
  DFF \mreg_reg[95]  ( .D(mreg[95]), .CLK(clk), .RST(rst), .I(g_init[95]), .Q(
        mreg[95]) );
  DFF \mreg_reg[94]  ( .D(mreg[94]), .CLK(clk), .RST(rst), .I(g_init[94]), .Q(
        mreg[94]) );
  DFF \mreg_reg[93]  ( .D(mreg[93]), .CLK(clk), .RST(rst), .I(g_init[93]), .Q(
        mreg[93]) );
  DFF \mreg_reg[92]  ( .D(mreg[92]), .CLK(clk), .RST(rst), .I(g_init[92]), .Q(
        mreg[92]) );
  DFF \mreg_reg[91]  ( .D(mreg[91]), .CLK(clk), .RST(rst), .I(g_init[91]), .Q(
        mreg[91]) );
  DFF \mreg_reg[90]  ( .D(mreg[90]), .CLK(clk), .RST(rst), .I(g_init[90]), .Q(
        mreg[90]) );
  DFF \mreg_reg[89]  ( .D(mreg[89]), .CLK(clk), .RST(rst), .I(g_init[89]), .Q(
        mreg[89]) );
  DFF \mreg_reg[88]  ( .D(mreg[88]), .CLK(clk), .RST(rst), .I(g_init[88]), .Q(
        mreg[88]) );
  DFF \mreg_reg[87]  ( .D(mreg[87]), .CLK(clk), .RST(rst), .I(g_init[87]), .Q(
        mreg[87]) );
  DFF \mreg_reg[86]  ( .D(mreg[86]), .CLK(clk), .RST(rst), .I(g_init[86]), .Q(
        mreg[86]) );
  DFF \mreg_reg[85]  ( .D(mreg[85]), .CLK(clk), .RST(rst), .I(g_init[85]), .Q(
        mreg[85]) );
  DFF \mreg_reg[84]  ( .D(mreg[84]), .CLK(clk), .RST(rst), .I(g_init[84]), .Q(
        mreg[84]) );
  DFF \mreg_reg[83]  ( .D(mreg[83]), .CLK(clk), .RST(rst), .I(g_init[83]), .Q(
        mreg[83]) );
  DFF \mreg_reg[82]  ( .D(mreg[82]), .CLK(clk), .RST(rst), .I(g_init[82]), .Q(
        mreg[82]) );
  DFF \mreg_reg[81]  ( .D(mreg[81]), .CLK(clk), .RST(rst), .I(g_init[81]), .Q(
        mreg[81]) );
  DFF \mreg_reg[80]  ( .D(mreg[80]), .CLK(clk), .RST(rst), .I(g_init[80]), .Q(
        mreg[80]) );
  DFF \mreg_reg[79]  ( .D(mreg[79]), .CLK(clk), .RST(rst), .I(g_init[79]), .Q(
        mreg[79]) );
  DFF \mreg_reg[78]  ( .D(mreg[78]), .CLK(clk), .RST(rst), .I(g_init[78]), .Q(
        mreg[78]) );
  DFF \mreg_reg[77]  ( .D(mreg[77]), .CLK(clk), .RST(rst), .I(g_init[77]), .Q(
        mreg[77]) );
  DFF \mreg_reg[76]  ( .D(mreg[76]), .CLK(clk), .RST(rst), .I(g_init[76]), .Q(
        mreg[76]) );
  DFF \mreg_reg[75]  ( .D(mreg[75]), .CLK(clk), .RST(rst), .I(g_init[75]), .Q(
        mreg[75]) );
  DFF \mreg_reg[74]  ( .D(mreg[74]), .CLK(clk), .RST(rst), .I(g_init[74]), .Q(
        mreg[74]) );
  DFF \mreg_reg[73]  ( .D(mreg[73]), .CLK(clk), .RST(rst), .I(g_init[73]), .Q(
        mreg[73]) );
  DFF \mreg_reg[72]  ( .D(mreg[72]), .CLK(clk), .RST(rst), .I(g_init[72]), .Q(
        mreg[72]) );
  DFF \mreg_reg[71]  ( .D(mreg[71]), .CLK(clk), .RST(rst), .I(g_init[71]), .Q(
        mreg[71]) );
  DFF \mreg_reg[70]  ( .D(mreg[70]), .CLK(clk), .RST(rst), .I(g_init[70]), .Q(
        mreg[70]) );
  DFF \mreg_reg[69]  ( .D(mreg[69]), .CLK(clk), .RST(rst), .I(g_init[69]), .Q(
        mreg[69]) );
  DFF \mreg_reg[68]  ( .D(mreg[68]), .CLK(clk), .RST(rst), .I(g_init[68]), .Q(
        mreg[68]) );
  DFF \mreg_reg[67]  ( .D(mreg[67]), .CLK(clk), .RST(rst), .I(g_init[67]), .Q(
        mreg[67]) );
  DFF \mreg_reg[66]  ( .D(mreg[66]), .CLK(clk), .RST(rst), .I(g_init[66]), .Q(
        mreg[66]) );
  DFF \mreg_reg[65]  ( .D(mreg[65]), .CLK(clk), .RST(rst), .I(g_init[65]), .Q(
        mreg[65]) );
  DFF \mreg_reg[64]  ( .D(mreg[64]), .CLK(clk), .RST(rst), .I(g_init[64]), .Q(
        mreg[64]) );
  DFF \mreg_reg[63]  ( .D(mreg[63]), .CLK(clk), .RST(rst), .I(g_init[63]), .Q(
        mreg[63]) );
  DFF \mreg_reg[62]  ( .D(mreg[62]), .CLK(clk), .RST(rst), .I(g_init[62]), .Q(
        mreg[62]) );
  DFF \mreg_reg[61]  ( .D(mreg[61]), .CLK(clk), .RST(rst), .I(g_init[61]), .Q(
        mreg[61]) );
  DFF \mreg_reg[60]  ( .D(mreg[60]), .CLK(clk), .RST(rst), .I(g_init[60]), .Q(
        mreg[60]) );
  DFF \mreg_reg[59]  ( .D(mreg[59]), .CLK(clk), .RST(rst), .I(g_init[59]), .Q(
        mreg[59]) );
  DFF \mreg_reg[58]  ( .D(mreg[58]), .CLK(clk), .RST(rst), .I(g_init[58]), .Q(
        mreg[58]) );
  DFF \mreg_reg[57]  ( .D(mreg[57]), .CLK(clk), .RST(rst), .I(g_init[57]), .Q(
        mreg[57]) );
  DFF \mreg_reg[56]  ( .D(mreg[56]), .CLK(clk), .RST(rst), .I(g_init[56]), .Q(
        mreg[56]) );
  DFF \mreg_reg[55]  ( .D(mreg[55]), .CLK(clk), .RST(rst), .I(g_init[55]), .Q(
        mreg[55]) );
  DFF \mreg_reg[54]  ( .D(mreg[54]), .CLK(clk), .RST(rst), .I(g_init[54]), .Q(
        mreg[54]) );
  DFF \mreg_reg[53]  ( .D(mreg[53]), .CLK(clk), .RST(rst), .I(g_init[53]), .Q(
        mreg[53]) );
  DFF \mreg_reg[52]  ( .D(mreg[52]), .CLK(clk), .RST(rst), .I(g_init[52]), .Q(
        mreg[52]) );
  DFF \mreg_reg[51]  ( .D(mreg[51]), .CLK(clk), .RST(rst), .I(g_init[51]), .Q(
        mreg[51]) );
  DFF \mreg_reg[50]  ( .D(mreg[50]), .CLK(clk), .RST(rst), .I(g_init[50]), .Q(
        mreg[50]) );
  DFF \mreg_reg[49]  ( .D(mreg[49]), .CLK(clk), .RST(rst), .I(g_init[49]), .Q(
        mreg[49]) );
  DFF \mreg_reg[48]  ( .D(mreg[48]), .CLK(clk), .RST(rst), .I(g_init[48]), .Q(
        mreg[48]) );
  DFF \mreg_reg[47]  ( .D(mreg[47]), .CLK(clk), .RST(rst), .I(g_init[47]), .Q(
        mreg[47]) );
  DFF \mreg_reg[46]  ( .D(mreg[46]), .CLK(clk), .RST(rst), .I(g_init[46]), .Q(
        mreg[46]) );
  DFF \mreg_reg[45]  ( .D(mreg[45]), .CLK(clk), .RST(rst), .I(g_init[45]), .Q(
        mreg[45]) );
  DFF \mreg_reg[44]  ( .D(mreg[44]), .CLK(clk), .RST(rst), .I(g_init[44]), .Q(
        mreg[44]) );
  DFF \mreg_reg[43]  ( .D(mreg[43]), .CLK(clk), .RST(rst), .I(g_init[43]), .Q(
        mreg[43]) );
  DFF \mreg_reg[42]  ( .D(mreg[42]), .CLK(clk), .RST(rst), .I(g_init[42]), .Q(
        mreg[42]) );
  DFF \mreg_reg[41]  ( .D(mreg[41]), .CLK(clk), .RST(rst), .I(g_init[41]), .Q(
        mreg[41]) );
  DFF \mreg_reg[40]  ( .D(mreg[40]), .CLK(clk), .RST(rst), .I(g_init[40]), .Q(
        mreg[40]) );
  DFF \mreg_reg[39]  ( .D(mreg[39]), .CLK(clk), .RST(rst), .I(g_init[39]), .Q(
        mreg[39]) );
  DFF \mreg_reg[38]  ( .D(mreg[38]), .CLK(clk), .RST(rst), .I(g_init[38]), .Q(
        mreg[38]) );
  DFF \mreg_reg[37]  ( .D(mreg[37]), .CLK(clk), .RST(rst), .I(g_init[37]), .Q(
        mreg[37]) );
  DFF \mreg_reg[36]  ( .D(mreg[36]), .CLK(clk), .RST(rst), .I(g_init[36]), .Q(
        mreg[36]) );
  DFF \mreg_reg[35]  ( .D(mreg[35]), .CLK(clk), .RST(rst), .I(g_init[35]), .Q(
        mreg[35]) );
  DFF \mreg_reg[34]  ( .D(mreg[34]), .CLK(clk), .RST(rst), .I(g_init[34]), .Q(
        mreg[34]) );
  DFF \mreg_reg[33]  ( .D(mreg[33]), .CLK(clk), .RST(rst), .I(g_init[33]), .Q(
        mreg[33]) );
  DFF \mreg_reg[32]  ( .D(mreg[32]), .CLK(clk), .RST(rst), .I(g_init[32]), .Q(
        mreg[32]) );
  DFF \mreg_reg[31]  ( .D(mreg[31]), .CLK(clk), .RST(rst), .I(g_init[31]), .Q(
        mreg[31]) );
  DFF \mreg_reg[30]  ( .D(mreg[30]), .CLK(clk), .RST(rst), .I(g_init[30]), .Q(
        mreg[30]) );
  DFF \mreg_reg[29]  ( .D(mreg[29]), .CLK(clk), .RST(rst), .I(g_init[29]), .Q(
        mreg[29]) );
  DFF \mreg_reg[28]  ( .D(mreg[28]), .CLK(clk), .RST(rst), .I(g_init[28]), .Q(
        mreg[28]) );
  DFF \mreg_reg[27]  ( .D(mreg[27]), .CLK(clk), .RST(rst), .I(g_init[27]), .Q(
        mreg[27]) );
  DFF \mreg_reg[26]  ( .D(mreg[26]), .CLK(clk), .RST(rst), .I(g_init[26]), .Q(
        mreg[26]) );
  DFF \mreg_reg[25]  ( .D(mreg[25]), .CLK(clk), .RST(rst), .I(g_init[25]), .Q(
        mreg[25]) );
  DFF \mreg_reg[24]  ( .D(mreg[24]), .CLK(clk), .RST(rst), .I(g_init[24]), .Q(
        mreg[24]) );
  DFF \mreg_reg[23]  ( .D(mreg[23]), .CLK(clk), .RST(rst), .I(g_init[23]), .Q(
        mreg[23]) );
  DFF \mreg_reg[22]  ( .D(mreg[22]), .CLK(clk), .RST(rst), .I(g_init[22]), .Q(
        mreg[22]) );
  DFF \mreg_reg[21]  ( .D(mreg[21]), .CLK(clk), .RST(rst), .I(g_init[21]), .Q(
        mreg[21]) );
  DFF \mreg_reg[20]  ( .D(mreg[20]), .CLK(clk), .RST(rst), .I(g_init[20]), .Q(
        mreg[20]) );
  DFF \mreg_reg[19]  ( .D(mreg[19]), .CLK(clk), .RST(rst), .I(g_init[19]), .Q(
        mreg[19]) );
  DFF \mreg_reg[18]  ( .D(mreg[18]), .CLK(clk), .RST(rst), .I(g_init[18]), .Q(
        mreg[18]) );
  DFF \mreg_reg[17]  ( .D(mreg[17]), .CLK(clk), .RST(rst), .I(g_init[17]), .Q(
        mreg[17]) );
  DFF \mreg_reg[16]  ( .D(mreg[16]), .CLK(clk), .RST(rst), .I(g_init[16]), .Q(
        mreg[16]) );
  DFF \mreg_reg[15]  ( .D(mreg[15]), .CLK(clk), .RST(rst), .I(g_init[15]), .Q(
        mreg[15]) );
  DFF \mreg_reg[14]  ( .D(mreg[14]), .CLK(clk), .RST(rst), .I(g_init[14]), .Q(
        mreg[14]) );
  DFF \mreg_reg[13]  ( .D(mreg[13]), .CLK(clk), .RST(rst), .I(g_init[13]), .Q(
        mreg[13]) );
  DFF \mreg_reg[12]  ( .D(mreg[12]), .CLK(clk), .RST(rst), .I(g_init[12]), .Q(
        mreg[12]) );
  DFF \mreg_reg[11]  ( .D(mreg[11]), .CLK(clk), .RST(rst), .I(g_init[11]), .Q(
        mreg[11]) );
  DFF \mreg_reg[10]  ( .D(mreg[10]), .CLK(clk), .RST(rst), .I(g_init[10]), .Q(
        mreg[10]) );
  DFF \mreg_reg[9]  ( .D(mreg[9]), .CLK(clk), .RST(rst), .I(g_init[9]), .Q(
        mreg[9]) );
  DFF \mreg_reg[8]  ( .D(mreg[8]), .CLK(clk), .RST(rst), .I(g_init[8]), .Q(
        mreg[8]) );
  DFF \mreg_reg[7]  ( .D(mreg[7]), .CLK(clk), .RST(rst), .I(g_init[7]), .Q(
        mreg[7]) );
  DFF \mreg_reg[6]  ( .D(mreg[6]), .CLK(clk), .RST(rst), .I(g_init[6]), .Q(
        mreg[6]) );
  DFF \mreg_reg[5]  ( .D(mreg[5]), .CLK(clk), .RST(rst), .I(g_init[5]), .Q(
        mreg[5]) );
  DFF \mreg_reg[4]  ( .D(mreg[4]), .CLK(clk), .RST(rst), .I(g_init[4]), .Q(
        mreg[4]) );
  DFF \mreg_reg[3]  ( .D(mreg[3]), .CLK(clk), .RST(rst), .I(g_init[3]), .Q(
        mreg[3]) );
  DFF \mreg_reg[2]  ( .D(mreg[2]), .CLK(clk), .RST(rst), .I(g_init[2]), .Q(
        mreg[2]) );
  DFF \mreg_reg[1]  ( .D(mreg[1]), .CLK(clk), .RST(rst), .I(g_init[1]), .Q(
        mreg[1]) );
  DFF \mreg_reg[0]  ( .D(mreg[0]), .CLK(clk), .RST(rst), .I(g_init[0]), .Q(
        mreg[0]) );
  DFF \creg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(g_init[0]), .Q(
        creg[0]) );
  DFF \creg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(g_init[1]), .Q(
        creg[1]) );
  DFF \creg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(g_init[2]), .Q(
        creg[2]) );
  DFF \creg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(g_init[3]), .Q(
        creg[3]) );
  DFF \creg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(g_init[4]), .Q(
        creg[4]) );
  DFF \creg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(g_init[5]), .Q(
        creg[5]) );
  DFF \creg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(g_init[6]), .Q(
        creg[6]) );
  DFF \creg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(g_init[7]), .Q(
        creg[7]) );
  DFF \creg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(g_init[8]), .Q(
        creg[8]) );
  DFF \creg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(g_init[9]), .Q(
        creg[9]) );
  DFF \creg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(g_init[10]), .Q(
        creg[10]) );
  DFF \creg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(g_init[11]), .Q(
        creg[11]) );
  DFF \creg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(g_init[12]), .Q(
        creg[12]) );
  DFF \creg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(g_init[13]), .Q(
        creg[13]) );
  DFF \creg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(g_init[14]), .Q(
        creg[14]) );
  DFF \creg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(g_init[15]), .Q(
        creg[15]) );
  DFF \creg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .I(g_init[16]), .Q(
        creg[16]) );
  DFF \creg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .I(g_init[17]), .Q(
        creg[17]) );
  DFF \creg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .I(g_init[18]), .Q(
        creg[18]) );
  DFF \creg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .I(g_init[19]), .Q(
        creg[19]) );
  DFF \creg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .I(g_init[20]), .Q(
        creg[20]) );
  DFF \creg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .I(g_init[21]), .Q(
        creg[21]) );
  DFF \creg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .I(g_init[22]), .Q(
        creg[22]) );
  DFF \creg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .I(g_init[23]), .Q(
        creg[23]) );
  DFF \creg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .I(g_init[24]), .Q(
        creg[24]) );
  DFF \creg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .I(g_init[25]), .Q(
        creg[25]) );
  DFF \creg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .I(g_init[26]), .Q(
        creg[26]) );
  DFF \creg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .I(g_init[27]), .Q(
        creg[27]) );
  DFF \creg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .I(g_init[28]), .Q(
        creg[28]) );
  DFF \creg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .I(g_init[29]), .Q(
        creg[29]) );
  DFF \creg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .I(g_init[30]), .Q(
        creg[30]) );
  DFF \creg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .I(g_init[31]), .Q(
        creg[31]) );
  DFF \creg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(rst), .I(g_init[32]), .Q(
        creg[32]) );
  DFF \creg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(rst), .I(g_init[33]), .Q(
        creg[33]) );
  DFF \creg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(rst), .I(g_init[34]), .Q(
        creg[34]) );
  DFF \creg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(rst), .I(g_init[35]), .Q(
        creg[35]) );
  DFF \creg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(rst), .I(g_init[36]), .Q(
        creg[36]) );
  DFF \creg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(rst), .I(g_init[37]), .Q(
        creg[37]) );
  DFF \creg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(rst), .I(g_init[38]), .Q(
        creg[38]) );
  DFF \creg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(rst), .I(g_init[39]), .Q(
        creg[39]) );
  DFF \creg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(rst), .I(g_init[40]), .Q(
        creg[40]) );
  DFF \creg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(rst), .I(g_init[41]), .Q(
        creg[41]) );
  DFF \creg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(rst), .I(g_init[42]), .Q(
        creg[42]) );
  DFF \creg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(rst), .I(g_init[43]), .Q(
        creg[43]) );
  DFF \creg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(rst), .I(g_init[44]), .Q(
        creg[44]) );
  DFF \creg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(rst), .I(g_init[45]), .Q(
        creg[45]) );
  DFF \creg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(rst), .I(g_init[46]), .Q(
        creg[46]) );
  DFF \creg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(rst), .I(g_init[47]), .Q(
        creg[47]) );
  DFF \creg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(rst), .I(g_init[48]), .Q(
        creg[48]) );
  DFF \creg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(rst), .I(g_init[49]), .Q(
        creg[49]) );
  DFF \creg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(rst), .I(g_init[50]), .Q(
        creg[50]) );
  DFF \creg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(rst), .I(g_init[51]), .Q(
        creg[51]) );
  DFF \creg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(rst), .I(g_init[52]), .Q(
        creg[52]) );
  DFF \creg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(rst), .I(g_init[53]), .Q(
        creg[53]) );
  DFF \creg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(rst), .I(g_init[54]), .Q(
        creg[54]) );
  DFF \creg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(rst), .I(g_init[55]), .Q(
        creg[55]) );
  DFF \creg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(rst), .I(g_init[56]), .Q(
        creg[56]) );
  DFF \creg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(rst), .I(g_init[57]), .Q(
        creg[57]) );
  DFF \creg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(rst), .I(g_init[58]), .Q(
        creg[58]) );
  DFF \creg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(rst), .I(g_init[59]), .Q(
        creg[59]) );
  DFF \creg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(rst), .I(g_init[60]), .Q(
        creg[60]) );
  DFF \creg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(rst), .I(g_init[61]), .Q(
        creg[61]) );
  DFF \creg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(rst), .I(g_init[62]), .Q(
        creg[62]) );
  DFF \creg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(rst), .I(g_init[63]), .Q(
        creg[63]) );
  DFF \creg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(rst), .I(g_init[64]), .Q(
        creg[64]) );
  DFF \creg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(rst), .I(g_init[65]), .Q(
        creg[65]) );
  DFF \creg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(rst), .I(g_init[66]), .Q(
        creg[66]) );
  DFF \creg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(rst), .I(g_init[67]), .Q(
        creg[67]) );
  DFF \creg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(rst), .I(g_init[68]), .Q(
        creg[68]) );
  DFF \creg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(rst), .I(g_init[69]), .Q(
        creg[69]) );
  DFF \creg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(rst), .I(g_init[70]), .Q(
        creg[70]) );
  DFF \creg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(rst), .I(g_init[71]), .Q(
        creg[71]) );
  DFF \creg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(rst), .I(g_init[72]), .Q(
        creg[72]) );
  DFF \creg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(rst), .I(g_init[73]), .Q(
        creg[73]) );
  DFF \creg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(rst), .I(g_init[74]), .Q(
        creg[74]) );
  DFF \creg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(rst), .I(g_init[75]), .Q(
        creg[75]) );
  DFF \creg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(rst), .I(g_init[76]), .Q(
        creg[76]) );
  DFF \creg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(rst), .I(g_init[77]), .Q(
        creg[77]) );
  DFF \creg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(rst), .I(g_init[78]), .Q(
        creg[78]) );
  DFF \creg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(rst), .I(g_init[79]), .Q(
        creg[79]) );
  DFF \creg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(rst), .I(g_init[80]), .Q(
        creg[80]) );
  DFF \creg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(rst), .I(g_init[81]), .Q(
        creg[81]) );
  DFF \creg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(rst), .I(g_init[82]), .Q(
        creg[82]) );
  DFF \creg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(rst), .I(g_init[83]), .Q(
        creg[83]) );
  DFF \creg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(rst), .I(g_init[84]), .Q(
        creg[84]) );
  DFF \creg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(rst), .I(g_init[85]), .Q(
        creg[85]) );
  DFF \creg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(rst), .I(g_init[86]), .Q(
        creg[86]) );
  DFF \creg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(rst), .I(g_init[87]), .Q(
        creg[87]) );
  DFF \creg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(rst), .I(g_init[88]), .Q(
        creg[88]) );
  DFF \creg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(rst), .I(g_init[89]), .Q(
        creg[89]) );
  DFF \creg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(rst), .I(g_init[90]), .Q(
        creg[90]) );
  DFF \creg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(rst), .I(g_init[91]), .Q(
        creg[91]) );
  DFF \creg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(rst), .I(g_init[92]), .Q(
        creg[92]) );
  DFF \creg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(rst), .I(g_init[93]), .Q(
        creg[93]) );
  DFF \creg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(rst), .I(g_init[94]), .Q(
        creg[94]) );
  DFF \creg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(rst), .I(g_init[95]), .Q(
        creg[95]) );
  DFF \creg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(rst), .I(g_init[96]), .Q(
        creg[96]) );
  DFF \creg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(rst), .I(g_init[97]), .Q(
        creg[97]) );
  DFF \creg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(rst), .I(g_init[98]), .Q(
        creg[98]) );
  DFF \creg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(rst), .I(g_init[99]), .Q(
        creg[99]) );
  DFF \creg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(rst), .I(g_init[100]), .Q(
        creg[100]) );
  DFF \creg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(rst), .I(g_init[101]), .Q(
        creg[101]) );
  DFF \creg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(rst), .I(g_init[102]), .Q(
        creg[102]) );
  DFF \creg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(rst), .I(g_init[103]), .Q(
        creg[103]) );
  DFF \creg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(rst), .I(g_init[104]), .Q(
        creg[104]) );
  DFF \creg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(rst), .I(g_init[105]), .Q(
        creg[105]) );
  DFF \creg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(rst), .I(g_init[106]), .Q(
        creg[106]) );
  DFF \creg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(rst), .I(g_init[107]), .Q(
        creg[107]) );
  DFF \creg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(rst), .I(g_init[108]), .Q(
        creg[108]) );
  DFF \creg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(rst), .I(g_init[109]), .Q(
        creg[109]) );
  DFF \creg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(rst), .I(g_init[110]), .Q(
        creg[110]) );
  DFF \creg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(rst), .I(g_init[111]), .Q(
        creg[111]) );
  DFF \creg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(rst), .I(g_init[112]), .Q(
        creg[112]) );
  DFF \creg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(rst), .I(g_init[113]), .Q(
        creg[113]) );
  DFF \creg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(rst), .I(g_init[114]), .Q(
        creg[114]) );
  DFF \creg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(rst), .I(g_init[115]), .Q(
        creg[115]) );
  DFF \creg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(rst), .I(g_init[116]), .Q(
        creg[116]) );
  DFF \creg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(rst), .I(g_init[117]), .Q(
        creg[117]) );
  DFF \creg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(rst), .I(g_init[118]), .Q(
        creg[118]) );
  DFF \creg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(rst), .I(g_init[119]), .Q(
        creg[119]) );
  DFF \creg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(rst), .I(g_init[120]), .Q(
        creg[120]) );
  DFF \creg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(rst), .I(g_init[121]), .Q(
        creg[121]) );
  DFF \creg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(rst), .I(g_init[122]), .Q(
        creg[122]) );
  DFF \creg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(rst), .I(g_init[123]), .Q(
        creg[123]) );
  DFF \creg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(rst), .I(g_init[124]), .Q(
        creg[124]) );
  DFF \creg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(rst), .I(g_init[125]), .Q(
        creg[125]) );
  DFF \creg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(rst), .I(g_init[126]), .Q(
        creg[126]) );
  DFF \creg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(rst), .I(g_init[127]), .Q(
        creg[127]) );
  DFF \creg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(rst), .I(g_init[128]), .Q(
        creg[128]) );
  DFF \creg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(rst), .I(g_init[129]), .Q(
        creg[129]) );
  DFF \creg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(rst), .I(g_init[130]), .Q(
        creg[130]) );
  DFF \creg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(rst), .I(g_init[131]), .Q(
        creg[131]) );
  DFF \creg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(rst), .I(g_init[132]), .Q(
        creg[132]) );
  DFF \creg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(rst), .I(g_init[133]), .Q(
        creg[133]) );
  DFF \creg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(rst), .I(g_init[134]), .Q(
        creg[134]) );
  DFF \creg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(rst), .I(g_init[135]), .Q(
        creg[135]) );
  DFF \creg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(rst), .I(g_init[136]), .Q(
        creg[136]) );
  DFF \creg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(rst), .I(g_init[137]), .Q(
        creg[137]) );
  DFF \creg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(rst), .I(g_init[138]), .Q(
        creg[138]) );
  DFF \creg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(rst), .I(g_init[139]), .Q(
        creg[139]) );
  DFF \creg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(rst), .I(g_init[140]), .Q(
        creg[140]) );
  DFF \creg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(rst), .I(g_init[141]), .Q(
        creg[141]) );
  DFF \creg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(rst), .I(g_init[142]), .Q(
        creg[142]) );
  DFF \creg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(rst), .I(g_init[143]), .Q(
        creg[143]) );
  DFF \creg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(rst), .I(g_init[144]), .Q(
        creg[144]) );
  DFF \creg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(rst), .I(g_init[145]), .Q(
        creg[145]) );
  DFF \creg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(rst), .I(g_init[146]), .Q(
        creg[146]) );
  DFF \creg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(rst), .I(g_init[147]), .Q(
        creg[147]) );
  DFF \creg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(rst), .I(g_init[148]), .Q(
        creg[148]) );
  DFF \creg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(rst), .I(g_init[149]), .Q(
        creg[149]) );
  DFF \creg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(rst), .I(g_init[150]), .Q(
        creg[150]) );
  DFF \creg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(rst), .I(g_init[151]), .Q(
        creg[151]) );
  DFF \creg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(rst), .I(g_init[152]), .Q(
        creg[152]) );
  DFF \creg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(rst), .I(g_init[153]), .Q(
        creg[153]) );
  DFF \creg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(rst), .I(g_init[154]), .Q(
        creg[154]) );
  DFF \creg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(rst), .I(g_init[155]), .Q(
        creg[155]) );
  DFF \creg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(rst), .I(g_init[156]), .Q(
        creg[156]) );
  DFF \creg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(rst), .I(g_init[157]), .Q(
        creg[157]) );
  DFF \creg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(rst), .I(g_init[158]), .Q(
        creg[158]) );
  DFF \creg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(rst), .I(g_init[159]), .Q(
        creg[159]) );
  DFF \creg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(rst), .I(g_init[160]), .Q(
        creg[160]) );
  DFF \creg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(rst), .I(g_init[161]), .Q(
        creg[161]) );
  DFF \creg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(rst), .I(g_init[162]), .Q(
        creg[162]) );
  DFF \creg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(rst), .I(g_init[163]), .Q(
        creg[163]) );
  DFF \creg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(rst), .I(g_init[164]), .Q(
        creg[164]) );
  DFF \creg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(rst), .I(g_init[165]), .Q(
        creg[165]) );
  DFF \creg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(rst), .I(g_init[166]), .Q(
        creg[166]) );
  DFF \creg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(rst), .I(g_init[167]), .Q(
        creg[167]) );
  DFF \creg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(rst), .I(g_init[168]), .Q(
        creg[168]) );
  DFF \creg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(rst), .I(g_init[169]), .Q(
        creg[169]) );
  DFF \creg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(rst), .I(g_init[170]), .Q(
        creg[170]) );
  DFF \creg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(rst), .I(g_init[171]), .Q(
        creg[171]) );
  DFF \creg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(rst), .I(g_init[172]), .Q(
        creg[172]) );
  DFF \creg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(rst), .I(g_init[173]), .Q(
        creg[173]) );
  DFF \creg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(rst), .I(g_init[174]), .Q(
        creg[174]) );
  DFF \creg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(rst), .I(g_init[175]), .Q(
        creg[175]) );
  DFF \creg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(rst), .I(g_init[176]), .Q(
        creg[176]) );
  DFF \creg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(rst), .I(g_init[177]), .Q(
        creg[177]) );
  DFF \creg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(rst), .I(g_init[178]), .Q(
        creg[178]) );
  DFF \creg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(rst), .I(g_init[179]), .Q(
        creg[179]) );
  DFF \creg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(rst), .I(g_init[180]), .Q(
        creg[180]) );
  DFF \creg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(rst), .I(g_init[181]), .Q(
        creg[181]) );
  DFF \creg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(rst), .I(g_init[182]), .Q(
        creg[182]) );
  DFF \creg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(rst), .I(g_init[183]), .Q(
        creg[183]) );
  DFF \creg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(rst), .I(g_init[184]), .Q(
        creg[184]) );
  DFF \creg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(rst), .I(g_init[185]), .Q(
        creg[185]) );
  DFF \creg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(rst), .I(g_init[186]), .Q(
        creg[186]) );
  DFF \creg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(rst), .I(g_init[187]), .Q(
        creg[187]) );
  DFF \creg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(rst), .I(g_init[188]), .Q(
        creg[188]) );
  DFF \creg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(rst), .I(g_init[189]), .Q(
        creg[189]) );
  DFF \creg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(rst), .I(g_init[190]), .Q(
        creg[190]) );
  DFF \creg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(rst), .I(g_init[191]), .Q(
        creg[191]) );
  DFF \creg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(rst), .I(g_init[192]), .Q(
        creg[192]) );
  DFF \creg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(rst), .I(g_init[193]), .Q(
        creg[193]) );
  DFF \creg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(rst), .I(g_init[194]), .Q(
        creg[194]) );
  DFF \creg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(rst), .I(g_init[195]), .Q(
        creg[195]) );
  DFF \creg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(rst), .I(g_init[196]), .Q(
        creg[196]) );
  DFF \creg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(rst), .I(g_init[197]), .Q(
        creg[197]) );
  DFF \creg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(rst), .I(g_init[198]), .Q(
        creg[198]) );
  DFF \creg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(rst), .I(g_init[199]), .Q(
        creg[199]) );
  DFF \creg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(rst), .I(g_init[200]), .Q(
        creg[200]) );
  DFF \creg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(rst), .I(g_init[201]), .Q(
        creg[201]) );
  DFF \creg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(rst), .I(g_init[202]), .Q(
        creg[202]) );
  DFF \creg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(rst), .I(g_init[203]), .Q(
        creg[203]) );
  DFF \creg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(rst), .I(g_init[204]), .Q(
        creg[204]) );
  DFF \creg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(rst), .I(g_init[205]), .Q(
        creg[205]) );
  DFF \creg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(rst), .I(g_init[206]), .Q(
        creg[206]) );
  DFF \creg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(rst), .I(g_init[207]), .Q(
        creg[207]) );
  DFF \creg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(rst), .I(g_init[208]), .Q(
        creg[208]) );
  DFF \creg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(rst), .I(g_init[209]), .Q(
        creg[209]) );
  DFF \creg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(rst), .I(g_init[210]), .Q(
        creg[210]) );
  DFF \creg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(rst), .I(g_init[211]), .Q(
        creg[211]) );
  DFF \creg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(rst), .I(g_init[212]), .Q(
        creg[212]) );
  DFF \creg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(rst), .I(g_init[213]), .Q(
        creg[213]) );
  DFF \creg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(rst), .I(g_init[214]), .Q(
        creg[214]) );
  DFF \creg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(rst), .I(g_init[215]), .Q(
        creg[215]) );
  DFF \creg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(rst), .I(g_init[216]), .Q(
        creg[216]) );
  DFF \creg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(rst), .I(g_init[217]), .Q(
        creg[217]) );
  DFF \creg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(rst), .I(g_init[218]), .Q(
        creg[218]) );
  DFF \creg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(rst), .I(g_init[219]), .Q(
        creg[219]) );
  DFF \creg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(rst), .I(g_init[220]), .Q(
        creg[220]) );
  DFF \creg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(rst), .I(g_init[221]), .Q(
        creg[221]) );
  DFF \creg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(rst), .I(g_init[222]), .Q(
        creg[222]) );
  DFF \creg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(rst), .I(g_init[223]), .Q(
        creg[223]) );
  DFF \creg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(rst), .I(g_init[224]), .Q(
        creg[224]) );
  DFF \creg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(rst), .I(g_init[225]), .Q(
        creg[225]) );
  DFF \creg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(rst), .I(g_init[226]), .Q(
        creg[226]) );
  DFF \creg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(rst), .I(g_init[227]), .Q(
        creg[227]) );
  DFF \creg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(rst), .I(g_init[228]), .Q(
        creg[228]) );
  DFF \creg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(rst), .I(g_init[229]), .Q(
        creg[229]) );
  DFF \creg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(rst), .I(g_init[230]), .Q(
        creg[230]) );
  DFF \creg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(rst), .I(g_init[231]), .Q(
        creg[231]) );
  DFF \creg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(rst), .I(g_init[232]), .Q(
        creg[232]) );
  DFF \creg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(rst), .I(g_init[233]), .Q(
        creg[233]) );
  DFF \creg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(rst), .I(g_init[234]), .Q(
        creg[234]) );
  DFF \creg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(rst), .I(g_init[235]), .Q(
        creg[235]) );
  DFF \creg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(rst), .I(g_init[236]), .Q(
        creg[236]) );
  DFF \creg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(rst), .I(g_init[237]), .Q(
        creg[237]) );
  DFF \creg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(rst), .I(g_init[238]), .Q(
        creg[238]) );
  DFF \creg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(rst), .I(g_init[239]), .Q(
        creg[239]) );
  DFF \creg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(rst), .I(g_init[240]), .Q(
        creg[240]) );
  DFF \creg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(rst), .I(g_init[241]), .Q(
        creg[241]) );
  DFF \creg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(rst), .I(g_init[242]), .Q(
        creg[242]) );
  DFF \creg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(rst), .I(g_init[243]), .Q(
        creg[243]) );
  DFF \creg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(rst), .I(g_init[244]), .Q(
        creg[244]) );
  DFF \creg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(rst), .I(g_init[245]), .Q(
        creg[245]) );
  DFF \creg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(rst), .I(g_init[246]), .Q(
        creg[246]) );
  DFF \creg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(rst), .I(g_init[247]), .Q(
        creg[247]) );
  DFF \creg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(rst), .I(g_init[248]), .Q(
        creg[248]) );
  DFF \creg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(rst), .I(g_init[249]), .Q(
        creg[249]) );
  DFF \creg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(rst), .I(g_init[250]), .Q(
        creg[250]) );
  DFF \creg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(rst), .I(g_init[251]), .Q(
        creg[251]) );
  DFF \creg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(rst), .I(g_init[252]), .Q(
        creg[252]) );
  DFF \creg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(rst), .I(g_init[253]), .Q(
        creg[253]) );
  DFF \creg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(rst), .I(g_init[254]), .Q(
        creg[254]) );
  DFF \creg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(rst), .I(g_init[255]), .Q(
        creg[255]) );
  DFF \creg_reg[256]  ( .D(o[256]), .CLK(clk), .RST(rst), .I(g_init[256]), .Q(
        creg[256]) );
  DFF \creg_reg[257]  ( .D(o[257]), .CLK(clk), .RST(rst), .I(g_init[257]), .Q(
        creg[257]) );
  DFF \creg_reg[258]  ( .D(o[258]), .CLK(clk), .RST(rst), .I(g_init[258]), .Q(
        creg[258]) );
  DFF \creg_reg[259]  ( .D(o[259]), .CLK(clk), .RST(rst), .I(g_init[259]), .Q(
        creg[259]) );
  DFF \creg_reg[260]  ( .D(o[260]), .CLK(clk), .RST(rst), .I(g_init[260]), .Q(
        creg[260]) );
  DFF \creg_reg[261]  ( .D(o[261]), .CLK(clk), .RST(rst), .I(g_init[261]), .Q(
        creg[261]) );
  DFF \creg_reg[262]  ( .D(o[262]), .CLK(clk), .RST(rst), .I(g_init[262]), .Q(
        creg[262]) );
  DFF \creg_reg[263]  ( .D(o[263]), .CLK(clk), .RST(rst), .I(g_init[263]), .Q(
        creg[263]) );
  DFF \creg_reg[264]  ( .D(o[264]), .CLK(clk), .RST(rst), .I(g_init[264]), .Q(
        creg[264]) );
  DFF \creg_reg[265]  ( .D(o[265]), .CLK(clk), .RST(rst), .I(g_init[265]), .Q(
        creg[265]) );
  DFF \creg_reg[266]  ( .D(o[266]), .CLK(clk), .RST(rst), .I(g_init[266]), .Q(
        creg[266]) );
  DFF \creg_reg[267]  ( .D(o[267]), .CLK(clk), .RST(rst), .I(g_init[267]), .Q(
        creg[267]) );
  DFF \creg_reg[268]  ( .D(o[268]), .CLK(clk), .RST(rst), .I(g_init[268]), .Q(
        creg[268]) );
  DFF \creg_reg[269]  ( .D(o[269]), .CLK(clk), .RST(rst), .I(g_init[269]), .Q(
        creg[269]) );
  DFF \creg_reg[270]  ( .D(o[270]), .CLK(clk), .RST(rst), .I(g_init[270]), .Q(
        creg[270]) );
  DFF \creg_reg[271]  ( .D(o[271]), .CLK(clk), .RST(rst), .I(g_init[271]), .Q(
        creg[271]) );
  DFF \creg_reg[272]  ( .D(o[272]), .CLK(clk), .RST(rst), .I(g_init[272]), .Q(
        creg[272]) );
  DFF \creg_reg[273]  ( .D(o[273]), .CLK(clk), .RST(rst), .I(g_init[273]), .Q(
        creg[273]) );
  DFF \creg_reg[274]  ( .D(o[274]), .CLK(clk), .RST(rst), .I(g_init[274]), .Q(
        creg[274]) );
  DFF \creg_reg[275]  ( .D(o[275]), .CLK(clk), .RST(rst), .I(g_init[275]), .Q(
        creg[275]) );
  DFF \creg_reg[276]  ( .D(o[276]), .CLK(clk), .RST(rst), .I(g_init[276]), .Q(
        creg[276]) );
  DFF \creg_reg[277]  ( .D(o[277]), .CLK(clk), .RST(rst), .I(g_init[277]), .Q(
        creg[277]) );
  DFF \creg_reg[278]  ( .D(o[278]), .CLK(clk), .RST(rst), .I(g_init[278]), .Q(
        creg[278]) );
  DFF \creg_reg[279]  ( .D(o[279]), .CLK(clk), .RST(rst), .I(g_init[279]), .Q(
        creg[279]) );
  DFF \creg_reg[280]  ( .D(o[280]), .CLK(clk), .RST(rst), .I(g_init[280]), .Q(
        creg[280]) );
  DFF \creg_reg[281]  ( .D(o[281]), .CLK(clk), .RST(rst), .I(g_init[281]), .Q(
        creg[281]) );
  DFF \creg_reg[282]  ( .D(o[282]), .CLK(clk), .RST(rst), .I(g_init[282]), .Q(
        creg[282]) );
  DFF \creg_reg[283]  ( .D(o[283]), .CLK(clk), .RST(rst), .I(g_init[283]), .Q(
        creg[283]) );
  DFF \creg_reg[284]  ( .D(o[284]), .CLK(clk), .RST(rst), .I(g_init[284]), .Q(
        creg[284]) );
  DFF \creg_reg[285]  ( .D(o[285]), .CLK(clk), .RST(rst), .I(g_init[285]), .Q(
        creg[285]) );
  DFF \creg_reg[286]  ( .D(o[286]), .CLK(clk), .RST(rst), .I(g_init[286]), .Q(
        creg[286]) );
  DFF \creg_reg[287]  ( .D(o[287]), .CLK(clk), .RST(rst), .I(g_init[287]), .Q(
        creg[287]) );
  DFF \creg_reg[288]  ( .D(o[288]), .CLK(clk), .RST(rst), .I(g_init[288]), .Q(
        creg[288]) );
  DFF \creg_reg[289]  ( .D(o[289]), .CLK(clk), .RST(rst), .I(g_init[289]), .Q(
        creg[289]) );
  DFF \creg_reg[290]  ( .D(o[290]), .CLK(clk), .RST(rst), .I(g_init[290]), .Q(
        creg[290]) );
  DFF \creg_reg[291]  ( .D(o[291]), .CLK(clk), .RST(rst), .I(g_init[291]), .Q(
        creg[291]) );
  DFF \creg_reg[292]  ( .D(o[292]), .CLK(clk), .RST(rst), .I(g_init[292]), .Q(
        creg[292]) );
  DFF \creg_reg[293]  ( .D(o[293]), .CLK(clk), .RST(rst), .I(g_init[293]), .Q(
        creg[293]) );
  DFF \creg_reg[294]  ( .D(o[294]), .CLK(clk), .RST(rst), .I(g_init[294]), .Q(
        creg[294]) );
  DFF \creg_reg[295]  ( .D(o[295]), .CLK(clk), .RST(rst), .I(g_init[295]), .Q(
        creg[295]) );
  DFF \creg_reg[296]  ( .D(o[296]), .CLK(clk), .RST(rst), .I(g_init[296]), .Q(
        creg[296]) );
  DFF \creg_reg[297]  ( .D(o[297]), .CLK(clk), .RST(rst), .I(g_init[297]), .Q(
        creg[297]) );
  DFF \creg_reg[298]  ( .D(o[298]), .CLK(clk), .RST(rst), .I(g_init[298]), .Q(
        creg[298]) );
  DFF \creg_reg[299]  ( .D(o[299]), .CLK(clk), .RST(rst), .I(g_init[299]), .Q(
        creg[299]) );
  DFF \creg_reg[300]  ( .D(o[300]), .CLK(clk), .RST(rst), .I(g_init[300]), .Q(
        creg[300]) );
  DFF \creg_reg[301]  ( .D(o[301]), .CLK(clk), .RST(rst), .I(g_init[301]), .Q(
        creg[301]) );
  DFF \creg_reg[302]  ( .D(o[302]), .CLK(clk), .RST(rst), .I(g_init[302]), .Q(
        creg[302]) );
  DFF \creg_reg[303]  ( .D(o[303]), .CLK(clk), .RST(rst), .I(g_init[303]), .Q(
        creg[303]) );
  DFF \creg_reg[304]  ( .D(o[304]), .CLK(clk), .RST(rst), .I(g_init[304]), .Q(
        creg[304]) );
  DFF \creg_reg[305]  ( .D(o[305]), .CLK(clk), .RST(rst), .I(g_init[305]), .Q(
        creg[305]) );
  DFF \creg_reg[306]  ( .D(o[306]), .CLK(clk), .RST(rst), .I(g_init[306]), .Q(
        creg[306]) );
  DFF \creg_reg[307]  ( .D(o[307]), .CLK(clk), .RST(rst), .I(g_init[307]), .Q(
        creg[307]) );
  DFF \creg_reg[308]  ( .D(o[308]), .CLK(clk), .RST(rst), .I(g_init[308]), .Q(
        creg[308]) );
  DFF \creg_reg[309]  ( .D(o[309]), .CLK(clk), .RST(rst), .I(g_init[309]), .Q(
        creg[309]) );
  DFF \creg_reg[310]  ( .D(o[310]), .CLK(clk), .RST(rst), .I(g_init[310]), .Q(
        creg[310]) );
  DFF \creg_reg[311]  ( .D(o[311]), .CLK(clk), .RST(rst), .I(g_init[311]), .Q(
        creg[311]) );
  DFF \creg_reg[312]  ( .D(o[312]), .CLK(clk), .RST(rst), .I(g_init[312]), .Q(
        creg[312]) );
  DFF \creg_reg[313]  ( .D(o[313]), .CLK(clk), .RST(rst), .I(g_init[313]), .Q(
        creg[313]) );
  DFF \creg_reg[314]  ( .D(o[314]), .CLK(clk), .RST(rst), .I(g_init[314]), .Q(
        creg[314]) );
  DFF \creg_reg[315]  ( .D(o[315]), .CLK(clk), .RST(rst), .I(g_init[315]), .Q(
        creg[315]) );
  DFF \creg_reg[316]  ( .D(o[316]), .CLK(clk), .RST(rst), .I(g_init[316]), .Q(
        creg[316]) );
  DFF \creg_reg[317]  ( .D(o[317]), .CLK(clk), .RST(rst), .I(g_init[317]), .Q(
        creg[317]) );
  DFF \creg_reg[318]  ( .D(o[318]), .CLK(clk), .RST(rst), .I(g_init[318]), .Q(
        creg[318]) );
  DFF \creg_reg[319]  ( .D(o[319]), .CLK(clk), .RST(rst), .I(g_init[319]), .Q(
        creg[319]) );
  DFF \creg_reg[320]  ( .D(o[320]), .CLK(clk), .RST(rst), .I(g_init[320]), .Q(
        creg[320]) );
  DFF \creg_reg[321]  ( .D(o[321]), .CLK(clk), .RST(rst), .I(g_init[321]), .Q(
        creg[321]) );
  DFF \creg_reg[322]  ( .D(o[322]), .CLK(clk), .RST(rst), .I(g_init[322]), .Q(
        creg[322]) );
  DFF \creg_reg[323]  ( .D(o[323]), .CLK(clk), .RST(rst), .I(g_init[323]), .Q(
        creg[323]) );
  DFF \creg_reg[324]  ( .D(o[324]), .CLK(clk), .RST(rst), .I(g_init[324]), .Q(
        creg[324]) );
  DFF \creg_reg[325]  ( .D(o[325]), .CLK(clk), .RST(rst), .I(g_init[325]), .Q(
        creg[325]) );
  DFF \creg_reg[326]  ( .D(o[326]), .CLK(clk), .RST(rst), .I(g_init[326]), .Q(
        creg[326]) );
  DFF \creg_reg[327]  ( .D(o[327]), .CLK(clk), .RST(rst), .I(g_init[327]), .Q(
        creg[327]) );
  DFF \creg_reg[328]  ( .D(o[328]), .CLK(clk), .RST(rst), .I(g_init[328]), .Q(
        creg[328]) );
  DFF \creg_reg[329]  ( .D(o[329]), .CLK(clk), .RST(rst), .I(g_init[329]), .Q(
        creg[329]) );
  DFF \creg_reg[330]  ( .D(o[330]), .CLK(clk), .RST(rst), .I(g_init[330]), .Q(
        creg[330]) );
  DFF \creg_reg[331]  ( .D(o[331]), .CLK(clk), .RST(rst), .I(g_init[331]), .Q(
        creg[331]) );
  DFF \creg_reg[332]  ( .D(o[332]), .CLK(clk), .RST(rst), .I(g_init[332]), .Q(
        creg[332]) );
  DFF \creg_reg[333]  ( .D(o[333]), .CLK(clk), .RST(rst), .I(g_init[333]), .Q(
        creg[333]) );
  DFF \creg_reg[334]  ( .D(o[334]), .CLK(clk), .RST(rst), .I(g_init[334]), .Q(
        creg[334]) );
  DFF \creg_reg[335]  ( .D(o[335]), .CLK(clk), .RST(rst), .I(g_init[335]), .Q(
        creg[335]) );
  DFF \creg_reg[336]  ( .D(o[336]), .CLK(clk), .RST(rst), .I(g_init[336]), .Q(
        creg[336]) );
  DFF \creg_reg[337]  ( .D(o[337]), .CLK(clk), .RST(rst), .I(g_init[337]), .Q(
        creg[337]) );
  DFF \creg_reg[338]  ( .D(o[338]), .CLK(clk), .RST(rst), .I(g_init[338]), .Q(
        creg[338]) );
  DFF \creg_reg[339]  ( .D(o[339]), .CLK(clk), .RST(rst), .I(g_init[339]), .Q(
        creg[339]) );
  DFF \creg_reg[340]  ( .D(o[340]), .CLK(clk), .RST(rst), .I(g_init[340]), .Q(
        creg[340]) );
  DFF \creg_reg[341]  ( .D(o[341]), .CLK(clk), .RST(rst), .I(g_init[341]), .Q(
        creg[341]) );
  DFF \creg_reg[342]  ( .D(o[342]), .CLK(clk), .RST(rst), .I(g_init[342]), .Q(
        creg[342]) );
  DFF \creg_reg[343]  ( .D(o[343]), .CLK(clk), .RST(rst), .I(g_init[343]), .Q(
        creg[343]) );
  DFF \creg_reg[344]  ( .D(o[344]), .CLK(clk), .RST(rst), .I(g_init[344]), .Q(
        creg[344]) );
  DFF \creg_reg[345]  ( .D(o[345]), .CLK(clk), .RST(rst), .I(g_init[345]), .Q(
        creg[345]) );
  DFF \creg_reg[346]  ( .D(o[346]), .CLK(clk), .RST(rst), .I(g_init[346]), .Q(
        creg[346]) );
  DFF \creg_reg[347]  ( .D(o[347]), .CLK(clk), .RST(rst), .I(g_init[347]), .Q(
        creg[347]) );
  DFF \creg_reg[348]  ( .D(o[348]), .CLK(clk), .RST(rst), .I(g_init[348]), .Q(
        creg[348]) );
  DFF \creg_reg[349]  ( .D(o[349]), .CLK(clk), .RST(rst), .I(g_init[349]), .Q(
        creg[349]) );
  DFF \creg_reg[350]  ( .D(o[350]), .CLK(clk), .RST(rst), .I(g_init[350]), .Q(
        creg[350]) );
  DFF \creg_reg[351]  ( .D(o[351]), .CLK(clk), .RST(rst), .I(g_init[351]), .Q(
        creg[351]) );
  DFF \creg_reg[352]  ( .D(o[352]), .CLK(clk), .RST(rst), .I(g_init[352]), .Q(
        creg[352]) );
  DFF \creg_reg[353]  ( .D(o[353]), .CLK(clk), .RST(rst), .I(g_init[353]), .Q(
        creg[353]) );
  DFF \creg_reg[354]  ( .D(o[354]), .CLK(clk), .RST(rst), .I(g_init[354]), .Q(
        creg[354]) );
  DFF \creg_reg[355]  ( .D(o[355]), .CLK(clk), .RST(rst), .I(g_init[355]), .Q(
        creg[355]) );
  DFF \creg_reg[356]  ( .D(o[356]), .CLK(clk), .RST(rst), .I(g_init[356]), .Q(
        creg[356]) );
  DFF \creg_reg[357]  ( .D(o[357]), .CLK(clk), .RST(rst), .I(g_init[357]), .Q(
        creg[357]) );
  DFF \creg_reg[358]  ( .D(o[358]), .CLK(clk), .RST(rst), .I(g_init[358]), .Q(
        creg[358]) );
  DFF \creg_reg[359]  ( .D(o[359]), .CLK(clk), .RST(rst), .I(g_init[359]), .Q(
        creg[359]) );
  DFF \creg_reg[360]  ( .D(o[360]), .CLK(clk), .RST(rst), .I(g_init[360]), .Q(
        creg[360]) );
  DFF \creg_reg[361]  ( .D(o[361]), .CLK(clk), .RST(rst), .I(g_init[361]), .Q(
        creg[361]) );
  DFF \creg_reg[362]  ( .D(o[362]), .CLK(clk), .RST(rst), .I(g_init[362]), .Q(
        creg[362]) );
  DFF \creg_reg[363]  ( .D(o[363]), .CLK(clk), .RST(rst), .I(g_init[363]), .Q(
        creg[363]) );
  DFF \creg_reg[364]  ( .D(o[364]), .CLK(clk), .RST(rst), .I(g_init[364]), .Q(
        creg[364]) );
  DFF \creg_reg[365]  ( .D(o[365]), .CLK(clk), .RST(rst), .I(g_init[365]), .Q(
        creg[365]) );
  DFF \creg_reg[366]  ( .D(o[366]), .CLK(clk), .RST(rst), .I(g_init[366]), .Q(
        creg[366]) );
  DFF \creg_reg[367]  ( .D(o[367]), .CLK(clk), .RST(rst), .I(g_init[367]), .Q(
        creg[367]) );
  DFF \creg_reg[368]  ( .D(o[368]), .CLK(clk), .RST(rst), .I(g_init[368]), .Q(
        creg[368]) );
  DFF \creg_reg[369]  ( .D(o[369]), .CLK(clk), .RST(rst), .I(g_init[369]), .Q(
        creg[369]) );
  DFF \creg_reg[370]  ( .D(o[370]), .CLK(clk), .RST(rst), .I(g_init[370]), .Q(
        creg[370]) );
  DFF \creg_reg[371]  ( .D(o[371]), .CLK(clk), .RST(rst), .I(g_init[371]), .Q(
        creg[371]) );
  DFF \creg_reg[372]  ( .D(o[372]), .CLK(clk), .RST(rst), .I(g_init[372]), .Q(
        creg[372]) );
  DFF \creg_reg[373]  ( .D(o[373]), .CLK(clk), .RST(rst), .I(g_init[373]), .Q(
        creg[373]) );
  DFF \creg_reg[374]  ( .D(o[374]), .CLK(clk), .RST(rst), .I(g_init[374]), .Q(
        creg[374]) );
  DFF \creg_reg[375]  ( .D(o[375]), .CLK(clk), .RST(rst), .I(g_init[375]), .Q(
        creg[375]) );
  DFF \creg_reg[376]  ( .D(o[376]), .CLK(clk), .RST(rst), .I(g_init[376]), .Q(
        creg[376]) );
  DFF \creg_reg[377]  ( .D(o[377]), .CLK(clk), .RST(rst), .I(g_init[377]), .Q(
        creg[377]) );
  DFF \creg_reg[378]  ( .D(o[378]), .CLK(clk), .RST(rst), .I(g_init[378]), .Q(
        creg[378]) );
  DFF \creg_reg[379]  ( .D(o[379]), .CLK(clk), .RST(rst), .I(g_init[379]), .Q(
        creg[379]) );
  DFF \creg_reg[380]  ( .D(o[380]), .CLK(clk), .RST(rst), .I(g_init[380]), .Q(
        creg[380]) );
  DFF \creg_reg[381]  ( .D(o[381]), .CLK(clk), .RST(rst), .I(g_init[381]), .Q(
        creg[381]) );
  DFF \creg_reg[382]  ( .D(o[382]), .CLK(clk), .RST(rst), .I(g_init[382]), .Q(
        creg[382]) );
  DFF \creg_reg[383]  ( .D(o[383]), .CLK(clk), .RST(rst), .I(g_init[383]), .Q(
        creg[383]) );
  DFF \creg_reg[384]  ( .D(o[384]), .CLK(clk), .RST(rst), .I(g_init[384]), .Q(
        creg[384]) );
  DFF \creg_reg[385]  ( .D(o[385]), .CLK(clk), .RST(rst), .I(g_init[385]), .Q(
        creg[385]) );
  DFF \creg_reg[386]  ( .D(o[386]), .CLK(clk), .RST(rst), .I(g_init[386]), .Q(
        creg[386]) );
  DFF \creg_reg[387]  ( .D(o[387]), .CLK(clk), .RST(rst), .I(g_init[387]), .Q(
        creg[387]) );
  DFF \creg_reg[388]  ( .D(o[388]), .CLK(clk), .RST(rst), .I(g_init[388]), .Q(
        creg[388]) );
  DFF \creg_reg[389]  ( .D(o[389]), .CLK(clk), .RST(rst), .I(g_init[389]), .Q(
        creg[389]) );
  DFF \creg_reg[390]  ( .D(o[390]), .CLK(clk), .RST(rst), .I(g_init[390]), .Q(
        creg[390]) );
  DFF \creg_reg[391]  ( .D(o[391]), .CLK(clk), .RST(rst), .I(g_init[391]), .Q(
        creg[391]) );
  DFF \creg_reg[392]  ( .D(o[392]), .CLK(clk), .RST(rst), .I(g_init[392]), .Q(
        creg[392]) );
  DFF \creg_reg[393]  ( .D(o[393]), .CLK(clk), .RST(rst), .I(g_init[393]), .Q(
        creg[393]) );
  DFF \creg_reg[394]  ( .D(o[394]), .CLK(clk), .RST(rst), .I(g_init[394]), .Q(
        creg[394]) );
  DFF \creg_reg[395]  ( .D(o[395]), .CLK(clk), .RST(rst), .I(g_init[395]), .Q(
        creg[395]) );
  DFF \creg_reg[396]  ( .D(o[396]), .CLK(clk), .RST(rst), .I(g_init[396]), .Q(
        creg[396]) );
  DFF \creg_reg[397]  ( .D(o[397]), .CLK(clk), .RST(rst), .I(g_init[397]), .Q(
        creg[397]) );
  DFF \creg_reg[398]  ( .D(o[398]), .CLK(clk), .RST(rst), .I(g_init[398]), .Q(
        creg[398]) );
  DFF \creg_reg[399]  ( .D(o[399]), .CLK(clk), .RST(rst), .I(g_init[399]), .Q(
        creg[399]) );
  DFF \creg_reg[400]  ( .D(o[400]), .CLK(clk), .RST(rst), .I(g_init[400]), .Q(
        creg[400]) );
  DFF \creg_reg[401]  ( .D(o[401]), .CLK(clk), .RST(rst), .I(g_init[401]), .Q(
        creg[401]) );
  DFF \creg_reg[402]  ( .D(o[402]), .CLK(clk), .RST(rst), .I(g_init[402]), .Q(
        creg[402]) );
  DFF \creg_reg[403]  ( .D(o[403]), .CLK(clk), .RST(rst), .I(g_init[403]), .Q(
        creg[403]) );
  DFF \creg_reg[404]  ( .D(o[404]), .CLK(clk), .RST(rst), .I(g_init[404]), .Q(
        creg[404]) );
  DFF \creg_reg[405]  ( .D(o[405]), .CLK(clk), .RST(rst), .I(g_init[405]), .Q(
        creg[405]) );
  DFF \creg_reg[406]  ( .D(o[406]), .CLK(clk), .RST(rst), .I(g_init[406]), .Q(
        creg[406]) );
  DFF \creg_reg[407]  ( .D(o[407]), .CLK(clk), .RST(rst), .I(g_init[407]), .Q(
        creg[407]) );
  DFF \creg_reg[408]  ( .D(o[408]), .CLK(clk), .RST(rst), .I(g_init[408]), .Q(
        creg[408]) );
  DFF \creg_reg[409]  ( .D(o[409]), .CLK(clk), .RST(rst), .I(g_init[409]), .Q(
        creg[409]) );
  DFF \creg_reg[410]  ( .D(o[410]), .CLK(clk), .RST(rst), .I(g_init[410]), .Q(
        creg[410]) );
  DFF \creg_reg[411]  ( .D(o[411]), .CLK(clk), .RST(rst), .I(g_init[411]), .Q(
        creg[411]) );
  DFF \creg_reg[412]  ( .D(o[412]), .CLK(clk), .RST(rst), .I(g_init[412]), .Q(
        creg[412]) );
  DFF \creg_reg[413]  ( .D(o[413]), .CLK(clk), .RST(rst), .I(g_init[413]), .Q(
        creg[413]) );
  DFF \creg_reg[414]  ( .D(o[414]), .CLK(clk), .RST(rst), .I(g_init[414]), .Q(
        creg[414]) );
  DFF \creg_reg[415]  ( .D(o[415]), .CLK(clk), .RST(rst), .I(g_init[415]), .Q(
        creg[415]) );
  DFF \creg_reg[416]  ( .D(o[416]), .CLK(clk), .RST(rst), .I(g_init[416]), .Q(
        creg[416]) );
  DFF \creg_reg[417]  ( .D(o[417]), .CLK(clk), .RST(rst), .I(g_init[417]), .Q(
        creg[417]) );
  DFF \creg_reg[418]  ( .D(o[418]), .CLK(clk), .RST(rst), .I(g_init[418]), .Q(
        creg[418]) );
  DFF \creg_reg[419]  ( .D(o[419]), .CLK(clk), .RST(rst), .I(g_init[419]), .Q(
        creg[419]) );
  DFF \creg_reg[420]  ( .D(o[420]), .CLK(clk), .RST(rst), .I(g_init[420]), .Q(
        creg[420]) );
  DFF \creg_reg[421]  ( .D(o[421]), .CLK(clk), .RST(rst), .I(g_init[421]), .Q(
        creg[421]) );
  DFF \creg_reg[422]  ( .D(o[422]), .CLK(clk), .RST(rst), .I(g_init[422]), .Q(
        creg[422]) );
  DFF \creg_reg[423]  ( .D(o[423]), .CLK(clk), .RST(rst), .I(g_init[423]), .Q(
        creg[423]) );
  DFF \creg_reg[424]  ( .D(o[424]), .CLK(clk), .RST(rst), .I(g_init[424]), .Q(
        creg[424]) );
  DFF \creg_reg[425]  ( .D(o[425]), .CLK(clk), .RST(rst), .I(g_init[425]), .Q(
        creg[425]) );
  DFF \creg_reg[426]  ( .D(o[426]), .CLK(clk), .RST(rst), .I(g_init[426]), .Q(
        creg[426]) );
  DFF \creg_reg[427]  ( .D(o[427]), .CLK(clk), .RST(rst), .I(g_init[427]), .Q(
        creg[427]) );
  DFF \creg_reg[428]  ( .D(o[428]), .CLK(clk), .RST(rst), .I(g_init[428]), .Q(
        creg[428]) );
  DFF \creg_reg[429]  ( .D(o[429]), .CLK(clk), .RST(rst), .I(g_init[429]), .Q(
        creg[429]) );
  DFF \creg_reg[430]  ( .D(o[430]), .CLK(clk), .RST(rst), .I(g_init[430]), .Q(
        creg[430]) );
  DFF \creg_reg[431]  ( .D(o[431]), .CLK(clk), .RST(rst), .I(g_init[431]), .Q(
        creg[431]) );
  DFF \creg_reg[432]  ( .D(o[432]), .CLK(clk), .RST(rst), .I(g_init[432]), .Q(
        creg[432]) );
  DFF \creg_reg[433]  ( .D(o[433]), .CLK(clk), .RST(rst), .I(g_init[433]), .Q(
        creg[433]) );
  DFF \creg_reg[434]  ( .D(o[434]), .CLK(clk), .RST(rst), .I(g_init[434]), .Q(
        creg[434]) );
  DFF \creg_reg[435]  ( .D(o[435]), .CLK(clk), .RST(rst), .I(g_init[435]), .Q(
        creg[435]) );
  DFF \creg_reg[436]  ( .D(o[436]), .CLK(clk), .RST(rst), .I(g_init[436]), .Q(
        creg[436]) );
  DFF \creg_reg[437]  ( .D(o[437]), .CLK(clk), .RST(rst), .I(g_init[437]), .Q(
        creg[437]) );
  DFF \creg_reg[438]  ( .D(o[438]), .CLK(clk), .RST(rst), .I(g_init[438]), .Q(
        creg[438]) );
  DFF \creg_reg[439]  ( .D(o[439]), .CLK(clk), .RST(rst), .I(g_init[439]), .Q(
        creg[439]) );
  DFF \creg_reg[440]  ( .D(o[440]), .CLK(clk), .RST(rst), .I(g_init[440]), .Q(
        creg[440]) );
  DFF \creg_reg[441]  ( .D(o[441]), .CLK(clk), .RST(rst), .I(g_init[441]), .Q(
        creg[441]) );
  DFF \creg_reg[442]  ( .D(o[442]), .CLK(clk), .RST(rst), .I(g_init[442]), .Q(
        creg[442]) );
  DFF \creg_reg[443]  ( .D(o[443]), .CLK(clk), .RST(rst), .I(g_init[443]), .Q(
        creg[443]) );
  DFF \creg_reg[444]  ( .D(o[444]), .CLK(clk), .RST(rst), .I(g_init[444]), .Q(
        creg[444]) );
  DFF \creg_reg[445]  ( .D(o[445]), .CLK(clk), .RST(rst), .I(g_init[445]), .Q(
        creg[445]) );
  DFF \creg_reg[446]  ( .D(o[446]), .CLK(clk), .RST(rst), .I(g_init[446]), .Q(
        creg[446]) );
  DFF \creg_reg[447]  ( .D(o[447]), .CLK(clk), .RST(rst), .I(g_init[447]), .Q(
        creg[447]) );
  DFF \creg_reg[448]  ( .D(o[448]), .CLK(clk), .RST(rst), .I(g_init[448]), .Q(
        creg[448]) );
  DFF \creg_reg[449]  ( .D(o[449]), .CLK(clk), .RST(rst), .I(g_init[449]), .Q(
        creg[449]) );
  DFF \creg_reg[450]  ( .D(o[450]), .CLK(clk), .RST(rst), .I(g_init[450]), .Q(
        creg[450]) );
  DFF \creg_reg[451]  ( .D(o[451]), .CLK(clk), .RST(rst), .I(g_init[451]), .Q(
        creg[451]) );
  DFF \creg_reg[452]  ( .D(o[452]), .CLK(clk), .RST(rst), .I(g_init[452]), .Q(
        creg[452]) );
  DFF \creg_reg[453]  ( .D(o[453]), .CLK(clk), .RST(rst), .I(g_init[453]), .Q(
        creg[453]) );
  DFF \creg_reg[454]  ( .D(o[454]), .CLK(clk), .RST(rst), .I(g_init[454]), .Q(
        creg[454]) );
  DFF \creg_reg[455]  ( .D(o[455]), .CLK(clk), .RST(rst), .I(g_init[455]), .Q(
        creg[455]) );
  DFF \creg_reg[456]  ( .D(o[456]), .CLK(clk), .RST(rst), .I(g_init[456]), .Q(
        creg[456]) );
  DFF \creg_reg[457]  ( .D(o[457]), .CLK(clk), .RST(rst), .I(g_init[457]), .Q(
        creg[457]) );
  DFF \creg_reg[458]  ( .D(o[458]), .CLK(clk), .RST(rst), .I(g_init[458]), .Q(
        creg[458]) );
  DFF \creg_reg[459]  ( .D(o[459]), .CLK(clk), .RST(rst), .I(g_init[459]), .Q(
        creg[459]) );
  DFF \creg_reg[460]  ( .D(o[460]), .CLK(clk), .RST(rst), .I(g_init[460]), .Q(
        creg[460]) );
  DFF \creg_reg[461]  ( .D(o[461]), .CLK(clk), .RST(rst), .I(g_init[461]), .Q(
        creg[461]) );
  DFF \creg_reg[462]  ( .D(o[462]), .CLK(clk), .RST(rst), .I(g_init[462]), .Q(
        creg[462]) );
  DFF \creg_reg[463]  ( .D(o[463]), .CLK(clk), .RST(rst), .I(g_init[463]), .Q(
        creg[463]) );
  DFF \creg_reg[464]  ( .D(o[464]), .CLK(clk), .RST(rst), .I(g_init[464]), .Q(
        creg[464]) );
  DFF \creg_reg[465]  ( .D(o[465]), .CLK(clk), .RST(rst), .I(g_init[465]), .Q(
        creg[465]) );
  DFF \creg_reg[466]  ( .D(o[466]), .CLK(clk), .RST(rst), .I(g_init[466]), .Q(
        creg[466]) );
  DFF \creg_reg[467]  ( .D(o[467]), .CLK(clk), .RST(rst), .I(g_init[467]), .Q(
        creg[467]) );
  DFF \creg_reg[468]  ( .D(o[468]), .CLK(clk), .RST(rst), .I(g_init[468]), .Q(
        creg[468]) );
  DFF \creg_reg[469]  ( .D(o[469]), .CLK(clk), .RST(rst), .I(g_init[469]), .Q(
        creg[469]) );
  DFF \creg_reg[470]  ( .D(o[470]), .CLK(clk), .RST(rst), .I(g_init[470]), .Q(
        creg[470]) );
  DFF \creg_reg[471]  ( .D(o[471]), .CLK(clk), .RST(rst), .I(g_init[471]), .Q(
        creg[471]) );
  DFF \creg_reg[472]  ( .D(o[472]), .CLK(clk), .RST(rst), .I(g_init[472]), .Q(
        creg[472]) );
  DFF \creg_reg[473]  ( .D(o[473]), .CLK(clk), .RST(rst), .I(g_init[473]), .Q(
        creg[473]) );
  DFF \creg_reg[474]  ( .D(o[474]), .CLK(clk), .RST(rst), .I(g_init[474]), .Q(
        creg[474]) );
  DFF \creg_reg[475]  ( .D(o[475]), .CLK(clk), .RST(rst), .I(g_init[475]), .Q(
        creg[475]) );
  DFF \creg_reg[476]  ( .D(o[476]), .CLK(clk), .RST(rst), .I(g_init[476]), .Q(
        creg[476]) );
  DFF \creg_reg[477]  ( .D(o[477]), .CLK(clk), .RST(rst), .I(g_init[477]), .Q(
        creg[477]) );
  DFF \creg_reg[478]  ( .D(o[478]), .CLK(clk), .RST(rst), .I(g_init[478]), .Q(
        creg[478]) );
  DFF \creg_reg[479]  ( .D(o[479]), .CLK(clk), .RST(rst), .I(g_init[479]), .Q(
        creg[479]) );
  DFF \creg_reg[480]  ( .D(o[480]), .CLK(clk), .RST(rst), .I(g_init[480]), .Q(
        creg[480]) );
  DFF \creg_reg[481]  ( .D(o[481]), .CLK(clk), .RST(rst), .I(g_init[481]), .Q(
        creg[481]) );
  DFF \creg_reg[482]  ( .D(o[482]), .CLK(clk), .RST(rst), .I(g_init[482]), .Q(
        creg[482]) );
  DFF \creg_reg[483]  ( .D(o[483]), .CLK(clk), .RST(rst), .I(g_init[483]), .Q(
        creg[483]) );
  DFF \creg_reg[484]  ( .D(o[484]), .CLK(clk), .RST(rst), .I(g_init[484]), .Q(
        creg[484]) );
  DFF \creg_reg[485]  ( .D(o[485]), .CLK(clk), .RST(rst), .I(g_init[485]), .Q(
        creg[485]) );
  DFF \creg_reg[486]  ( .D(o[486]), .CLK(clk), .RST(rst), .I(g_init[486]), .Q(
        creg[486]) );
  DFF \creg_reg[487]  ( .D(o[487]), .CLK(clk), .RST(rst), .I(g_init[487]), .Q(
        creg[487]) );
  DFF \creg_reg[488]  ( .D(o[488]), .CLK(clk), .RST(rst), .I(g_init[488]), .Q(
        creg[488]) );
  DFF \creg_reg[489]  ( .D(o[489]), .CLK(clk), .RST(rst), .I(g_init[489]), .Q(
        creg[489]) );
  DFF \creg_reg[490]  ( .D(o[490]), .CLK(clk), .RST(rst), .I(g_init[490]), .Q(
        creg[490]) );
  DFF \creg_reg[491]  ( .D(o[491]), .CLK(clk), .RST(rst), .I(g_init[491]), .Q(
        creg[491]) );
  DFF \creg_reg[492]  ( .D(o[492]), .CLK(clk), .RST(rst), .I(g_init[492]), .Q(
        creg[492]) );
  DFF \creg_reg[493]  ( .D(o[493]), .CLK(clk), .RST(rst), .I(g_init[493]), .Q(
        creg[493]) );
  DFF \creg_reg[494]  ( .D(o[494]), .CLK(clk), .RST(rst), .I(g_init[494]), .Q(
        creg[494]) );
  DFF \creg_reg[495]  ( .D(o[495]), .CLK(clk), .RST(rst), .I(g_init[495]), .Q(
        creg[495]) );
  DFF \creg_reg[496]  ( .D(o[496]), .CLK(clk), .RST(rst), .I(g_init[496]), .Q(
        creg[496]) );
  DFF \creg_reg[497]  ( .D(o[497]), .CLK(clk), .RST(rst), .I(g_init[497]), .Q(
        creg[497]) );
  DFF \creg_reg[498]  ( .D(o[498]), .CLK(clk), .RST(rst), .I(g_init[498]), .Q(
        creg[498]) );
  DFF \creg_reg[499]  ( .D(o[499]), .CLK(clk), .RST(rst), .I(g_init[499]), .Q(
        creg[499]) );
  DFF \creg_reg[500]  ( .D(o[500]), .CLK(clk), .RST(rst), .I(g_init[500]), .Q(
        creg[500]) );
  DFF \creg_reg[501]  ( .D(o[501]), .CLK(clk), .RST(rst), .I(g_init[501]), .Q(
        creg[501]) );
  DFF \creg_reg[502]  ( .D(o[502]), .CLK(clk), .RST(rst), .I(g_init[502]), .Q(
        creg[502]) );
  DFF \creg_reg[503]  ( .D(o[503]), .CLK(clk), .RST(rst), .I(g_init[503]), .Q(
        creg[503]) );
  DFF \creg_reg[504]  ( .D(o[504]), .CLK(clk), .RST(rst), .I(g_init[504]), .Q(
        creg[504]) );
  DFF \creg_reg[505]  ( .D(o[505]), .CLK(clk), .RST(rst), .I(g_init[505]), .Q(
        creg[505]) );
  DFF \creg_reg[506]  ( .D(o[506]), .CLK(clk), .RST(rst), .I(g_init[506]), .Q(
        creg[506]) );
  DFF \creg_reg[507]  ( .D(o[507]), .CLK(clk), .RST(rst), .I(g_init[507]), .Q(
        creg[507]) );
  DFF \creg_reg[508]  ( .D(o[508]), .CLK(clk), .RST(rst), .I(g_init[508]), .Q(
        creg[508]) );
  DFF \creg_reg[509]  ( .D(o[509]), .CLK(clk), .RST(rst), .I(g_init[509]), .Q(
        creg[509]) );
  DFF \creg_reg[510]  ( .D(o[510]), .CLK(clk), .RST(rst), .I(g_init[510]), .Q(
        creg[510]) );
  DFF \creg_reg[511]  ( .D(o[511]), .CLK(clk), .RST(rst), .I(g_init[511]), .Q(
        creg[511]) );
  DFF \creg_reg[512]  ( .D(o[512]), .CLK(clk), .RST(rst), .I(g_init[512]), .Q(
        creg[512]) );
  DFF \creg_reg[513]  ( .D(o[513]), .CLK(clk), .RST(rst), .I(g_init[513]), .Q(
        creg[513]) );
  DFF \creg_reg[514]  ( .D(o[514]), .CLK(clk), .RST(rst), .I(g_init[514]), .Q(
        creg[514]) );
  DFF \creg_reg[515]  ( .D(o[515]), .CLK(clk), .RST(rst), .I(g_init[515]), .Q(
        creg[515]) );
  DFF \creg_reg[516]  ( .D(o[516]), .CLK(clk), .RST(rst), .I(g_init[516]), .Q(
        creg[516]) );
  DFF \creg_reg[517]  ( .D(o[517]), .CLK(clk), .RST(rst), .I(g_init[517]), .Q(
        creg[517]) );
  DFF \creg_reg[518]  ( .D(o[518]), .CLK(clk), .RST(rst), .I(g_init[518]), .Q(
        creg[518]) );
  DFF \creg_reg[519]  ( .D(o[519]), .CLK(clk), .RST(rst), .I(g_init[519]), .Q(
        creg[519]) );
  DFF \creg_reg[520]  ( .D(o[520]), .CLK(clk), .RST(rst), .I(g_init[520]), .Q(
        creg[520]) );
  DFF \creg_reg[521]  ( .D(o[521]), .CLK(clk), .RST(rst), .I(g_init[521]), .Q(
        creg[521]) );
  DFF \creg_reg[522]  ( .D(o[522]), .CLK(clk), .RST(rst), .I(g_init[522]), .Q(
        creg[522]) );
  DFF \creg_reg[523]  ( .D(o[523]), .CLK(clk), .RST(rst), .I(g_init[523]), .Q(
        creg[523]) );
  DFF \creg_reg[524]  ( .D(o[524]), .CLK(clk), .RST(rst), .I(g_init[524]), .Q(
        creg[524]) );
  DFF \creg_reg[525]  ( .D(o[525]), .CLK(clk), .RST(rst), .I(g_init[525]), .Q(
        creg[525]) );
  DFF \creg_reg[526]  ( .D(o[526]), .CLK(clk), .RST(rst), .I(g_init[526]), .Q(
        creg[526]) );
  DFF \creg_reg[527]  ( .D(o[527]), .CLK(clk), .RST(rst), .I(g_init[527]), .Q(
        creg[527]) );
  DFF \creg_reg[528]  ( .D(o[528]), .CLK(clk), .RST(rst), .I(g_init[528]), .Q(
        creg[528]) );
  DFF \creg_reg[529]  ( .D(o[529]), .CLK(clk), .RST(rst), .I(g_init[529]), .Q(
        creg[529]) );
  DFF \creg_reg[530]  ( .D(o[530]), .CLK(clk), .RST(rst), .I(g_init[530]), .Q(
        creg[530]) );
  DFF \creg_reg[531]  ( .D(o[531]), .CLK(clk), .RST(rst), .I(g_init[531]), .Q(
        creg[531]) );
  DFF \creg_reg[532]  ( .D(o[532]), .CLK(clk), .RST(rst), .I(g_init[532]), .Q(
        creg[532]) );
  DFF \creg_reg[533]  ( .D(o[533]), .CLK(clk), .RST(rst), .I(g_init[533]), .Q(
        creg[533]) );
  DFF \creg_reg[534]  ( .D(o[534]), .CLK(clk), .RST(rst), .I(g_init[534]), .Q(
        creg[534]) );
  DFF \creg_reg[535]  ( .D(o[535]), .CLK(clk), .RST(rst), .I(g_init[535]), .Q(
        creg[535]) );
  DFF \creg_reg[536]  ( .D(o[536]), .CLK(clk), .RST(rst), .I(g_init[536]), .Q(
        creg[536]) );
  DFF \creg_reg[537]  ( .D(o[537]), .CLK(clk), .RST(rst), .I(g_init[537]), .Q(
        creg[537]) );
  DFF \creg_reg[538]  ( .D(o[538]), .CLK(clk), .RST(rst), .I(g_init[538]), .Q(
        creg[538]) );
  DFF \creg_reg[539]  ( .D(o[539]), .CLK(clk), .RST(rst), .I(g_init[539]), .Q(
        creg[539]) );
  DFF \creg_reg[540]  ( .D(o[540]), .CLK(clk), .RST(rst), .I(g_init[540]), .Q(
        creg[540]) );
  DFF \creg_reg[541]  ( .D(o[541]), .CLK(clk), .RST(rst), .I(g_init[541]), .Q(
        creg[541]) );
  DFF \creg_reg[542]  ( .D(o[542]), .CLK(clk), .RST(rst), .I(g_init[542]), .Q(
        creg[542]) );
  DFF \creg_reg[543]  ( .D(o[543]), .CLK(clk), .RST(rst), .I(g_init[543]), .Q(
        creg[543]) );
  DFF \creg_reg[544]  ( .D(o[544]), .CLK(clk), .RST(rst), .I(g_init[544]), .Q(
        creg[544]) );
  DFF \creg_reg[545]  ( .D(o[545]), .CLK(clk), .RST(rst), .I(g_init[545]), .Q(
        creg[545]) );
  DFF \creg_reg[546]  ( .D(o[546]), .CLK(clk), .RST(rst), .I(g_init[546]), .Q(
        creg[546]) );
  DFF \creg_reg[547]  ( .D(o[547]), .CLK(clk), .RST(rst), .I(g_init[547]), .Q(
        creg[547]) );
  DFF \creg_reg[548]  ( .D(o[548]), .CLK(clk), .RST(rst), .I(g_init[548]), .Q(
        creg[548]) );
  DFF \creg_reg[549]  ( .D(o[549]), .CLK(clk), .RST(rst), .I(g_init[549]), .Q(
        creg[549]) );
  DFF \creg_reg[550]  ( .D(o[550]), .CLK(clk), .RST(rst), .I(g_init[550]), .Q(
        creg[550]) );
  DFF \creg_reg[551]  ( .D(o[551]), .CLK(clk), .RST(rst), .I(g_init[551]), .Q(
        creg[551]) );
  DFF \creg_reg[552]  ( .D(o[552]), .CLK(clk), .RST(rst), .I(g_init[552]), .Q(
        creg[552]) );
  DFF \creg_reg[553]  ( .D(o[553]), .CLK(clk), .RST(rst), .I(g_init[553]), .Q(
        creg[553]) );
  DFF \creg_reg[554]  ( .D(o[554]), .CLK(clk), .RST(rst), .I(g_init[554]), .Q(
        creg[554]) );
  DFF \creg_reg[555]  ( .D(o[555]), .CLK(clk), .RST(rst), .I(g_init[555]), .Q(
        creg[555]) );
  DFF \creg_reg[556]  ( .D(o[556]), .CLK(clk), .RST(rst), .I(g_init[556]), .Q(
        creg[556]) );
  DFF \creg_reg[557]  ( .D(o[557]), .CLK(clk), .RST(rst), .I(g_init[557]), .Q(
        creg[557]) );
  DFF \creg_reg[558]  ( .D(o[558]), .CLK(clk), .RST(rst), .I(g_init[558]), .Q(
        creg[558]) );
  DFF \creg_reg[559]  ( .D(o[559]), .CLK(clk), .RST(rst), .I(g_init[559]), .Q(
        creg[559]) );
  DFF \creg_reg[560]  ( .D(o[560]), .CLK(clk), .RST(rst), .I(g_init[560]), .Q(
        creg[560]) );
  DFF \creg_reg[561]  ( .D(o[561]), .CLK(clk), .RST(rst), .I(g_init[561]), .Q(
        creg[561]) );
  DFF \creg_reg[562]  ( .D(o[562]), .CLK(clk), .RST(rst), .I(g_init[562]), .Q(
        creg[562]) );
  DFF \creg_reg[563]  ( .D(o[563]), .CLK(clk), .RST(rst), .I(g_init[563]), .Q(
        creg[563]) );
  DFF \creg_reg[564]  ( .D(o[564]), .CLK(clk), .RST(rst), .I(g_init[564]), .Q(
        creg[564]) );
  DFF \creg_reg[565]  ( .D(o[565]), .CLK(clk), .RST(rst), .I(g_init[565]), .Q(
        creg[565]) );
  DFF \creg_reg[566]  ( .D(o[566]), .CLK(clk), .RST(rst), .I(g_init[566]), .Q(
        creg[566]) );
  DFF \creg_reg[567]  ( .D(o[567]), .CLK(clk), .RST(rst), .I(g_init[567]), .Q(
        creg[567]) );
  DFF \creg_reg[568]  ( .D(o[568]), .CLK(clk), .RST(rst), .I(g_init[568]), .Q(
        creg[568]) );
  DFF \creg_reg[569]  ( .D(o[569]), .CLK(clk), .RST(rst), .I(g_init[569]), .Q(
        creg[569]) );
  DFF \creg_reg[570]  ( .D(o[570]), .CLK(clk), .RST(rst), .I(g_init[570]), .Q(
        creg[570]) );
  DFF \creg_reg[571]  ( .D(o[571]), .CLK(clk), .RST(rst), .I(g_init[571]), .Q(
        creg[571]) );
  DFF \creg_reg[572]  ( .D(o[572]), .CLK(clk), .RST(rst), .I(g_init[572]), .Q(
        creg[572]) );
  DFF \creg_reg[573]  ( .D(o[573]), .CLK(clk), .RST(rst), .I(g_init[573]), .Q(
        creg[573]) );
  DFF \creg_reg[574]  ( .D(o[574]), .CLK(clk), .RST(rst), .I(g_init[574]), .Q(
        creg[574]) );
  DFF \creg_reg[575]  ( .D(o[575]), .CLK(clk), .RST(rst), .I(g_init[575]), .Q(
        creg[575]) );
  DFF \creg_reg[576]  ( .D(o[576]), .CLK(clk), .RST(rst), .I(g_init[576]), .Q(
        creg[576]) );
  DFF \creg_reg[577]  ( .D(o[577]), .CLK(clk), .RST(rst), .I(g_init[577]), .Q(
        creg[577]) );
  DFF \creg_reg[578]  ( .D(o[578]), .CLK(clk), .RST(rst), .I(g_init[578]), .Q(
        creg[578]) );
  DFF \creg_reg[579]  ( .D(o[579]), .CLK(clk), .RST(rst), .I(g_init[579]), .Q(
        creg[579]) );
  DFF \creg_reg[580]  ( .D(o[580]), .CLK(clk), .RST(rst), .I(g_init[580]), .Q(
        creg[580]) );
  DFF \creg_reg[581]  ( .D(o[581]), .CLK(clk), .RST(rst), .I(g_init[581]), .Q(
        creg[581]) );
  DFF \creg_reg[582]  ( .D(o[582]), .CLK(clk), .RST(rst), .I(g_init[582]), .Q(
        creg[582]) );
  DFF \creg_reg[583]  ( .D(o[583]), .CLK(clk), .RST(rst), .I(g_init[583]), .Q(
        creg[583]) );
  DFF \creg_reg[584]  ( .D(o[584]), .CLK(clk), .RST(rst), .I(g_init[584]), .Q(
        creg[584]) );
  DFF \creg_reg[585]  ( .D(o[585]), .CLK(clk), .RST(rst), .I(g_init[585]), .Q(
        creg[585]) );
  DFF \creg_reg[586]  ( .D(o[586]), .CLK(clk), .RST(rst), .I(g_init[586]), .Q(
        creg[586]) );
  DFF \creg_reg[587]  ( .D(o[587]), .CLK(clk), .RST(rst), .I(g_init[587]), .Q(
        creg[587]) );
  DFF \creg_reg[588]  ( .D(o[588]), .CLK(clk), .RST(rst), .I(g_init[588]), .Q(
        creg[588]) );
  DFF \creg_reg[589]  ( .D(o[589]), .CLK(clk), .RST(rst), .I(g_init[589]), .Q(
        creg[589]) );
  DFF \creg_reg[590]  ( .D(o[590]), .CLK(clk), .RST(rst), .I(g_init[590]), .Q(
        creg[590]) );
  DFF \creg_reg[591]  ( .D(o[591]), .CLK(clk), .RST(rst), .I(g_init[591]), .Q(
        creg[591]) );
  DFF \creg_reg[592]  ( .D(o[592]), .CLK(clk), .RST(rst), .I(g_init[592]), .Q(
        creg[592]) );
  DFF \creg_reg[593]  ( .D(o[593]), .CLK(clk), .RST(rst), .I(g_init[593]), .Q(
        creg[593]) );
  DFF \creg_reg[594]  ( .D(o[594]), .CLK(clk), .RST(rst), .I(g_init[594]), .Q(
        creg[594]) );
  DFF \creg_reg[595]  ( .D(o[595]), .CLK(clk), .RST(rst), .I(g_init[595]), .Q(
        creg[595]) );
  DFF \creg_reg[596]  ( .D(o[596]), .CLK(clk), .RST(rst), .I(g_init[596]), .Q(
        creg[596]) );
  DFF \creg_reg[597]  ( .D(o[597]), .CLK(clk), .RST(rst), .I(g_init[597]), .Q(
        creg[597]) );
  DFF \creg_reg[598]  ( .D(o[598]), .CLK(clk), .RST(rst), .I(g_init[598]), .Q(
        creg[598]) );
  DFF \creg_reg[599]  ( .D(o[599]), .CLK(clk), .RST(rst), .I(g_init[599]), .Q(
        creg[599]) );
  DFF \creg_reg[600]  ( .D(o[600]), .CLK(clk), .RST(rst), .I(g_init[600]), .Q(
        creg[600]) );
  DFF \creg_reg[601]  ( .D(o[601]), .CLK(clk), .RST(rst), .I(g_init[601]), .Q(
        creg[601]) );
  DFF \creg_reg[602]  ( .D(o[602]), .CLK(clk), .RST(rst), .I(g_init[602]), .Q(
        creg[602]) );
  DFF \creg_reg[603]  ( .D(o[603]), .CLK(clk), .RST(rst), .I(g_init[603]), .Q(
        creg[603]) );
  DFF \creg_reg[604]  ( .D(o[604]), .CLK(clk), .RST(rst), .I(g_init[604]), .Q(
        creg[604]) );
  DFF \creg_reg[605]  ( .D(o[605]), .CLK(clk), .RST(rst), .I(g_init[605]), .Q(
        creg[605]) );
  DFF \creg_reg[606]  ( .D(o[606]), .CLK(clk), .RST(rst), .I(g_init[606]), .Q(
        creg[606]) );
  DFF \creg_reg[607]  ( .D(o[607]), .CLK(clk), .RST(rst), .I(g_init[607]), .Q(
        creg[607]) );
  DFF \creg_reg[608]  ( .D(o[608]), .CLK(clk), .RST(rst), .I(g_init[608]), .Q(
        creg[608]) );
  DFF \creg_reg[609]  ( .D(o[609]), .CLK(clk), .RST(rst), .I(g_init[609]), .Q(
        creg[609]) );
  DFF \creg_reg[610]  ( .D(o[610]), .CLK(clk), .RST(rst), .I(g_init[610]), .Q(
        creg[610]) );
  DFF \creg_reg[611]  ( .D(o[611]), .CLK(clk), .RST(rst), .I(g_init[611]), .Q(
        creg[611]) );
  DFF \creg_reg[612]  ( .D(o[612]), .CLK(clk), .RST(rst), .I(g_init[612]), .Q(
        creg[612]) );
  DFF \creg_reg[613]  ( .D(o[613]), .CLK(clk), .RST(rst), .I(g_init[613]), .Q(
        creg[613]) );
  DFF \creg_reg[614]  ( .D(o[614]), .CLK(clk), .RST(rst), .I(g_init[614]), .Q(
        creg[614]) );
  DFF \creg_reg[615]  ( .D(o[615]), .CLK(clk), .RST(rst), .I(g_init[615]), .Q(
        creg[615]) );
  DFF \creg_reg[616]  ( .D(o[616]), .CLK(clk), .RST(rst), .I(g_init[616]), .Q(
        creg[616]) );
  DFF \creg_reg[617]  ( .D(o[617]), .CLK(clk), .RST(rst), .I(g_init[617]), .Q(
        creg[617]) );
  DFF \creg_reg[618]  ( .D(o[618]), .CLK(clk), .RST(rst), .I(g_init[618]), .Q(
        creg[618]) );
  DFF \creg_reg[619]  ( .D(o[619]), .CLK(clk), .RST(rst), .I(g_init[619]), .Q(
        creg[619]) );
  DFF \creg_reg[620]  ( .D(o[620]), .CLK(clk), .RST(rst), .I(g_init[620]), .Q(
        creg[620]) );
  DFF \creg_reg[621]  ( .D(o[621]), .CLK(clk), .RST(rst), .I(g_init[621]), .Q(
        creg[621]) );
  DFF \creg_reg[622]  ( .D(o[622]), .CLK(clk), .RST(rst), .I(g_init[622]), .Q(
        creg[622]) );
  DFF \creg_reg[623]  ( .D(o[623]), .CLK(clk), .RST(rst), .I(g_init[623]), .Q(
        creg[623]) );
  DFF \creg_reg[624]  ( .D(o[624]), .CLK(clk), .RST(rst), .I(g_init[624]), .Q(
        creg[624]) );
  DFF \creg_reg[625]  ( .D(o[625]), .CLK(clk), .RST(rst), .I(g_init[625]), .Q(
        creg[625]) );
  DFF \creg_reg[626]  ( .D(o[626]), .CLK(clk), .RST(rst), .I(g_init[626]), .Q(
        creg[626]) );
  DFF \creg_reg[627]  ( .D(o[627]), .CLK(clk), .RST(rst), .I(g_init[627]), .Q(
        creg[627]) );
  DFF \creg_reg[628]  ( .D(o[628]), .CLK(clk), .RST(rst), .I(g_init[628]), .Q(
        creg[628]) );
  DFF \creg_reg[629]  ( .D(o[629]), .CLK(clk), .RST(rst), .I(g_init[629]), .Q(
        creg[629]) );
  DFF \creg_reg[630]  ( .D(o[630]), .CLK(clk), .RST(rst), .I(g_init[630]), .Q(
        creg[630]) );
  DFF \creg_reg[631]  ( .D(o[631]), .CLK(clk), .RST(rst), .I(g_init[631]), .Q(
        creg[631]) );
  DFF \creg_reg[632]  ( .D(o[632]), .CLK(clk), .RST(rst), .I(g_init[632]), .Q(
        creg[632]) );
  DFF \creg_reg[633]  ( .D(o[633]), .CLK(clk), .RST(rst), .I(g_init[633]), .Q(
        creg[633]) );
  DFF \creg_reg[634]  ( .D(o[634]), .CLK(clk), .RST(rst), .I(g_init[634]), .Q(
        creg[634]) );
  DFF \creg_reg[635]  ( .D(o[635]), .CLK(clk), .RST(rst), .I(g_init[635]), .Q(
        creg[635]) );
  DFF \creg_reg[636]  ( .D(o[636]), .CLK(clk), .RST(rst), .I(g_init[636]), .Q(
        creg[636]) );
  DFF \creg_reg[637]  ( .D(o[637]), .CLK(clk), .RST(rst), .I(g_init[637]), .Q(
        creg[637]) );
  DFF \creg_reg[638]  ( .D(o[638]), .CLK(clk), .RST(rst), .I(g_init[638]), .Q(
        creg[638]) );
  DFF \creg_reg[639]  ( .D(o[639]), .CLK(clk), .RST(rst), .I(g_init[639]), .Q(
        creg[639]) );
  DFF \creg_reg[640]  ( .D(o[640]), .CLK(clk), .RST(rst), .I(g_init[640]), .Q(
        creg[640]) );
  DFF \creg_reg[641]  ( .D(o[641]), .CLK(clk), .RST(rst), .I(g_init[641]), .Q(
        creg[641]) );
  DFF \creg_reg[642]  ( .D(o[642]), .CLK(clk), .RST(rst), .I(g_init[642]), .Q(
        creg[642]) );
  DFF \creg_reg[643]  ( .D(o[643]), .CLK(clk), .RST(rst), .I(g_init[643]), .Q(
        creg[643]) );
  DFF \creg_reg[644]  ( .D(o[644]), .CLK(clk), .RST(rst), .I(g_init[644]), .Q(
        creg[644]) );
  DFF \creg_reg[645]  ( .D(o[645]), .CLK(clk), .RST(rst), .I(g_init[645]), .Q(
        creg[645]) );
  DFF \creg_reg[646]  ( .D(o[646]), .CLK(clk), .RST(rst), .I(g_init[646]), .Q(
        creg[646]) );
  DFF \creg_reg[647]  ( .D(o[647]), .CLK(clk), .RST(rst), .I(g_init[647]), .Q(
        creg[647]) );
  DFF \creg_reg[648]  ( .D(o[648]), .CLK(clk), .RST(rst), .I(g_init[648]), .Q(
        creg[648]) );
  DFF \creg_reg[649]  ( .D(o[649]), .CLK(clk), .RST(rst), .I(g_init[649]), .Q(
        creg[649]) );
  DFF \creg_reg[650]  ( .D(o[650]), .CLK(clk), .RST(rst), .I(g_init[650]), .Q(
        creg[650]) );
  DFF \creg_reg[651]  ( .D(o[651]), .CLK(clk), .RST(rst), .I(g_init[651]), .Q(
        creg[651]) );
  DFF \creg_reg[652]  ( .D(o[652]), .CLK(clk), .RST(rst), .I(g_init[652]), .Q(
        creg[652]) );
  DFF \creg_reg[653]  ( .D(o[653]), .CLK(clk), .RST(rst), .I(g_init[653]), .Q(
        creg[653]) );
  DFF \creg_reg[654]  ( .D(o[654]), .CLK(clk), .RST(rst), .I(g_init[654]), .Q(
        creg[654]) );
  DFF \creg_reg[655]  ( .D(o[655]), .CLK(clk), .RST(rst), .I(g_init[655]), .Q(
        creg[655]) );
  DFF \creg_reg[656]  ( .D(o[656]), .CLK(clk), .RST(rst), .I(g_init[656]), .Q(
        creg[656]) );
  DFF \creg_reg[657]  ( .D(o[657]), .CLK(clk), .RST(rst), .I(g_init[657]), .Q(
        creg[657]) );
  DFF \creg_reg[658]  ( .D(o[658]), .CLK(clk), .RST(rst), .I(g_init[658]), .Q(
        creg[658]) );
  DFF \creg_reg[659]  ( .D(o[659]), .CLK(clk), .RST(rst), .I(g_init[659]), .Q(
        creg[659]) );
  DFF \creg_reg[660]  ( .D(o[660]), .CLK(clk), .RST(rst), .I(g_init[660]), .Q(
        creg[660]) );
  DFF \creg_reg[661]  ( .D(o[661]), .CLK(clk), .RST(rst), .I(g_init[661]), .Q(
        creg[661]) );
  DFF \creg_reg[662]  ( .D(o[662]), .CLK(clk), .RST(rst), .I(g_init[662]), .Q(
        creg[662]) );
  DFF \creg_reg[663]  ( .D(o[663]), .CLK(clk), .RST(rst), .I(g_init[663]), .Q(
        creg[663]) );
  DFF \creg_reg[664]  ( .D(o[664]), .CLK(clk), .RST(rst), .I(g_init[664]), .Q(
        creg[664]) );
  DFF \creg_reg[665]  ( .D(o[665]), .CLK(clk), .RST(rst), .I(g_init[665]), .Q(
        creg[665]) );
  DFF \creg_reg[666]  ( .D(o[666]), .CLK(clk), .RST(rst), .I(g_init[666]), .Q(
        creg[666]) );
  DFF \creg_reg[667]  ( .D(o[667]), .CLK(clk), .RST(rst), .I(g_init[667]), .Q(
        creg[667]) );
  DFF \creg_reg[668]  ( .D(o[668]), .CLK(clk), .RST(rst), .I(g_init[668]), .Q(
        creg[668]) );
  DFF \creg_reg[669]  ( .D(o[669]), .CLK(clk), .RST(rst), .I(g_init[669]), .Q(
        creg[669]) );
  DFF \creg_reg[670]  ( .D(o[670]), .CLK(clk), .RST(rst), .I(g_init[670]), .Q(
        creg[670]) );
  DFF \creg_reg[671]  ( .D(o[671]), .CLK(clk), .RST(rst), .I(g_init[671]), .Q(
        creg[671]) );
  DFF \creg_reg[672]  ( .D(o[672]), .CLK(clk), .RST(rst), .I(g_init[672]), .Q(
        creg[672]) );
  DFF \creg_reg[673]  ( .D(o[673]), .CLK(clk), .RST(rst), .I(g_init[673]), .Q(
        creg[673]) );
  DFF \creg_reg[674]  ( .D(o[674]), .CLK(clk), .RST(rst), .I(g_init[674]), .Q(
        creg[674]) );
  DFF \creg_reg[675]  ( .D(o[675]), .CLK(clk), .RST(rst), .I(g_init[675]), .Q(
        creg[675]) );
  DFF \creg_reg[676]  ( .D(o[676]), .CLK(clk), .RST(rst), .I(g_init[676]), .Q(
        creg[676]) );
  DFF \creg_reg[677]  ( .D(o[677]), .CLK(clk), .RST(rst), .I(g_init[677]), .Q(
        creg[677]) );
  DFF \creg_reg[678]  ( .D(o[678]), .CLK(clk), .RST(rst), .I(g_init[678]), .Q(
        creg[678]) );
  DFF \creg_reg[679]  ( .D(o[679]), .CLK(clk), .RST(rst), .I(g_init[679]), .Q(
        creg[679]) );
  DFF \creg_reg[680]  ( .D(o[680]), .CLK(clk), .RST(rst), .I(g_init[680]), .Q(
        creg[680]) );
  DFF \creg_reg[681]  ( .D(o[681]), .CLK(clk), .RST(rst), .I(g_init[681]), .Q(
        creg[681]) );
  DFF \creg_reg[682]  ( .D(o[682]), .CLK(clk), .RST(rst), .I(g_init[682]), .Q(
        creg[682]) );
  DFF \creg_reg[683]  ( .D(o[683]), .CLK(clk), .RST(rst), .I(g_init[683]), .Q(
        creg[683]) );
  DFF \creg_reg[684]  ( .D(o[684]), .CLK(clk), .RST(rst), .I(g_init[684]), .Q(
        creg[684]) );
  DFF \creg_reg[685]  ( .D(o[685]), .CLK(clk), .RST(rst), .I(g_init[685]), .Q(
        creg[685]) );
  DFF \creg_reg[686]  ( .D(o[686]), .CLK(clk), .RST(rst), .I(g_init[686]), .Q(
        creg[686]) );
  DFF \creg_reg[687]  ( .D(o[687]), .CLK(clk), .RST(rst), .I(g_init[687]), .Q(
        creg[687]) );
  DFF \creg_reg[688]  ( .D(o[688]), .CLK(clk), .RST(rst), .I(g_init[688]), .Q(
        creg[688]) );
  DFF \creg_reg[689]  ( .D(o[689]), .CLK(clk), .RST(rst), .I(g_init[689]), .Q(
        creg[689]) );
  DFF \creg_reg[690]  ( .D(o[690]), .CLK(clk), .RST(rst), .I(g_init[690]), .Q(
        creg[690]) );
  DFF \creg_reg[691]  ( .D(o[691]), .CLK(clk), .RST(rst), .I(g_init[691]), .Q(
        creg[691]) );
  DFF \creg_reg[692]  ( .D(o[692]), .CLK(clk), .RST(rst), .I(g_init[692]), .Q(
        creg[692]) );
  DFF \creg_reg[693]  ( .D(o[693]), .CLK(clk), .RST(rst), .I(g_init[693]), .Q(
        creg[693]) );
  DFF \creg_reg[694]  ( .D(o[694]), .CLK(clk), .RST(rst), .I(g_init[694]), .Q(
        creg[694]) );
  DFF \creg_reg[695]  ( .D(o[695]), .CLK(clk), .RST(rst), .I(g_init[695]), .Q(
        creg[695]) );
  DFF \creg_reg[696]  ( .D(o[696]), .CLK(clk), .RST(rst), .I(g_init[696]), .Q(
        creg[696]) );
  DFF \creg_reg[697]  ( .D(o[697]), .CLK(clk), .RST(rst), .I(g_init[697]), .Q(
        creg[697]) );
  DFF \creg_reg[698]  ( .D(o[698]), .CLK(clk), .RST(rst), .I(g_init[698]), .Q(
        creg[698]) );
  DFF \creg_reg[699]  ( .D(o[699]), .CLK(clk), .RST(rst), .I(g_init[699]), .Q(
        creg[699]) );
  DFF \creg_reg[700]  ( .D(o[700]), .CLK(clk), .RST(rst), .I(g_init[700]), .Q(
        creg[700]) );
  DFF \creg_reg[701]  ( .D(o[701]), .CLK(clk), .RST(rst), .I(g_init[701]), .Q(
        creg[701]) );
  DFF \creg_reg[702]  ( .D(o[702]), .CLK(clk), .RST(rst), .I(g_init[702]), .Q(
        creg[702]) );
  DFF \creg_reg[703]  ( .D(o[703]), .CLK(clk), .RST(rst), .I(g_init[703]), .Q(
        creg[703]) );
  DFF \creg_reg[704]  ( .D(o[704]), .CLK(clk), .RST(rst), .I(g_init[704]), .Q(
        creg[704]) );
  DFF \creg_reg[705]  ( .D(o[705]), .CLK(clk), .RST(rst), .I(g_init[705]), .Q(
        creg[705]) );
  DFF \creg_reg[706]  ( .D(o[706]), .CLK(clk), .RST(rst), .I(g_init[706]), .Q(
        creg[706]) );
  DFF \creg_reg[707]  ( .D(o[707]), .CLK(clk), .RST(rst), .I(g_init[707]), .Q(
        creg[707]) );
  DFF \creg_reg[708]  ( .D(o[708]), .CLK(clk), .RST(rst), .I(g_init[708]), .Q(
        creg[708]) );
  DFF \creg_reg[709]  ( .D(o[709]), .CLK(clk), .RST(rst), .I(g_init[709]), .Q(
        creg[709]) );
  DFF \creg_reg[710]  ( .D(o[710]), .CLK(clk), .RST(rst), .I(g_init[710]), .Q(
        creg[710]) );
  DFF \creg_reg[711]  ( .D(o[711]), .CLK(clk), .RST(rst), .I(g_init[711]), .Q(
        creg[711]) );
  DFF \creg_reg[712]  ( .D(o[712]), .CLK(clk), .RST(rst), .I(g_init[712]), .Q(
        creg[712]) );
  DFF \creg_reg[713]  ( .D(o[713]), .CLK(clk), .RST(rst), .I(g_init[713]), .Q(
        creg[713]) );
  DFF \creg_reg[714]  ( .D(o[714]), .CLK(clk), .RST(rst), .I(g_init[714]), .Q(
        creg[714]) );
  DFF \creg_reg[715]  ( .D(o[715]), .CLK(clk), .RST(rst), .I(g_init[715]), .Q(
        creg[715]) );
  DFF \creg_reg[716]  ( .D(o[716]), .CLK(clk), .RST(rst), .I(g_init[716]), .Q(
        creg[716]) );
  DFF \creg_reg[717]  ( .D(o[717]), .CLK(clk), .RST(rst), .I(g_init[717]), .Q(
        creg[717]) );
  DFF \creg_reg[718]  ( .D(o[718]), .CLK(clk), .RST(rst), .I(g_init[718]), .Q(
        creg[718]) );
  DFF \creg_reg[719]  ( .D(o[719]), .CLK(clk), .RST(rst), .I(g_init[719]), .Q(
        creg[719]) );
  DFF \creg_reg[720]  ( .D(o[720]), .CLK(clk), .RST(rst), .I(g_init[720]), .Q(
        creg[720]) );
  DFF \creg_reg[721]  ( .D(o[721]), .CLK(clk), .RST(rst), .I(g_init[721]), .Q(
        creg[721]) );
  DFF \creg_reg[722]  ( .D(o[722]), .CLK(clk), .RST(rst), .I(g_init[722]), .Q(
        creg[722]) );
  DFF \creg_reg[723]  ( .D(o[723]), .CLK(clk), .RST(rst), .I(g_init[723]), .Q(
        creg[723]) );
  DFF \creg_reg[724]  ( .D(o[724]), .CLK(clk), .RST(rst), .I(g_init[724]), .Q(
        creg[724]) );
  DFF \creg_reg[725]  ( .D(o[725]), .CLK(clk), .RST(rst), .I(g_init[725]), .Q(
        creg[725]) );
  DFF \creg_reg[726]  ( .D(o[726]), .CLK(clk), .RST(rst), .I(g_init[726]), .Q(
        creg[726]) );
  DFF \creg_reg[727]  ( .D(o[727]), .CLK(clk), .RST(rst), .I(g_init[727]), .Q(
        creg[727]) );
  DFF \creg_reg[728]  ( .D(o[728]), .CLK(clk), .RST(rst), .I(g_init[728]), .Q(
        creg[728]) );
  DFF \creg_reg[729]  ( .D(o[729]), .CLK(clk), .RST(rst), .I(g_init[729]), .Q(
        creg[729]) );
  DFF \creg_reg[730]  ( .D(o[730]), .CLK(clk), .RST(rst), .I(g_init[730]), .Q(
        creg[730]) );
  DFF \creg_reg[731]  ( .D(o[731]), .CLK(clk), .RST(rst), .I(g_init[731]), .Q(
        creg[731]) );
  DFF \creg_reg[732]  ( .D(o[732]), .CLK(clk), .RST(rst), .I(g_init[732]), .Q(
        creg[732]) );
  DFF \creg_reg[733]  ( .D(o[733]), .CLK(clk), .RST(rst), .I(g_init[733]), .Q(
        creg[733]) );
  DFF \creg_reg[734]  ( .D(o[734]), .CLK(clk), .RST(rst), .I(g_init[734]), .Q(
        creg[734]) );
  DFF \creg_reg[735]  ( .D(o[735]), .CLK(clk), .RST(rst), .I(g_init[735]), .Q(
        creg[735]) );
  DFF \creg_reg[736]  ( .D(o[736]), .CLK(clk), .RST(rst), .I(g_init[736]), .Q(
        creg[736]) );
  DFF \creg_reg[737]  ( .D(o[737]), .CLK(clk), .RST(rst), .I(g_init[737]), .Q(
        creg[737]) );
  DFF \creg_reg[738]  ( .D(o[738]), .CLK(clk), .RST(rst), .I(g_init[738]), .Q(
        creg[738]) );
  DFF \creg_reg[739]  ( .D(o[739]), .CLK(clk), .RST(rst), .I(g_init[739]), .Q(
        creg[739]) );
  DFF \creg_reg[740]  ( .D(o[740]), .CLK(clk), .RST(rst), .I(g_init[740]), .Q(
        creg[740]) );
  DFF \creg_reg[741]  ( .D(o[741]), .CLK(clk), .RST(rst), .I(g_init[741]), .Q(
        creg[741]) );
  DFF \creg_reg[742]  ( .D(o[742]), .CLK(clk), .RST(rst), .I(g_init[742]), .Q(
        creg[742]) );
  DFF \creg_reg[743]  ( .D(o[743]), .CLK(clk), .RST(rst), .I(g_init[743]), .Q(
        creg[743]) );
  DFF \creg_reg[744]  ( .D(o[744]), .CLK(clk), .RST(rst), .I(g_init[744]), .Q(
        creg[744]) );
  DFF \creg_reg[745]  ( .D(o[745]), .CLK(clk), .RST(rst), .I(g_init[745]), .Q(
        creg[745]) );
  DFF \creg_reg[746]  ( .D(o[746]), .CLK(clk), .RST(rst), .I(g_init[746]), .Q(
        creg[746]) );
  DFF \creg_reg[747]  ( .D(o[747]), .CLK(clk), .RST(rst), .I(g_init[747]), .Q(
        creg[747]) );
  DFF \creg_reg[748]  ( .D(o[748]), .CLK(clk), .RST(rst), .I(g_init[748]), .Q(
        creg[748]) );
  DFF \creg_reg[749]  ( .D(o[749]), .CLK(clk), .RST(rst), .I(g_init[749]), .Q(
        creg[749]) );
  DFF \creg_reg[750]  ( .D(o[750]), .CLK(clk), .RST(rst), .I(g_init[750]), .Q(
        creg[750]) );
  DFF \creg_reg[751]  ( .D(o[751]), .CLK(clk), .RST(rst), .I(g_init[751]), .Q(
        creg[751]) );
  DFF \creg_reg[752]  ( .D(o[752]), .CLK(clk), .RST(rst), .I(g_init[752]), .Q(
        creg[752]) );
  DFF \creg_reg[753]  ( .D(o[753]), .CLK(clk), .RST(rst), .I(g_init[753]), .Q(
        creg[753]) );
  DFF \creg_reg[754]  ( .D(o[754]), .CLK(clk), .RST(rst), .I(g_init[754]), .Q(
        creg[754]) );
  DFF \creg_reg[755]  ( .D(o[755]), .CLK(clk), .RST(rst), .I(g_init[755]), .Q(
        creg[755]) );
  DFF \creg_reg[756]  ( .D(o[756]), .CLK(clk), .RST(rst), .I(g_init[756]), .Q(
        creg[756]) );
  DFF \creg_reg[757]  ( .D(o[757]), .CLK(clk), .RST(rst), .I(g_init[757]), .Q(
        creg[757]) );
  DFF \creg_reg[758]  ( .D(o[758]), .CLK(clk), .RST(rst), .I(g_init[758]), .Q(
        creg[758]) );
  DFF \creg_reg[759]  ( .D(o[759]), .CLK(clk), .RST(rst), .I(g_init[759]), .Q(
        creg[759]) );
  DFF \creg_reg[760]  ( .D(o[760]), .CLK(clk), .RST(rst), .I(g_init[760]), .Q(
        creg[760]) );
  DFF \creg_reg[761]  ( .D(o[761]), .CLK(clk), .RST(rst), .I(g_init[761]), .Q(
        creg[761]) );
  DFF \creg_reg[762]  ( .D(o[762]), .CLK(clk), .RST(rst), .I(g_init[762]), .Q(
        creg[762]) );
  DFF \creg_reg[763]  ( .D(o[763]), .CLK(clk), .RST(rst), .I(g_init[763]), .Q(
        creg[763]) );
  DFF \creg_reg[764]  ( .D(o[764]), .CLK(clk), .RST(rst), .I(g_init[764]), .Q(
        creg[764]) );
  DFF \creg_reg[765]  ( .D(o[765]), .CLK(clk), .RST(rst), .I(g_init[765]), .Q(
        creg[765]) );
  DFF \creg_reg[766]  ( .D(o[766]), .CLK(clk), .RST(rst), .I(g_init[766]), .Q(
        creg[766]) );
  DFF \creg_reg[767]  ( .D(o[767]), .CLK(clk), .RST(rst), .I(g_init[767]), .Q(
        creg[767]) );
  DFF \creg_reg[768]  ( .D(o[768]), .CLK(clk), .RST(rst), .I(g_init[768]), .Q(
        creg[768]) );
  DFF \creg_reg[769]  ( .D(o[769]), .CLK(clk), .RST(rst), .I(g_init[769]), .Q(
        creg[769]) );
  DFF \creg_reg[770]  ( .D(o[770]), .CLK(clk), .RST(rst), .I(g_init[770]), .Q(
        creg[770]) );
  DFF \creg_reg[771]  ( .D(o[771]), .CLK(clk), .RST(rst), .I(g_init[771]), .Q(
        creg[771]) );
  DFF \creg_reg[772]  ( .D(o[772]), .CLK(clk), .RST(rst), .I(g_init[772]), .Q(
        creg[772]) );
  DFF \creg_reg[773]  ( .D(o[773]), .CLK(clk), .RST(rst), .I(g_init[773]), .Q(
        creg[773]) );
  DFF \creg_reg[774]  ( .D(o[774]), .CLK(clk), .RST(rst), .I(g_init[774]), .Q(
        creg[774]) );
  DFF \creg_reg[775]  ( .D(o[775]), .CLK(clk), .RST(rst), .I(g_init[775]), .Q(
        creg[775]) );
  DFF \creg_reg[776]  ( .D(o[776]), .CLK(clk), .RST(rst), .I(g_init[776]), .Q(
        creg[776]) );
  DFF \creg_reg[777]  ( .D(o[777]), .CLK(clk), .RST(rst), .I(g_init[777]), .Q(
        creg[777]) );
  DFF \creg_reg[778]  ( .D(o[778]), .CLK(clk), .RST(rst), .I(g_init[778]), .Q(
        creg[778]) );
  DFF \creg_reg[779]  ( .D(o[779]), .CLK(clk), .RST(rst), .I(g_init[779]), .Q(
        creg[779]) );
  DFF \creg_reg[780]  ( .D(o[780]), .CLK(clk), .RST(rst), .I(g_init[780]), .Q(
        creg[780]) );
  DFF \creg_reg[781]  ( .D(o[781]), .CLK(clk), .RST(rst), .I(g_init[781]), .Q(
        creg[781]) );
  DFF \creg_reg[782]  ( .D(o[782]), .CLK(clk), .RST(rst), .I(g_init[782]), .Q(
        creg[782]) );
  DFF \creg_reg[783]  ( .D(o[783]), .CLK(clk), .RST(rst), .I(g_init[783]), .Q(
        creg[783]) );
  DFF \creg_reg[784]  ( .D(o[784]), .CLK(clk), .RST(rst), .I(g_init[784]), .Q(
        creg[784]) );
  DFF \creg_reg[785]  ( .D(o[785]), .CLK(clk), .RST(rst), .I(g_init[785]), .Q(
        creg[785]) );
  DFF \creg_reg[786]  ( .D(o[786]), .CLK(clk), .RST(rst), .I(g_init[786]), .Q(
        creg[786]) );
  DFF \creg_reg[787]  ( .D(o[787]), .CLK(clk), .RST(rst), .I(g_init[787]), .Q(
        creg[787]) );
  DFF \creg_reg[788]  ( .D(o[788]), .CLK(clk), .RST(rst), .I(g_init[788]), .Q(
        creg[788]) );
  DFF \creg_reg[789]  ( .D(o[789]), .CLK(clk), .RST(rst), .I(g_init[789]), .Q(
        creg[789]) );
  DFF \creg_reg[790]  ( .D(o[790]), .CLK(clk), .RST(rst), .I(g_init[790]), .Q(
        creg[790]) );
  DFF \creg_reg[791]  ( .D(o[791]), .CLK(clk), .RST(rst), .I(g_init[791]), .Q(
        creg[791]) );
  DFF \creg_reg[792]  ( .D(o[792]), .CLK(clk), .RST(rst), .I(g_init[792]), .Q(
        creg[792]) );
  DFF \creg_reg[793]  ( .D(o[793]), .CLK(clk), .RST(rst), .I(g_init[793]), .Q(
        creg[793]) );
  DFF \creg_reg[794]  ( .D(o[794]), .CLK(clk), .RST(rst), .I(g_init[794]), .Q(
        creg[794]) );
  DFF \creg_reg[795]  ( .D(o[795]), .CLK(clk), .RST(rst), .I(g_init[795]), .Q(
        creg[795]) );
  DFF \creg_reg[796]  ( .D(o[796]), .CLK(clk), .RST(rst), .I(g_init[796]), .Q(
        creg[796]) );
  DFF \creg_reg[797]  ( .D(o[797]), .CLK(clk), .RST(rst), .I(g_init[797]), .Q(
        creg[797]) );
  DFF \creg_reg[798]  ( .D(o[798]), .CLK(clk), .RST(rst), .I(g_init[798]), .Q(
        creg[798]) );
  DFF \creg_reg[799]  ( .D(o[799]), .CLK(clk), .RST(rst), .I(g_init[799]), .Q(
        creg[799]) );
  DFF \creg_reg[800]  ( .D(o[800]), .CLK(clk), .RST(rst), .I(g_init[800]), .Q(
        creg[800]) );
  DFF \creg_reg[801]  ( .D(o[801]), .CLK(clk), .RST(rst), .I(g_init[801]), .Q(
        creg[801]) );
  DFF \creg_reg[802]  ( .D(o[802]), .CLK(clk), .RST(rst), .I(g_init[802]), .Q(
        creg[802]) );
  DFF \creg_reg[803]  ( .D(o[803]), .CLK(clk), .RST(rst), .I(g_init[803]), .Q(
        creg[803]) );
  DFF \creg_reg[804]  ( .D(o[804]), .CLK(clk), .RST(rst), .I(g_init[804]), .Q(
        creg[804]) );
  DFF \creg_reg[805]  ( .D(o[805]), .CLK(clk), .RST(rst), .I(g_init[805]), .Q(
        creg[805]) );
  DFF \creg_reg[806]  ( .D(o[806]), .CLK(clk), .RST(rst), .I(g_init[806]), .Q(
        creg[806]) );
  DFF \creg_reg[807]  ( .D(o[807]), .CLK(clk), .RST(rst), .I(g_init[807]), .Q(
        creg[807]) );
  DFF \creg_reg[808]  ( .D(o[808]), .CLK(clk), .RST(rst), .I(g_init[808]), .Q(
        creg[808]) );
  DFF \creg_reg[809]  ( .D(o[809]), .CLK(clk), .RST(rst), .I(g_init[809]), .Q(
        creg[809]) );
  DFF \creg_reg[810]  ( .D(o[810]), .CLK(clk), .RST(rst), .I(g_init[810]), .Q(
        creg[810]) );
  DFF \creg_reg[811]  ( .D(o[811]), .CLK(clk), .RST(rst), .I(g_init[811]), .Q(
        creg[811]) );
  DFF \creg_reg[812]  ( .D(o[812]), .CLK(clk), .RST(rst), .I(g_init[812]), .Q(
        creg[812]) );
  DFF \creg_reg[813]  ( .D(o[813]), .CLK(clk), .RST(rst), .I(g_init[813]), .Q(
        creg[813]) );
  DFF \creg_reg[814]  ( .D(o[814]), .CLK(clk), .RST(rst), .I(g_init[814]), .Q(
        creg[814]) );
  DFF \creg_reg[815]  ( .D(o[815]), .CLK(clk), .RST(rst), .I(g_init[815]), .Q(
        creg[815]) );
  DFF \creg_reg[816]  ( .D(o[816]), .CLK(clk), .RST(rst), .I(g_init[816]), .Q(
        creg[816]) );
  DFF \creg_reg[817]  ( .D(o[817]), .CLK(clk), .RST(rst), .I(g_init[817]), .Q(
        creg[817]) );
  DFF \creg_reg[818]  ( .D(o[818]), .CLK(clk), .RST(rst), .I(g_init[818]), .Q(
        creg[818]) );
  DFF \creg_reg[819]  ( .D(o[819]), .CLK(clk), .RST(rst), .I(g_init[819]), .Q(
        creg[819]) );
  DFF \creg_reg[820]  ( .D(o[820]), .CLK(clk), .RST(rst), .I(g_init[820]), .Q(
        creg[820]) );
  DFF \creg_reg[821]  ( .D(o[821]), .CLK(clk), .RST(rst), .I(g_init[821]), .Q(
        creg[821]) );
  DFF \creg_reg[822]  ( .D(o[822]), .CLK(clk), .RST(rst), .I(g_init[822]), .Q(
        creg[822]) );
  DFF \creg_reg[823]  ( .D(o[823]), .CLK(clk), .RST(rst), .I(g_init[823]), .Q(
        creg[823]) );
  DFF \creg_reg[824]  ( .D(o[824]), .CLK(clk), .RST(rst), .I(g_init[824]), .Q(
        creg[824]) );
  DFF \creg_reg[825]  ( .D(o[825]), .CLK(clk), .RST(rst), .I(g_init[825]), .Q(
        creg[825]) );
  DFF \creg_reg[826]  ( .D(o[826]), .CLK(clk), .RST(rst), .I(g_init[826]), .Q(
        creg[826]) );
  DFF \creg_reg[827]  ( .D(o[827]), .CLK(clk), .RST(rst), .I(g_init[827]), .Q(
        creg[827]) );
  DFF \creg_reg[828]  ( .D(o[828]), .CLK(clk), .RST(rst), .I(g_init[828]), .Q(
        creg[828]) );
  DFF \creg_reg[829]  ( .D(o[829]), .CLK(clk), .RST(rst), .I(g_init[829]), .Q(
        creg[829]) );
  DFF \creg_reg[830]  ( .D(o[830]), .CLK(clk), .RST(rst), .I(g_init[830]), .Q(
        creg[830]) );
  DFF \creg_reg[831]  ( .D(o[831]), .CLK(clk), .RST(rst), .I(g_init[831]), .Q(
        creg[831]) );
  DFF \creg_reg[832]  ( .D(o[832]), .CLK(clk), .RST(rst), .I(g_init[832]), .Q(
        creg[832]) );
  DFF \creg_reg[833]  ( .D(o[833]), .CLK(clk), .RST(rst), .I(g_init[833]), .Q(
        creg[833]) );
  DFF \creg_reg[834]  ( .D(o[834]), .CLK(clk), .RST(rst), .I(g_init[834]), .Q(
        creg[834]) );
  DFF \creg_reg[835]  ( .D(o[835]), .CLK(clk), .RST(rst), .I(g_init[835]), .Q(
        creg[835]) );
  DFF \creg_reg[836]  ( .D(o[836]), .CLK(clk), .RST(rst), .I(g_init[836]), .Q(
        creg[836]) );
  DFF \creg_reg[837]  ( .D(o[837]), .CLK(clk), .RST(rst), .I(g_init[837]), .Q(
        creg[837]) );
  DFF \creg_reg[838]  ( .D(o[838]), .CLK(clk), .RST(rst), .I(g_init[838]), .Q(
        creg[838]) );
  DFF \creg_reg[839]  ( .D(o[839]), .CLK(clk), .RST(rst), .I(g_init[839]), .Q(
        creg[839]) );
  DFF \creg_reg[840]  ( .D(o[840]), .CLK(clk), .RST(rst), .I(g_init[840]), .Q(
        creg[840]) );
  DFF \creg_reg[841]  ( .D(o[841]), .CLK(clk), .RST(rst), .I(g_init[841]), .Q(
        creg[841]) );
  DFF \creg_reg[842]  ( .D(o[842]), .CLK(clk), .RST(rst), .I(g_init[842]), .Q(
        creg[842]) );
  DFF \creg_reg[843]  ( .D(o[843]), .CLK(clk), .RST(rst), .I(g_init[843]), .Q(
        creg[843]) );
  DFF \creg_reg[844]  ( .D(o[844]), .CLK(clk), .RST(rst), .I(g_init[844]), .Q(
        creg[844]) );
  DFF \creg_reg[845]  ( .D(o[845]), .CLK(clk), .RST(rst), .I(g_init[845]), .Q(
        creg[845]) );
  DFF \creg_reg[846]  ( .D(o[846]), .CLK(clk), .RST(rst), .I(g_init[846]), .Q(
        creg[846]) );
  DFF \creg_reg[847]  ( .D(o[847]), .CLK(clk), .RST(rst), .I(g_init[847]), .Q(
        creg[847]) );
  DFF \creg_reg[848]  ( .D(o[848]), .CLK(clk), .RST(rst), .I(g_init[848]), .Q(
        creg[848]) );
  DFF \creg_reg[849]  ( .D(o[849]), .CLK(clk), .RST(rst), .I(g_init[849]), .Q(
        creg[849]) );
  DFF \creg_reg[850]  ( .D(o[850]), .CLK(clk), .RST(rst), .I(g_init[850]), .Q(
        creg[850]) );
  DFF \creg_reg[851]  ( .D(o[851]), .CLK(clk), .RST(rst), .I(g_init[851]), .Q(
        creg[851]) );
  DFF \creg_reg[852]  ( .D(o[852]), .CLK(clk), .RST(rst), .I(g_init[852]), .Q(
        creg[852]) );
  DFF \creg_reg[853]  ( .D(o[853]), .CLK(clk), .RST(rst), .I(g_init[853]), .Q(
        creg[853]) );
  DFF \creg_reg[854]  ( .D(o[854]), .CLK(clk), .RST(rst), .I(g_init[854]), .Q(
        creg[854]) );
  DFF \creg_reg[855]  ( .D(o[855]), .CLK(clk), .RST(rst), .I(g_init[855]), .Q(
        creg[855]) );
  DFF \creg_reg[856]  ( .D(o[856]), .CLK(clk), .RST(rst), .I(g_init[856]), .Q(
        creg[856]) );
  DFF \creg_reg[857]  ( .D(o[857]), .CLK(clk), .RST(rst), .I(g_init[857]), .Q(
        creg[857]) );
  DFF \creg_reg[858]  ( .D(o[858]), .CLK(clk), .RST(rst), .I(g_init[858]), .Q(
        creg[858]) );
  DFF \creg_reg[859]  ( .D(o[859]), .CLK(clk), .RST(rst), .I(g_init[859]), .Q(
        creg[859]) );
  DFF \creg_reg[860]  ( .D(o[860]), .CLK(clk), .RST(rst), .I(g_init[860]), .Q(
        creg[860]) );
  DFF \creg_reg[861]  ( .D(o[861]), .CLK(clk), .RST(rst), .I(g_init[861]), .Q(
        creg[861]) );
  DFF \creg_reg[862]  ( .D(o[862]), .CLK(clk), .RST(rst), .I(g_init[862]), .Q(
        creg[862]) );
  DFF \creg_reg[863]  ( .D(o[863]), .CLK(clk), .RST(rst), .I(g_init[863]), .Q(
        creg[863]) );
  DFF \creg_reg[864]  ( .D(o[864]), .CLK(clk), .RST(rst), .I(g_init[864]), .Q(
        creg[864]) );
  DFF \creg_reg[865]  ( .D(o[865]), .CLK(clk), .RST(rst), .I(g_init[865]), .Q(
        creg[865]) );
  DFF \creg_reg[866]  ( .D(o[866]), .CLK(clk), .RST(rst), .I(g_init[866]), .Q(
        creg[866]) );
  DFF \creg_reg[867]  ( .D(o[867]), .CLK(clk), .RST(rst), .I(g_init[867]), .Q(
        creg[867]) );
  DFF \creg_reg[868]  ( .D(o[868]), .CLK(clk), .RST(rst), .I(g_init[868]), .Q(
        creg[868]) );
  DFF \creg_reg[869]  ( .D(o[869]), .CLK(clk), .RST(rst), .I(g_init[869]), .Q(
        creg[869]) );
  DFF \creg_reg[870]  ( .D(o[870]), .CLK(clk), .RST(rst), .I(g_init[870]), .Q(
        creg[870]) );
  DFF \creg_reg[871]  ( .D(o[871]), .CLK(clk), .RST(rst), .I(g_init[871]), .Q(
        creg[871]) );
  DFF \creg_reg[872]  ( .D(o[872]), .CLK(clk), .RST(rst), .I(g_init[872]), .Q(
        creg[872]) );
  DFF \creg_reg[873]  ( .D(o[873]), .CLK(clk), .RST(rst), .I(g_init[873]), .Q(
        creg[873]) );
  DFF \creg_reg[874]  ( .D(o[874]), .CLK(clk), .RST(rst), .I(g_init[874]), .Q(
        creg[874]) );
  DFF \creg_reg[875]  ( .D(o[875]), .CLK(clk), .RST(rst), .I(g_init[875]), .Q(
        creg[875]) );
  DFF \creg_reg[876]  ( .D(o[876]), .CLK(clk), .RST(rst), .I(g_init[876]), .Q(
        creg[876]) );
  DFF \creg_reg[877]  ( .D(o[877]), .CLK(clk), .RST(rst), .I(g_init[877]), .Q(
        creg[877]) );
  DFF \creg_reg[878]  ( .D(o[878]), .CLK(clk), .RST(rst), .I(g_init[878]), .Q(
        creg[878]) );
  DFF \creg_reg[879]  ( .D(o[879]), .CLK(clk), .RST(rst), .I(g_init[879]), .Q(
        creg[879]) );
  DFF \creg_reg[880]  ( .D(o[880]), .CLK(clk), .RST(rst), .I(g_init[880]), .Q(
        creg[880]) );
  DFF \creg_reg[881]  ( .D(o[881]), .CLK(clk), .RST(rst), .I(g_init[881]), .Q(
        creg[881]) );
  DFF \creg_reg[882]  ( .D(o[882]), .CLK(clk), .RST(rst), .I(g_init[882]), .Q(
        creg[882]) );
  DFF \creg_reg[883]  ( .D(o[883]), .CLK(clk), .RST(rst), .I(g_init[883]), .Q(
        creg[883]) );
  DFF \creg_reg[884]  ( .D(o[884]), .CLK(clk), .RST(rst), .I(g_init[884]), .Q(
        creg[884]) );
  DFF \creg_reg[885]  ( .D(o[885]), .CLK(clk), .RST(rst), .I(g_init[885]), .Q(
        creg[885]) );
  DFF \creg_reg[886]  ( .D(o[886]), .CLK(clk), .RST(rst), .I(g_init[886]), .Q(
        creg[886]) );
  DFF \creg_reg[887]  ( .D(o[887]), .CLK(clk), .RST(rst), .I(g_init[887]), .Q(
        creg[887]) );
  DFF \creg_reg[888]  ( .D(o[888]), .CLK(clk), .RST(rst), .I(g_init[888]), .Q(
        creg[888]) );
  DFF \creg_reg[889]  ( .D(o[889]), .CLK(clk), .RST(rst), .I(g_init[889]), .Q(
        creg[889]) );
  DFF \creg_reg[890]  ( .D(o[890]), .CLK(clk), .RST(rst), .I(g_init[890]), .Q(
        creg[890]) );
  DFF \creg_reg[891]  ( .D(o[891]), .CLK(clk), .RST(rst), .I(g_init[891]), .Q(
        creg[891]) );
  DFF \creg_reg[892]  ( .D(o[892]), .CLK(clk), .RST(rst), .I(g_init[892]), .Q(
        creg[892]) );
  DFF \creg_reg[893]  ( .D(o[893]), .CLK(clk), .RST(rst), .I(g_init[893]), .Q(
        creg[893]) );
  DFF \creg_reg[894]  ( .D(o[894]), .CLK(clk), .RST(rst), .I(g_init[894]), .Q(
        creg[894]) );
  DFF \creg_reg[895]  ( .D(o[895]), .CLK(clk), .RST(rst), .I(g_init[895]), .Q(
        creg[895]) );
  DFF \creg_reg[896]  ( .D(o[896]), .CLK(clk), .RST(rst), .I(g_init[896]), .Q(
        creg[896]) );
  DFF \creg_reg[897]  ( .D(o[897]), .CLK(clk), .RST(rst), .I(g_init[897]), .Q(
        creg[897]) );
  DFF \creg_reg[898]  ( .D(o[898]), .CLK(clk), .RST(rst), .I(g_init[898]), .Q(
        creg[898]) );
  DFF \creg_reg[899]  ( .D(o[899]), .CLK(clk), .RST(rst), .I(g_init[899]), .Q(
        creg[899]) );
  DFF \creg_reg[900]  ( .D(o[900]), .CLK(clk), .RST(rst), .I(g_init[900]), .Q(
        creg[900]) );
  DFF \creg_reg[901]  ( .D(o[901]), .CLK(clk), .RST(rst), .I(g_init[901]), .Q(
        creg[901]) );
  DFF \creg_reg[902]  ( .D(o[902]), .CLK(clk), .RST(rst), .I(g_init[902]), .Q(
        creg[902]) );
  DFF \creg_reg[903]  ( .D(o[903]), .CLK(clk), .RST(rst), .I(g_init[903]), .Q(
        creg[903]) );
  DFF \creg_reg[904]  ( .D(o[904]), .CLK(clk), .RST(rst), .I(g_init[904]), .Q(
        creg[904]) );
  DFF \creg_reg[905]  ( .D(o[905]), .CLK(clk), .RST(rst), .I(g_init[905]), .Q(
        creg[905]) );
  DFF \creg_reg[906]  ( .D(o[906]), .CLK(clk), .RST(rst), .I(g_init[906]), .Q(
        creg[906]) );
  DFF \creg_reg[907]  ( .D(o[907]), .CLK(clk), .RST(rst), .I(g_init[907]), .Q(
        creg[907]) );
  DFF \creg_reg[908]  ( .D(o[908]), .CLK(clk), .RST(rst), .I(g_init[908]), .Q(
        creg[908]) );
  DFF \creg_reg[909]  ( .D(o[909]), .CLK(clk), .RST(rst), .I(g_init[909]), .Q(
        creg[909]) );
  DFF \creg_reg[910]  ( .D(o[910]), .CLK(clk), .RST(rst), .I(g_init[910]), .Q(
        creg[910]) );
  DFF \creg_reg[911]  ( .D(o[911]), .CLK(clk), .RST(rst), .I(g_init[911]), .Q(
        creg[911]) );
  DFF \creg_reg[912]  ( .D(o[912]), .CLK(clk), .RST(rst), .I(g_init[912]), .Q(
        creg[912]) );
  DFF \creg_reg[913]  ( .D(o[913]), .CLK(clk), .RST(rst), .I(g_init[913]), .Q(
        creg[913]) );
  DFF \creg_reg[914]  ( .D(o[914]), .CLK(clk), .RST(rst), .I(g_init[914]), .Q(
        creg[914]) );
  DFF \creg_reg[915]  ( .D(o[915]), .CLK(clk), .RST(rst), .I(g_init[915]), .Q(
        creg[915]) );
  DFF \creg_reg[916]  ( .D(o[916]), .CLK(clk), .RST(rst), .I(g_init[916]), .Q(
        creg[916]) );
  DFF \creg_reg[917]  ( .D(o[917]), .CLK(clk), .RST(rst), .I(g_init[917]), .Q(
        creg[917]) );
  DFF \creg_reg[918]  ( .D(o[918]), .CLK(clk), .RST(rst), .I(g_init[918]), .Q(
        creg[918]) );
  DFF \creg_reg[919]  ( .D(o[919]), .CLK(clk), .RST(rst), .I(g_init[919]), .Q(
        creg[919]) );
  DFF \creg_reg[920]  ( .D(o[920]), .CLK(clk), .RST(rst), .I(g_init[920]), .Q(
        creg[920]) );
  DFF \creg_reg[921]  ( .D(o[921]), .CLK(clk), .RST(rst), .I(g_init[921]), .Q(
        creg[921]) );
  DFF \creg_reg[922]  ( .D(o[922]), .CLK(clk), .RST(rst), .I(g_init[922]), .Q(
        creg[922]) );
  DFF \creg_reg[923]  ( .D(o[923]), .CLK(clk), .RST(rst), .I(g_init[923]), .Q(
        creg[923]) );
  DFF \creg_reg[924]  ( .D(o[924]), .CLK(clk), .RST(rst), .I(g_init[924]), .Q(
        creg[924]) );
  DFF \creg_reg[925]  ( .D(o[925]), .CLK(clk), .RST(rst), .I(g_init[925]), .Q(
        creg[925]) );
  DFF \creg_reg[926]  ( .D(o[926]), .CLK(clk), .RST(rst), .I(g_init[926]), .Q(
        creg[926]) );
  DFF \creg_reg[927]  ( .D(o[927]), .CLK(clk), .RST(rst), .I(g_init[927]), .Q(
        creg[927]) );
  DFF \creg_reg[928]  ( .D(o[928]), .CLK(clk), .RST(rst), .I(g_init[928]), .Q(
        creg[928]) );
  DFF \creg_reg[929]  ( .D(o[929]), .CLK(clk), .RST(rst), .I(g_init[929]), .Q(
        creg[929]) );
  DFF \creg_reg[930]  ( .D(o[930]), .CLK(clk), .RST(rst), .I(g_init[930]), .Q(
        creg[930]) );
  DFF \creg_reg[931]  ( .D(o[931]), .CLK(clk), .RST(rst), .I(g_init[931]), .Q(
        creg[931]) );
  DFF \creg_reg[932]  ( .D(o[932]), .CLK(clk), .RST(rst), .I(g_init[932]), .Q(
        creg[932]) );
  DFF \creg_reg[933]  ( .D(o[933]), .CLK(clk), .RST(rst), .I(g_init[933]), .Q(
        creg[933]) );
  DFF \creg_reg[934]  ( .D(o[934]), .CLK(clk), .RST(rst), .I(g_init[934]), .Q(
        creg[934]) );
  DFF \creg_reg[935]  ( .D(o[935]), .CLK(clk), .RST(rst), .I(g_init[935]), .Q(
        creg[935]) );
  DFF \creg_reg[936]  ( .D(o[936]), .CLK(clk), .RST(rst), .I(g_init[936]), .Q(
        creg[936]) );
  DFF \creg_reg[937]  ( .D(o[937]), .CLK(clk), .RST(rst), .I(g_init[937]), .Q(
        creg[937]) );
  DFF \creg_reg[938]  ( .D(o[938]), .CLK(clk), .RST(rst), .I(g_init[938]), .Q(
        creg[938]) );
  DFF \creg_reg[939]  ( .D(o[939]), .CLK(clk), .RST(rst), .I(g_init[939]), .Q(
        creg[939]) );
  DFF \creg_reg[940]  ( .D(o[940]), .CLK(clk), .RST(rst), .I(g_init[940]), .Q(
        creg[940]) );
  DFF \creg_reg[941]  ( .D(o[941]), .CLK(clk), .RST(rst), .I(g_init[941]), .Q(
        creg[941]) );
  DFF \creg_reg[942]  ( .D(o[942]), .CLK(clk), .RST(rst), .I(g_init[942]), .Q(
        creg[942]) );
  DFF \creg_reg[943]  ( .D(o[943]), .CLK(clk), .RST(rst), .I(g_init[943]), .Q(
        creg[943]) );
  DFF \creg_reg[944]  ( .D(o[944]), .CLK(clk), .RST(rst), .I(g_init[944]), .Q(
        creg[944]) );
  DFF \creg_reg[945]  ( .D(o[945]), .CLK(clk), .RST(rst), .I(g_init[945]), .Q(
        creg[945]) );
  DFF \creg_reg[946]  ( .D(o[946]), .CLK(clk), .RST(rst), .I(g_init[946]), .Q(
        creg[946]) );
  DFF \creg_reg[947]  ( .D(o[947]), .CLK(clk), .RST(rst), .I(g_init[947]), .Q(
        creg[947]) );
  DFF \creg_reg[948]  ( .D(o[948]), .CLK(clk), .RST(rst), .I(g_init[948]), .Q(
        creg[948]) );
  DFF \creg_reg[949]  ( .D(o[949]), .CLK(clk), .RST(rst), .I(g_init[949]), .Q(
        creg[949]) );
  DFF \creg_reg[950]  ( .D(o[950]), .CLK(clk), .RST(rst), .I(g_init[950]), .Q(
        creg[950]) );
  DFF \creg_reg[951]  ( .D(o[951]), .CLK(clk), .RST(rst), .I(g_init[951]), .Q(
        creg[951]) );
  DFF \creg_reg[952]  ( .D(o[952]), .CLK(clk), .RST(rst), .I(g_init[952]), .Q(
        creg[952]) );
  DFF \creg_reg[953]  ( .D(o[953]), .CLK(clk), .RST(rst), .I(g_init[953]), .Q(
        creg[953]) );
  DFF \creg_reg[954]  ( .D(o[954]), .CLK(clk), .RST(rst), .I(g_init[954]), .Q(
        creg[954]) );
  DFF \creg_reg[955]  ( .D(o[955]), .CLK(clk), .RST(rst), .I(g_init[955]), .Q(
        creg[955]) );
  DFF \creg_reg[956]  ( .D(o[956]), .CLK(clk), .RST(rst), .I(g_init[956]), .Q(
        creg[956]) );
  DFF \creg_reg[957]  ( .D(o[957]), .CLK(clk), .RST(rst), .I(g_init[957]), .Q(
        creg[957]) );
  DFF \creg_reg[958]  ( .D(o[958]), .CLK(clk), .RST(rst), .I(g_init[958]), .Q(
        creg[958]) );
  DFF \creg_reg[959]  ( .D(o[959]), .CLK(clk), .RST(rst), .I(g_init[959]), .Q(
        creg[959]) );
  DFF \creg_reg[960]  ( .D(o[960]), .CLK(clk), .RST(rst), .I(g_init[960]), .Q(
        creg[960]) );
  DFF \creg_reg[961]  ( .D(o[961]), .CLK(clk), .RST(rst), .I(g_init[961]), .Q(
        creg[961]) );
  DFF \creg_reg[962]  ( .D(o[962]), .CLK(clk), .RST(rst), .I(g_init[962]), .Q(
        creg[962]) );
  DFF \creg_reg[963]  ( .D(o[963]), .CLK(clk), .RST(rst), .I(g_init[963]), .Q(
        creg[963]) );
  DFF \creg_reg[964]  ( .D(o[964]), .CLK(clk), .RST(rst), .I(g_init[964]), .Q(
        creg[964]) );
  DFF \creg_reg[965]  ( .D(o[965]), .CLK(clk), .RST(rst), .I(g_init[965]), .Q(
        creg[965]) );
  DFF \creg_reg[966]  ( .D(o[966]), .CLK(clk), .RST(rst), .I(g_init[966]), .Q(
        creg[966]) );
  DFF \creg_reg[967]  ( .D(o[967]), .CLK(clk), .RST(rst), .I(g_init[967]), .Q(
        creg[967]) );
  DFF \creg_reg[968]  ( .D(o[968]), .CLK(clk), .RST(rst), .I(g_init[968]), .Q(
        creg[968]) );
  DFF \creg_reg[969]  ( .D(o[969]), .CLK(clk), .RST(rst), .I(g_init[969]), .Q(
        creg[969]) );
  DFF \creg_reg[970]  ( .D(o[970]), .CLK(clk), .RST(rst), .I(g_init[970]), .Q(
        creg[970]) );
  DFF \creg_reg[971]  ( .D(o[971]), .CLK(clk), .RST(rst), .I(g_init[971]), .Q(
        creg[971]) );
  DFF \creg_reg[972]  ( .D(o[972]), .CLK(clk), .RST(rst), .I(g_init[972]), .Q(
        creg[972]) );
  DFF \creg_reg[973]  ( .D(o[973]), .CLK(clk), .RST(rst), .I(g_init[973]), .Q(
        creg[973]) );
  DFF \creg_reg[974]  ( .D(o[974]), .CLK(clk), .RST(rst), .I(g_init[974]), .Q(
        creg[974]) );
  DFF \creg_reg[975]  ( .D(o[975]), .CLK(clk), .RST(rst), .I(g_init[975]), .Q(
        creg[975]) );
  DFF \creg_reg[976]  ( .D(o[976]), .CLK(clk), .RST(rst), .I(g_init[976]), .Q(
        creg[976]) );
  DFF \creg_reg[977]  ( .D(o[977]), .CLK(clk), .RST(rst), .I(g_init[977]), .Q(
        creg[977]) );
  DFF \creg_reg[978]  ( .D(o[978]), .CLK(clk), .RST(rst), .I(g_init[978]), .Q(
        creg[978]) );
  DFF \creg_reg[979]  ( .D(o[979]), .CLK(clk), .RST(rst), .I(g_init[979]), .Q(
        creg[979]) );
  DFF \creg_reg[980]  ( .D(o[980]), .CLK(clk), .RST(rst), .I(g_init[980]), .Q(
        creg[980]) );
  DFF \creg_reg[981]  ( .D(o[981]), .CLK(clk), .RST(rst), .I(g_init[981]), .Q(
        creg[981]) );
  DFF \creg_reg[982]  ( .D(o[982]), .CLK(clk), .RST(rst), .I(g_init[982]), .Q(
        creg[982]) );
  DFF \creg_reg[983]  ( .D(o[983]), .CLK(clk), .RST(rst), .I(g_init[983]), .Q(
        creg[983]) );
  DFF \creg_reg[984]  ( .D(o[984]), .CLK(clk), .RST(rst), .I(g_init[984]), .Q(
        creg[984]) );
  DFF \creg_reg[985]  ( .D(o[985]), .CLK(clk), .RST(rst), .I(g_init[985]), .Q(
        creg[985]) );
  DFF \creg_reg[986]  ( .D(o[986]), .CLK(clk), .RST(rst), .I(g_init[986]), .Q(
        creg[986]) );
  DFF \creg_reg[987]  ( .D(o[987]), .CLK(clk), .RST(rst), .I(g_init[987]), .Q(
        creg[987]) );
  DFF \creg_reg[988]  ( .D(o[988]), .CLK(clk), .RST(rst), .I(g_init[988]), .Q(
        creg[988]) );
  DFF \creg_reg[989]  ( .D(o[989]), .CLK(clk), .RST(rst), .I(g_init[989]), .Q(
        creg[989]) );
  DFF \creg_reg[990]  ( .D(o[990]), .CLK(clk), .RST(rst), .I(g_init[990]), .Q(
        creg[990]) );
  DFF \creg_reg[991]  ( .D(o[991]), .CLK(clk), .RST(rst), .I(g_init[991]), .Q(
        creg[991]) );
  DFF \creg_reg[992]  ( .D(o[992]), .CLK(clk), .RST(rst), .I(g_init[992]), .Q(
        creg[992]) );
  DFF \creg_reg[993]  ( .D(o[993]), .CLK(clk), .RST(rst), .I(g_init[993]), .Q(
        creg[993]) );
  DFF \creg_reg[994]  ( .D(o[994]), .CLK(clk), .RST(rst), .I(g_init[994]), .Q(
        creg[994]) );
  DFF \creg_reg[995]  ( .D(o[995]), .CLK(clk), .RST(rst), .I(g_init[995]), .Q(
        creg[995]) );
  DFF \creg_reg[996]  ( .D(o[996]), .CLK(clk), .RST(rst), .I(g_init[996]), .Q(
        creg[996]) );
  DFF \creg_reg[997]  ( .D(o[997]), .CLK(clk), .RST(rst), .I(g_init[997]), .Q(
        creg[997]) );
  DFF \creg_reg[998]  ( .D(o[998]), .CLK(clk), .RST(rst), .I(g_init[998]), .Q(
        creg[998]) );
  DFF \creg_reg[999]  ( .D(o[999]), .CLK(clk), .RST(rst), .I(g_init[999]), .Q(
        creg[999]) );
  DFF \creg_reg[1000]  ( .D(o[1000]), .CLK(clk), .RST(rst), .I(g_init[1000]), 
        .Q(creg[1000]) );
  DFF \creg_reg[1001]  ( .D(o[1001]), .CLK(clk), .RST(rst), .I(g_init[1001]), 
        .Q(creg[1001]) );
  DFF \creg_reg[1002]  ( .D(o[1002]), .CLK(clk), .RST(rst), .I(g_init[1002]), 
        .Q(creg[1002]) );
  DFF \creg_reg[1003]  ( .D(o[1003]), .CLK(clk), .RST(rst), .I(g_init[1003]), 
        .Q(creg[1003]) );
  DFF \creg_reg[1004]  ( .D(o[1004]), .CLK(clk), .RST(rst), .I(g_init[1004]), 
        .Q(creg[1004]) );
  DFF \creg_reg[1005]  ( .D(o[1005]), .CLK(clk), .RST(rst), .I(g_init[1005]), 
        .Q(creg[1005]) );
  DFF \creg_reg[1006]  ( .D(o[1006]), .CLK(clk), .RST(rst), .I(g_init[1006]), 
        .Q(creg[1006]) );
  DFF \creg_reg[1007]  ( .D(o[1007]), .CLK(clk), .RST(rst), .I(g_init[1007]), 
        .Q(creg[1007]) );
  DFF \creg_reg[1008]  ( .D(o[1008]), .CLK(clk), .RST(rst), .I(g_init[1008]), 
        .Q(creg[1008]) );
  DFF \creg_reg[1009]  ( .D(o[1009]), .CLK(clk), .RST(rst), .I(g_init[1009]), 
        .Q(creg[1009]) );
  DFF \creg_reg[1010]  ( .D(o[1010]), .CLK(clk), .RST(rst), .I(g_init[1010]), 
        .Q(creg[1010]) );
  DFF \creg_reg[1011]  ( .D(o[1011]), .CLK(clk), .RST(rst), .I(g_init[1011]), 
        .Q(creg[1011]) );
  DFF \creg_reg[1012]  ( .D(o[1012]), .CLK(clk), .RST(rst), .I(g_init[1012]), 
        .Q(creg[1012]) );
  DFF \creg_reg[1013]  ( .D(o[1013]), .CLK(clk), .RST(rst), .I(g_init[1013]), 
        .Q(creg[1013]) );
  DFF \creg_reg[1014]  ( .D(o[1014]), .CLK(clk), .RST(rst), .I(g_init[1014]), 
        .Q(creg[1014]) );
  DFF \creg_reg[1015]  ( .D(o[1015]), .CLK(clk), .RST(rst), .I(g_init[1015]), 
        .Q(creg[1015]) );
  DFF \creg_reg[1016]  ( .D(o[1016]), .CLK(clk), .RST(rst), .I(g_init[1016]), 
        .Q(creg[1016]) );
  DFF \creg_reg[1017]  ( .D(o[1017]), .CLK(clk), .RST(rst), .I(g_init[1017]), 
        .Q(creg[1017]) );
  DFF \creg_reg[1018]  ( .D(o[1018]), .CLK(clk), .RST(rst), .I(g_init[1018]), 
        .Q(creg[1018]) );
  DFF \creg_reg[1019]  ( .D(o[1019]), .CLK(clk), .RST(rst), .I(g_init[1019]), 
        .Q(creg[1019]) );
  DFF \creg_reg[1020]  ( .D(o[1020]), .CLK(clk), .RST(rst), .I(g_init[1020]), 
        .Q(creg[1020]) );
  DFF \creg_reg[1021]  ( .D(o[1021]), .CLK(clk), .RST(rst), .I(g_init[1021]), 
        .Q(creg[1021]) );
  DFF \creg_reg[1022]  ( .D(o[1022]), .CLK(clk), .RST(rst), .I(g_init[1022]), 
        .Q(creg[1022]) );
  DFF \creg_reg[1023]  ( .D(o[1023]), .CLK(clk), .RST(rst), .I(g_init[1023]), 
        .Q(creg[1023]) );
  DFF \modmult_1/zreg_reg[1024]  ( .D(\modmult_1/N1027 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1024] ) );
  DFF \modmult_1/zreg_reg[1023]  ( .D(\modmult_1/N1026 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1023] ) );
  DFF \modmult_1/zreg_reg[1022]  ( .D(\modmult_1/N1025 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1022] ) );
  DFF \modmult_1/zreg_reg[1021]  ( .D(\modmult_1/N1024 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1021] ) );
  DFF \modmult_1/zreg_reg[1020]  ( .D(\modmult_1/N1023 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1020] ) );
  DFF \modmult_1/zreg_reg[1019]  ( .D(\modmult_1/N1022 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1019] ) );
  DFF \modmult_1/zreg_reg[1018]  ( .D(\modmult_1/N1021 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1018] ) );
  DFF \modmult_1/zreg_reg[1017]  ( .D(\modmult_1/N1020 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1017] ) );
  DFF \modmult_1/zreg_reg[1016]  ( .D(\modmult_1/N1019 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1016] ) );
  DFF \modmult_1/zreg_reg[1015]  ( .D(\modmult_1/N1018 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1015] ) );
  DFF \modmult_1/zreg_reg[1014]  ( .D(\modmult_1/N1017 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1014] ) );
  DFF \modmult_1/zreg_reg[1013]  ( .D(\modmult_1/N1016 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1013] ) );
  DFF \modmult_1/zreg_reg[1012]  ( .D(\modmult_1/N1015 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1012] ) );
  DFF \modmult_1/zreg_reg[1011]  ( .D(\modmult_1/N1014 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1011] ) );
  DFF \modmult_1/zreg_reg[1010]  ( .D(\modmult_1/N1013 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1010] ) );
  DFF \modmult_1/zreg_reg[1009]  ( .D(\modmult_1/N1012 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1009] ) );
  DFF \modmult_1/zreg_reg[1008]  ( .D(\modmult_1/N1011 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1008] ) );
  DFF \modmult_1/zreg_reg[1007]  ( .D(\modmult_1/N1010 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1007] ) );
  DFF \modmult_1/zreg_reg[1006]  ( .D(\modmult_1/N1009 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1006] ) );
  DFF \modmult_1/zreg_reg[1005]  ( .D(\modmult_1/N1008 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1005] ) );
  DFF \modmult_1/zreg_reg[1004]  ( .D(\modmult_1/N1007 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1004] ) );
  DFF \modmult_1/zreg_reg[1003]  ( .D(\modmult_1/N1006 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1003] ) );
  DFF \modmult_1/zreg_reg[1002]  ( .D(\modmult_1/N1005 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1002] ) );
  DFF \modmult_1/zreg_reg[1001]  ( .D(\modmult_1/N1004 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1001] ) );
  DFF \modmult_1/zreg_reg[1000]  ( .D(\modmult_1/N1003 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][1000] ) );
  DFF \modmult_1/zreg_reg[999]  ( .D(\modmult_1/N1002 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][999] ) );
  DFF \modmult_1/zreg_reg[998]  ( .D(\modmult_1/N1001 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][998] ) );
  DFF \modmult_1/zreg_reg[997]  ( .D(\modmult_1/N1000 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][997] ) );
  DFF \modmult_1/zreg_reg[996]  ( .D(\modmult_1/N999 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][996] ) );
  DFF \modmult_1/zreg_reg[995]  ( .D(\modmult_1/N998 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][995] ) );
  DFF \modmult_1/zreg_reg[994]  ( .D(\modmult_1/N997 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][994] ) );
  DFF \modmult_1/zreg_reg[993]  ( .D(\modmult_1/N996 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][993] ) );
  DFF \modmult_1/zreg_reg[992]  ( .D(\modmult_1/N995 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][992] ) );
  DFF \modmult_1/zreg_reg[991]  ( .D(\modmult_1/N994 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][991] ) );
  DFF \modmult_1/zreg_reg[990]  ( .D(\modmult_1/N993 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][990] ) );
  DFF \modmult_1/zreg_reg[989]  ( .D(\modmult_1/N992 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][989] ) );
  DFF \modmult_1/zreg_reg[988]  ( .D(\modmult_1/N991 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][988] ) );
  DFF \modmult_1/zreg_reg[987]  ( .D(\modmult_1/N990 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][987] ) );
  DFF \modmult_1/zreg_reg[986]  ( .D(\modmult_1/N989 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][986] ) );
  DFF \modmult_1/zreg_reg[985]  ( .D(\modmult_1/N988 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][985] ) );
  DFF \modmult_1/zreg_reg[984]  ( .D(\modmult_1/N987 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][984] ) );
  DFF \modmult_1/zreg_reg[983]  ( .D(\modmult_1/N986 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][983] ) );
  DFF \modmult_1/zreg_reg[982]  ( .D(\modmult_1/N985 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][982] ) );
  DFF \modmult_1/zreg_reg[981]  ( .D(\modmult_1/N984 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][981] ) );
  DFF \modmult_1/zreg_reg[980]  ( .D(\modmult_1/N983 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][980] ) );
  DFF \modmult_1/zreg_reg[979]  ( .D(\modmult_1/N982 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][979] ) );
  DFF \modmult_1/zreg_reg[978]  ( .D(\modmult_1/N981 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][978] ) );
  DFF \modmult_1/zreg_reg[977]  ( .D(\modmult_1/N980 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][977] ) );
  DFF \modmult_1/zreg_reg[976]  ( .D(\modmult_1/N979 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][976] ) );
  DFF \modmult_1/zreg_reg[975]  ( .D(\modmult_1/N978 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][975] ) );
  DFF \modmult_1/zreg_reg[974]  ( .D(\modmult_1/N977 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][974] ) );
  DFF \modmult_1/zreg_reg[973]  ( .D(\modmult_1/N976 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][973] ) );
  DFF \modmult_1/zreg_reg[972]  ( .D(\modmult_1/N975 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][972] ) );
  DFF \modmult_1/zreg_reg[971]  ( .D(\modmult_1/N974 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][971] ) );
  DFF \modmult_1/zreg_reg[970]  ( .D(\modmult_1/N973 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][970] ) );
  DFF \modmult_1/zreg_reg[969]  ( .D(\modmult_1/N972 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][969] ) );
  DFF \modmult_1/zreg_reg[968]  ( .D(\modmult_1/N971 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][968] ) );
  DFF \modmult_1/zreg_reg[967]  ( .D(\modmult_1/N970 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][967] ) );
  DFF \modmult_1/zreg_reg[966]  ( .D(\modmult_1/N969 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][966] ) );
  DFF \modmult_1/zreg_reg[965]  ( .D(\modmult_1/N968 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][965] ) );
  DFF \modmult_1/zreg_reg[964]  ( .D(\modmult_1/N967 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][964] ) );
  DFF \modmult_1/zreg_reg[963]  ( .D(\modmult_1/N966 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][963] ) );
  DFF \modmult_1/zreg_reg[962]  ( .D(\modmult_1/N965 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][962] ) );
  DFF \modmult_1/zreg_reg[961]  ( .D(\modmult_1/N964 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][961] ) );
  DFF \modmult_1/zreg_reg[960]  ( .D(\modmult_1/N963 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][960] ) );
  DFF \modmult_1/zreg_reg[959]  ( .D(\modmult_1/N962 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][959] ) );
  DFF \modmult_1/zreg_reg[958]  ( .D(\modmult_1/N961 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][958] ) );
  DFF \modmult_1/zreg_reg[957]  ( .D(\modmult_1/N960 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][957] ) );
  DFF \modmult_1/zreg_reg[956]  ( .D(\modmult_1/N959 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][956] ) );
  DFF \modmult_1/zreg_reg[955]  ( .D(\modmult_1/N958 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][955] ) );
  DFF \modmult_1/zreg_reg[954]  ( .D(\modmult_1/N957 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][954] ) );
  DFF \modmult_1/zreg_reg[953]  ( .D(\modmult_1/N956 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][953] ) );
  DFF \modmult_1/zreg_reg[952]  ( .D(\modmult_1/N955 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][952] ) );
  DFF \modmult_1/zreg_reg[951]  ( .D(\modmult_1/N954 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][951] ) );
  DFF \modmult_1/zreg_reg[950]  ( .D(\modmult_1/N953 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][950] ) );
  DFF \modmult_1/zreg_reg[949]  ( .D(\modmult_1/N952 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][949] ) );
  DFF \modmult_1/zreg_reg[948]  ( .D(\modmult_1/N951 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][948] ) );
  DFF \modmult_1/zreg_reg[947]  ( .D(\modmult_1/N950 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][947] ) );
  DFF \modmult_1/zreg_reg[946]  ( .D(\modmult_1/N949 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][946] ) );
  DFF \modmult_1/zreg_reg[945]  ( .D(\modmult_1/N948 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][945] ) );
  DFF \modmult_1/zreg_reg[944]  ( .D(\modmult_1/N947 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][944] ) );
  DFF \modmult_1/zreg_reg[943]  ( .D(\modmult_1/N946 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][943] ) );
  DFF \modmult_1/zreg_reg[942]  ( .D(\modmult_1/N945 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][942] ) );
  DFF \modmult_1/zreg_reg[941]  ( .D(\modmult_1/N944 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][941] ) );
  DFF \modmult_1/zreg_reg[940]  ( .D(\modmult_1/N943 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][940] ) );
  DFF \modmult_1/zreg_reg[939]  ( .D(\modmult_1/N942 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][939] ) );
  DFF \modmult_1/zreg_reg[938]  ( .D(\modmult_1/N941 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][938] ) );
  DFF \modmult_1/zreg_reg[937]  ( .D(\modmult_1/N940 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][937] ) );
  DFF \modmult_1/zreg_reg[936]  ( .D(\modmult_1/N939 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][936] ) );
  DFF \modmult_1/zreg_reg[935]  ( .D(\modmult_1/N938 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][935] ) );
  DFF \modmult_1/zreg_reg[934]  ( .D(\modmult_1/N937 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][934] ) );
  DFF \modmult_1/zreg_reg[933]  ( .D(\modmult_1/N936 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][933] ) );
  DFF \modmult_1/zreg_reg[932]  ( .D(\modmult_1/N935 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][932] ) );
  DFF \modmult_1/zreg_reg[931]  ( .D(\modmult_1/N934 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][931] ) );
  DFF \modmult_1/zreg_reg[930]  ( .D(\modmult_1/N933 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][930] ) );
  DFF \modmult_1/zreg_reg[929]  ( .D(\modmult_1/N932 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][929] ) );
  DFF \modmult_1/zreg_reg[928]  ( .D(\modmult_1/N931 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][928] ) );
  DFF \modmult_1/zreg_reg[927]  ( .D(\modmult_1/N930 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][927] ) );
  DFF \modmult_1/zreg_reg[926]  ( .D(\modmult_1/N929 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][926] ) );
  DFF \modmult_1/zreg_reg[925]  ( .D(\modmult_1/N928 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][925] ) );
  DFF \modmult_1/zreg_reg[924]  ( .D(\modmult_1/N927 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][924] ) );
  DFF \modmult_1/zreg_reg[923]  ( .D(\modmult_1/N926 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][923] ) );
  DFF \modmult_1/zreg_reg[922]  ( .D(\modmult_1/N925 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][922] ) );
  DFF \modmult_1/zreg_reg[921]  ( .D(\modmult_1/N924 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][921] ) );
  DFF \modmult_1/zreg_reg[920]  ( .D(\modmult_1/N923 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][920] ) );
  DFF \modmult_1/zreg_reg[919]  ( .D(\modmult_1/N922 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][919] ) );
  DFF \modmult_1/zreg_reg[918]  ( .D(\modmult_1/N921 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][918] ) );
  DFF \modmult_1/zreg_reg[917]  ( .D(\modmult_1/N920 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][917] ) );
  DFF \modmult_1/zreg_reg[916]  ( .D(\modmult_1/N919 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][916] ) );
  DFF \modmult_1/zreg_reg[915]  ( .D(\modmult_1/N918 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][915] ) );
  DFF \modmult_1/zreg_reg[914]  ( .D(\modmult_1/N917 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][914] ) );
  DFF \modmult_1/zreg_reg[913]  ( .D(\modmult_1/N916 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][913] ) );
  DFF \modmult_1/zreg_reg[912]  ( .D(\modmult_1/N915 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][912] ) );
  DFF \modmult_1/zreg_reg[911]  ( .D(\modmult_1/N914 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][911] ) );
  DFF \modmult_1/zreg_reg[910]  ( .D(\modmult_1/N913 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][910] ) );
  DFF \modmult_1/zreg_reg[909]  ( .D(\modmult_1/N912 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][909] ) );
  DFF \modmult_1/zreg_reg[908]  ( .D(\modmult_1/N911 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][908] ) );
  DFF \modmult_1/zreg_reg[907]  ( .D(\modmult_1/N910 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][907] ) );
  DFF \modmult_1/zreg_reg[906]  ( .D(\modmult_1/N909 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][906] ) );
  DFF \modmult_1/zreg_reg[905]  ( .D(\modmult_1/N908 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][905] ) );
  DFF \modmult_1/zreg_reg[904]  ( .D(\modmult_1/N907 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][904] ) );
  DFF \modmult_1/zreg_reg[903]  ( .D(\modmult_1/N906 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][903] ) );
  DFF \modmult_1/zreg_reg[902]  ( .D(\modmult_1/N905 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][902] ) );
  DFF \modmult_1/zreg_reg[901]  ( .D(\modmult_1/N904 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][901] ) );
  DFF \modmult_1/zreg_reg[900]  ( .D(\modmult_1/N903 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][900] ) );
  DFF \modmult_1/zreg_reg[899]  ( .D(\modmult_1/N902 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][899] ) );
  DFF \modmult_1/zreg_reg[898]  ( .D(\modmult_1/N901 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][898] ) );
  DFF \modmult_1/zreg_reg[897]  ( .D(\modmult_1/N900 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][897] ) );
  DFF \modmult_1/zreg_reg[896]  ( .D(\modmult_1/N899 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][896] ) );
  DFF \modmult_1/zreg_reg[895]  ( .D(\modmult_1/N898 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][895] ) );
  DFF \modmult_1/zreg_reg[894]  ( .D(\modmult_1/N897 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][894] ) );
  DFF \modmult_1/zreg_reg[893]  ( .D(\modmult_1/N896 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][893] ) );
  DFF \modmult_1/zreg_reg[892]  ( .D(\modmult_1/N895 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][892] ) );
  DFF \modmult_1/zreg_reg[891]  ( .D(\modmult_1/N894 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][891] ) );
  DFF \modmult_1/zreg_reg[890]  ( .D(\modmult_1/N893 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][890] ) );
  DFF \modmult_1/zreg_reg[889]  ( .D(\modmult_1/N892 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][889] ) );
  DFF \modmult_1/zreg_reg[888]  ( .D(\modmult_1/N891 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][888] ) );
  DFF \modmult_1/zreg_reg[887]  ( .D(\modmult_1/N890 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][887] ) );
  DFF \modmult_1/zreg_reg[886]  ( .D(\modmult_1/N889 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][886] ) );
  DFF \modmult_1/zreg_reg[885]  ( .D(\modmult_1/N888 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][885] ) );
  DFF \modmult_1/zreg_reg[884]  ( .D(\modmult_1/N887 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][884] ) );
  DFF \modmult_1/zreg_reg[883]  ( .D(\modmult_1/N886 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][883] ) );
  DFF \modmult_1/zreg_reg[882]  ( .D(\modmult_1/N885 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][882] ) );
  DFF \modmult_1/zreg_reg[881]  ( .D(\modmult_1/N884 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][881] ) );
  DFF \modmult_1/zreg_reg[880]  ( .D(\modmult_1/N883 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][880] ) );
  DFF \modmult_1/zreg_reg[879]  ( .D(\modmult_1/N882 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][879] ) );
  DFF \modmult_1/zreg_reg[878]  ( .D(\modmult_1/N881 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][878] ) );
  DFF \modmult_1/zreg_reg[877]  ( .D(\modmult_1/N880 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][877] ) );
  DFF \modmult_1/zreg_reg[876]  ( .D(\modmult_1/N879 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][876] ) );
  DFF \modmult_1/zreg_reg[875]  ( .D(\modmult_1/N878 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][875] ) );
  DFF \modmult_1/zreg_reg[874]  ( .D(\modmult_1/N877 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][874] ) );
  DFF \modmult_1/zreg_reg[873]  ( .D(\modmult_1/N876 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][873] ) );
  DFF \modmult_1/zreg_reg[872]  ( .D(\modmult_1/N875 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][872] ) );
  DFF \modmult_1/zreg_reg[871]  ( .D(\modmult_1/N874 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][871] ) );
  DFF \modmult_1/zreg_reg[870]  ( .D(\modmult_1/N873 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][870] ) );
  DFF \modmult_1/zreg_reg[869]  ( .D(\modmult_1/N872 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][869] ) );
  DFF \modmult_1/zreg_reg[868]  ( .D(\modmult_1/N871 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][868] ) );
  DFF \modmult_1/zreg_reg[867]  ( .D(\modmult_1/N870 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][867] ) );
  DFF \modmult_1/zreg_reg[866]  ( .D(\modmult_1/N869 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][866] ) );
  DFF \modmult_1/zreg_reg[865]  ( .D(\modmult_1/N868 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][865] ) );
  DFF \modmult_1/zreg_reg[864]  ( .D(\modmult_1/N867 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][864] ) );
  DFF \modmult_1/zreg_reg[863]  ( .D(\modmult_1/N866 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][863] ) );
  DFF \modmult_1/zreg_reg[862]  ( .D(\modmult_1/N865 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][862] ) );
  DFF \modmult_1/zreg_reg[861]  ( .D(\modmult_1/N864 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][861] ) );
  DFF \modmult_1/zreg_reg[860]  ( .D(\modmult_1/N863 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][860] ) );
  DFF \modmult_1/zreg_reg[859]  ( .D(\modmult_1/N862 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][859] ) );
  DFF \modmult_1/zreg_reg[858]  ( .D(\modmult_1/N861 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][858] ) );
  DFF \modmult_1/zreg_reg[857]  ( .D(\modmult_1/N860 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][857] ) );
  DFF \modmult_1/zreg_reg[856]  ( .D(\modmult_1/N859 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][856] ) );
  DFF \modmult_1/zreg_reg[855]  ( .D(\modmult_1/N858 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][855] ) );
  DFF \modmult_1/zreg_reg[854]  ( .D(\modmult_1/N857 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][854] ) );
  DFF \modmult_1/zreg_reg[853]  ( .D(\modmult_1/N856 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][853] ) );
  DFF \modmult_1/zreg_reg[852]  ( .D(\modmult_1/N855 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][852] ) );
  DFF \modmult_1/zreg_reg[851]  ( .D(\modmult_1/N854 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][851] ) );
  DFF \modmult_1/zreg_reg[850]  ( .D(\modmult_1/N853 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][850] ) );
  DFF \modmult_1/zreg_reg[849]  ( .D(\modmult_1/N852 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][849] ) );
  DFF \modmult_1/zreg_reg[848]  ( .D(\modmult_1/N851 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][848] ) );
  DFF \modmult_1/zreg_reg[847]  ( .D(\modmult_1/N850 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][847] ) );
  DFF \modmult_1/zreg_reg[846]  ( .D(\modmult_1/N849 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][846] ) );
  DFF \modmult_1/zreg_reg[845]  ( .D(\modmult_1/N848 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][845] ) );
  DFF \modmult_1/zreg_reg[844]  ( .D(\modmult_1/N847 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][844] ) );
  DFF \modmult_1/zreg_reg[843]  ( .D(\modmult_1/N846 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][843] ) );
  DFF \modmult_1/zreg_reg[842]  ( .D(\modmult_1/N845 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][842] ) );
  DFF \modmult_1/zreg_reg[841]  ( .D(\modmult_1/N844 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][841] ) );
  DFF \modmult_1/zreg_reg[840]  ( .D(\modmult_1/N843 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][840] ) );
  DFF \modmult_1/zreg_reg[839]  ( .D(\modmult_1/N842 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][839] ) );
  DFF \modmult_1/zreg_reg[838]  ( .D(\modmult_1/N841 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][838] ) );
  DFF \modmult_1/zreg_reg[837]  ( .D(\modmult_1/N840 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][837] ) );
  DFF \modmult_1/zreg_reg[836]  ( .D(\modmult_1/N839 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][836] ) );
  DFF \modmult_1/zreg_reg[835]  ( .D(\modmult_1/N838 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][835] ) );
  DFF \modmult_1/zreg_reg[834]  ( .D(\modmult_1/N837 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][834] ) );
  DFF \modmult_1/zreg_reg[833]  ( .D(\modmult_1/N836 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][833] ) );
  DFF \modmult_1/zreg_reg[832]  ( .D(\modmult_1/N835 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][832] ) );
  DFF \modmult_1/zreg_reg[831]  ( .D(\modmult_1/N834 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][831] ) );
  DFF \modmult_1/zreg_reg[830]  ( .D(\modmult_1/N833 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][830] ) );
  DFF \modmult_1/zreg_reg[829]  ( .D(\modmult_1/N832 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][829] ) );
  DFF \modmult_1/zreg_reg[828]  ( .D(\modmult_1/N831 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][828] ) );
  DFF \modmult_1/zreg_reg[827]  ( .D(\modmult_1/N830 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][827] ) );
  DFF \modmult_1/zreg_reg[826]  ( .D(\modmult_1/N829 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][826] ) );
  DFF \modmult_1/zreg_reg[825]  ( .D(\modmult_1/N828 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][825] ) );
  DFF \modmult_1/zreg_reg[824]  ( .D(\modmult_1/N827 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][824] ) );
  DFF \modmult_1/zreg_reg[823]  ( .D(\modmult_1/N826 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][823] ) );
  DFF \modmult_1/zreg_reg[822]  ( .D(\modmult_1/N825 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][822] ) );
  DFF \modmult_1/zreg_reg[821]  ( .D(\modmult_1/N824 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][821] ) );
  DFF \modmult_1/zreg_reg[820]  ( .D(\modmult_1/N823 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][820] ) );
  DFF \modmult_1/zreg_reg[819]  ( .D(\modmult_1/N822 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][819] ) );
  DFF \modmult_1/zreg_reg[818]  ( .D(\modmult_1/N821 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][818] ) );
  DFF \modmult_1/zreg_reg[817]  ( .D(\modmult_1/N820 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][817] ) );
  DFF \modmult_1/zreg_reg[816]  ( .D(\modmult_1/N819 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][816] ) );
  DFF \modmult_1/zreg_reg[815]  ( .D(\modmult_1/N818 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][815] ) );
  DFF \modmult_1/zreg_reg[814]  ( .D(\modmult_1/N817 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][814] ) );
  DFF \modmult_1/zreg_reg[813]  ( .D(\modmult_1/N816 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][813] ) );
  DFF \modmult_1/zreg_reg[812]  ( .D(\modmult_1/N815 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][812] ) );
  DFF \modmult_1/zreg_reg[811]  ( .D(\modmult_1/N814 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][811] ) );
  DFF \modmult_1/zreg_reg[810]  ( .D(\modmult_1/N813 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][810] ) );
  DFF \modmult_1/zreg_reg[809]  ( .D(\modmult_1/N812 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][809] ) );
  DFF \modmult_1/zreg_reg[808]  ( .D(\modmult_1/N811 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][808] ) );
  DFF \modmult_1/zreg_reg[807]  ( .D(\modmult_1/N810 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][807] ) );
  DFF \modmult_1/zreg_reg[806]  ( .D(\modmult_1/N809 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][806] ) );
  DFF \modmult_1/zreg_reg[805]  ( .D(\modmult_1/N808 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][805] ) );
  DFF \modmult_1/zreg_reg[804]  ( .D(\modmult_1/N807 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][804] ) );
  DFF \modmult_1/zreg_reg[803]  ( .D(\modmult_1/N806 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][803] ) );
  DFF \modmult_1/zreg_reg[802]  ( .D(\modmult_1/N805 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][802] ) );
  DFF \modmult_1/zreg_reg[801]  ( .D(\modmult_1/N804 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][801] ) );
  DFF \modmult_1/zreg_reg[800]  ( .D(\modmult_1/N803 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][800] ) );
  DFF \modmult_1/zreg_reg[799]  ( .D(\modmult_1/N802 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][799] ) );
  DFF \modmult_1/zreg_reg[798]  ( .D(\modmult_1/N801 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][798] ) );
  DFF \modmult_1/zreg_reg[797]  ( .D(\modmult_1/N800 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][797] ) );
  DFF \modmult_1/zreg_reg[796]  ( .D(\modmult_1/N799 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][796] ) );
  DFF \modmult_1/zreg_reg[795]  ( .D(\modmult_1/N798 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][795] ) );
  DFF \modmult_1/zreg_reg[794]  ( .D(\modmult_1/N797 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][794] ) );
  DFF \modmult_1/zreg_reg[793]  ( .D(\modmult_1/N796 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][793] ) );
  DFF \modmult_1/zreg_reg[792]  ( .D(\modmult_1/N795 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][792] ) );
  DFF \modmult_1/zreg_reg[791]  ( .D(\modmult_1/N794 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][791] ) );
  DFF \modmult_1/zreg_reg[790]  ( .D(\modmult_1/N793 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][790] ) );
  DFF \modmult_1/zreg_reg[789]  ( .D(\modmult_1/N792 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][789] ) );
  DFF \modmult_1/zreg_reg[788]  ( .D(\modmult_1/N791 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][788] ) );
  DFF \modmult_1/zreg_reg[787]  ( .D(\modmult_1/N790 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][787] ) );
  DFF \modmult_1/zreg_reg[786]  ( .D(\modmult_1/N789 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][786] ) );
  DFF \modmult_1/zreg_reg[785]  ( .D(\modmult_1/N788 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][785] ) );
  DFF \modmult_1/zreg_reg[784]  ( .D(\modmult_1/N787 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][784] ) );
  DFF \modmult_1/zreg_reg[783]  ( .D(\modmult_1/N786 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][783] ) );
  DFF \modmult_1/zreg_reg[782]  ( .D(\modmult_1/N785 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][782] ) );
  DFF \modmult_1/zreg_reg[781]  ( .D(\modmult_1/N784 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][781] ) );
  DFF \modmult_1/zreg_reg[780]  ( .D(\modmult_1/N783 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][780] ) );
  DFF \modmult_1/zreg_reg[779]  ( .D(\modmult_1/N782 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][779] ) );
  DFF \modmult_1/zreg_reg[778]  ( .D(\modmult_1/N781 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][778] ) );
  DFF \modmult_1/zreg_reg[777]  ( .D(\modmult_1/N780 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][777] ) );
  DFF \modmult_1/zreg_reg[776]  ( .D(\modmult_1/N779 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][776] ) );
  DFF \modmult_1/zreg_reg[775]  ( .D(\modmult_1/N778 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][775] ) );
  DFF \modmult_1/zreg_reg[774]  ( .D(\modmult_1/N777 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][774] ) );
  DFF \modmult_1/zreg_reg[773]  ( .D(\modmult_1/N776 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][773] ) );
  DFF \modmult_1/zreg_reg[772]  ( .D(\modmult_1/N775 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][772] ) );
  DFF \modmult_1/zreg_reg[771]  ( .D(\modmult_1/N774 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][771] ) );
  DFF \modmult_1/zreg_reg[770]  ( .D(\modmult_1/N773 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][770] ) );
  DFF \modmult_1/zreg_reg[769]  ( .D(\modmult_1/N772 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][769] ) );
  DFF \modmult_1/zreg_reg[768]  ( .D(\modmult_1/N771 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][768] ) );
  DFF \modmult_1/zreg_reg[767]  ( .D(\modmult_1/N770 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][767] ) );
  DFF \modmult_1/zreg_reg[766]  ( .D(\modmult_1/N769 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][766] ) );
  DFF \modmult_1/zreg_reg[765]  ( .D(\modmult_1/N768 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][765] ) );
  DFF \modmult_1/zreg_reg[764]  ( .D(\modmult_1/N767 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][764] ) );
  DFF \modmult_1/zreg_reg[763]  ( .D(\modmult_1/N766 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][763] ) );
  DFF \modmult_1/zreg_reg[762]  ( .D(\modmult_1/N765 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][762] ) );
  DFF \modmult_1/zreg_reg[761]  ( .D(\modmult_1/N764 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][761] ) );
  DFF \modmult_1/zreg_reg[760]  ( .D(\modmult_1/N763 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][760] ) );
  DFF \modmult_1/zreg_reg[759]  ( .D(\modmult_1/N762 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][759] ) );
  DFF \modmult_1/zreg_reg[758]  ( .D(\modmult_1/N761 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][758] ) );
  DFF \modmult_1/zreg_reg[757]  ( .D(\modmult_1/N760 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][757] ) );
  DFF \modmult_1/zreg_reg[756]  ( .D(\modmult_1/N759 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][756] ) );
  DFF \modmult_1/zreg_reg[755]  ( .D(\modmult_1/N758 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][755] ) );
  DFF \modmult_1/zreg_reg[754]  ( .D(\modmult_1/N757 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][754] ) );
  DFF \modmult_1/zreg_reg[753]  ( .D(\modmult_1/N756 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][753] ) );
  DFF \modmult_1/zreg_reg[752]  ( .D(\modmult_1/N755 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][752] ) );
  DFF \modmult_1/zreg_reg[751]  ( .D(\modmult_1/N754 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][751] ) );
  DFF \modmult_1/zreg_reg[750]  ( .D(\modmult_1/N753 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][750] ) );
  DFF \modmult_1/zreg_reg[749]  ( .D(\modmult_1/N752 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][749] ) );
  DFF \modmult_1/zreg_reg[748]  ( .D(\modmult_1/N751 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][748] ) );
  DFF \modmult_1/zreg_reg[747]  ( .D(\modmult_1/N750 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][747] ) );
  DFF \modmult_1/zreg_reg[746]  ( .D(\modmult_1/N749 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][746] ) );
  DFF \modmult_1/zreg_reg[745]  ( .D(\modmult_1/N748 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][745] ) );
  DFF \modmult_1/zreg_reg[744]  ( .D(\modmult_1/N747 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][744] ) );
  DFF \modmult_1/zreg_reg[743]  ( .D(\modmult_1/N746 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][743] ) );
  DFF \modmult_1/zreg_reg[742]  ( .D(\modmult_1/N745 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][742] ) );
  DFF \modmult_1/zreg_reg[741]  ( .D(\modmult_1/N744 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][741] ) );
  DFF \modmult_1/zreg_reg[740]  ( .D(\modmult_1/N743 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][740] ) );
  DFF \modmult_1/zreg_reg[739]  ( .D(\modmult_1/N742 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][739] ) );
  DFF \modmult_1/zreg_reg[738]  ( .D(\modmult_1/N741 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][738] ) );
  DFF \modmult_1/zreg_reg[737]  ( .D(\modmult_1/N740 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][737] ) );
  DFF \modmult_1/zreg_reg[736]  ( .D(\modmult_1/N739 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][736] ) );
  DFF \modmult_1/zreg_reg[735]  ( .D(\modmult_1/N738 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][735] ) );
  DFF \modmult_1/zreg_reg[734]  ( .D(\modmult_1/N737 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][734] ) );
  DFF \modmult_1/zreg_reg[733]  ( .D(\modmult_1/N736 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][733] ) );
  DFF \modmult_1/zreg_reg[732]  ( .D(\modmult_1/N735 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][732] ) );
  DFF \modmult_1/zreg_reg[731]  ( .D(\modmult_1/N734 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][731] ) );
  DFF \modmult_1/zreg_reg[730]  ( .D(\modmult_1/N733 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][730] ) );
  DFF \modmult_1/zreg_reg[729]  ( .D(\modmult_1/N732 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][729] ) );
  DFF \modmult_1/zreg_reg[728]  ( .D(\modmult_1/N731 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][728] ) );
  DFF \modmult_1/zreg_reg[727]  ( .D(\modmult_1/N730 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][727] ) );
  DFF \modmult_1/zreg_reg[726]  ( .D(\modmult_1/N729 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][726] ) );
  DFF \modmult_1/zreg_reg[725]  ( .D(\modmult_1/N728 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][725] ) );
  DFF \modmult_1/zreg_reg[724]  ( .D(\modmult_1/N727 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][724] ) );
  DFF \modmult_1/zreg_reg[723]  ( .D(\modmult_1/N726 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][723] ) );
  DFF \modmult_1/zreg_reg[722]  ( .D(\modmult_1/N725 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][722] ) );
  DFF \modmult_1/zreg_reg[721]  ( .D(\modmult_1/N724 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][721] ) );
  DFF \modmult_1/zreg_reg[720]  ( .D(\modmult_1/N723 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][720] ) );
  DFF \modmult_1/zreg_reg[719]  ( .D(\modmult_1/N722 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][719] ) );
  DFF \modmult_1/zreg_reg[718]  ( .D(\modmult_1/N721 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][718] ) );
  DFF \modmult_1/zreg_reg[717]  ( .D(\modmult_1/N720 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][717] ) );
  DFF \modmult_1/zreg_reg[716]  ( .D(\modmult_1/N719 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][716] ) );
  DFF \modmult_1/zreg_reg[715]  ( .D(\modmult_1/N718 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][715] ) );
  DFF \modmult_1/zreg_reg[714]  ( .D(\modmult_1/N717 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][714] ) );
  DFF \modmult_1/zreg_reg[713]  ( .D(\modmult_1/N716 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][713] ) );
  DFF \modmult_1/zreg_reg[712]  ( .D(\modmult_1/N715 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][712] ) );
  DFF \modmult_1/zreg_reg[711]  ( .D(\modmult_1/N714 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][711] ) );
  DFF \modmult_1/zreg_reg[710]  ( .D(\modmult_1/N713 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][710] ) );
  DFF \modmult_1/zreg_reg[709]  ( .D(\modmult_1/N712 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][709] ) );
  DFF \modmult_1/zreg_reg[708]  ( .D(\modmult_1/N711 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][708] ) );
  DFF \modmult_1/zreg_reg[707]  ( .D(\modmult_1/N710 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][707] ) );
  DFF \modmult_1/zreg_reg[706]  ( .D(\modmult_1/N709 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][706] ) );
  DFF \modmult_1/zreg_reg[705]  ( .D(\modmult_1/N708 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][705] ) );
  DFF \modmult_1/zreg_reg[704]  ( .D(\modmult_1/N707 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][704] ) );
  DFF \modmult_1/zreg_reg[703]  ( .D(\modmult_1/N706 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][703] ) );
  DFF \modmult_1/zreg_reg[702]  ( .D(\modmult_1/N705 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][702] ) );
  DFF \modmult_1/zreg_reg[701]  ( .D(\modmult_1/N704 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][701] ) );
  DFF \modmult_1/zreg_reg[700]  ( .D(\modmult_1/N703 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][700] ) );
  DFF \modmult_1/zreg_reg[699]  ( .D(\modmult_1/N702 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][699] ) );
  DFF \modmult_1/zreg_reg[698]  ( .D(\modmult_1/N701 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][698] ) );
  DFF \modmult_1/zreg_reg[697]  ( .D(\modmult_1/N700 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][697] ) );
  DFF \modmult_1/zreg_reg[696]  ( .D(\modmult_1/N699 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][696] ) );
  DFF \modmult_1/zreg_reg[695]  ( .D(\modmult_1/N698 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][695] ) );
  DFF \modmult_1/zreg_reg[694]  ( .D(\modmult_1/N697 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][694] ) );
  DFF \modmult_1/zreg_reg[693]  ( .D(\modmult_1/N696 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][693] ) );
  DFF \modmult_1/zreg_reg[692]  ( .D(\modmult_1/N695 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][692] ) );
  DFF \modmult_1/zreg_reg[691]  ( .D(\modmult_1/N694 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][691] ) );
  DFF \modmult_1/zreg_reg[690]  ( .D(\modmult_1/N693 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][690] ) );
  DFF \modmult_1/zreg_reg[689]  ( .D(\modmult_1/N692 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][689] ) );
  DFF \modmult_1/zreg_reg[688]  ( .D(\modmult_1/N691 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][688] ) );
  DFF \modmult_1/zreg_reg[687]  ( .D(\modmult_1/N690 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][687] ) );
  DFF \modmult_1/zreg_reg[686]  ( .D(\modmult_1/N689 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][686] ) );
  DFF \modmult_1/zreg_reg[685]  ( .D(\modmult_1/N688 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][685] ) );
  DFF \modmult_1/zreg_reg[684]  ( .D(\modmult_1/N687 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][684] ) );
  DFF \modmult_1/zreg_reg[683]  ( .D(\modmult_1/N686 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][683] ) );
  DFF \modmult_1/zreg_reg[682]  ( .D(\modmult_1/N685 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][682] ) );
  DFF \modmult_1/zreg_reg[681]  ( .D(\modmult_1/N684 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][681] ) );
  DFF \modmult_1/zreg_reg[680]  ( .D(\modmult_1/N683 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][680] ) );
  DFF \modmult_1/zreg_reg[679]  ( .D(\modmult_1/N682 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][679] ) );
  DFF \modmult_1/zreg_reg[678]  ( .D(\modmult_1/N681 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][678] ) );
  DFF \modmult_1/zreg_reg[677]  ( .D(\modmult_1/N680 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][677] ) );
  DFF \modmult_1/zreg_reg[676]  ( .D(\modmult_1/N679 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][676] ) );
  DFF \modmult_1/zreg_reg[675]  ( .D(\modmult_1/N678 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][675] ) );
  DFF \modmult_1/zreg_reg[674]  ( .D(\modmult_1/N677 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][674] ) );
  DFF \modmult_1/zreg_reg[673]  ( .D(\modmult_1/N676 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][673] ) );
  DFF \modmult_1/zreg_reg[672]  ( .D(\modmult_1/N675 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][672] ) );
  DFF \modmult_1/zreg_reg[671]  ( .D(\modmult_1/N674 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][671] ) );
  DFF \modmult_1/zreg_reg[670]  ( .D(\modmult_1/N673 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][670] ) );
  DFF \modmult_1/zreg_reg[669]  ( .D(\modmult_1/N672 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][669] ) );
  DFF \modmult_1/zreg_reg[668]  ( .D(\modmult_1/N671 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][668] ) );
  DFF \modmult_1/zreg_reg[667]  ( .D(\modmult_1/N670 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][667] ) );
  DFF \modmult_1/zreg_reg[666]  ( .D(\modmult_1/N669 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][666] ) );
  DFF \modmult_1/zreg_reg[665]  ( .D(\modmult_1/N668 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][665] ) );
  DFF \modmult_1/zreg_reg[664]  ( .D(\modmult_1/N667 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][664] ) );
  DFF \modmult_1/zreg_reg[663]  ( .D(\modmult_1/N666 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][663] ) );
  DFF \modmult_1/zreg_reg[662]  ( .D(\modmult_1/N665 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][662] ) );
  DFF \modmult_1/zreg_reg[661]  ( .D(\modmult_1/N664 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][661] ) );
  DFF \modmult_1/zreg_reg[660]  ( .D(\modmult_1/N663 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][660] ) );
  DFF \modmult_1/zreg_reg[659]  ( .D(\modmult_1/N662 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][659] ) );
  DFF \modmult_1/zreg_reg[658]  ( .D(\modmult_1/N661 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][658] ) );
  DFF \modmult_1/zreg_reg[657]  ( .D(\modmult_1/N660 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][657] ) );
  DFF \modmult_1/zreg_reg[656]  ( .D(\modmult_1/N659 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][656] ) );
  DFF \modmult_1/zreg_reg[655]  ( .D(\modmult_1/N658 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][655] ) );
  DFF \modmult_1/zreg_reg[654]  ( .D(\modmult_1/N657 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][654] ) );
  DFF \modmult_1/zreg_reg[653]  ( .D(\modmult_1/N656 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][653] ) );
  DFF \modmult_1/zreg_reg[652]  ( .D(\modmult_1/N655 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][652] ) );
  DFF \modmult_1/zreg_reg[651]  ( .D(\modmult_1/N654 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][651] ) );
  DFF \modmult_1/zreg_reg[650]  ( .D(\modmult_1/N653 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][650] ) );
  DFF \modmult_1/zreg_reg[649]  ( .D(\modmult_1/N652 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][649] ) );
  DFF \modmult_1/zreg_reg[648]  ( .D(\modmult_1/N651 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][648] ) );
  DFF \modmult_1/zreg_reg[647]  ( .D(\modmult_1/N650 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][647] ) );
  DFF \modmult_1/zreg_reg[646]  ( .D(\modmult_1/N649 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][646] ) );
  DFF \modmult_1/zreg_reg[645]  ( .D(\modmult_1/N648 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][645] ) );
  DFF \modmult_1/zreg_reg[644]  ( .D(\modmult_1/N647 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][644] ) );
  DFF \modmult_1/zreg_reg[643]  ( .D(\modmult_1/N646 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][643] ) );
  DFF \modmult_1/zreg_reg[642]  ( .D(\modmult_1/N645 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][642] ) );
  DFF \modmult_1/zreg_reg[641]  ( .D(\modmult_1/N644 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][641] ) );
  DFF \modmult_1/zreg_reg[640]  ( .D(\modmult_1/N643 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][640] ) );
  DFF \modmult_1/zreg_reg[639]  ( .D(\modmult_1/N642 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][639] ) );
  DFF \modmult_1/zreg_reg[638]  ( .D(\modmult_1/N641 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][638] ) );
  DFF \modmult_1/zreg_reg[637]  ( .D(\modmult_1/N640 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][637] ) );
  DFF \modmult_1/zreg_reg[636]  ( .D(\modmult_1/N639 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][636] ) );
  DFF \modmult_1/zreg_reg[635]  ( .D(\modmult_1/N638 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][635] ) );
  DFF \modmult_1/zreg_reg[634]  ( .D(\modmult_1/N637 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][634] ) );
  DFF \modmult_1/zreg_reg[633]  ( .D(\modmult_1/N636 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][633] ) );
  DFF \modmult_1/zreg_reg[632]  ( .D(\modmult_1/N635 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][632] ) );
  DFF \modmult_1/zreg_reg[631]  ( .D(\modmult_1/N634 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][631] ) );
  DFF \modmult_1/zreg_reg[630]  ( .D(\modmult_1/N633 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][630] ) );
  DFF \modmult_1/zreg_reg[629]  ( .D(\modmult_1/N632 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][629] ) );
  DFF \modmult_1/zreg_reg[628]  ( .D(\modmult_1/N631 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][628] ) );
  DFF \modmult_1/zreg_reg[627]  ( .D(\modmult_1/N630 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][627] ) );
  DFF \modmult_1/zreg_reg[626]  ( .D(\modmult_1/N629 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][626] ) );
  DFF \modmult_1/zreg_reg[625]  ( .D(\modmult_1/N628 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][625] ) );
  DFF \modmult_1/zreg_reg[624]  ( .D(\modmult_1/N627 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][624] ) );
  DFF \modmult_1/zreg_reg[623]  ( .D(\modmult_1/N626 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][623] ) );
  DFF \modmult_1/zreg_reg[622]  ( .D(\modmult_1/N625 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][622] ) );
  DFF \modmult_1/zreg_reg[621]  ( .D(\modmult_1/N624 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][621] ) );
  DFF \modmult_1/zreg_reg[620]  ( .D(\modmult_1/N623 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][620] ) );
  DFF \modmult_1/zreg_reg[619]  ( .D(\modmult_1/N622 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][619] ) );
  DFF \modmult_1/zreg_reg[618]  ( .D(\modmult_1/N621 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][618] ) );
  DFF \modmult_1/zreg_reg[617]  ( .D(\modmult_1/N620 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][617] ) );
  DFF \modmult_1/zreg_reg[616]  ( .D(\modmult_1/N619 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][616] ) );
  DFF \modmult_1/zreg_reg[615]  ( .D(\modmult_1/N618 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][615] ) );
  DFF \modmult_1/zreg_reg[614]  ( .D(\modmult_1/N617 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][614] ) );
  DFF \modmult_1/zreg_reg[613]  ( .D(\modmult_1/N616 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][613] ) );
  DFF \modmult_1/zreg_reg[612]  ( .D(\modmult_1/N615 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][612] ) );
  DFF \modmult_1/zreg_reg[611]  ( .D(\modmult_1/N614 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][611] ) );
  DFF \modmult_1/zreg_reg[610]  ( .D(\modmult_1/N613 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][610] ) );
  DFF \modmult_1/zreg_reg[609]  ( .D(\modmult_1/N612 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][609] ) );
  DFF \modmult_1/zreg_reg[608]  ( .D(\modmult_1/N611 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][608] ) );
  DFF \modmult_1/zreg_reg[607]  ( .D(\modmult_1/N610 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][607] ) );
  DFF \modmult_1/zreg_reg[606]  ( .D(\modmult_1/N609 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][606] ) );
  DFF \modmult_1/zreg_reg[605]  ( .D(\modmult_1/N608 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][605] ) );
  DFF \modmult_1/zreg_reg[604]  ( .D(\modmult_1/N607 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][604] ) );
  DFF \modmult_1/zreg_reg[603]  ( .D(\modmult_1/N606 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][603] ) );
  DFF \modmult_1/zreg_reg[602]  ( .D(\modmult_1/N605 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][602] ) );
  DFF \modmult_1/zreg_reg[601]  ( .D(\modmult_1/N604 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][601] ) );
  DFF \modmult_1/zreg_reg[600]  ( .D(\modmult_1/N603 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][600] ) );
  DFF \modmult_1/zreg_reg[599]  ( .D(\modmult_1/N602 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][599] ) );
  DFF \modmult_1/zreg_reg[598]  ( .D(\modmult_1/N601 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][598] ) );
  DFF \modmult_1/zreg_reg[597]  ( .D(\modmult_1/N600 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][597] ) );
  DFF \modmult_1/zreg_reg[596]  ( .D(\modmult_1/N599 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][596] ) );
  DFF \modmult_1/zreg_reg[595]  ( .D(\modmult_1/N598 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][595] ) );
  DFF \modmult_1/zreg_reg[594]  ( .D(\modmult_1/N597 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][594] ) );
  DFF \modmult_1/zreg_reg[593]  ( .D(\modmult_1/N596 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][593] ) );
  DFF \modmult_1/zreg_reg[592]  ( .D(\modmult_1/N595 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][592] ) );
  DFF \modmult_1/zreg_reg[591]  ( .D(\modmult_1/N594 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][591] ) );
  DFF \modmult_1/zreg_reg[590]  ( .D(\modmult_1/N593 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][590] ) );
  DFF \modmult_1/zreg_reg[589]  ( .D(\modmult_1/N592 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][589] ) );
  DFF \modmult_1/zreg_reg[588]  ( .D(\modmult_1/N591 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][588] ) );
  DFF \modmult_1/zreg_reg[587]  ( .D(\modmult_1/N590 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][587] ) );
  DFF \modmult_1/zreg_reg[586]  ( .D(\modmult_1/N589 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][586] ) );
  DFF \modmult_1/zreg_reg[585]  ( .D(\modmult_1/N588 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][585] ) );
  DFF \modmult_1/zreg_reg[584]  ( .D(\modmult_1/N587 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][584] ) );
  DFF \modmult_1/zreg_reg[583]  ( .D(\modmult_1/N586 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][583] ) );
  DFF \modmult_1/zreg_reg[582]  ( .D(\modmult_1/N585 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][582] ) );
  DFF \modmult_1/zreg_reg[581]  ( .D(\modmult_1/N584 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][581] ) );
  DFF \modmult_1/zreg_reg[580]  ( .D(\modmult_1/N583 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][580] ) );
  DFF \modmult_1/zreg_reg[579]  ( .D(\modmult_1/N582 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][579] ) );
  DFF \modmult_1/zreg_reg[578]  ( .D(\modmult_1/N581 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][578] ) );
  DFF \modmult_1/zreg_reg[577]  ( .D(\modmult_1/N580 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][577] ) );
  DFF \modmult_1/zreg_reg[576]  ( .D(\modmult_1/N579 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][576] ) );
  DFF \modmult_1/zreg_reg[575]  ( .D(\modmult_1/N578 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][575] ) );
  DFF \modmult_1/zreg_reg[574]  ( .D(\modmult_1/N577 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][574] ) );
  DFF \modmult_1/zreg_reg[573]  ( .D(\modmult_1/N576 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][573] ) );
  DFF \modmult_1/zreg_reg[572]  ( .D(\modmult_1/N575 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][572] ) );
  DFF \modmult_1/zreg_reg[571]  ( .D(\modmult_1/N574 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][571] ) );
  DFF \modmult_1/zreg_reg[570]  ( .D(\modmult_1/N573 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][570] ) );
  DFF \modmult_1/zreg_reg[569]  ( .D(\modmult_1/N572 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][569] ) );
  DFF \modmult_1/zreg_reg[568]  ( .D(\modmult_1/N571 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][568] ) );
  DFF \modmult_1/zreg_reg[567]  ( .D(\modmult_1/N570 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][567] ) );
  DFF \modmult_1/zreg_reg[566]  ( .D(\modmult_1/N569 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][566] ) );
  DFF \modmult_1/zreg_reg[565]  ( .D(\modmult_1/N568 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][565] ) );
  DFF \modmult_1/zreg_reg[564]  ( .D(\modmult_1/N567 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][564] ) );
  DFF \modmult_1/zreg_reg[563]  ( .D(\modmult_1/N566 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][563] ) );
  DFF \modmult_1/zreg_reg[562]  ( .D(\modmult_1/N565 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][562] ) );
  DFF \modmult_1/zreg_reg[561]  ( .D(\modmult_1/N564 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][561] ) );
  DFF \modmult_1/zreg_reg[560]  ( .D(\modmult_1/N563 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][560] ) );
  DFF \modmult_1/zreg_reg[559]  ( .D(\modmult_1/N562 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][559] ) );
  DFF \modmult_1/zreg_reg[558]  ( .D(\modmult_1/N561 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][558] ) );
  DFF \modmult_1/zreg_reg[557]  ( .D(\modmult_1/N560 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][557] ) );
  DFF \modmult_1/zreg_reg[556]  ( .D(\modmult_1/N559 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][556] ) );
  DFF \modmult_1/zreg_reg[555]  ( .D(\modmult_1/N558 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][555] ) );
  DFF \modmult_1/zreg_reg[554]  ( .D(\modmult_1/N557 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][554] ) );
  DFF \modmult_1/zreg_reg[553]  ( .D(\modmult_1/N556 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][553] ) );
  DFF \modmult_1/zreg_reg[552]  ( .D(\modmult_1/N555 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][552] ) );
  DFF \modmult_1/zreg_reg[551]  ( .D(\modmult_1/N554 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][551] ) );
  DFF \modmult_1/zreg_reg[550]  ( .D(\modmult_1/N553 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][550] ) );
  DFF \modmult_1/zreg_reg[549]  ( .D(\modmult_1/N552 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][549] ) );
  DFF \modmult_1/zreg_reg[548]  ( .D(\modmult_1/N551 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][548] ) );
  DFF \modmult_1/zreg_reg[547]  ( .D(\modmult_1/N550 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][547] ) );
  DFF \modmult_1/zreg_reg[546]  ( .D(\modmult_1/N549 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][546] ) );
  DFF \modmult_1/zreg_reg[545]  ( .D(\modmult_1/N548 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][545] ) );
  DFF \modmult_1/zreg_reg[544]  ( .D(\modmult_1/N547 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][544] ) );
  DFF \modmult_1/zreg_reg[543]  ( .D(\modmult_1/N546 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][543] ) );
  DFF \modmult_1/zreg_reg[542]  ( .D(\modmult_1/N545 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][542] ) );
  DFF \modmult_1/zreg_reg[541]  ( .D(\modmult_1/N544 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][541] ) );
  DFF \modmult_1/zreg_reg[540]  ( .D(\modmult_1/N543 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][540] ) );
  DFF \modmult_1/zreg_reg[539]  ( .D(\modmult_1/N542 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][539] ) );
  DFF \modmult_1/zreg_reg[538]  ( .D(\modmult_1/N541 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][538] ) );
  DFF \modmult_1/zreg_reg[537]  ( .D(\modmult_1/N540 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][537] ) );
  DFF \modmult_1/zreg_reg[536]  ( .D(\modmult_1/N539 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][536] ) );
  DFF \modmult_1/zreg_reg[535]  ( .D(\modmult_1/N538 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][535] ) );
  DFF \modmult_1/zreg_reg[534]  ( .D(\modmult_1/N537 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][534] ) );
  DFF \modmult_1/zreg_reg[533]  ( .D(\modmult_1/N536 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][533] ) );
  DFF \modmult_1/zreg_reg[532]  ( .D(\modmult_1/N535 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][532] ) );
  DFF \modmult_1/zreg_reg[531]  ( .D(\modmult_1/N534 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][531] ) );
  DFF \modmult_1/zreg_reg[530]  ( .D(\modmult_1/N533 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][530] ) );
  DFF \modmult_1/zreg_reg[529]  ( .D(\modmult_1/N532 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][529] ) );
  DFF \modmult_1/zreg_reg[528]  ( .D(\modmult_1/N531 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][528] ) );
  DFF \modmult_1/zreg_reg[527]  ( .D(\modmult_1/N530 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][527] ) );
  DFF \modmult_1/zreg_reg[526]  ( .D(\modmult_1/N529 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][526] ) );
  DFF \modmult_1/zreg_reg[525]  ( .D(\modmult_1/N528 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][525] ) );
  DFF \modmult_1/zreg_reg[524]  ( .D(\modmult_1/N527 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][524] ) );
  DFF \modmult_1/zreg_reg[523]  ( .D(\modmult_1/N526 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][523] ) );
  DFF \modmult_1/zreg_reg[522]  ( .D(\modmult_1/N525 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][522] ) );
  DFF \modmult_1/zreg_reg[521]  ( .D(\modmult_1/N524 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][521] ) );
  DFF \modmult_1/zreg_reg[520]  ( .D(\modmult_1/N523 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][520] ) );
  DFF \modmult_1/zreg_reg[519]  ( .D(\modmult_1/N522 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][519] ) );
  DFF \modmult_1/zreg_reg[518]  ( .D(\modmult_1/N521 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][518] ) );
  DFF \modmult_1/zreg_reg[517]  ( .D(\modmult_1/N520 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][517] ) );
  DFF \modmult_1/zreg_reg[516]  ( .D(\modmult_1/N519 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][516] ) );
  DFF \modmult_1/zreg_reg[515]  ( .D(\modmult_1/N518 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][515] ) );
  DFF \modmult_1/zreg_reg[514]  ( .D(\modmult_1/N517 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][514] ) );
  DFF \modmult_1/zreg_reg[513]  ( .D(\modmult_1/N516 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][513] ) );
  DFF \modmult_1/zreg_reg[512]  ( .D(\modmult_1/N515 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][512] ) );
  DFF \modmult_1/zreg_reg[511]  ( .D(\modmult_1/N514 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][511] ) );
  DFF \modmult_1/zreg_reg[510]  ( .D(\modmult_1/N513 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][510] ) );
  DFF \modmult_1/zreg_reg[509]  ( .D(\modmult_1/N512 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][509] ) );
  DFF \modmult_1/zreg_reg[508]  ( .D(\modmult_1/N511 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][508] ) );
  DFF \modmult_1/zreg_reg[507]  ( .D(\modmult_1/N510 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][507] ) );
  DFF \modmult_1/zreg_reg[506]  ( .D(\modmult_1/N509 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][506] ) );
  DFF \modmult_1/zreg_reg[505]  ( .D(\modmult_1/N508 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][505] ) );
  DFF \modmult_1/zreg_reg[504]  ( .D(\modmult_1/N507 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][504] ) );
  DFF \modmult_1/zreg_reg[503]  ( .D(\modmult_1/N506 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][503] ) );
  DFF \modmult_1/zreg_reg[502]  ( .D(\modmult_1/N505 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][502] ) );
  DFF \modmult_1/zreg_reg[501]  ( .D(\modmult_1/N504 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][501] ) );
  DFF \modmult_1/zreg_reg[500]  ( .D(\modmult_1/N503 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][500] ) );
  DFF \modmult_1/zreg_reg[499]  ( .D(\modmult_1/N502 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][499] ) );
  DFF \modmult_1/zreg_reg[498]  ( .D(\modmult_1/N501 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][498] ) );
  DFF \modmult_1/zreg_reg[497]  ( .D(\modmult_1/N500 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][497] ) );
  DFF \modmult_1/zreg_reg[496]  ( .D(\modmult_1/N499 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][496] ) );
  DFF \modmult_1/zreg_reg[495]  ( .D(\modmult_1/N498 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][495] ) );
  DFF \modmult_1/zreg_reg[494]  ( .D(\modmult_1/N497 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][494] ) );
  DFF \modmult_1/zreg_reg[493]  ( .D(\modmult_1/N496 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][493] ) );
  DFF \modmult_1/zreg_reg[492]  ( .D(\modmult_1/N495 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][492] ) );
  DFF \modmult_1/zreg_reg[491]  ( .D(\modmult_1/N494 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][491] ) );
  DFF \modmult_1/zreg_reg[490]  ( .D(\modmult_1/N493 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][490] ) );
  DFF \modmult_1/zreg_reg[489]  ( .D(\modmult_1/N492 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][489] ) );
  DFF \modmult_1/zreg_reg[488]  ( .D(\modmult_1/N491 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][488] ) );
  DFF \modmult_1/zreg_reg[487]  ( .D(\modmult_1/N490 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][487] ) );
  DFF \modmult_1/zreg_reg[486]  ( .D(\modmult_1/N489 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][486] ) );
  DFF \modmult_1/zreg_reg[485]  ( .D(\modmult_1/N488 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][485] ) );
  DFF \modmult_1/zreg_reg[484]  ( .D(\modmult_1/N487 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][484] ) );
  DFF \modmult_1/zreg_reg[483]  ( .D(\modmult_1/N486 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][483] ) );
  DFF \modmult_1/zreg_reg[482]  ( .D(\modmult_1/N485 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][482] ) );
  DFF \modmult_1/zreg_reg[481]  ( .D(\modmult_1/N484 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][481] ) );
  DFF \modmult_1/zreg_reg[480]  ( .D(\modmult_1/N483 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][480] ) );
  DFF \modmult_1/zreg_reg[479]  ( .D(\modmult_1/N482 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][479] ) );
  DFF \modmult_1/zreg_reg[478]  ( .D(\modmult_1/N481 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][478] ) );
  DFF \modmult_1/zreg_reg[477]  ( .D(\modmult_1/N480 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][477] ) );
  DFF \modmult_1/zreg_reg[476]  ( .D(\modmult_1/N479 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][476] ) );
  DFF \modmult_1/zreg_reg[475]  ( .D(\modmult_1/N478 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][475] ) );
  DFF \modmult_1/zreg_reg[474]  ( .D(\modmult_1/N477 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][474] ) );
  DFF \modmult_1/zreg_reg[473]  ( .D(\modmult_1/N476 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][473] ) );
  DFF \modmult_1/zreg_reg[472]  ( .D(\modmult_1/N475 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][472] ) );
  DFF \modmult_1/zreg_reg[471]  ( .D(\modmult_1/N474 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][471] ) );
  DFF \modmult_1/zreg_reg[470]  ( .D(\modmult_1/N473 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][470] ) );
  DFF \modmult_1/zreg_reg[469]  ( .D(\modmult_1/N472 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][469] ) );
  DFF \modmult_1/zreg_reg[468]  ( .D(\modmult_1/N471 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][468] ) );
  DFF \modmult_1/zreg_reg[467]  ( .D(\modmult_1/N470 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][467] ) );
  DFF \modmult_1/zreg_reg[466]  ( .D(\modmult_1/N469 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][466] ) );
  DFF \modmult_1/zreg_reg[465]  ( .D(\modmult_1/N468 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][465] ) );
  DFF \modmult_1/zreg_reg[464]  ( .D(\modmult_1/N467 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][464] ) );
  DFF \modmult_1/zreg_reg[463]  ( .D(\modmult_1/N466 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][463] ) );
  DFF \modmult_1/zreg_reg[462]  ( .D(\modmult_1/N465 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][462] ) );
  DFF \modmult_1/zreg_reg[461]  ( .D(\modmult_1/N464 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][461] ) );
  DFF \modmult_1/zreg_reg[460]  ( .D(\modmult_1/N463 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][460] ) );
  DFF \modmult_1/zreg_reg[459]  ( .D(\modmult_1/N462 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][459] ) );
  DFF \modmult_1/zreg_reg[458]  ( .D(\modmult_1/N461 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][458] ) );
  DFF \modmult_1/zreg_reg[457]  ( .D(\modmult_1/N460 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][457] ) );
  DFF \modmult_1/zreg_reg[456]  ( .D(\modmult_1/N459 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][456] ) );
  DFF \modmult_1/zreg_reg[455]  ( .D(\modmult_1/N458 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][455] ) );
  DFF \modmult_1/zreg_reg[454]  ( .D(\modmult_1/N457 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][454] ) );
  DFF \modmult_1/zreg_reg[453]  ( .D(\modmult_1/N456 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][453] ) );
  DFF \modmult_1/zreg_reg[452]  ( .D(\modmult_1/N455 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][452] ) );
  DFF \modmult_1/zreg_reg[451]  ( .D(\modmult_1/N454 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][451] ) );
  DFF \modmult_1/zreg_reg[450]  ( .D(\modmult_1/N453 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][450] ) );
  DFF \modmult_1/zreg_reg[449]  ( .D(\modmult_1/N452 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][449] ) );
  DFF \modmult_1/zreg_reg[448]  ( .D(\modmult_1/N451 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][448] ) );
  DFF \modmult_1/zreg_reg[447]  ( .D(\modmult_1/N450 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][447] ) );
  DFF \modmult_1/zreg_reg[446]  ( .D(\modmult_1/N449 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][446] ) );
  DFF \modmult_1/zreg_reg[445]  ( .D(\modmult_1/N448 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][445] ) );
  DFF \modmult_1/zreg_reg[444]  ( .D(\modmult_1/N447 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][444] ) );
  DFF \modmult_1/zreg_reg[443]  ( .D(\modmult_1/N446 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][443] ) );
  DFF \modmult_1/zreg_reg[442]  ( .D(\modmult_1/N445 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][442] ) );
  DFF \modmult_1/zreg_reg[441]  ( .D(\modmult_1/N444 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][441] ) );
  DFF \modmult_1/zreg_reg[440]  ( .D(\modmult_1/N443 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][440] ) );
  DFF \modmult_1/zreg_reg[439]  ( .D(\modmult_1/N442 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][439] ) );
  DFF \modmult_1/zreg_reg[438]  ( .D(\modmult_1/N441 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][438] ) );
  DFF \modmult_1/zreg_reg[437]  ( .D(\modmult_1/N440 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][437] ) );
  DFF \modmult_1/zreg_reg[436]  ( .D(\modmult_1/N439 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][436] ) );
  DFF \modmult_1/zreg_reg[435]  ( .D(\modmult_1/N438 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][435] ) );
  DFF \modmult_1/zreg_reg[434]  ( .D(\modmult_1/N437 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][434] ) );
  DFF \modmult_1/zreg_reg[433]  ( .D(\modmult_1/N436 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][433] ) );
  DFF \modmult_1/zreg_reg[432]  ( .D(\modmult_1/N435 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][432] ) );
  DFF \modmult_1/zreg_reg[431]  ( .D(\modmult_1/N434 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][431] ) );
  DFF \modmult_1/zreg_reg[430]  ( .D(\modmult_1/N433 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][430] ) );
  DFF \modmult_1/zreg_reg[429]  ( .D(\modmult_1/N432 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][429] ) );
  DFF \modmult_1/zreg_reg[428]  ( .D(\modmult_1/N431 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][428] ) );
  DFF \modmult_1/zreg_reg[427]  ( .D(\modmult_1/N430 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][427] ) );
  DFF \modmult_1/zreg_reg[426]  ( .D(\modmult_1/N429 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][426] ) );
  DFF \modmult_1/zreg_reg[425]  ( .D(\modmult_1/N428 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][425] ) );
  DFF \modmult_1/zreg_reg[424]  ( .D(\modmult_1/N427 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][424] ) );
  DFF \modmult_1/zreg_reg[423]  ( .D(\modmult_1/N426 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][423] ) );
  DFF \modmult_1/zreg_reg[422]  ( .D(\modmult_1/N425 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][422] ) );
  DFF \modmult_1/zreg_reg[421]  ( .D(\modmult_1/N424 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][421] ) );
  DFF \modmult_1/zreg_reg[420]  ( .D(\modmult_1/N423 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][420] ) );
  DFF \modmult_1/zreg_reg[419]  ( .D(\modmult_1/N422 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][419] ) );
  DFF \modmult_1/zreg_reg[418]  ( .D(\modmult_1/N421 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][418] ) );
  DFF \modmult_1/zreg_reg[417]  ( .D(\modmult_1/N420 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][417] ) );
  DFF \modmult_1/zreg_reg[416]  ( .D(\modmult_1/N419 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][416] ) );
  DFF \modmult_1/zreg_reg[415]  ( .D(\modmult_1/N418 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][415] ) );
  DFF \modmult_1/zreg_reg[414]  ( .D(\modmult_1/N417 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][414] ) );
  DFF \modmult_1/zreg_reg[413]  ( .D(\modmult_1/N416 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][413] ) );
  DFF \modmult_1/zreg_reg[412]  ( .D(\modmult_1/N415 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][412] ) );
  DFF \modmult_1/zreg_reg[411]  ( .D(\modmult_1/N414 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][411] ) );
  DFF \modmult_1/zreg_reg[410]  ( .D(\modmult_1/N413 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][410] ) );
  DFF \modmult_1/zreg_reg[409]  ( .D(\modmult_1/N412 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][409] ) );
  DFF \modmult_1/zreg_reg[408]  ( .D(\modmult_1/N411 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][408] ) );
  DFF \modmult_1/zreg_reg[407]  ( .D(\modmult_1/N410 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][407] ) );
  DFF \modmult_1/zreg_reg[406]  ( .D(\modmult_1/N409 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][406] ) );
  DFF \modmult_1/zreg_reg[405]  ( .D(\modmult_1/N408 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][405] ) );
  DFF \modmult_1/zreg_reg[404]  ( .D(\modmult_1/N407 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][404] ) );
  DFF \modmult_1/zreg_reg[403]  ( .D(\modmult_1/N406 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][403] ) );
  DFF \modmult_1/zreg_reg[402]  ( .D(\modmult_1/N405 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][402] ) );
  DFF \modmult_1/zreg_reg[401]  ( .D(\modmult_1/N404 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][401] ) );
  DFF \modmult_1/zreg_reg[400]  ( .D(\modmult_1/N403 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][400] ) );
  DFF \modmult_1/zreg_reg[399]  ( .D(\modmult_1/N402 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][399] ) );
  DFF \modmult_1/zreg_reg[398]  ( .D(\modmult_1/N401 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][398] ) );
  DFF \modmult_1/zreg_reg[397]  ( .D(\modmult_1/N400 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][397] ) );
  DFF \modmult_1/zreg_reg[396]  ( .D(\modmult_1/N399 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][396] ) );
  DFF \modmult_1/zreg_reg[395]  ( .D(\modmult_1/N398 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][395] ) );
  DFF \modmult_1/zreg_reg[394]  ( .D(\modmult_1/N397 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][394] ) );
  DFF \modmult_1/zreg_reg[393]  ( .D(\modmult_1/N396 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][393] ) );
  DFF \modmult_1/zreg_reg[392]  ( .D(\modmult_1/N395 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][392] ) );
  DFF \modmult_1/zreg_reg[391]  ( .D(\modmult_1/N394 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][391] ) );
  DFF \modmult_1/zreg_reg[390]  ( .D(\modmult_1/N393 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][390] ) );
  DFF \modmult_1/zreg_reg[389]  ( .D(\modmult_1/N392 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][389] ) );
  DFF \modmult_1/zreg_reg[388]  ( .D(\modmult_1/N391 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][388] ) );
  DFF \modmult_1/zreg_reg[387]  ( .D(\modmult_1/N390 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][387] ) );
  DFF \modmult_1/zreg_reg[386]  ( .D(\modmult_1/N389 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][386] ) );
  DFF \modmult_1/zreg_reg[385]  ( .D(\modmult_1/N388 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][385] ) );
  DFF \modmult_1/zreg_reg[384]  ( .D(\modmult_1/N387 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][384] ) );
  DFF \modmult_1/zreg_reg[383]  ( .D(\modmult_1/N386 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][383] ) );
  DFF \modmult_1/zreg_reg[382]  ( .D(\modmult_1/N385 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][382] ) );
  DFF \modmult_1/zreg_reg[381]  ( .D(\modmult_1/N384 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][381] ) );
  DFF \modmult_1/zreg_reg[380]  ( .D(\modmult_1/N383 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][380] ) );
  DFF \modmult_1/zreg_reg[379]  ( .D(\modmult_1/N382 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][379] ) );
  DFF \modmult_1/zreg_reg[378]  ( .D(\modmult_1/N381 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][378] ) );
  DFF \modmult_1/zreg_reg[377]  ( .D(\modmult_1/N380 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][377] ) );
  DFF \modmult_1/zreg_reg[376]  ( .D(\modmult_1/N379 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][376] ) );
  DFF \modmult_1/zreg_reg[375]  ( .D(\modmult_1/N378 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][375] ) );
  DFF \modmult_1/zreg_reg[374]  ( .D(\modmult_1/N377 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][374] ) );
  DFF \modmult_1/zreg_reg[373]  ( .D(\modmult_1/N376 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][373] ) );
  DFF \modmult_1/zreg_reg[372]  ( .D(\modmult_1/N375 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][372] ) );
  DFF \modmult_1/zreg_reg[371]  ( .D(\modmult_1/N374 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][371] ) );
  DFF \modmult_1/zreg_reg[370]  ( .D(\modmult_1/N373 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][370] ) );
  DFF \modmult_1/zreg_reg[369]  ( .D(\modmult_1/N372 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][369] ) );
  DFF \modmult_1/zreg_reg[368]  ( .D(\modmult_1/N371 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][368] ) );
  DFF \modmult_1/zreg_reg[367]  ( .D(\modmult_1/N370 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][367] ) );
  DFF \modmult_1/zreg_reg[366]  ( .D(\modmult_1/N369 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][366] ) );
  DFF \modmult_1/zreg_reg[365]  ( .D(\modmult_1/N368 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][365] ) );
  DFF \modmult_1/zreg_reg[364]  ( .D(\modmult_1/N367 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][364] ) );
  DFF \modmult_1/zreg_reg[363]  ( .D(\modmult_1/N366 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][363] ) );
  DFF \modmult_1/zreg_reg[362]  ( .D(\modmult_1/N365 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][362] ) );
  DFF \modmult_1/zreg_reg[361]  ( .D(\modmult_1/N364 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][361] ) );
  DFF \modmult_1/zreg_reg[360]  ( .D(\modmult_1/N363 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][360] ) );
  DFF \modmult_1/zreg_reg[359]  ( .D(\modmult_1/N362 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][359] ) );
  DFF \modmult_1/zreg_reg[358]  ( .D(\modmult_1/N361 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][358] ) );
  DFF \modmult_1/zreg_reg[357]  ( .D(\modmult_1/N360 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][357] ) );
  DFF \modmult_1/zreg_reg[356]  ( .D(\modmult_1/N359 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][356] ) );
  DFF \modmult_1/zreg_reg[355]  ( .D(\modmult_1/N358 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][355] ) );
  DFF \modmult_1/zreg_reg[354]  ( .D(\modmult_1/N357 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][354] ) );
  DFF \modmult_1/zreg_reg[353]  ( .D(\modmult_1/N356 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][353] ) );
  DFF \modmult_1/zreg_reg[352]  ( .D(\modmult_1/N355 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][352] ) );
  DFF \modmult_1/zreg_reg[351]  ( .D(\modmult_1/N354 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][351] ) );
  DFF \modmult_1/zreg_reg[350]  ( .D(\modmult_1/N353 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][350] ) );
  DFF \modmult_1/zreg_reg[349]  ( .D(\modmult_1/N352 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][349] ) );
  DFF \modmult_1/zreg_reg[348]  ( .D(\modmult_1/N351 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][348] ) );
  DFF \modmult_1/zreg_reg[347]  ( .D(\modmult_1/N350 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][347] ) );
  DFF \modmult_1/zreg_reg[346]  ( .D(\modmult_1/N349 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][346] ) );
  DFF \modmult_1/zreg_reg[345]  ( .D(\modmult_1/N348 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][345] ) );
  DFF \modmult_1/zreg_reg[344]  ( .D(\modmult_1/N347 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][344] ) );
  DFF \modmult_1/zreg_reg[343]  ( .D(\modmult_1/N346 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][343] ) );
  DFF \modmult_1/zreg_reg[342]  ( .D(\modmult_1/N345 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][342] ) );
  DFF \modmult_1/zreg_reg[341]  ( .D(\modmult_1/N344 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][341] ) );
  DFF \modmult_1/zreg_reg[340]  ( .D(\modmult_1/N343 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][340] ) );
  DFF \modmult_1/zreg_reg[339]  ( .D(\modmult_1/N342 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][339] ) );
  DFF \modmult_1/zreg_reg[338]  ( .D(\modmult_1/N341 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][338] ) );
  DFF \modmult_1/zreg_reg[337]  ( .D(\modmult_1/N340 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][337] ) );
  DFF \modmult_1/zreg_reg[336]  ( .D(\modmult_1/N339 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][336] ) );
  DFF \modmult_1/zreg_reg[335]  ( .D(\modmult_1/N338 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][335] ) );
  DFF \modmult_1/zreg_reg[334]  ( .D(\modmult_1/N337 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][334] ) );
  DFF \modmult_1/zreg_reg[333]  ( .D(\modmult_1/N336 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][333] ) );
  DFF \modmult_1/zreg_reg[332]  ( .D(\modmult_1/N335 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][332] ) );
  DFF \modmult_1/zreg_reg[331]  ( .D(\modmult_1/N334 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][331] ) );
  DFF \modmult_1/zreg_reg[330]  ( .D(\modmult_1/N333 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][330] ) );
  DFF \modmult_1/zreg_reg[329]  ( .D(\modmult_1/N332 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][329] ) );
  DFF \modmult_1/zreg_reg[328]  ( .D(\modmult_1/N331 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][328] ) );
  DFF \modmult_1/zreg_reg[327]  ( .D(\modmult_1/N330 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][327] ) );
  DFF \modmult_1/zreg_reg[326]  ( .D(\modmult_1/N329 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][326] ) );
  DFF \modmult_1/zreg_reg[325]  ( .D(\modmult_1/N328 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][325] ) );
  DFF \modmult_1/zreg_reg[324]  ( .D(\modmult_1/N327 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][324] ) );
  DFF \modmult_1/zreg_reg[323]  ( .D(\modmult_1/N326 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][323] ) );
  DFF \modmult_1/zreg_reg[322]  ( .D(\modmult_1/N325 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][322] ) );
  DFF \modmult_1/zreg_reg[321]  ( .D(\modmult_1/N324 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][321] ) );
  DFF \modmult_1/zreg_reg[320]  ( .D(\modmult_1/N323 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][320] ) );
  DFF \modmult_1/zreg_reg[319]  ( .D(\modmult_1/N322 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][319] ) );
  DFF \modmult_1/zreg_reg[318]  ( .D(\modmult_1/N321 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][318] ) );
  DFF \modmult_1/zreg_reg[317]  ( .D(\modmult_1/N320 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][317] ) );
  DFF \modmult_1/zreg_reg[316]  ( .D(\modmult_1/N319 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][316] ) );
  DFF \modmult_1/zreg_reg[315]  ( .D(\modmult_1/N318 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][315] ) );
  DFF \modmult_1/zreg_reg[314]  ( .D(\modmult_1/N317 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][314] ) );
  DFF \modmult_1/zreg_reg[313]  ( .D(\modmult_1/N316 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][313] ) );
  DFF \modmult_1/zreg_reg[312]  ( .D(\modmult_1/N315 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][312] ) );
  DFF \modmult_1/zreg_reg[311]  ( .D(\modmult_1/N314 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][311] ) );
  DFF \modmult_1/zreg_reg[310]  ( .D(\modmult_1/N313 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][310] ) );
  DFF \modmult_1/zreg_reg[309]  ( .D(\modmult_1/N312 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][309] ) );
  DFF \modmult_1/zreg_reg[308]  ( .D(\modmult_1/N311 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][308] ) );
  DFF \modmult_1/zreg_reg[307]  ( .D(\modmult_1/N310 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][307] ) );
  DFF \modmult_1/zreg_reg[306]  ( .D(\modmult_1/N309 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][306] ) );
  DFF \modmult_1/zreg_reg[305]  ( .D(\modmult_1/N308 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][305] ) );
  DFF \modmult_1/zreg_reg[304]  ( .D(\modmult_1/N307 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][304] ) );
  DFF \modmult_1/zreg_reg[303]  ( .D(\modmult_1/N306 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][303] ) );
  DFF \modmult_1/zreg_reg[302]  ( .D(\modmult_1/N305 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][302] ) );
  DFF \modmult_1/zreg_reg[301]  ( .D(\modmult_1/N304 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][301] ) );
  DFF \modmult_1/zreg_reg[300]  ( .D(\modmult_1/N303 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][300] ) );
  DFF \modmult_1/zreg_reg[299]  ( .D(\modmult_1/N302 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][299] ) );
  DFF \modmult_1/zreg_reg[298]  ( .D(\modmult_1/N301 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][298] ) );
  DFF \modmult_1/zreg_reg[297]  ( .D(\modmult_1/N300 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][297] ) );
  DFF \modmult_1/zreg_reg[296]  ( .D(\modmult_1/N299 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][296] ) );
  DFF \modmult_1/zreg_reg[295]  ( .D(\modmult_1/N298 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][295] ) );
  DFF \modmult_1/zreg_reg[294]  ( .D(\modmult_1/N297 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][294] ) );
  DFF \modmult_1/zreg_reg[293]  ( .D(\modmult_1/N296 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][293] ) );
  DFF \modmult_1/zreg_reg[292]  ( .D(\modmult_1/N295 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][292] ) );
  DFF \modmult_1/zreg_reg[291]  ( .D(\modmult_1/N294 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][291] ) );
  DFF \modmult_1/zreg_reg[290]  ( .D(\modmult_1/N293 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][290] ) );
  DFF \modmult_1/zreg_reg[289]  ( .D(\modmult_1/N292 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][289] ) );
  DFF \modmult_1/zreg_reg[288]  ( .D(\modmult_1/N291 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][288] ) );
  DFF \modmult_1/zreg_reg[287]  ( .D(\modmult_1/N290 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][287] ) );
  DFF \modmult_1/zreg_reg[286]  ( .D(\modmult_1/N289 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][286] ) );
  DFF \modmult_1/zreg_reg[285]  ( .D(\modmult_1/N288 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][285] ) );
  DFF \modmult_1/zreg_reg[284]  ( .D(\modmult_1/N287 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][284] ) );
  DFF \modmult_1/zreg_reg[283]  ( .D(\modmult_1/N286 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][283] ) );
  DFF \modmult_1/zreg_reg[282]  ( .D(\modmult_1/N285 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][282] ) );
  DFF \modmult_1/zreg_reg[281]  ( .D(\modmult_1/N284 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][281] ) );
  DFF \modmult_1/zreg_reg[280]  ( .D(\modmult_1/N283 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][280] ) );
  DFF \modmult_1/zreg_reg[279]  ( .D(\modmult_1/N282 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][279] ) );
  DFF \modmult_1/zreg_reg[278]  ( .D(\modmult_1/N281 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][278] ) );
  DFF \modmult_1/zreg_reg[277]  ( .D(\modmult_1/N280 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][277] ) );
  DFF \modmult_1/zreg_reg[276]  ( .D(\modmult_1/N279 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][276] ) );
  DFF \modmult_1/zreg_reg[275]  ( .D(\modmult_1/N278 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][275] ) );
  DFF \modmult_1/zreg_reg[274]  ( .D(\modmult_1/N277 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][274] ) );
  DFF \modmult_1/zreg_reg[273]  ( .D(\modmult_1/N276 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][273] ) );
  DFF \modmult_1/zreg_reg[272]  ( .D(\modmult_1/N275 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][272] ) );
  DFF \modmult_1/zreg_reg[271]  ( .D(\modmult_1/N274 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][271] ) );
  DFF \modmult_1/zreg_reg[270]  ( .D(\modmult_1/N273 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][270] ) );
  DFF \modmult_1/zreg_reg[269]  ( .D(\modmult_1/N272 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][269] ) );
  DFF \modmult_1/zreg_reg[268]  ( .D(\modmult_1/N271 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][268] ) );
  DFF \modmult_1/zreg_reg[267]  ( .D(\modmult_1/N270 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][267] ) );
  DFF \modmult_1/zreg_reg[266]  ( .D(\modmult_1/N269 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][266] ) );
  DFF \modmult_1/zreg_reg[265]  ( .D(\modmult_1/N268 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][265] ) );
  DFF \modmult_1/zreg_reg[264]  ( .D(\modmult_1/N267 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][264] ) );
  DFF \modmult_1/zreg_reg[263]  ( .D(\modmult_1/N266 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][263] ) );
  DFF \modmult_1/zreg_reg[262]  ( .D(\modmult_1/N265 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][262] ) );
  DFF \modmult_1/zreg_reg[261]  ( .D(\modmult_1/N264 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][261] ) );
  DFF \modmult_1/zreg_reg[260]  ( .D(\modmult_1/N263 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][260] ) );
  DFF \modmult_1/zreg_reg[259]  ( .D(\modmult_1/N262 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][259] ) );
  DFF \modmult_1/zreg_reg[258]  ( .D(\modmult_1/N261 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][258] ) );
  DFF \modmult_1/zreg_reg[257]  ( .D(\modmult_1/N260 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][257] ) );
  DFF \modmult_1/zreg_reg[256]  ( .D(\modmult_1/N259 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][256] ) );
  DFF \modmult_1/zreg_reg[255]  ( .D(\modmult_1/N258 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][255] ) );
  DFF \modmult_1/zreg_reg[254]  ( .D(\modmult_1/N257 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][254] ) );
  DFF \modmult_1/zreg_reg[253]  ( .D(\modmult_1/N256 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][253] ) );
  DFF \modmult_1/zreg_reg[252]  ( .D(\modmult_1/N255 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][252] ) );
  DFF \modmult_1/zreg_reg[251]  ( .D(\modmult_1/N254 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][251] ) );
  DFF \modmult_1/zreg_reg[250]  ( .D(\modmult_1/N253 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][250] ) );
  DFF \modmult_1/zreg_reg[249]  ( .D(\modmult_1/N252 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][249] ) );
  DFF \modmult_1/zreg_reg[248]  ( .D(\modmult_1/N251 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][248] ) );
  DFF \modmult_1/zreg_reg[247]  ( .D(\modmult_1/N250 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][247] ) );
  DFF \modmult_1/zreg_reg[246]  ( .D(\modmult_1/N249 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][246] ) );
  DFF \modmult_1/zreg_reg[245]  ( .D(\modmult_1/N248 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][245] ) );
  DFF \modmult_1/zreg_reg[244]  ( .D(\modmult_1/N247 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][244] ) );
  DFF \modmult_1/zreg_reg[243]  ( .D(\modmult_1/N246 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][243] ) );
  DFF \modmult_1/zreg_reg[242]  ( .D(\modmult_1/N245 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][242] ) );
  DFF \modmult_1/zreg_reg[241]  ( .D(\modmult_1/N244 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][241] ) );
  DFF \modmult_1/zreg_reg[240]  ( .D(\modmult_1/N243 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][240] ) );
  DFF \modmult_1/zreg_reg[239]  ( .D(\modmult_1/N242 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][239] ) );
  DFF \modmult_1/zreg_reg[238]  ( .D(\modmult_1/N241 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][238] ) );
  DFF \modmult_1/zreg_reg[237]  ( .D(\modmult_1/N240 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][237] ) );
  DFF \modmult_1/zreg_reg[236]  ( .D(\modmult_1/N239 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][236] ) );
  DFF \modmult_1/zreg_reg[235]  ( .D(\modmult_1/N238 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][235] ) );
  DFF \modmult_1/zreg_reg[234]  ( .D(\modmult_1/N237 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][234] ) );
  DFF \modmult_1/zreg_reg[233]  ( .D(\modmult_1/N236 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][233] ) );
  DFF \modmult_1/zreg_reg[232]  ( .D(\modmult_1/N235 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][232] ) );
  DFF \modmult_1/zreg_reg[231]  ( .D(\modmult_1/N234 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][231] ) );
  DFF \modmult_1/zreg_reg[230]  ( .D(\modmult_1/N233 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][230] ) );
  DFF \modmult_1/zreg_reg[229]  ( .D(\modmult_1/N232 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][229] ) );
  DFF \modmult_1/zreg_reg[228]  ( .D(\modmult_1/N231 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][228] ) );
  DFF \modmult_1/zreg_reg[227]  ( .D(\modmult_1/N230 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][227] ) );
  DFF \modmult_1/zreg_reg[226]  ( .D(\modmult_1/N229 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][226] ) );
  DFF \modmult_1/zreg_reg[225]  ( .D(\modmult_1/N228 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][225] ) );
  DFF \modmult_1/zreg_reg[224]  ( .D(\modmult_1/N227 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][224] ) );
  DFF \modmult_1/zreg_reg[223]  ( .D(\modmult_1/N226 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][223] ) );
  DFF \modmult_1/zreg_reg[222]  ( .D(\modmult_1/N225 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][222] ) );
  DFF \modmult_1/zreg_reg[221]  ( .D(\modmult_1/N224 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][221] ) );
  DFF \modmult_1/zreg_reg[220]  ( .D(\modmult_1/N223 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][220] ) );
  DFF \modmult_1/zreg_reg[219]  ( .D(\modmult_1/N222 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][219] ) );
  DFF \modmult_1/zreg_reg[218]  ( .D(\modmult_1/N221 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][218] ) );
  DFF \modmult_1/zreg_reg[217]  ( .D(\modmult_1/N220 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][217] ) );
  DFF \modmult_1/zreg_reg[216]  ( .D(\modmult_1/N219 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][216] ) );
  DFF \modmult_1/zreg_reg[215]  ( .D(\modmult_1/N218 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][215] ) );
  DFF \modmult_1/zreg_reg[214]  ( .D(\modmult_1/N217 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][214] ) );
  DFF \modmult_1/zreg_reg[213]  ( .D(\modmult_1/N216 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][213] ) );
  DFF \modmult_1/zreg_reg[212]  ( .D(\modmult_1/N215 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][212] ) );
  DFF \modmult_1/zreg_reg[211]  ( .D(\modmult_1/N214 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][211] ) );
  DFF \modmult_1/zreg_reg[210]  ( .D(\modmult_1/N213 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][210] ) );
  DFF \modmult_1/zreg_reg[209]  ( .D(\modmult_1/N212 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][209] ) );
  DFF \modmult_1/zreg_reg[208]  ( .D(\modmult_1/N211 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][208] ) );
  DFF \modmult_1/zreg_reg[207]  ( .D(\modmult_1/N210 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][207] ) );
  DFF \modmult_1/zreg_reg[206]  ( .D(\modmult_1/N209 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][206] ) );
  DFF \modmult_1/zreg_reg[205]  ( .D(\modmult_1/N208 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][205] ) );
  DFF \modmult_1/zreg_reg[204]  ( .D(\modmult_1/N207 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][204] ) );
  DFF \modmult_1/zreg_reg[203]  ( .D(\modmult_1/N206 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][203] ) );
  DFF \modmult_1/zreg_reg[202]  ( .D(\modmult_1/N205 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][202] ) );
  DFF \modmult_1/zreg_reg[201]  ( .D(\modmult_1/N204 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][201] ) );
  DFF \modmult_1/zreg_reg[200]  ( .D(\modmult_1/N203 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][200] ) );
  DFF \modmult_1/zreg_reg[199]  ( .D(\modmult_1/N202 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][199] ) );
  DFF \modmult_1/zreg_reg[198]  ( .D(\modmult_1/N201 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][198] ) );
  DFF \modmult_1/zreg_reg[197]  ( .D(\modmult_1/N200 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][197] ) );
  DFF \modmult_1/zreg_reg[196]  ( .D(\modmult_1/N199 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][196] ) );
  DFF \modmult_1/zreg_reg[195]  ( .D(\modmult_1/N198 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][195] ) );
  DFF \modmult_1/zreg_reg[194]  ( .D(\modmult_1/N197 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][194] ) );
  DFF \modmult_1/zreg_reg[193]  ( .D(\modmult_1/N196 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][193] ) );
  DFF \modmult_1/zreg_reg[192]  ( .D(\modmult_1/N195 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][192] ) );
  DFF \modmult_1/zreg_reg[191]  ( .D(\modmult_1/N194 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][191] ) );
  DFF \modmult_1/zreg_reg[190]  ( .D(\modmult_1/N193 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][190] ) );
  DFF \modmult_1/zreg_reg[189]  ( .D(\modmult_1/N192 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][189] ) );
  DFF \modmult_1/zreg_reg[188]  ( .D(\modmult_1/N191 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][188] ) );
  DFF \modmult_1/zreg_reg[187]  ( .D(\modmult_1/N190 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][187] ) );
  DFF \modmult_1/zreg_reg[186]  ( .D(\modmult_1/N189 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][186] ) );
  DFF \modmult_1/zreg_reg[185]  ( .D(\modmult_1/N188 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][185] ) );
  DFF \modmult_1/zreg_reg[184]  ( .D(\modmult_1/N187 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][184] ) );
  DFF \modmult_1/zreg_reg[183]  ( .D(\modmult_1/N186 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][183] ) );
  DFF \modmult_1/zreg_reg[182]  ( .D(\modmult_1/N185 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][182] ) );
  DFF \modmult_1/zreg_reg[181]  ( .D(\modmult_1/N184 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][181] ) );
  DFF \modmult_1/zreg_reg[180]  ( .D(\modmult_1/N183 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][180] ) );
  DFF \modmult_1/zreg_reg[179]  ( .D(\modmult_1/N182 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][179] ) );
  DFF \modmult_1/zreg_reg[178]  ( .D(\modmult_1/N181 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][178] ) );
  DFF \modmult_1/zreg_reg[177]  ( .D(\modmult_1/N180 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][177] ) );
  DFF \modmult_1/zreg_reg[176]  ( .D(\modmult_1/N179 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][176] ) );
  DFF \modmult_1/zreg_reg[175]  ( .D(\modmult_1/N178 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][175] ) );
  DFF \modmult_1/zreg_reg[174]  ( .D(\modmult_1/N177 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][174] ) );
  DFF \modmult_1/zreg_reg[173]  ( .D(\modmult_1/N176 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][173] ) );
  DFF \modmult_1/zreg_reg[172]  ( .D(\modmult_1/N175 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][172] ) );
  DFF \modmult_1/zreg_reg[171]  ( .D(\modmult_1/N174 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][171] ) );
  DFF \modmult_1/zreg_reg[170]  ( .D(\modmult_1/N173 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][170] ) );
  DFF \modmult_1/zreg_reg[169]  ( .D(\modmult_1/N172 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][169] ) );
  DFF \modmult_1/zreg_reg[168]  ( .D(\modmult_1/N171 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][168] ) );
  DFF \modmult_1/zreg_reg[167]  ( .D(\modmult_1/N170 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][167] ) );
  DFF \modmult_1/zreg_reg[166]  ( .D(\modmult_1/N169 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][166] ) );
  DFF \modmult_1/zreg_reg[165]  ( .D(\modmult_1/N168 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][165] ) );
  DFF \modmult_1/zreg_reg[164]  ( .D(\modmult_1/N167 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][164] ) );
  DFF \modmult_1/zreg_reg[163]  ( .D(\modmult_1/N166 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][163] ) );
  DFF \modmult_1/zreg_reg[162]  ( .D(\modmult_1/N165 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][162] ) );
  DFF \modmult_1/zreg_reg[161]  ( .D(\modmult_1/N164 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][161] ) );
  DFF \modmult_1/zreg_reg[160]  ( .D(\modmult_1/N163 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][160] ) );
  DFF \modmult_1/zreg_reg[159]  ( .D(\modmult_1/N162 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][159] ) );
  DFF \modmult_1/zreg_reg[158]  ( .D(\modmult_1/N161 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][158] ) );
  DFF \modmult_1/zreg_reg[157]  ( .D(\modmult_1/N160 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][157] ) );
  DFF \modmult_1/zreg_reg[156]  ( .D(\modmult_1/N159 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][156] ) );
  DFF \modmult_1/zreg_reg[155]  ( .D(\modmult_1/N158 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][155] ) );
  DFF \modmult_1/zreg_reg[154]  ( .D(\modmult_1/N157 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][154] ) );
  DFF \modmult_1/zreg_reg[153]  ( .D(\modmult_1/N156 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][153] ) );
  DFF \modmult_1/zreg_reg[152]  ( .D(\modmult_1/N155 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][152] ) );
  DFF \modmult_1/zreg_reg[151]  ( .D(\modmult_1/N154 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][151] ) );
  DFF \modmult_1/zreg_reg[150]  ( .D(\modmult_1/N153 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][150] ) );
  DFF \modmult_1/zreg_reg[149]  ( .D(\modmult_1/N152 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][149] ) );
  DFF \modmult_1/zreg_reg[148]  ( .D(\modmult_1/N151 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][148] ) );
  DFF \modmult_1/zreg_reg[147]  ( .D(\modmult_1/N150 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][147] ) );
  DFF \modmult_1/zreg_reg[146]  ( .D(\modmult_1/N149 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][146] ) );
  DFF \modmult_1/zreg_reg[145]  ( .D(\modmult_1/N148 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][145] ) );
  DFF \modmult_1/zreg_reg[144]  ( .D(\modmult_1/N147 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][144] ) );
  DFF \modmult_1/zreg_reg[143]  ( .D(\modmult_1/N146 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][143] ) );
  DFF \modmult_1/zreg_reg[142]  ( .D(\modmult_1/N145 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][142] ) );
  DFF \modmult_1/zreg_reg[141]  ( .D(\modmult_1/N144 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][141] ) );
  DFF \modmult_1/zreg_reg[140]  ( .D(\modmult_1/N143 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][140] ) );
  DFF \modmult_1/zreg_reg[139]  ( .D(\modmult_1/N142 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][139] ) );
  DFF \modmult_1/zreg_reg[138]  ( .D(\modmult_1/N141 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][138] ) );
  DFF \modmult_1/zreg_reg[137]  ( .D(\modmult_1/N140 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][137] ) );
  DFF \modmult_1/zreg_reg[136]  ( .D(\modmult_1/N139 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][136] ) );
  DFF \modmult_1/zreg_reg[135]  ( .D(\modmult_1/N138 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][135] ) );
  DFF \modmult_1/zreg_reg[134]  ( .D(\modmult_1/N137 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][134] ) );
  DFF \modmult_1/zreg_reg[133]  ( .D(\modmult_1/N136 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][133] ) );
  DFF \modmult_1/zreg_reg[132]  ( .D(\modmult_1/N135 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][132] ) );
  DFF \modmult_1/zreg_reg[131]  ( .D(\modmult_1/N134 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][131] ) );
  DFF \modmult_1/zreg_reg[130]  ( .D(\modmult_1/N133 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][130] ) );
  DFF \modmult_1/zreg_reg[129]  ( .D(\modmult_1/N132 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][129] ) );
  DFF \modmult_1/zreg_reg[128]  ( .D(\modmult_1/N131 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][128] ) );
  DFF \modmult_1/zreg_reg[127]  ( .D(\modmult_1/N130 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][127] ) );
  DFF \modmult_1/zreg_reg[126]  ( .D(\modmult_1/N129 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][126] ) );
  DFF \modmult_1/zreg_reg[125]  ( .D(\modmult_1/N128 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][125] ) );
  DFF \modmult_1/zreg_reg[124]  ( .D(\modmult_1/N127 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][124] ) );
  DFF \modmult_1/zreg_reg[123]  ( .D(\modmult_1/N126 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][123] ) );
  DFF \modmult_1/zreg_reg[122]  ( .D(\modmult_1/N125 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][122] ) );
  DFF \modmult_1/zreg_reg[121]  ( .D(\modmult_1/N124 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][121] ) );
  DFF \modmult_1/zreg_reg[120]  ( .D(\modmult_1/N123 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][120] ) );
  DFF \modmult_1/zreg_reg[119]  ( .D(\modmult_1/N122 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][119] ) );
  DFF \modmult_1/zreg_reg[118]  ( .D(\modmult_1/N121 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][118] ) );
  DFF \modmult_1/zreg_reg[117]  ( .D(\modmult_1/N120 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][117] ) );
  DFF \modmult_1/zreg_reg[116]  ( .D(\modmult_1/N119 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][116] ) );
  DFF \modmult_1/zreg_reg[115]  ( .D(\modmult_1/N118 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][115] ) );
  DFF \modmult_1/zreg_reg[114]  ( .D(\modmult_1/N117 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][114] ) );
  DFF \modmult_1/zreg_reg[113]  ( .D(\modmult_1/N116 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][113] ) );
  DFF \modmult_1/zreg_reg[112]  ( .D(\modmult_1/N115 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][112] ) );
  DFF \modmult_1/zreg_reg[111]  ( .D(\modmult_1/N114 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][111] ) );
  DFF \modmult_1/zreg_reg[110]  ( .D(\modmult_1/N113 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][110] ) );
  DFF \modmult_1/zreg_reg[109]  ( .D(\modmult_1/N112 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][109] ) );
  DFF \modmult_1/zreg_reg[108]  ( .D(\modmult_1/N111 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][108] ) );
  DFF \modmult_1/zreg_reg[107]  ( .D(\modmult_1/N110 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][107] ) );
  DFF \modmult_1/zreg_reg[106]  ( .D(\modmult_1/N109 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][106] ) );
  DFF \modmult_1/zreg_reg[105]  ( .D(\modmult_1/N108 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][105] ) );
  DFF \modmult_1/zreg_reg[104]  ( .D(\modmult_1/N107 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][104] ) );
  DFF \modmult_1/zreg_reg[103]  ( .D(\modmult_1/N106 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][103] ) );
  DFF \modmult_1/zreg_reg[102]  ( .D(\modmult_1/N105 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][102] ) );
  DFF \modmult_1/zreg_reg[101]  ( .D(\modmult_1/N104 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][101] ) );
  DFF \modmult_1/zreg_reg[100]  ( .D(\modmult_1/N103 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][100] ) );
  DFF \modmult_1/zreg_reg[99]  ( .D(\modmult_1/N102 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][99] ) );
  DFF \modmult_1/zreg_reg[98]  ( .D(\modmult_1/N101 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][98] ) );
  DFF \modmult_1/zreg_reg[97]  ( .D(\modmult_1/N100 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][97] ) );
  DFF \modmult_1/zreg_reg[96]  ( .D(\modmult_1/N99 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][96] ) );
  DFF \modmult_1/zreg_reg[95]  ( .D(\modmult_1/N98 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][95] ) );
  DFF \modmult_1/zreg_reg[94]  ( .D(\modmult_1/N97 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][94] ) );
  DFF \modmult_1/zreg_reg[93]  ( .D(\modmult_1/N96 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][93] ) );
  DFF \modmult_1/zreg_reg[92]  ( .D(\modmult_1/N95 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][92] ) );
  DFF \modmult_1/zreg_reg[91]  ( .D(\modmult_1/N94 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][91] ) );
  DFF \modmult_1/zreg_reg[90]  ( .D(\modmult_1/N93 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][90] ) );
  DFF \modmult_1/zreg_reg[89]  ( .D(\modmult_1/N92 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][89] ) );
  DFF \modmult_1/zreg_reg[88]  ( .D(\modmult_1/N91 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][88] ) );
  DFF \modmult_1/zreg_reg[87]  ( .D(\modmult_1/N90 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][87] ) );
  DFF \modmult_1/zreg_reg[86]  ( .D(\modmult_1/N89 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][86] ) );
  DFF \modmult_1/zreg_reg[85]  ( .D(\modmult_1/N88 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][85] ) );
  DFF \modmult_1/zreg_reg[84]  ( .D(\modmult_1/N87 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][84] ) );
  DFF \modmult_1/zreg_reg[83]  ( .D(\modmult_1/N86 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][83] ) );
  DFF \modmult_1/zreg_reg[82]  ( .D(\modmult_1/N85 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][82] ) );
  DFF \modmult_1/zreg_reg[81]  ( .D(\modmult_1/N84 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][81] ) );
  DFF \modmult_1/zreg_reg[80]  ( .D(\modmult_1/N83 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][80] ) );
  DFF \modmult_1/zreg_reg[79]  ( .D(\modmult_1/N82 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][79] ) );
  DFF \modmult_1/zreg_reg[78]  ( .D(\modmult_1/N81 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][78] ) );
  DFF \modmult_1/zreg_reg[77]  ( .D(\modmult_1/N80 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][77] ) );
  DFF \modmult_1/zreg_reg[76]  ( .D(\modmult_1/N79 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][76] ) );
  DFF \modmult_1/zreg_reg[75]  ( .D(\modmult_1/N78 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][75] ) );
  DFF \modmult_1/zreg_reg[74]  ( .D(\modmult_1/N77 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][74] ) );
  DFF \modmult_1/zreg_reg[73]  ( .D(\modmult_1/N76 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][73] ) );
  DFF \modmult_1/zreg_reg[72]  ( .D(\modmult_1/N75 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][72] ) );
  DFF \modmult_1/zreg_reg[71]  ( .D(\modmult_1/N74 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][71] ) );
  DFF \modmult_1/zreg_reg[70]  ( .D(\modmult_1/N73 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][70] ) );
  DFF \modmult_1/zreg_reg[69]  ( .D(\modmult_1/N72 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][69] ) );
  DFF \modmult_1/zreg_reg[68]  ( .D(\modmult_1/N71 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][68] ) );
  DFF \modmult_1/zreg_reg[67]  ( .D(\modmult_1/N70 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][67] ) );
  DFF \modmult_1/zreg_reg[66]  ( .D(\modmult_1/N69 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][66] ) );
  DFF \modmult_1/zreg_reg[65]  ( .D(\modmult_1/N68 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][65] ) );
  DFF \modmult_1/zreg_reg[64]  ( .D(\modmult_1/N67 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][64] ) );
  DFF \modmult_1/zreg_reg[63]  ( .D(\modmult_1/N66 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][63] ) );
  DFF \modmult_1/zreg_reg[62]  ( .D(\modmult_1/N65 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][62] ) );
  DFF \modmult_1/zreg_reg[61]  ( .D(\modmult_1/N64 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][61] ) );
  DFF \modmult_1/zreg_reg[60]  ( .D(\modmult_1/N63 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][60] ) );
  DFF \modmult_1/zreg_reg[59]  ( .D(\modmult_1/N62 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][59] ) );
  DFF \modmult_1/zreg_reg[58]  ( .D(\modmult_1/N61 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][58] ) );
  DFF \modmult_1/zreg_reg[57]  ( .D(\modmult_1/N60 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][57] ) );
  DFF \modmult_1/zreg_reg[56]  ( .D(\modmult_1/N59 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][56] ) );
  DFF \modmult_1/zreg_reg[55]  ( .D(\modmult_1/N58 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][55] ) );
  DFF \modmult_1/zreg_reg[54]  ( .D(\modmult_1/N57 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][54] ) );
  DFF \modmult_1/zreg_reg[53]  ( .D(\modmult_1/N56 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][53] ) );
  DFF \modmult_1/zreg_reg[52]  ( .D(\modmult_1/N55 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][52] ) );
  DFF \modmult_1/zreg_reg[51]  ( .D(\modmult_1/N54 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][51] ) );
  DFF \modmult_1/zreg_reg[50]  ( .D(\modmult_1/N53 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][50] ) );
  DFF \modmult_1/zreg_reg[49]  ( .D(\modmult_1/N52 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][49] ) );
  DFF \modmult_1/zreg_reg[48]  ( .D(\modmult_1/N51 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][48] ) );
  DFF \modmult_1/zreg_reg[47]  ( .D(\modmult_1/N50 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][47] ) );
  DFF \modmult_1/zreg_reg[46]  ( .D(\modmult_1/N49 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][46] ) );
  DFF \modmult_1/zreg_reg[45]  ( .D(\modmult_1/N48 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][45] ) );
  DFF \modmult_1/zreg_reg[44]  ( .D(\modmult_1/N47 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][44] ) );
  DFF \modmult_1/zreg_reg[43]  ( .D(\modmult_1/N46 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][43] ) );
  DFF \modmult_1/zreg_reg[42]  ( .D(\modmult_1/N45 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][42] ) );
  DFF \modmult_1/zreg_reg[41]  ( .D(\modmult_1/N44 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][41] ) );
  DFF \modmult_1/zreg_reg[40]  ( .D(\modmult_1/N43 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][40] ) );
  DFF \modmult_1/zreg_reg[39]  ( .D(\modmult_1/N42 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][39] ) );
  DFF \modmult_1/zreg_reg[38]  ( .D(\modmult_1/N41 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][38] ) );
  DFF \modmult_1/zreg_reg[37]  ( .D(\modmult_1/N40 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][37] ) );
  DFF \modmult_1/zreg_reg[36]  ( .D(\modmult_1/N39 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][36] ) );
  DFF \modmult_1/zreg_reg[35]  ( .D(\modmult_1/N38 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][35] ) );
  DFF \modmult_1/zreg_reg[34]  ( .D(\modmult_1/N37 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][34] ) );
  DFF \modmult_1/zreg_reg[33]  ( .D(\modmult_1/N36 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][33] ) );
  DFF \modmult_1/zreg_reg[32]  ( .D(\modmult_1/N35 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][32] ) );
  DFF \modmult_1/zreg_reg[31]  ( .D(\modmult_1/N34 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][31] ) );
  DFF \modmult_1/zreg_reg[30]  ( .D(\modmult_1/N33 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][30] ) );
  DFF \modmult_1/zreg_reg[29]  ( .D(\modmult_1/N32 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][29] ) );
  DFF \modmult_1/zreg_reg[28]  ( .D(\modmult_1/N31 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][28] ) );
  DFF \modmult_1/zreg_reg[27]  ( .D(\modmult_1/N30 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][27] ) );
  DFF \modmult_1/zreg_reg[26]  ( .D(\modmult_1/N29 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][26] ) );
  DFF \modmult_1/zreg_reg[25]  ( .D(\modmult_1/N28 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][25] ) );
  DFF \modmult_1/zreg_reg[24]  ( .D(\modmult_1/N27 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][24] ) );
  DFF \modmult_1/zreg_reg[23]  ( .D(\modmult_1/N26 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][23] ) );
  DFF \modmult_1/zreg_reg[22]  ( .D(\modmult_1/N25 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][22] ) );
  DFF \modmult_1/zreg_reg[21]  ( .D(\modmult_1/N24 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][21] ) );
  DFF \modmult_1/zreg_reg[20]  ( .D(\modmult_1/N23 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][20] ) );
  DFF \modmult_1/zreg_reg[19]  ( .D(\modmult_1/N22 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][19] ) );
  DFF \modmult_1/zreg_reg[18]  ( .D(\modmult_1/N21 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][18] ) );
  DFF \modmult_1/zreg_reg[17]  ( .D(\modmult_1/N20 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][17] ) );
  DFF \modmult_1/zreg_reg[16]  ( .D(\modmult_1/N19 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][16] ) );
  DFF \modmult_1/zreg_reg[15]  ( .D(\modmult_1/N18 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][15] ) );
  DFF \modmult_1/zreg_reg[14]  ( .D(\modmult_1/N17 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][14] ) );
  DFF \modmult_1/zreg_reg[13]  ( .D(\modmult_1/N16 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][13] ) );
  DFF \modmult_1/zreg_reg[12]  ( .D(\modmult_1/N15 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][12] ) );
  DFF \modmult_1/zreg_reg[11]  ( .D(\modmult_1/N14 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][11] ) );
  DFF \modmult_1/zreg_reg[10]  ( .D(\modmult_1/N13 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/zin[0][10] ) );
  DFF \modmult_1/zreg_reg[9]  ( .D(\modmult_1/N12 ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\modmult_1/zin[0][9] ) );
  DFF \modmult_1/zreg_reg[8]  ( .D(\modmult_1/N11 ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\modmult_1/zin[0][8] ) );
  DFF \modmult_1/zreg_reg[7]  ( .D(\modmult_1/N10 ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\modmult_1/zin[0][7] ) );
  DFF \modmult_1/zreg_reg[6]  ( .D(\modmult_1/N9 ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\modmult_1/zin[0][6] ) );
  DFF \modmult_1/zreg_reg[5]  ( .D(\modmult_1/N8 ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\modmult_1/zin[0][5] ) );
  DFF \modmult_1/zreg_reg[4]  ( .D(\modmult_1/N7 ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\modmult_1/zin[0][4] ) );
  DFF \modmult_1/zreg_reg[3]  ( .D(\modmult_1/N6 ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\modmult_1/zin[0][3] ) );
  DFF \modmult_1/zreg_reg[2]  ( .D(\modmult_1/N5 ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\modmult_1/zin[0][2] ) );
  DFF \modmult_1/zreg_reg[1]  ( .D(\modmult_1/N4 ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\modmult_1/zin[0][1] ) );
  DFF \modmult_1/zreg_reg[0]  ( .D(\modmult_1/N3 ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\modmult_1/zin[0][0] ) );
  DFF \modmult_1/xreg_reg[1023]  ( .D(\modmult_1/N2052 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1023] ) );
  DFF \modmult_1/xreg_reg[1022]  ( .D(\modmult_1/N2051 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1022] ) );
  DFF \modmult_1/xreg_reg[1021]  ( .D(\modmult_1/N2050 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1021] ) );
  DFF \modmult_1/xreg_reg[1020]  ( .D(\modmult_1/N2049 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1020] ) );
  DFF \modmult_1/xreg_reg[1019]  ( .D(\modmult_1/N2048 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1019] ) );
  DFF \modmult_1/xreg_reg[1018]  ( .D(\modmult_1/N2047 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1018] ) );
  DFF \modmult_1/xreg_reg[1017]  ( .D(\modmult_1/N2046 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1017] ) );
  DFF \modmult_1/xreg_reg[1016]  ( .D(\modmult_1/N2045 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1016] ) );
  DFF \modmult_1/xreg_reg[1015]  ( .D(\modmult_1/N2044 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1015] ) );
  DFF \modmult_1/xreg_reg[1014]  ( .D(\modmult_1/N2043 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1014] ) );
  DFF \modmult_1/xreg_reg[1013]  ( .D(\modmult_1/N2042 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1013] ) );
  DFF \modmult_1/xreg_reg[1012]  ( .D(\modmult_1/N2041 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1012] ) );
  DFF \modmult_1/xreg_reg[1011]  ( .D(\modmult_1/N2040 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1011] ) );
  DFF \modmult_1/xreg_reg[1010]  ( .D(\modmult_1/N2039 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1010] ) );
  DFF \modmult_1/xreg_reg[1009]  ( .D(\modmult_1/N2038 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1009] ) );
  DFF \modmult_1/xreg_reg[1008]  ( .D(\modmult_1/N2037 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1008] ) );
  DFF \modmult_1/xreg_reg[1007]  ( .D(\modmult_1/N2036 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1007] ) );
  DFF \modmult_1/xreg_reg[1006]  ( .D(\modmult_1/N2035 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1006] ) );
  DFF \modmult_1/xreg_reg[1005]  ( .D(\modmult_1/N2034 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1005] ) );
  DFF \modmult_1/xreg_reg[1004]  ( .D(\modmult_1/N2033 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1004] ) );
  DFF \modmult_1/xreg_reg[1003]  ( .D(\modmult_1/N2032 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1003] ) );
  DFF \modmult_1/xreg_reg[1002]  ( .D(\modmult_1/N2031 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1002] ) );
  DFF \modmult_1/xreg_reg[1001]  ( .D(\modmult_1/N2030 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1001] ) );
  DFF \modmult_1/xreg_reg[1000]  ( .D(\modmult_1/N2029 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1000] ) );
  DFF \modmult_1/xreg_reg[999]  ( .D(\modmult_1/N2028 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[999] ) );
  DFF \modmult_1/xreg_reg[998]  ( .D(\modmult_1/N2027 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[998] ) );
  DFF \modmult_1/xreg_reg[997]  ( .D(\modmult_1/N2026 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[997] ) );
  DFF \modmult_1/xreg_reg[996]  ( .D(\modmult_1/N2025 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[996] ) );
  DFF \modmult_1/xreg_reg[995]  ( .D(\modmult_1/N2024 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[995] ) );
  DFF \modmult_1/xreg_reg[994]  ( .D(\modmult_1/N2023 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[994] ) );
  DFF \modmult_1/xreg_reg[993]  ( .D(\modmult_1/N2022 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[993] ) );
  DFF \modmult_1/xreg_reg[992]  ( .D(\modmult_1/N2021 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[992] ) );
  DFF \modmult_1/xreg_reg[991]  ( .D(\modmult_1/N2020 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[991] ) );
  DFF \modmult_1/xreg_reg[990]  ( .D(\modmult_1/N2019 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[990] ) );
  DFF \modmult_1/xreg_reg[989]  ( .D(\modmult_1/N2018 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[989] ) );
  DFF \modmult_1/xreg_reg[988]  ( .D(\modmult_1/N2017 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[988] ) );
  DFF \modmult_1/xreg_reg[987]  ( .D(\modmult_1/N2016 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[987] ) );
  DFF \modmult_1/xreg_reg[986]  ( .D(\modmult_1/N2015 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[986] ) );
  DFF \modmult_1/xreg_reg[985]  ( .D(\modmult_1/N2014 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[985] ) );
  DFF \modmult_1/xreg_reg[984]  ( .D(\modmult_1/N2013 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[984] ) );
  DFF \modmult_1/xreg_reg[983]  ( .D(\modmult_1/N2012 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[983] ) );
  DFF \modmult_1/xreg_reg[982]  ( .D(\modmult_1/N2011 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[982] ) );
  DFF \modmult_1/xreg_reg[981]  ( .D(\modmult_1/N2010 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[981] ) );
  DFF \modmult_1/xreg_reg[980]  ( .D(\modmult_1/N2009 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[980] ) );
  DFF \modmult_1/xreg_reg[979]  ( .D(\modmult_1/N2008 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[979] ) );
  DFF \modmult_1/xreg_reg[978]  ( .D(\modmult_1/N2007 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[978] ) );
  DFF \modmult_1/xreg_reg[977]  ( .D(\modmult_1/N2006 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[977] ) );
  DFF \modmult_1/xreg_reg[976]  ( .D(\modmult_1/N2005 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[976] ) );
  DFF \modmult_1/xreg_reg[975]  ( .D(\modmult_1/N2004 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[975] ) );
  DFF \modmult_1/xreg_reg[974]  ( .D(\modmult_1/N2003 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[974] ) );
  DFF \modmult_1/xreg_reg[973]  ( .D(\modmult_1/N2002 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[973] ) );
  DFF \modmult_1/xreg_reg[972]  ( .D(\modmult_1/N2001 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[972] ) );
  DFF \modmult_1/xreg_reg[971]  ( .D(\modmult_1/N2000 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[971] ) );
  DFF \modmult_1/xreg_reg[970]  ( .D(\modmult_1/N1999 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[970] ) );
  DFF \modmult_1/xreg_reg[969]  ( .D(\modmult_1/N1998 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[969] ) );
  DFF \modmult_1/xreg_reg[968]  ( .D(\modmult_1/N1997 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[968] ) );
  DFF \modmult_1/xreg_reg[967]  ( .D(\modmult_1/N1996 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[967] ) );
  DFF \modmult_1/xreg_reg[966]  ( .D(\modmult_1/N1995 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[966] ) );
  DFF \modmult_1/xreg_reg[965]  ( .D(\modmult_1/N1994 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[965] ) );
  DFF \modmult_1/xreg_reg[964]  ( .D(\modmult_1/N1993 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[964] ) );
  DFF \modmult_1/xreg_reg[963]  ( .D(\modmult_1/N1992 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[963] ) );
  DFF \modmult_1/xreg_reg[962]  ( .D(\modmult_1/N1991 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[962] ) );
  DFF \modmult_1/xreg_reg[961]  ( .D(\modmult_1/N1990 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[961] ) );
  DFF \modmult_1/xreg_reg[960]  ( .D(\modmult_1/N1989 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[960] ) );
  DFF \modmult_1/xreg_reg[959]  ( .D(\modmult_1/N1988 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[959] ) );
  DFF \modmult_1/xreg_reg[958]  ( .D(\modmult_1/N1987 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[958] ) );
  DFF \modmult_1/xreg_reg[957]  ( .D(\modmult_1/N1986 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[957] ) );
  DFF \modmult_1/xreg_reg[956]  ( .D(\modmult_1/N1985 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[956] ) );
  DFF \modmult_1/xreg_reg[955]  ( .D(\modmult_1/N1984 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[955] ) );
  DFF \modmult_1/xreg_reg[954]  ( .D(\modmult_1/N1983 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[954] ) );
  DFF \modmult_1/xreg_reg[953]  ( .D(\modmult_1/N1982 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[953] ) );
  DFF \modmult_1/xreg_reg[952]  ( .D(\modmult_1/N1981 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[952] ) );
  DFF \modmult_1/xreg_reg[951]  ( .D(\modmult_1/N1980 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[951] ) );
  DFF \modmult_1/xreg_reg[950]  ( .D(\modmult_1/N1979 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[950] ) );
  DFF \modmult_1/xreg_reg[949]  ( .D(\modmult_1/N1978 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[949] ) );
  DFF \modmult_1/xreg_reg[948]  ( .D(\modmult_1/N1977 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[948] ) );
  DFF \modmult_1/xreg_reg[947]  ( .D(\modmult_1/N1976 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[947] ) );
  DFF \modmult_1/xreg_reg[946]  ( .D(\modmult_1/N1975 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[946] ) );
  DFF \modmult_1/xreg_reg[945]  ( .D(\modmult_1/N1974 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[945] ) );
  DFF \modmult_1/xreg_reg[944]  ( .D(\modmult_1/N1973 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[944] ) );
  DFF \modmult_1/xreg_reg[943]  ( .D(\modmult_1/N1972 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[943] ) );
  DFF \modmult_1/xreg_reg[942]  ( .D(\modmult_1/N1971 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[942] ) );
  DFF \modmult_1/xreg_reg[941]  ( .D(\modmult_1/N1970 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[941] ) );
  DFF \modmult_1/xreg_reg[940]  ( .D(\modmult_1/N1969 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[940] ) );
  DFF \modmult_1/xreg_reg[939]  ( .D(\modmult_1/N1968 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[939] ) );
  DFF \modmult_1/xreg_reg[938]  ( .D(\modmult_1/N1967 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[938] ) );
  DFF \modmult_1/xreg_reg[937]  ( .D(\modmult_1/N1966 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[937] ) );
  DFF \modmult_1/xreg_reg[936]  ( .D(\modmult_1/N1965 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[936] ) );
  DFF \modmult_1/xreg_reg[935]  ( .D(\modmult_1/N1964 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[935] ) );
  DFF \modmult_1/xreg_reg[934]  ( .D(\modmult_1/N1963 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[934] ) );
  DFF \modmult_1/xreg_reg[933]  ( .D(\modmult_1/N1962 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[933] ) );
  DFF \modmult_1/xreg_reg[932]  ( .D(\modmult_1/N1961 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[932] ) );
  DFF \modmult_1/xreg_reg[931]  ( .D(\modmult_1/N1960 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[931] ) );
  DFF \modmult_1/xreg_reg[930]  ( .D(\modmult_1/N1959 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[930] ) );
  DFF \modmult_1/xreg_reg[929]  ( .D(\modmult_1/N1958 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[929] ) );
  DFF \modmult_1/xreg_reg[928]  ( .D(\modmult_1/N1957 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[928] ) );
  DFF \modmult_1/xreg_reg[927]  ( .D(\modmult_1/N1956 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[927] ) );
  DFF \modmult_1/xreg_reg[926]  ( .D(\modmult_1/N1955 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[926] ) );
  DFF \modmult_1/xreg_reg[925]  ( .D(\modmult_1/N1954 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[925] ) );
  DFF \modmult_1/xreg_reg[924]  ( .D(\modmult_1/N1953 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[924] ) );
  DFF \modmult_1/xreg_reg[923]  ( .D(\modmult_1/N1952 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[923] ) );
  DFF \modmult_1/xreg_reg[922]  ( .D(\modmult_1/N1951 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[922] ) );
  DFF \modmult_1/xreg_reg[921]  ( .D(\modmult_1/N1950 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[921] ) );
  DFF \modmult_1/xreg_reg[920]  ( .D(\modmult_1/N1949 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[920] ) );
  DFF \modmult_1/xreg_reg[919]  ( .D(\modmult_1/N1948 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[919] ) );
  DFF \modmult_1/xreg_reg[918]  ( .D(\modmult_1/N1947 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[918] ) );
  DFF \modmult_1/xreg_reg[917]  ( .D(\modmult_1/N1946 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[917] ) );
  DFF \modmult_1/xreg_reg[916]  ( .D(\modmult_1/N1945 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[916] ) );
  DFF \modmult_1/xreg_reg[915]  ( .D(\modmult_1/N1944 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[915] ) );
  DFF \modmult_1/xreg_reg[914]  ( .D(\modmult_1/N1943 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[914] ) );
  DFF \modmult_1/xreg_reg[913]  ( .D(\modmult_1/N1942 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[913] ) );
  DFF \modmult_1/xreg_reg[912]  ( .D(\modmult_1/N1941 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[912] ) );
  DFF \modmult_1/xreg_reg[911]  ( .D(\modmult_1/N1940 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[911] ) );
  DFF \modmult_1/xreg_reg[910]  ( .D(\modmult_1/N1939 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[910] ) );
  DFF \modmult_1/xreg_reg[909]  ( .D(\modmult_1/N1938 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[909] ) );
  DFF \modmult_1/xreg_reg[908]  ( .D(\modmult_1/N1937 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[908] ) );
  DFF \modmult_1/xreg_reg[907]  ( .D(\modmult_1/N1936 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[907] ) );
  DFF \modmult_1/xreg_reg[906]  ( .D(\modmult_1/N1935 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[906] ) );
  DFF \modmult_1/xreg_reg[905]  ( .D(\modmult_1/N1934 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[905] ) );
  DFF \modmult_1/xreg_reg[904]  ( .D(\modmult_1/N1933 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[904] ) );
  DFF \modmult_1/xreg_reg[903]  ( .D(\modmult_1/N1932 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[903] ) );
  DFF \modmult_1/xreg_reg[902]  ( .D(\modmult_1/N1931 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[902] ) );
  DFF \modmult_1/xreg_reg[901]  ( .D(\modmult_1/N1930 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[901] ) );
  DFF \modmult_1/xreg_reg[900]  ( .D(\modmult_1/N1929 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[900] ) );
  DFF \modmult_1/xreg_reg[899]  ( .D(\modmult_1/N1928 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[899] ) );
  DFF \modmult_1/xreg_reg[898]  ( .D(\modmult_1/N1927 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[898] ) );
  DFF \modmult_1/xreg_reg[897]  ( .D(\modmult_1/N1926 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[897] ) );
  DFF \modmult_1/xreg_reg[896]  ( .D(\modmult_1/N1925 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[896] ) );
  DFF \modmult_1/xreg_reg[895]  ( .D(\modmult_1/N1924 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[895] ) );
  DFF \modmult_1/xreg_reg[894]  ( .D(\modmult_1/N1923 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[894] ) );
  DFF \modmult_1/xreg_reg[893]  ( .D(\modmult_1/N1922 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[893] ) );
  DFF \modmult_1/xreg_reg[892]  ( .D(\modmult_1/N1921 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[892] ) );
  DFF \modmult_1/xreg_reg[891]  ( .D(\modmult_1/N1920 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[891] ) );
  DFF \modmult_1/xreg_reg[890]  ( .D(\modmult_1/N1919 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[890] ) );
  DFF \modmult_1/xreg_reg[889]  ( .D(\modmult_1/N1918 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[889] ) );
  DFF \modmult_1/xreg_reg[888]  ( .D(\modmult_1/N1917 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[888] ) );
  DFF \modmult_1/xreg_reg[887]  ( .D(\modmult_1/N1916 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[887] ) );
  DFF \modmult_1/xreg_reg[886]  ( .D(\modmult_1/N1915 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[886] ) );
  DFF \modmult_1/xreg_reg[885]  ( .D(\modmult_1/N1914 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[885] ) );
  DFF \modmult_1/xreg_reg[884]  ( .D(\modmult_1/N1913 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[884] ) );
  DFF \modmult_1/xreg_reg[883]  ( .D(\modmult_1/N1912 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[883] ) );
  DFF \modmult_1/xreg_reg[882]  ( .D(\modmult_1/N1911 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[882] ) );
  DFF \modmult_1/xreg_reg[881]  ( .D(\modmult_1/N1910 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[881] ) );
  DFF \modmult_1/xreg_reg[880]  ( .D(\modmult_1/N1909 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[880] ) );
  DFF \modmult_1/xreg_reg[879]  ( .D(\modmult_1/N1908 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[879] ) );
  DFF \modmult_1/xreg_reg[878]  ( .D(\modmult_1/N1907 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[878] ) );
  DFF \modmult_1/xreg_reg[877]  ( .D(\modmult_1/N1906 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[877] ) );
  DFF \modmult_1/xreg_reg[876]  ( .D(\modmult_1/N1905 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[876] ) );
  DFF \modmult_1/xreg_reg[875]  ( .D(\modmult_1/N1904 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[875] ) );
  DFF \modmult_1/xreg_reg[874]  ( .D(\modmult_1/N1903 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[874] ) );
  DFF \modmult_1/xreg_reg[873]  ( .D(\modmult_1/N1902 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[873] ) );
  DFF \modmult_1/xreg_reg[872]  ( .D(\modmult_1/N1901 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[872] ) );
  DFF \modmult_1/xreg_reg[871]  ( .D(\modmult_1/N1900 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[871] ) );
  DFF \modmult_1/xreg_reg[870]  ( .D(\modmult_1/N1899 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[870] ) );
  DFF \modmult_1/xreg_reg[869]  ( .D(\modmult_1/N1898 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[869] ) );
  DFF \modmult_1/xreg_reg[868]  ( .D(\modmult_1/N1897 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[868] ) );
  DFF \modmult_1/xreg_reg[867]  ( .D(\modmult_1/N1896 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[867] ) );
  DFF \modmult_1/xreg_reg[866]  ( .D(\modmult_1/N1895 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[866] ) );
  DFF \modmult_1/xreg_reg[865]  ( .D(\modmult_1/N1894 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[865] ) );
  DFF \modmult_1/xreg_reg[864]  ( .D(\modmult_1/N1893 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[864] ) );
  DFF \modmult_1/xreg_reg[863]  ( .D(\modmult_1/N1892 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[863] ) );
  DFF \modmult_1/xreg_reg[862]  ( .D(\modmult_1/N1891 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[862] ) );
  DFF \modmult_1/xreg_reg[861]  ( .D(\modmult_1/N1890 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[861] ) );
  DFF \modmult_1/xreg_reg[860]  ( .D(\modmult_1/N1889 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[860] ) );
  DFF \modmult_1/xreg_reg[859]  ( .D(\modmult_1/N1888 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[859] ) );
  DFF \modmult_1/xreg_reg[858]  ( .D(\modmult_1/N1887 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[858] ) );
  DFF \modmult_1/xreg_reg[857]  ( .D(\modmult_1/N1886 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[857] ) );
  DFF \modmult_1/xreg_reg[856]  ( .D(\modmult_1/N1885 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[856] ) );
  DFF \modmult_1/xreg_reg[855]  ( .D(\modmult_1/N1884 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[855] ) );
  DFF \modmult_1/xreg_reg[854]  ( .D(\modmult_1/N1883 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[854] ) );
  DFF \modmult_1/xreg_reg[853]  ( .D(\modmult_1/N1882 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[853] ) );
  DFF \modmult_1/xreg_reg[852]  ( .D(\modmult_1/N1881 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[852] ) );
  DFF \modmult_1/xreg_reg[851]  ( .D(\modmult_1/N1880 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[851] ) );
  DFF \modmult_1/xreg_reg[850]  ( .D(\modmult_1/N1879 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[850] ) );
  DFF \modmult_1/xreg_reg[849]  ( .D(\modmult_1/N1878 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[849] ) );
  DFF \modmult_1/xreg_reg[848]  ( .D(\modmult_1/N1877 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[848] ) );
  DFF \modmult_1/xreg_reg[847]  ( .D(\modmult_1/N1876 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[847] ) );
  DFF \modmult_1/xreg_reg[846]  ( .D(\modmult_1/N1875 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[846] ) );
  DFF \modmult_1/xreg_reg[845]  ( .D(\modmult_1/N1874 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[845] ) );
  DFF \modmult_1/xreg_reg[844]  ( .D(\modmult_1/N1873 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[844] ) );
  DFF \modmult_1/xreg_reg[843]  ( .D(\modmult_1/N1872 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[843] ) );
  DFF \modmult_1/xreg_reg[842]  ( .D(\modmult_1/N1871 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[842] ) );
  DFF \modmult_1/xreg_reg[841]  ( .D(\modmult_1/N1870 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[841] ) );
  DFF \modmult_1/xreg_reg[840]  ( .D(\modmult_1/N1869 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[840] ) );
  DFF \modmult_1/xreg_reg[839]  ( .D(\modmult_1/N1868 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[839] ) );
  DFF \modmult_1/xreg_reg[838]  ( .D(\modmult_1/N1867 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[838] ) );
  DFF \modmult_1/xreg_reg[837]  ( .D(\modmult_1/N1866 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[837] ) );
  DFF \modmult_1/xreg_reg[836]  ( .D(\modmult_1/N1865 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[836] ) );
  DFF \modmult_1/xreg_reg[835]  ( .D(\modmult_1/N1864 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[835] ) );
  DFF \modmult_1/xreg_reg[834]  ( .D(\modmult_1/N1863 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[834] ) );
  DFF \modmult_1/xreg_reg[833]  ( .D(\modmult_1/N1862 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[833] ) );
  DFF \modmult_1/xreg_reg[832]  ( .D(\modmult_1/N1861 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[832] ) );
  DFF \modmult_1/xreg_reg[831]  ( .D(\modmult_1/N1860 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[831] ) );
  DFF \modmult_1/xreg_reg[830]  ( .D(\modmult_1/N1859 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[830] ) );
  DFF \modmult_1/xreg_reg[829]  ( .D(\modmult_1/N1858 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[829] ) );
  DFF \modmult_1/xreg_reg[828]  ( .D(\modmult_1/N1857 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[828] ) );
  DFF \modmult_1/xreg_reg[827]  ( .D(\modmult_1/N1856 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[827] ) );
  DFF \modmult_1/xreg_reg[826]  ( .D(\modmult_1/N1855 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[826] ) );
  DFF \modmult_1/xreg_reg[825]  ( .D(\modmult_1/N1854 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[825] ) );
  DFF \modmult_1/xreg_reg[824]  ( .D(\modmult_1/N1853 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[824] ) );
  DFF \modmult_1/xreg_reg[823]  ( .D(\modmult_1/N1852 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[823] ) );
  DFF \modmult_1/xreg_reg[822]  ( .D(\modmult_1/N1851 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[822] ) );
  DFF \modmult_1/xreg_reg[821]  ( .D(\modmult_1/N1850 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[821] ) );
  DFF \modmult_1/xreg_reg[820]  ( .D(\modmult_1/N1849 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[820] ) );
  DFF \modmult_1/xreg_reg[819]  ( .D(\modmult_1/N1848 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[819] ) );
  DFF \modmult_1/xreg_reg[818]  ( .D(\modmult_1/N1847 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[818] ) );
  DFF \modmult_1/xreg_reg[817]  ( .D(\modmult_1/N1846 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[817] ) );
  DFF \modmult_1/xreg_reg[816]  ( .D(\modmult_1/N1845 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[816] ) );
  DFF \modmult_1/xreg_reg[815]  ( .D(\modmult_1/N1844 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[815] ) );
  DFF \modmult_1/xreg_reg[814]  ( .D(\modmult_1/N1843 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[814] ) );
  DFF \modmult_1/xreg_reg[813]  ( .D(\modmult_1/N1842 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[813] ) );
  DFF \modmult_1/xreg_reg[812]  ( .D(\modmult_1/N1841 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[812] ) );
  DFF \modmult_1/xreg_reg[811]  ( .D(\modmult_1/N1840 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[811] ) );
  DFF \modmult_1/xreg_reg[810]  ( .D(\modmult_1/N1839 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[810] ) );
  DFF \modmult_1/xreg_reg[809]  ( .D(\modmult_1/N1838 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[809] ) );
  DFF \modmult_1/xreg_reg[808]  ( .D(\modmult_1/N1837 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[808] ) );
  DFF \modmult_1/xreg_reg[807]  ( .D(\modmult_1/N1836 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[807] ) );
  DFF \modmult_1/xreg_reg[806]  ( .D(\modmult_1/N1835 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[806] ) );
  DFF \modmult_1/xreg_reg[805]  ( .D(\modmult_1/N1834 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[805] ) );
  DFF \modmult_1/xreg_reg[804]  ( .D(\modmult_1/N1833 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[804] ) );
  DFF \modmult_1/xreg_reg[803]  ( .D(\modmult_1/N1832 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[803] ) );
  DFF \modmult_1/xreg_reg[802]  ( .D(\modmult_1/N1831 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[802] ) );
  DFF \modmult_1/xreg_reg[801]  ( .D(\modmult_1/N1830 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[801] ) );
  DFF \modmult_1/xreg_reg[800]  ( .D(\modmult_1/N1829 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[800] ) );
  DFF \modmult_1/xreg_reg[799]  ( .D(\modmult_1/N1828 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[799] ) );
  DFF \modmult_1/xreg_reg[798]  ( .D(\modmult_1/N1827 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[798] ) );
  DFF \modmult_1/xreg_reg[797]  ( .D(\modmult_1/N1826 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[797] ) );
  DFF \modmult_1/xreg_reg[796]  ( .D(\modmult_1/N1825 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[796] ) );
  DFF \modmult_1/xreg_reg[795]  ( .D(\modmult_1/N1824 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[795] ) );
  DFF \modmult_1/xreg_reg[794]  ( .D(\modmult_1/N1823 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[794] ) );
  DFF \modmult_1/xreg_reg[793]  ( .D(\modmult_1/N1822 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[793] ) );
  DFF \modmult_1/xreg_reg[792]  ( .D(\modmult_1/N1821 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[792] ) );
  DFF \modmult_1/xreg_reg[791]  ( .D(\modmult_1/N1820 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[791] ) );
  DFF \modmult_1/xreg_reg[790]  ( .D(\modmult_1/N1819 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[790] ) );
  DFF \modmult_1/xreg_reg[789]  ( .D(\modmult_1/N1818 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[789] ) );
  DFF \modmult_1/xreg_reg[788]  ( .D(\modmult_1/N1817 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[788] ) );
  DFF \modmult_1/xreg_reg[787]  ( .D(\modmult_1/N1816 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[787] ) );
  DFF \modmult_1/xreg_reg[786]  ( .D(\modmult_1/N1815 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[786] ) );
  DFF \modmult_1/xreg_reg[785]  ( .D(\modmult_1/N1814 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[785] ) );
  DFF \modmult_1/xreg_reg[784]  ( .D(\modmult_1/N1813 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[784] ) );
  DFF \modmult_1/xreg_reg[783]  ( .D(\modmult_1/N1812 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[783] ) );
  DFF \modmult_1/xreg_reg[782]  ( .D(\modmult_1/N1811 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[782] ) );
  DFF \modmult_1/xreg_reg[781]  ( .D(\modmult_1/N1810 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[781] ) );
  DFF \modmult_1/xreg_reg[780]  ( .D(\modmult_1/N1809 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[780] ) );
  DFF \modmult_1/xreg_reg[779]  ( .D(\modmult_1/N1808 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[779] ) );
  DFF \modmult_1/xreg_reg[778]  ( .D(\modmult_1/N1807 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[778] ) );
  DFF \modmult_1/xreg_reg[777]  ( .D(\modmult_1/N1806 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[777] ) );
  DFF \modmult_1/xreg_reg[776]  ( .D(\modmult_1/N1805 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[776] ) );
  DFF \modmult_1/xreg_reg[775]  ( .D(\modmult_1/N1804 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[775] ) );
  DFF \modmult_1/xreg_reg[774]  ( .D(\modmult_1/N1803 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[774] ) );
  DFF \modmult_1/xreg_reg[773]  ( .D(\modmult_1/N1802 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[773] ) );
  DFF \modmult_1/xreg_reg[772]  ( .D(\modmult_1/N1801 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[772] ) );
  DFF \modmult_1/xreg_reg[771]  ( .D(\modmult_1/N1800 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[771] ) );
  DFF \modmult_1/xreg_reg[770]  ( .D(\modmult_1/N1799 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[770] ) );
  DFF \modmult_1/xreg_reg[769]  ( .D(\modmult_1/N1798 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[769] ) );
  DFF \modmult_1/xreg_reg[768]  ( .D(\modmult_1/N1797 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[768] ) );
  DFF \modmult_1/xreg_reg[767]  ( .D(\modmult_1/N1796 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[767] ) );
  DFF \modmult_1/xreg_reg[766]  ( .D(\modmult_1/N1795 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[766] ) );
  DFF \modmult_1/xreg_reg[765]  ( .D(\modmult_1/N1794 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[765] ) );
  DFF \modmult_1/xreg_reg[764]  ( .D(\modmult_1/N1793 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[764] ) );
  DFF \modmult_1/xreg_reg[763]  ( .D(\modmult_1/N1792 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[763] ) );
  DFF \modmult_1/xreg_reg[762]  ( .D(\modmult_1/N1791 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[762] ) );
  DFF \modmult_1/xreg_reg[761]  ( .D(\modmult_1/N1790 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[761] ) );
  DFF \modmult_1/xreg_reg[760]  ( .D(\modmult_1/N1789 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[760] ) );
  DFF \modmult_1/xreg_reg[759]  ( .D(\modmult_1/N1788 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[759] ) );
  DFF \modmult_1/xreg_reg[758]  ( .D(\modmult_1/N1787 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[758] ) );
  DFF \modmult_1/xreg_reg[757]  ( .D(\modmult_1/N1786 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[757] ) );
  DFF \modmult_1/xreg_reg[756]  ( .D(\modmult_1/N1785 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[756] ) );
  DFF \modmult_1/xreg_reg[755]  ( .D(\modmult_1/N1784 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[755] ) );
  DFF \modmult_1/xreg_reg[754]  ( .D(\modmult_1/N1783 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[754] ) );
  DFF \modmult_1/xreg_reg[753]  ( .D(\modmult_1/N1782 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[753] ) );
  DFF \modmult_1/xreg_reg[752]  ( .D(\modmult_1/N1781 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[752] ) );
  DFF \modmult_1/xreg_reg[751]  ( .D(\modmult_1/N1780 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[751] ) );
  DFF \modmult_1/xreg_reg[750]  ( .D(\modmult_1/N1779 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[750] ) );
  DFF \modmult_1/xreg_reg[749]  ( .D(\modmult_1/N1778 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[749] ) );
  DFF \modmult_1/xreg_reg[748]  ( .D(\modmult_1/N1777 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[748] ) );
  DFF \modmult_1/xreg_reg[747]  ( .D(\modmult_1/N1776 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[747] ) );
  DFF \modmult_1/xreg_reg[746]  ( .D(\modmult_1/N1775 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[746] ) );
  DFF \modmult_1/xreg_reg[745]  ( .D(\modmult_1/N1774 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[745] ) );
  DFF \modmult_1/xreg_reg[744]  ( .D(\modmult_1/N1773 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[744] ) );
  DFF \modmult_1/xreg_reg[743]  ( .D(\modmult_1/N1772 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[743] ) );
  DFF \modmult_1/xreg_reg[742]  ( .D(\modmult_1/N1771 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[742] ) );
  DFF \modmult_1/xreg_reg[741]  ( .D(\modmult_1/N1770 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[741] ) );
  DFF \modmult_1/xreg_reg[740]  ( .D(\modmult_1/N1769 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[740] ) );
  DFF \modmult_1/xreg_reg[739]  ( .D(\modmult_1/N1768 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[739] ) );
  DFF \modmult_1/xreg_reg[738]  ( .D(\modmult_1/N1767 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[738] ) );
  DFF \modmult_1/xreg_reg[737]  ( .D(\modmult_1/N1766 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[737] ) );
  DFF \modmult_1/xreg_reg[736]  ( .D(\modmult_1/N1765 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[736] ) );
  DFF \modmult_1/xreg_reg[735]  ( .D(\modmult_1/N1764 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[735] ) );
  DFF \modmult_1/xreg_reg[734]  ( .D(\modmult_1/N1763 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[734] ) );
  DFF \modmult_1/xreg_reg[733]  ( .D(\modmult_1/N1762 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[733] ) );
  DFF \modmult_1/xreg_reg[732]  ( .D(\modmult_1/N1761 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[732] ) );
  DFF \modmult_1/xreg_reg[731]  ( .D(\modmult_1/N1760 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[731] ) );
  DFF \modmult_1/xreg_reg[730]  ( .D(\modmult_1/N1759 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[730] ) );
  DFF \modmult_1/xreg_reg[729]  ( .D(\modmult_1/N1758 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[729] ) );
  DFF \modmult_1/xreg_reg[728]  ( .D(\modmult_1/N1757 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[728] ) );
  DFF \modmult_1/xreg_reg[727]  ( .D(\modmult_1/N1756 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[727] ) );
  DFF \modmult_1/xreg_reg[726]  ( .D(\modmult_1/N1755 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[726] ) );
  DFF \modmult_1/xreg_reg[725]  ( .D(\modmult_1/N1754 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[725] ) );
  DFF \modmult_1/xreg_reg[724]  ( .D(\modmult_1/N1753 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[724] ) );
  DFF \modmult_1/xreg_reg[723]  ( .D(\modmult_1/N1752 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[723] ) );
  DFF \modmult_1/xreg_reg[722]  ( .D(\modmult_1/N1751 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[722] ) );
  DFF \modmult_1/xreg_reg[721]  ( .D(\modmult_1/N1750 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[721] ) );
  DFF \modmult_1/xreg_reg[720]  ( .D(\modmult_1/N1749 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[720] ) );
  DFF \modmult_1/xreg_reg[719]  ( .D(\modmult_1/N1748 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[719] ) );
  DFF \modmult_1/xreg_reg[718]  ( .D(\modmult_1/N1747 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[718] ) );
  DFF \modmult_1/xreg_reg[717]  ( .D(\modmult_1/N1746 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[717] ) );
  DFF \modmult_1/xreg_reg[716]  ( .D(\modmult_1/N1745 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[716] ) );
  DFF \modmult_1/xreg_reg[715]  ( .D(\modmult_1/N1744 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[715] ) );
  DFF \modmult_1/xreg_reg[714]  ( .D(\modmult_1/N1743 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[714] ) );
  DFF \modmult_1/xreg_reg[713]  ( .D(\modmult_1/N1742 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[713] ) );
  DFF \modmult_1/xreg_reg[712]  ( .D(\modmult_1/N1741 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[712] ) );
  DFF \modmult_1/xreg_reg[711]  ( .D(\modmult_1/N1740 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[711] ) );
  DFF \modmult_1/xreg_reg[710]  ( .D(\modmult_1/N1739 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[710] ) );
  DFF \modmult_1/xreg_reg[709]  ( .D(\modmult_1/N1738 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[709] ) );
  DFF \modmult_1/xreg_reg[708]  ( .D(\modmult_1/N1737 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[708] ) );
  DFF \modmult_1/xreg_reg[707]  ( .D(\modmult_1/N1736 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[707] ) );
  DFF \modmult_1/xreg_reg[706]  ( .D(\modmult_1/N1735 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[706] ) );
  DFF \modmult_1/xreg_reg[705]  ( .D(\modmult_1/N1734 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[705] ) );
  DFF \modmult_1/xreg_reg[704]  ( .D(\modmult_1/N1733 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[704] ) );
  DFF \modmult_1/xreg_reg[703]  ( .D(\modmult_1/N1732 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[703] ) );
  DFF \modmult_1/xreg_reg[702]  ( .D(\modmult_1/N1731 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[702] ) );
  DFF \modmult_1/xreg_reg[701]  ( .D(\modmult_1/N1730 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[701] ) );
  DFF \modmult_1/xreg_reg[700]  ( .D(\modmult_1/N1729 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[700] ) );
  DFF \modmult_1/xreg_reg[699]  ( .D(\modmult_1/N1728 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[699] ) );
  DFF \modmult_1/xreg_reg[698]  ( .D(\modmult_1/N1727 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[698] ) );
  DFF \modmult_1/xreg_reg[697]  ( .D(\modmult_1/N1726 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[697] ) );
  DFF \modmult_1/xreg_reg[696]  ( .D(\modmult_1/N1725 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[696] ) );
  DFF \modmult_1/xreg_reg[695]  ( .D(\modmult_1/N1724 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[695] ) );
  DFF \modmult_1/xreg_reg[694]  ( .D(\modmult_1/N1723 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[694] ) );
  DFF \modmult_1/xreg_reg[693]  ( .D(\modmult_1/N1722 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[693] ) );
  DFF \modmult_1/xreg_reg[692]  ( .D(\modmult_1/N1721 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[692] ) );
  DFF \modmult_1/xreg_reg[691]  ( .D(\modmult_1/N1720 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[691] ) );
  DFF \modmult_1/xreg_reg[690]  ( .D(\modmult_1/N1719 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[690] ) );
  DFF \modmult_1/xreg_reg[689]  ( .D(\modmult_1/N1718 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[689] ) );
  DFF \modmult_1/xreg_reg[688]  ( .D(\modmult_1/N1717 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[688] ) );
  DFF \modmult_1/xreg_reg[687]  ( .D(\modmult_1/N1716 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[687] ) );
  DFF \modmult_1/xreg_reg[686]  ( .D(\modmult_1/N1715 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[686] ) );
  DFF \modmult_1/xreg_reg[685]  ( .D(\modmult_1/N1714 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[685] ) );
  DFF \modmult_1/xreg_reg[684]  ( .D(\modmult_1/N1713 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[684] ) );
  DFF \modmult_1/xreg_reg[683]  ( .D(\modmult_1/N1712 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[683] ) );
  DFF \modmult_1/xreg_reg[682]  ( .D(\modmult_1/N1711 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[682] ) );
  DFF \modmult_1/xreg_reg[681]  ( .D(\modmult_1/N1710 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[681] ) );
  DFF \modmult_1/xreg_reg[680]  ( .D(\modmult_1/N1709 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[680] ) );
  DFF \modmult_1/xreg_reg[679]  ( .D(\modmult_1/N1708 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[679] ) );
  DFF \modmult_1/xreg_reg[678]  ( .D(\modmult_1/N1707 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[678] ) );
  DFF \modmult_1/xreg_reg[677]  ( .D(\modmult_1/N1706 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[677] ) );
  DFF \modmult_1/xreg_reg[676]  ( .D(\modmult_1/N1705 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[676] ) );
  DFF \modmult_1/xreg_reg[675]  ( .D(\modmult_1/N1704 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[675] ) );
  DFF \modmult_1/xreg_reg[674]  ( .D(\modmult_1/N1703 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[674] ) );
  DFF \modmult_1/xreg_reg[673]  ( .D(\modmult_1/N1702 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[673] ) );
  DFF \modmult_1/xreg_reg[672]  ( .D(\modmult_1/N1701 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[672] ) );
  DFF \modmult_1/xreg_reg[671]  ( .D(\modmult_1/N1700 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[671] ) );
  DFF \modmult_1/xreg_reg[670]  ( .D(\modmult_1/N1699 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[670] ) );
  DFF \modmult_1/xreg_reg[669]  ( .D(\modmult_1/N1698 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[669] ) );
  DFF \modmult_1/xreg_reg[668]  ( .D(\modmult_1/N1697 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[668] ) );
  DFF \modmult_1/xreg_reg[667]  ( .D(\modmult_1/N1696 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[667] ) );
  DFF \modmult_1/xreg_reg[666]  ( .D(\modmult_1/N1695 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[666] ) );
  DFF \modmult_1/xreg_reg[665]  ( .D(\modmult_1/N1694 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[665] ) );
  DFF \modmult_1/xreg_reg[664]  ( .D(\modmult_1/N1693 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[664] ) );
  DFF \modmult_1/xreg_reg[663]  ( .D(\modmult_1/N1692 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[663] ) );
  DFF \modmult_1/xreg_reg[662]  ( .D(\modmult_1/N1691 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[662] ) );
  DFF \modmult_1/xreg_reg[661]  ( .D(\modmult_1/N1690 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[661] ) );
  DFF \modmult_1/xreg_reg[660]  ( .D(\modmult_1/N1689 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[660] ) );
  DFF \modmult_1/xreg_reg[659]  ( .D(\modmult_1/N1688 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[659] ) );
  DFF \modmult_1/xreg_reg[658]  ( .D(\modmult_1/N1687 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[658] ) );
  DFF \modmult_1/xreg_reg[657]  ( .D(\modmult_1/N1686 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[657] ) );
  DFF \modmult_1/xreg_reg[656]  ( .D(\modmult_1/N1685 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[656] ) );
  DFF \modmult_1/xreg_reg[655]  ( .D(\modmult_1/N1684 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[655] ) );
  DFF \modmult_1/xreg_reg[654]  ( .D(\modmult_1/N1683 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[654] ) );
  DFF \modmult_1/xreg_reg[653]  ( .D(\modmult_1/N1682 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[653] ) );
  DFF \modmult_1/xreg_reg[652]  ( .D(\modmult_1/N1681 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[652] ) );
  DFF \modmult_1/xreg_reg[651]  ( .D(\modmult_1/N1680 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[651] ) );
  DFF \modmult_1/xreg_reg[650]  ( .D(\modmult_1/N1679 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[650] ) );
  DFF \modmult_1/xreg_reg[649]  ( .D(\modmult_1/N1678 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[649] ) );
  DFF \modmult_1/xreg_reg[648]  ( .D(\modmult_1/N1677 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[648] ) );
  DFF \modmult_1/xreg_reg[647]  ( .D(\modmult_1/N1676 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[647] ) );
  DFF \modmult_1/xreg_reg[646]  ( .D(\modmult_1/N1675 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[646] ) );
  DFF \modmult_1/xreg_reg[645]  ( .D(\modmult_1/N1674 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[645] ) );
  DFF \modmult_1/xreg_reg[644]  ( .D(\modmult_1/N1673 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[644] ) );
  DFF \modmult_1/xreg_reg[643]  ( .D(\modmult_1/N1672 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[643] ) );
  DFF \modmult_1/xreg_reg[642]  ( .D(\modmult_1/N1671 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[642] ) );
  DFF \modmult_1/xreg_reg[641]  ( .D(\modmult_1/N1670 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[641] ) );
  DFF \modmult_1/xreg_reg[640]  ( .D(\modmult_1/N1669 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[640] ) );
  DFF \modmult_1/xreg_reg[639]  ( .D(\modmult_1/N1668 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[639] ) );
  DFF \modmult_1/xreg_reg[638]  ( .D(\modmult_1/N1667 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[638] ) );
  DFF \modmult_1/xreg_reg[637]  ( .D(\modmult_1/N1666 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[637] ) );
  DFF \modmult_1/xreg_reg[636]  ( .D(\modmult_1/N1665 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[636] ) );
  DFF \modmult_1/xreg_reg[635]  ( .D(\modmult_1/N1664 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[635] ) );
  DFF \modmult_1/xreg_reg[634]  ( .D(\modmult_1/N1663 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[634] ) );
  DFF \modmult_1/xreg_reg[633]  ( .D(\modmult_1/N1662 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[633] ) );
  DFF \modmult_1/xreg_reg[632]  ( .D(\modmult_1/N1661 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[632] ) );
  DFF \modmult_1/xreg_reg[631]  ( .D(\modmult_1/N1660 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[631] ) );
  DFF \modmult_1/xreg_reg[630]  ( .D(\modmult_1/N1659 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[630] ) );
  DFF \modmult_1/xreg_reg[629]  ( .D(\modmult_1/N1658 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[629] ) );
  DFF \modmult_1/xreg_reg[628]  ( .D(\modmult_1/N1657 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[628] ) );
  DFF \modmult_1/xreg_reg[627]  ( .D(\modmult_1/N1656 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[627] ) );
  DFF \modmult_1/xreg_reg[626]  ( .D(\modmult_1/N1655 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[626] ) );
  DFF \modmult_1/xreg_reg[625]  ( .D(\modmult_1/N1654 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[625] ) );
  DFF \modmult_1/xreg_reg[624]  ( .D(\modmult_1/N1653 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[624] ) );
  DFF \modmult_1/xreg_reg[623]  ( .D(\modmult_1/N1652 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[623] ) );
  DFF \modmult_1/xreg_reg[622]  ( .D(\modmult_1/N1651 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[622] ) );
  DFF \modmult_1/xreg_reg[621]  ( .D(\modmult_1/N1650 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[621] ) );
  DFF \modmult_1/xreg_reg[620]  ( .D(\modmult_1/N1649 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[620] ) );
  DFF \modmult_1/xreg_reg[619]  ( .D(\modmult_1/N1648 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[619] ) );
  DFF \modmult_1/xreg_reg[618]  ( .D(\modmult_1/N1647 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[618] ) );
  DFF \modmult_1/xreg_reg[617]  ( .D(\modmult_1/N1646 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[617] ) );
  DFF \modmult_1/xreg_reg[616]  ( .D(\modmult_1/N1645 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[616] ) );
  DFF \modmult_1/xreg_reg[615]  ( .D(\modmult_1/N1644 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[615] ) );
  DFF \modmult_1/xreg_reg[614]  ( .D(\modmult_1/N1643 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[614] ) );
  DFF \modmult_1/xreg_reg[613]  ( .D(\modmult_1/N1642 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[613] ) );
  DFF \modmult_1/xreg_reg[612]  ( .D(\modmult_1/N1641 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[612] ) );
  DFF \modmult_1/xreg_reg[611]  ( .D(\modmult_1/N1640 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[611] ) );
  DFF \modmult_1/xreg_reg[610]  ( .D(\modmult_1/N1639 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[610] ) );
  DFF \modmult_1/xreg_reg[609]  ( .D(\modmult_1/N1638 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[609] ) );
  DFF \modmult_1/xreg_reg[608]  ( .D(\modmult_1/N1637 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[608] ) );
  DFF \modmult_1/xreg_reg[607]  ( .D(\modmult_1/N1636 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[607] ) );
  DFF \modmult_1/xreg_reg[606]  ( .D(\modmult_1/N1635 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[606] ) );
  DFF \modmult_1/xreg_reg[605]  ( .D(\modmult_1/N1634 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[605] ) );
  DFF \modmult_1/xreg_reg[604]  ( .D(\modmult_1/N1633 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[604] ) );
  DFF \modmult_1/xreg_reg[603]  ( .D(\modmult_1/N1632 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[603] ) );
  DFF \modmult_1/xreg_reg[602]  ( .D(\modmult_1/N1631 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[602] ) );
  DFF \modmult_1/xreg_reg[601]  ( .D(\modmult_1/N1630 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[601] ) );
  DFF \modmult_1/xreg_reg[600]  ( .D(\modmult_1/N1629 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[600] ) );
  DFF \modmult_1/xreg_reg[599]  ( .D(\modmult_1/N1628 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[599] ) );
  DFF \modmult_1/xreg_reg[598]  ( .D(\modmult_1/N1627 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[598] ) );
  DFF \modmult_1/xreg_reg[597]  ( .D(\modmult_1/N1626 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[597] ) );
  DFF \modmult_1/xreg_reg[596]  ( .D(\modmult_1/N1625 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[596] ) );
  DFF \modmult_1/xreg_reg[595]  ( .D(\modmult_1/N1624 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[595] ) );
  DFF \modmult_1/xreg_reg[594]  ( .D(\modmult_1/N1623 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[594] ) );
  DFF \modmult_1/xreg_reg[593]  ( .D(\modmult_1/N1622 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[593] ) );
  DFF \modmult_1/xreg_reg[592]  ( .D(\modmult_1/N1621 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[592] ) );
  DFF \modmult_1/xreg_reg[591]  ( .D(\modmult_1/N1620 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[591] ) );
  DFF \modmult_1/xreg_reg[590]  ( .D(\modmult_1/N1619 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[590] ) );
  DFF \modmult_1/xreg_reg[589]  ( .D(\modmult_1/N1618 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[589] ) );
  DFF \modmult_1/xreg_reg[588]  ( .D(\modmult_1/N1617 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[588] ) );
  DFF \modmult_1/xreg_reg[587]  ( .D(\modmult_1/N1616 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[587] ) );
  DFF \modmult_1/xreg_reg[586]  ( .D(\modmult_1/N1615 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[586] ) );
  DFF \modmult_1/xreg_reg[585]  ( .D(\modmult_1/N1614 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[585] ) );
  DFF \modmult_1/xreg_reg[584]  ( .D(\modmult_1/N1613 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[584] ) );
  DFF \modmult_1/xreg_reg[583]  ( .D(\modmult_1/N1612 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[583] ) );
  DFF \modmult_1/xreg_reg[582]  ( .D(\modmult_1/N1611 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[582] ) );
  DFF \modmult_1/xreg_reg[581]  ( .D(\modmult_1/N1610 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[581] ) );
  DFF \modmult_1/xreg_reg[580]  ( .D(\modmult_1/N1609 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[580] ) );
  DFF \modmult_1/xreg_reg[579]  ( .D(\modmult_1/N1608 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[579] ) );
  DFF \modmult_1/xreg_reg[578]  ( .D(\modmult_1/N1607 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[578] ) );
  DFF \modmult_1/xreg_reg[577]  ( .D(\modmult_1/N1606 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[577] ) );
  DFF \modmult_1/xreg_reg[576]  ( .D(\modmult_1/N1605 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[576] ) );
  DFF \modmult_1/xreg_reg[575]  ( .D(\modmult_1/N1604 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[575] ) );
  DFF \modmult_1/xreg_reg[574]  ( .D(\modmult_1/N1603 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[574] ) );
  DFF \modmult_1/xreg_reg[573]  ( .D(\modmult_1/N1602 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[573] ) );
  DFF \modmult_1/xreg_reg[572]  ( .D(\modmult_1/N1601 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[572] ) );
  DFF \modmult_1/xreg_reg[571]  ( .D(\modmult_1/N1600 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[571] ) );
  DFF \modmult_1/xreg_reg[570]  ( .D(\modmult_1/N1599 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[570] ) );
  DFF \modmult_1/xreg_reg[569]  ( .D(\modmult_1/N1598 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[569] ) );
  DFF \modmult_1/xreg_reg[568]  ( .D(\modmult_1/N1597 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[568] ) );
  DFF \modmult_1/xreg_reg[567]  ( .D(\modmult_1/N1596 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[567] ) );
  DFF \modmult_1/xreg_reg[566]  ( .D(\modmult_1/N1595 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[566] ) );
  DFF \modmult_1/xreg_reg[565]  ( .D(\modmult_1/N1594 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[565] ) );
  DFF \modmult_1/xreg_reg[564]  ( .D(\modmult_1/N1593 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[564] ) );
  DFF \modmult_1/xreg_reg[563]  ( .D(\modmult_1/N1592 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[563] ) );
  DFF \modmult_1/xreg_reg[562]  ( .D(\modmult_1/N1591 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[562] ) );
  DFF \modmult_1/xreg_reg[561]  ( .D(\modmult_1/N1590 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[561] ) );
  DFF \modmult_1/xreg_reg[560]  ( .D(\modmult_1/N1589 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[560] ) );
  DFF \modmult_1/xreg_reg[559]  ( .D(\modmult_1/N1588 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[559] ) );
  DFF \modmult_1/xreg_reg[558]  ( .D(\modmult_1/N1587 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[558] ) );
  DFF \modmult_1/xreg_reg[557]  ( .D(\modmult_1/N1586 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[557] ) );
  DFF \modmult_1/xreg_reg[556]  ( .D(\modmult_1/N1585 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[556] ) );
  DFF \modmult_1/xreg_reg[555]  ( .D(\modmult_1/N1584 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[555] ) );
  DFF \modmult_1/xreg_reg[554]  ( .D(\modmult_1/N1583 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[554] ) );
  DFF \modmult_1/xreg_reg[553]  ( .D(\modmult_1/N1582 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[553] ) );
  DFF \modmult_1/xreg_reg[552]  ( .D(\modmult_1/N1581 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[552] ) );
  DFF \modmult_1/xreg_reg[551]  ( .D(\modmult_1/N1580 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[551] ) );
  DFF \modmult_1/xreg_reg[550]  ( .D(\modmult_1/N1579 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[550] ) );
  DFF \modmult_1/xreg_reg[549]  ( .D(\modmult_1/N1578 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[549] ) );
  DFF \modmult_1/xreg_reg[548]  ( .D(\modmult_1/N1577 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[548] ) );
  DFF \modmult_1/xreg_reg[547]  ( .D(\modmult_1/N1576 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[547] ) );
  DFF \modmult_1/xreg_reg[546]  ( .D(\modmult_1/N1575 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[546] ) );
  DFF \modmult_1/xreg_reg[545]  ( .D(\modmult_1/N1574 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[545] ) );
  DFF \modmult_1/xreg_reg[544]  ( .D(\modmult_1/N1573 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[544] ) );
  DFF \modmult_1/xreg_reg[543]  ( .D(\modmult_1/N1572 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[543] ) );
  DFF \modmult_1/xreg_reg[542]  ( .D(\modmult_1/N1571 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[542] ) );
  DFF \modmult_1/xreg_reg[541]  ( .D(\modmult_1/N1570 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[541] ) );
  DFF \modmult_1/xreg_reg[540]  ( .D(\modmult_1/N1569 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[540] ) );
  DFF \modmult_1/xreg_reg[539]  ( .D(\modmult_1/N1568 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[539] ) );
  DFF \modmult_1/xreg_reg[538]  ( .D(\modmult_1/N1567 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[538] ) );
  DFF \modmult_1/xreg_reg[537]  ( .D(\modmult_1/N1566 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[537] ) );
  DFF \modmult_1/xreg_reg[536]  ( .D(\modmult_1/N1565 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[536] ) );
  DFF \modmult_1/xreg_reg[535]  ( .D(\modmult_1/N1564 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[535] ) );
  DFF \modmult_1/xreg_reg[534]  ( .D(\modmult_1/N1563 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[534] ) );
  DFF \modmult_1/xreg_reg[533]  ( .D(\modmult_1/N1562 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[533] ) );
  DFF \modmult_1/xreg_reg[532]  ( .D(\modmult_1/N1561 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[532] ) );
  DFF \modmult_1/xreg_reg[531]  ( .D(\modmult_1/N1560 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[531] ) );
  DFF \modmult_1/xreg_reg[530]  ( .D(\modmult_1/N1559 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[530] ) );
  DFF \modmult_1/xreg_reg[529]  ( .D(\modmult_1/N1558 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[529] ) );
  DFF \modmult_1/xreg_reg[528]  ( .D(\modmult_1/N1557 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[528] ) );
  DFF \modmult_1/xreg_reg[527]  ( .D(\modmult_1/N1556 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[527] ) );
  DFF \modmult_1/xreg_reg[526]  ( .D(\modmult_1/N1555 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[526] ) );
  DFF \modmult_1/xreg_reg[525]  ( .D(\modmult_1/N1554 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[525] ) );
  DFF \modmult_1/xreg_reg[524]  ( .D(\modmult_1/N1553 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[524] ) );
  DFF \modmult_1/xreg_reg[523]  ( .D(\modmult_1/N1552 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[523] ) );
  DFF \modmult_1/xreg_reg[522]  ( .D(\modmult_1/N1551 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[522] ) );
  DFF \modmult_1/xreg_reg[521]  ( .D(\modmult_1/N1550 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[521] ) );
  DFF \modmult_1/xreg_reg[520]  ( .D(\modmult_1/N1549 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[520] ) );
  DFF \modmult_1/xreg_reg[519]  ( .D(\modmult_1/N1548 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[519] ) );
  DFF \modmult_1/xreg_reg[518]  ( .D(\modmult_1/N1547 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[518] ) );
  DFF \modmult_1/xreg_reg[517]  ( .D(\modmult_1/N1546 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[517] ) );
  DFF \modmult_1/xreg_reg[516]  ( .D(\modmult_1/N1545 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[516] ) );
  DFF \modmult_1/xreg_reg[515]  ( .D(\modmult_1/N1544 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[515] ) );
  DFF \modmult_1/xreg_reg[514]  ( .D(\modmult_1/N1543 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[514] ) );
  DFF \modmult_1/xreg_reg[513]  ( .D(\modmult_1/N1542 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[513] ) );
  DFF \modmult_1/xreg_reg[512]  ( .D(\modmult_1/N1541 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[512] ) );
  DFF \modmult_1/xreg_reg[511]  ( .D(\modmult_1/N1540 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[511] ) );
  DFF \modmult_1/xreg_reg[510]  ( .D(\modmult_1/N1539 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[510] ) );
  DFF \modmult_1/xreg_reg[509]  ( .D(\modmult_1/N1538 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[509] ) );
  DFF \modmult_1/xreg_reg[508]  ( .D(\modmult_1/N1537 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[508] ) );
  DFF \modmult_1/xreg_reg[507]  ( .D(\modmult_1/N1536 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[507] ) );
  DFF \modmult_1/xreg_reg[506]  ( .D(\modmult_1/N1535 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[506] ) );
  DFF \modmult_1/xreg_reg[505]  ( .D(\modmult_1/N1534 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[505] ) );
  DFF \modmult_1/xreg_reg[504]  ( .D(\modmult_1/N1533 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[504] ) );
  DFF \modmult_1/xreg_reg[503]  ( .D(\modmult_1/N1532 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[503] ) );
  DFF \modmult_1/xreg_reg[502]  ( .D(\modmult_1/N1531 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[502] ) );
  DFF \modmult_1/xreg_reg[501]  ( .D(\modmult_1/N1530 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[501] ) );
  DFF \modmult_1/xreg_reg[500]  ( .D(\modmult_1/N1529 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[500] ) );
  DFF \modmult_1/xreg_reg[499]  ( .D(\modmult_1/N1528 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[499] ) );
  DFF \modmult_1/xreg_reg[498]  ( .D(\modmult_1/N1527 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[498] ) );
  DFF \modmult_1/xreg_reg[497]  ( .D(\modmult_1/N1526 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[497] ) );
  DFF \modmult_1/xreg_reg[496]  ( .D(\modmult_1/N1525 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[496] ) );
  DFF \modmult_1/xreg_reg[495]  ( .D(\modmult_1/N1524 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[495] ) );
  DFF \modmult_1/xreg_reg[494]  ( .D(\modmult_1/N1523 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[494] ) );
  DFF \modmult_1/xreg_reg[493]  ( .D(\modmult_1/N1522 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[493] ) );
  DFF \modmult_1/xreg_reg[492]  ( .D(\modmult_1/N1521 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[492] ) );
  DFF \modmult_1/xreg_reg[491]  ( .D(\modmult_1/N1520 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[491] ) );
  DFF \modmult_1/xreg_reg[490]  ( .D(\modmult_1/N1519 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[490] ) );
  DFF \modmult_1/xreg_reg[489]  ( .D(\modmult_1/N1518 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[489] ) );
  DFF \modmult_1/xreg_reg[488]  ( .D(\modmult_1/N1517 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[488] ) );
  DFF \modmult_1/xreg_reg[487]  ( .D(\modmult_1/N1516 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[487] ) );
  DFF \modmult_1/xreg_reg[486]  ( .D(\modmult_1/N1515 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[486] ) );
  DFF \modmult_1/xreg_reg[485]  ( .D(\modmult_1/N1514 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[485] ) );
  DFF \modmult_1/xreg_reg[484]  ( .D(\modmult_1/N1513 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[484] ) );
  DFF \modmult_1/xreg_reg[483]  ( .D(\modmult_1/N1512 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[483] ) );
  DFF \modmult_1/xreg_reg[482]  ( .D(\modmult_1/N1511 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[482] ) );
  DFF \modmult_1/xreg_reg[481]  ( .D(\modmult_1/N1510 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[481] ) );
  DFF \modmult_1/xreg_reg[480]  ( .D(\modmult_1/N1509 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[480] ) );
  DFF \modmult_1/xreg_reg[479]  ( .D(\modmult_1/N1508 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[479] ) );
  DFF \modmult_1/xreg_reg[478]  ( .D(\modmult_1/N1507 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[478] ) );
  DFF \modmult_1/xreg_reg[477]  ( .D(\modmult_1/N1506 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[477] ) );
  DFF \modmult_1/xreg_reg[476]  ( .D(\modmult_1/N1505 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[476] ) );
  DFF \modmult_1/xreg_reg[475]  ( .D(\modmult_1/N1504 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[475] ) );
  DFF \modmult_1/xreg_reg[474]  ( .D(\modmult_1/N1503 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[474] ) );
  DFF \modmult_1/xreg_reg[473]  ( .D(\modmult_1/N1502 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[473] ) );
  DFF \modmult_1/xreg_reg[472]  ( .D(\modmult_1/N1501 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[472] ) );
  DFF \modmult_1/xreg_reg[471]  ( .D(\modmult_1/N1500 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[471] ) );
  DFF \modmult_1/xreg_reg[470]  ( .D(\modmult_1/N1499 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[470] ) );
  DFF \modmult_1/xreg_reg[469]  ( .D(\modmult_1/N1498 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[469] ) );
  DFF \modmult_1/xreg_reg[468]  ( .D(\modmult_1/N1497 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[468] ) );
  DFF \modmult_1/xreg_reg[467]  ( .D(\modmult_1/N1496 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[467] ) );
  DFF \modmult_1/xreg_reg[466]  ( .D(\modmult_1/N1495 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[466] ) );
  DFF \modmult_1/xreg_reg[465]  ( .D(\modmult_1/N1494 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[465] ) );
  DFF \modmult_1/xreg_reg[464]  ( .D(\modmult_1/N1493 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[464] ) );
  DFF \modmult_1/xreg_reg[463]  ( .D(\modmult_1/N1492 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[463] ) );
  DFF \modmult_1/xreg_reg[462]  ( .D(\modmult_1/N1491 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[462] ) );
  DFF \modmult_1/xreg_reg[461]  ( .D(\modmult_1/N1490 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[461] ) );
  DFF \modmult_1/xreg_reg[460]  ( .D(\modmult_1/N1489 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[460] ) );
  DFF \modmult_1/xreg_reg[459]  ( .D(\modmult_1/N1488 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[459] ) );
  DFF \modmult_1/xreg_reg[458]  ( .D(\modmult_1/N1487 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[458] ) );
  DFF \modmult_1/xreg_reg[457]  ( .D(\modmult_1/N1486 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[457] ) );
  DFF \modmult_1/xreg_reg[456]  ( .D(\modmult_1/N1485 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[456] ) );
  DFF \modmult_1/xreg_reg[455]  ( .D(\modmult_1/N1484 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[455] ) );
  DFF \modmult_1/xreg_reg[454]  ( .D(\modmult_1/N1483 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[454] ) );
  DFF \modmult_1/xreg_reg[453]  ( .D(\modmult_1/N1482 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[453] ) );
  DFF \modmult_1/xreg_reg[452]  ( .D(\modmult_1/N1481 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[452] ) );
  DFF \modmult_1/xreg_reg[451]  ( .D(\modmult_1/N1480 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[451] ) );
  DFF \modmult_1/xreg_reg[450]  ( .D(\modmult_1/N1479 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[450] ) );
  DFF \modmult_1/xreg_reg[449]  ( .D(\modmult_1/N1478 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[449] ) );
  DFF \modmult_1/xreg_reg[448]  ( .D(\modmult_1/N1477 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[448] ) );
  DFF \modmult_1/xreg_reg[447]  ( .D(\modmult_1/N1476 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[447] ) );
  DFF \modmult_1/xreg_reg[446]  ( .D(\modmult_1/N1475 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[446] ) );
  DFF \modmult_1/xreg_reg[445]  ( .D(\modmult_1/N1474 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[445] ) );
  DFF \modmult_1/xreg_reg[444]  ( .D(\modmult_1/N1473 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[444] ) );
  DFF \modmult_1/xreg_reg[443]  ( .D(\modmult_1/N1472 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[443] ) );
  DFF \modmult_1/xreg_reg[442]  ( .D(\modmult_1/N1471 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[442] ) );
  DFF \modmult_1/xreg_reg[441]  ( .D(\modmult_1/N1470 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[441] ) );
  DFF \modmult_1/xreg_reg[440]  ( .D(\modmult_1/N1469 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[440] ) );
  DFF \modmult_1/xreg_reg[439]  ( .D(\modmult_1/N1468 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[439] ) );
  DFF \modmult_1/xreg_reg[438]  ( .D(\modmult_1/N1467 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[438] ) );
  DFF \modmult_1/xreg_reg[437]  ( .D(\modmult_1/N1466 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[437] ) );
  DFF \modmult_1/xreg_reg[436]  ( .D(\modmult_1/N1465 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[436] ) );
  DFF \modmult_1/xreg_reg[435]  ( .D(\modmult_1/N1464 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[435] ) );
  DFF \modmult_1/xreg_reg[434]  ( .D(\modmult_1/N1463 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[434] ) );
  DFF \modmult_1/xreg_reg[433]  ( .D(\modmult_1/N1462 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[433] ) );
  DFF \modmult_1/xreg_reg[432]  ( .D(\modmult_1/N1461 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[432] ) );
  DFF \modmult_1/xreg_reg[431]  ( .D(\modmult_1/N1460 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[431] ) );
  DFF \modmult_1/xreg_reg[430]  ( .D(\modmult_1/N1459 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[430] ) );
  DFF \modmult_1/xreg_reg[429]  ( .D(\modmult_1/N1458 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[429] ) );
  DFF \modmult_1/xreg_reg[428]  ( .D(\modmult_1/N1457 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[428] ) );
  DFF \modmult_1/xreg_reg[427]  ( .D(\modmult_1/N1456 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[427] ) );
  DFF \modmult_1/xreg_reg[426]  ( .D(\modmult_1/N1455 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[426] ) );
  DFF \modmult_1/xreg_reg[425]  ( .D(\modmult_1/N1454 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[425] ) );
  DFF \modmult_1/xreg_reg[424]  ( .D(\modmult_1/N1453 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[424] ) );
  DFF \modmult_1/xreg_reg[423]  ( .D(\modmult_1/N1452 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[423] ) );
  DFF \modmult_1/xreg_reg[422]  ( .D(\modmult_1/N1451 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[422] ) );
  DFF \modmult_1/xreg_reg[421]  ( .D(\modmult_1/N1450 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[421] ) );
  DFF \modmult_1/xreg_reg[420]  ( .D(\modmult_1/N1449 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[420] ) );
  DFF \modmult_1/xreg_reg[419]  ( .D(\modmult_1/N1448 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[419] ) );
  DFF \modmult_1/xreg_reg[418]  ( .D(\modmult_1/N1447 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[418] ) );
  DFF \modmult_1/xreg_reg[417]  ( .D(\modmult_1/N1446 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[417] ) );
  DFF \modmult_1/xreg_reg[416]  ( .D(\modmult_1/N1445 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[416] ) );
  DFF \modmult_1/xreg_reg[415]  ( .D(\modmult_1/N1444 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[415] ) );
  DFF \modmult_1/xreg_reg[414]  ( .D(\modmult_1/N1443 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[414] ) );
  DFF \modmult_1/xreg_reg[413]  ( .D(\modmult_1/N1442 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[413] ) );
  DFF \modmult_1/xreg_reg[412]  ( .D(\modmult_1/N1441 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[412] ) );
  DFF \modmult_1/xreg_reg[411]  ( .D(\modmult_1/N1440 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[411] ) );
  DFF \modmult_1/xreg_reg[410]  ( .D(\modmult_1/N1439 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[410] ) );
  DFF \modmult_1/xreg_reg[409]  ( .D(\modmult_1/N1438 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[409] ) );
  DFF \modmult_1/xreg_reg[408]  ( .D(\modmult_1/N1437 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[408] ) );
  DFF \modmult_1/xreg_reg[407]  ( .D(\modmult_1/N1436 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[407] ) );
  DFF \modmult_1/xreg_reg[406]  ( .D(\modmult_1/N1435 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[406] ) );
  DFF \modmult_1/xreg_reg[405]  ( .D(\modmult_1/N1434 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[405] ) );
  DFF \modmult_1/xreg_reg[404]  ( .D(\modmult_1/N1433 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[404] ) );
  DFF \modmult_1/xreg_reg[403]  ( .D(\modmult_1/N1432 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[403] ) );
  DFF \modmult_1/xreg_reg[402]  ( .D(\modmult_1/N1431 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[402] ) );
  DFF \modmult_1/xreg_reg[401]  ( .D(\modmult_1/N1430 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[401] ) );
  DFF \modmult_1/xreg_reg[400]  ( .D(\modmult_1/N1429 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[400] ) );
  DFF \modmult_1/xreg_reg[399]  ( .D(\modmult_1/N1428 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[399] ) );
  DFF \modmult_1/xreg_reg[398]  ( .D(\modmult_1/N1427 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[398] ) );
  DFF \modmult_1/xreg_reg[397]  ( .D(\modmult_1/N1426 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[397] ) );
  DFF \modmult_1/xreg_reg[396]  ( .D(\modmult_1/N1425 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[396] ) );
  DFF \modmult_1/xreg_reg[395]  ( .D(\modmult_1/N1424 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[395] ) );
  DFF \modmult_1/xreg_reg[394]  ( .D(\modmult_1/N1423 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[394] ) );
  DFF \modmult_1/xreg_reg[393]  ( .D(\modmult_1/N1422 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[393] ) );
  DFF \modmult_1/xreg_reg[392]  ( .D(\modmult_1/N1421 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[392] ) );
  DFF \modmult_1/xreg_reg[391]  ( .D(\modmult_1/N1420 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[391] ) );
  DFF \modmult_1/xreg_reg[390]  ( .D(\modmult_1/N1419 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[390] ) );
  DFF \modmult_1/xreg_reg[389]  ( .D(\modmult_1/N1418 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[389] ) );
  DFF \modmult_1/xreg_reg[388]  ( .D(\modmult_1/N1417 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[388] ) );
  DFF \modmult_1/xreg_reg[387]  ( .D(\modmult_1/N1416 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[387] ) );
  DFF \modmult_1/xreg_reg[386]  ( .D(\modmult_1/N1415 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[386] ) );
  DFF \modmult_1/xreg_reg[385]  ( .D(\modmult_1/N1414 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[385] ) );
  DFF \modmult_1/xreg_reg[384]  ( .D(\modmult_1/N1413 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[384] ) );
  DFF \modmult_1/xreg_reg[383]  ( .D(\modmult_1/N1412 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[383] ) );
  DFF \modmult_1/xreg_reg[382]  ( .D(\modmult_1/N1411 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[382] ) );
  DFF \modmult_1/xreg_reg[381]  ( .D(\modmult_1/N1410 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[381] ) );
  DFF \modmult_1/xreg_reg[380]  ( .D(\modmult_1/N1409 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[380] ) );
  DFF \modmult_1/xreg_reg[379]  ( .D(\modmult_1/N1408 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[379] ) );
  DFF \modmult_1/xreg_reg[378]  ( .D(\modmult_1/N1407 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[378] ) );
  DFF \modmult_1/xreg_reg[377]  ( .D(\modmult_1/N1406 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[377] ) );
  DFF \modmult_1/xreg_reg[376]  ( .D(\modmult_1/N1405 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[376] ) );
  DFF \modmult_1/xreg_reg[375]  ( .D(\modmult_1/N1404 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[375] ) );
  DFF \modmult_1/xreg_reg[374]  ( .D(\modmult_1/N1403 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[374] ) );
  DFF \modmult_1/xreg_reg[373]  ( .D(\modmult_1/N1402 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[373] ) );
  DFF \modmult_1/xreg_reg[372]  ( .D(\modmult_1/N1401 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[372] ) );
  DFF \modmult_1/xreg_reg[371]  ( .D(\modmult_1/N1400 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[371] ) );
  DFF \modmult_1/xreg_reg[370]  ( .D(\modmult_1/N1399 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[370] ) );
  DFF \modmult_1/xreg_reg[369]  ( .D(\modmult_1/N1398 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[369] ) );
  DFF \modmult_1/xreg_reg[368]  ( .D(\modmult_1/N1397 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[368] ) );
  DFF \modmult_1/xreg_reg[367]  ( .D(\modmult_1/N1396 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[367] ) );
  DFF \modmult_1/xreg_reg[366]  ( .D(\modmult_1/N1395 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[366] ) );
  DFF \modmult_1/xreg_reg[365]  ( .D(\modmult_1/N1394 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[365] ) );
  DFF \modmult_1/xreg_reg[364]  ( .D(\modmult_1/N1393 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[364] ) );
  DFF \modmult_1/xreg_reg[363]  ( .D(\modmult_1/N1392 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[363] ) );
  DFF \modmult_1/xreg_reg[362]  ( .D(\modmult_1/N1391 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[362] ) );
  DFF \modmult_1/xreg_reg[361]  ( .D(\modmult_1/N1390 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[361] ) );
  DFF \modmult_1/xreg_reg[360]  ( .D(\modmult_1/N1389 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[360] ) );
  DFF \modmult_1/xreg_reg[359]  ( .D(\modmult_1/N1388 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[359] ) );
  DFF \modmult_1/xreg_reg[358]  ( .D(\modmult_1/N1387 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[358] ) );
  DFF \modmult_1/xreg_reg[357]  ( .D(\modmult_1/N1386 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[357] ) );
  DFF \modmult_1/xreg_reg[356]  ( .D(\modmult_1/N1385 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[356] ) );
  DFF \modmult_1/xreg_reg[355]  ( .D(\modmult_1/N1384 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[355] ) );
  DFF \modmult_1/xreg_reg[354]  ( .D(\modmult_1/N1383 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[354] ) );
  DFF \modmult_1/xreg_reg[353]  ( .D(\modmult_1/N1382 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[353] ) );
  DFF \modmult_1/xreg_reg[352]  ( .D(\modmult_1/N1381 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[352] ) );
  DFF \modmult_1/xreg_reg[351]  ( .D(\modmult_1/N1380 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[351] ) );
  DFF \modmult_1/xreg_reg[350]  ( .D(\modmult_1/N1379 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[350] ) );
  DFF \modmult_1/xreg_reg[349]  ( .D(\modmult_1/N1378 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[349] ) );
  DFF \modmult_1/xreg_reg[348]  ( .D(\modmult_1/N1377 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[348] ) );
  DFF \modmult_1/xreg_reg[347]  ( .D(\modmult_1/N1376 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[347] ) );
  DFF \modmult_1/xreg_reg[346]  ( .D(\modmult_1/N1375 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[346] ) );
  DFF \modmult_1/xreg_reg[345]  ( .D(\modmult_1/N1374 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[345] ) );
  DFF \modmult_1/xreg_reg[344]  ( .D(\modmult_1/N1373 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[344] ) );
  DFF \modmult_1/xreg_reg[343]  ( .D(\modmult_1/N1372 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[343] ) );
  DFF \modmult_1/xreg_reg[342]  ( .D(\modmult_1/N1371 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[342] ) );
  DFF \modmult_1/xreg_reg[341]  ( .D(\modmult_1/N1370 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[341] ) );
  DFF \modmult_1/xreg_reg[340]  ( .D(\modmult_1/N1369 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[340] ) );
  DFF \modmult_1/xreg_reg[339]  ( .D(\modmult_1/N1368 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[339] ) );
  DFF \modmult_1/xreg_reg[338]  ( .D(\modmult_1/N1367 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[338] ) );
  DFF \modmult_1/xreg_reg[337]  ( .D(\modmult_1/N1366 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[337] ) );
  DFF \modmult_1/xreg_reg[336]  ( .D(\modmult_1/N1365 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[336] ) );
  DFF \modmult_1/xreg_reg[335]  ( .D(\modmult_1/N1364 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[335] ) );
  DFF \modmult_1/xreg_reg[334]  ( .D(\modmult_1/N1363 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[334] ) );
  DFF \modmult_1/xreg_reg[333]  ( .D(\modmult_1/N1362 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[333] ) );
  DFF \modmult_1/xreg_reg[332]  ( .D(\modmult_1/N1361 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[332] ) );
  DFF \modmult_1/xreg_reg[331]  ( .D(\modmult_1/N1360 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[331] ) );
  DFF \modmult_1/xreg_reg[330]  ( .D(\modmult_1/N1359 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[330] ) );
  DFF \modmult_1/xreg_reg[329]  ( .D(\modmult_1/N1358 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[329] ) );
  DFF \modmult_1/xreg_reg[328]  ( .D(\modmult_1/N1357 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[328] ) );
  DFF \modmult_1/xreg_reg[327]  ( .D(\modmult_1/N1356 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[327] ) );
  DFF \modmult_1/xreg_reg[326]  ( .D(\modmult_1/N1355 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[326] ) );
  DFF \modmult_1/xreg_reg[325]  ( .D(\modmult_1/N1354 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[325] ) );
  DFF \modmult_1/xreg_reg[324]  ( .D(\modmult_1/N1353 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[324] ) );
  DFF \modmult_1/xreg_reg[323]  ( .D(\modmult_1/N1352 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[323] ) );
  DFF \modmult_1/xreg_reg[322]  ( .D(\modmult_1/N1351 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[322] ) );
  DFF \modmult_1/xreg_reg[321]  ( .D(\modmult_1/N1350 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[321] ) );
  DFF \modmult_1/xreg_reg[320]  ( .D(\modmult_1/N1349 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[320] ) );
  DFF \modmult_1/xreg_reg[319]  ( .D(\modmult_1/N1348 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[319] ) );
  DFF \modmult_1/xreg_reg[318]  ( .D(\modmult_1/N1347 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[318] ) );
  DFF \modmult_1/xreg_reg[317]  ( .D(\modmult_1/N1346 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[317] ) );
  DFF \modmult_1/xreg_reg[316]  ( .D(\modmult_1/N1345 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[316] ) );
  DFF \modmult_1/xreg_reg[315]  ( .D(\modmult_1/N1344 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[315] ) );
  DFF \modmult_1/xreg_reg[314]  ( .D(\modmult_1/N1343 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[314] ) );
  DFF \modmult_1/xreg_reg[313]  ( .D(\modmult_1/N1342 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[313] ) );
  DFF \modmult_1/xreg_reg[312]  ( .D(\modmult_1/N1341 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[312] ) );
  DFF \modmult_1/xreg_reg[311]  ( .D(\modmult_1/N1340 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[311] ) );
  DFF \modmult_1/xreg_reg[310]  ( .D(\modmult_1/N1339 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[310] ) );
  DFF \modmult_1/xreg_reg[309]  ( .D(\modmult_1/N1338 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[309] ) );
  DFF \modmult_1/xreg_reg[308]  ( .D(\modmult_1/N1337 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[308] ) );
  DFF \modmult_1/xreg_reg[307]  ( .D(\modmult_1/N1336 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[307] ) );
  DFF \modmult_1/xreg_reg[306]  ( .D(\modmult_1/N1335 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[306] ) );
  DFF \modmult_1/xreg_reg[305]  ( .D(\modmult_1/N1334 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[305] ) );
  DFF \modmult_1/xreg_reg[304]  ( .D(\modmult_1/N1333 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[304] ) );
  DFF \modmult_1/xreg_reg[303]  ( .D(\modmult_1/N1332 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[303] ) );
  DFF \modmult_1/xreg_reg[302]  ( .D(\modmult_1/N1331 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[302] ) );
  DFF \modmult_1/xreg_reg[301]  ( .D(\modmult_1/N1330 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[301] ) );
  DFF \modmult_1/xreg_reg[300]  ( .D(\modmult_1/N1329 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[300] ) );
  DFF \modmult_1/xreg_reg[299]  ( .D(\modmult_1/N1328 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[299] ) );
  DFF \modmult_1/xreg_reg[298]  ( .D(\modmult_1/N1327 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[298] ) );
  DFF \modmult_1/xreg_reg[297]  ( .D(\modmult_1/N1326 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[297] ) );
  DFF \modmult_1/xreg_reg[296]  ( .D(\modmult_1/N1325 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[296] ) );
  DFF \modmult_1/xreg_reg[295]  ( .D(\modmult_1/N1324 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[295] ) );
  DFF \modmult_1/xreg_reg[294]  ( .D(\modmult_1/N1323 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[294] ) );
  DFF \modmult_1/xreg_reg[293]  ( .D(\modmult_1/N1322 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[293] ) );
  DFF \modmult_1/xreg_reg[292]  ( .D(\modmult_1/N1321 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[292] ) );
  DFF \modmult_1/xreg_reg[291]  ( .D(\modmult_1/N1320 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[291] ) );
  DFF \modmult_1/xreg_reg[290]  ( .D(\modmult_1/N1319 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[290] ) );
  DFF \modmult_1/xreg_reg[289]  ( .D(\modmult_1/N1318 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[289] ) );
  DFF \modmult_1/xreg_reg[288]  ( .D(\modmult_1/N1317 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[288] ) );
  DFF \modmult_1/xreg_reg[287]  ( .D(\modmult_1/N1316 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[287] ) );
  DFF \modmult_1/xreg_reg[286]  ( .D(\modmult_1/N1315 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[286] ) );
  DFF \modmult_1/xreg_reg[285]  ( .D(\modmult_1/N1314 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[285] ) );
  DFF \modmult_1/xreg_reg[284]  ( .D(\modmult_1/N1313 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[284] ) );
  DFF \modmult_1/xreg_reg[283]  ( .D(\modmult_1/N1312 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[283] ) );
  DFF \modmult_1/xreg_reg[282]  ( .D(\modmult_1/N1311 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[282] ) );
  DFF \modmult_1/xreg_reg[281]  ( .D(\modmult_1/N1310 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[281] ) );
  DFF \modmult_1/xreg_reg[280]  ( .D(\modmult_1/N1309 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[280] ) );
  DFF \modmult_1/xreg_reg[279]  ( .D(\modmult_1/N1308 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[279] ) );
  DFF \modmult_1/xreg_reg[278]  ( .D(\modmult_1/N1307 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[278] ) );
  DFF \modmult_1/xreg_reg[277]  ( .D(\modmult_1/N1306 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[277] ) );
  DFF \modmult_1/xreg_reg[276]  ( .D(\modmult_1/N1305 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[276] ) );
  DFF \modmult_1/xreg_reg[275]  ( .D(\modmult_1/N1304 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[275] ) );
  DFF \modmult_1/xreg_reg[274]  ( .D(\modmult_1/N1303 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[274] ) );
  DFF \modmult_1/xreg_reg[273]  ( .D(\modmult_1/N1302 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[273] ) );
  DFF \modmult_1/xreg_reg[272]  ( .D(\modmult_1/N1301 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[272] ) );
  DFF \modmult_1/xreg_reg[271]  ( .D(\modmult_1/N1300 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[271] ) );
  DFF \modmult_1/xreg_reg[270]  ( .D(\modmult_1/N1299 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[270] ) );
  DFF \modmult_1/xreg_reg[269]  ( .D(\modmult_1/N1298 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[269] ) );
  DFF \modmult_1/xreg_reg[268]  ( .D(\modmult_1/N1297 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[268] ) );
  DFF \modmult_1/xreg_reg[267]  ( .D(\modmult_1/N1296 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[267] ) );
  DFF \modmult_1/xreg_reg[266]  ( .D(\modmult_1/N1295 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[266] ) );
  DFF \modmult_1/xreg_reg[265]  ( .D(\modmult_1/N1294 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[265] ) );
  DFF \modmult_1/xreg_reg[264]  ( .D(\modmult_1/N1293 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[264] ) );
  DFF \modmult_1/xreg_reg[263]  ( .D(\modmult_1/N1292 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[263] ) );
  DFF \modmult_1/xreg_reg[262]  ( .D(\modmult_1/N1291 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[262] ) );
  DFF \modmult_1/xreg_reg[261]  ( .D(\modmult_1/N1290 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[261] ) );
  DFF \modmult_1/xreg_reg[260]  ( .D(\modmult_1/N1289 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[260] ) );
  DFF \modmult_1/xreg_reg[259]  ( .D(\modmult_1/N1288 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[259] ) );
  DFF \modmult_1/xreg_reg[258]  ( .D(\modmult_1/N1287 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[258] ) );
  DFF \modmult_1/xreg_reg[257]  ( .D(\modmult_1/N1286 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[257] ) );
  DFF \modmult_1/xreg_reg[256]  ( .D(\modmult_1/N1285 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[256] ) );
  DFF \modmult_1/xreg_reg[255]  ( .D(\modmult_1/N1284 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[255] ) );
  DFF \modmult_1/xreg_reg[254]  ( .D(\modmult_1/N1283 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[254] ) );
  DFF \modmult_1/xreg_reg[253]  ( .D(\modmult_1/N1282 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[253] ) );
  DFF \modmult_1/xreg_reg[252]  ( .D(\modmult_1/N1281 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[252] ) );
  DFF \modmult_1/xreg_reg[251]  ( .D(\modmult_1/N1280 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[251] ) );
  DFF \modmult_1/xreg_reg[250]  ( .D(\modmult_1/N1279 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[250] ) );
  DFF \modmult_1/xreg_reg[249]  ( .D(\modmult_1/N1278 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[249] ) );
  DFF \modmult_1/xreg_reg[248]  ( .D(\modmult_1/N1277 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[248] ) );
  DFF \modmult_1/xreg_reg[247]  ( .D(\modmult_1/N1276 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[247] ) );
  DFF \modmult_1/xreg_reg[246]  ( .D(\modmult_1/N1275 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[246] ) );
  DFF \modmult_1/xreg_reg[245]  ( .D(\modmult_1/N1274 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[245] ) );
  DFF \modmult_1/xreg_reg[244]  ( .D(\modmult_1/N1273 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[244] ) );
  DFF \modmult_1/xreg_reg[243]  ( .D(\modmult_1/N1272 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[243] ) );
  DFF \modmult_1/xreg_reg[242]  ( .D(\modmult_1/N1271 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[242] ) );
  DFF \modmult_1/xreg_reg[241]  ( .D(\modmult_1/N1270 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[241] ) );
  DFF \modmult_1/xreg_reg[240]  ( .D(\modmult_1/N1269 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[240] ) );
  DFF \modmult_1/xreg_reg[239]  ( .D(\modmult_1/N1268 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[239] ) );
  DFF \modmult_1/xreg_reg[238]  ( .D(\modmult_1/N1267 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[238] ) );
  DFF \modmult_1/xreg_reg[237]  ( .D(\modmult_1/N1266 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[237] ) );
  DFF \modmult_1/xreg_reg[236]  ( .D(\modmult_1/N1265 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[236] ) );
  DFF \modmult_1/xreg_reg[235]  ( .D(\modmult_1/N1264 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[235] ) );
  DFF \modmult_1/xreg_reg[234]  ( .D(\modmult_1/N1263 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[234] ) );
  DFF \modmult_1/xreg_reg[233]  ( .D(\modmult_1/N1262 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[233] ) );
  DFF \modmult_1/xreg_reg[232]  ( .D(\modmult_1/N1261 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[232] ) );
  DFF \modmult_1/xreg_reg[231]  ( .D(\modmult_1/N1260 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[231] ) );
  DFF \modmult_1/xreg_reg[230]  ( .D(\modmult_1/N1259 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[230] ) );
  DFF \modmult_1/xreg_reg[229]  ( .D(\modmult_1/N1258 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[229] ) );
  DFF \modmult_1/xreg_reg[228]  ( .D(\modmult_1/N1257 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[228] ) );
  DFF \modmult_1/xreg_reg[227]  ( .D(\modmult_1/N1256 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[227] ) );
  DFF \modmult_1/xreg_reg[226]  ( .D(\modmult_1/N1255 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[226] ) );
  DFF \modmult_1/xreg_reg[225]  ( .D(\modmult_1/N1254 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[225] ) );
  DFF \modmult_1/xreg_reg[224]  ( .D(\modmult_1/N1253 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[224] ) );
  DFF \modmult_1/xreg_reg[223]  ( .D(\modmult_1/N1252 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[223] ) );
  DFF \modmult_1/xreg_reg[222]  ( .D(\modmult_1/N1251 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[222] ) );
  DFF \modmult_1/xreg_reg[221]  ( .D(\modmult_1/N1250 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[221] ) );
  DFF \modmult_1/xreg_reg[220]  ( .D(\modmult_1/N1249 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[220] ) );
  DFF \modmult_1/xreg_reg[219]  ( .D(\modmult_1/N1248 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[219] ) );
  DFF \modmult_1/xreg_reg[218]  ( .D(\modmult_1/N1247 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[218] ) );
  DFF \modmult_1/xreg_reg[217]  ( .D(\modmult_1/N1246 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[217] ) );
  DFF \modmult_1/xreg_reg[216]  ( .D(\modmult_1/N1245 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[216] ) );
  DFF \modmult_1/xreg_reg[215]  ( .D(\modmult_1/N1244 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[215] ) );
  DFF \modmult_1/xreg_reg[214]  ( .D(\modmult_1/N1243 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[214] ) );
  DFF \modmult_1/xreg_reg[213]  ( .D(\modmult_1/N1242 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[213] ) );
  DFF \modmult_1/xreg_reg[212]  ( .D(\modmult_1/N1241 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[212] ) );
  DFF \modmult_1/xreg_reg[211]  ( .D(\modmult_1/N1240 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[211] ) );
  DFF \modmult_1/xreg_reg[210]  ( .D(\modmult_1/N1239 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[210] ) );
  DFF \modmult_1/xreg_reg[209]  ( .D(\modmult_1/N1238 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[209] ) );
  DFF \modmult_1/xreg_reg[208]  ( .D(\modmult_1/N1237 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[208] ) );
  DFF \modmult_1/xreg_reg[207]  ( .D(\modmult_1/N1236 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[207] ) );
  DFF \modmult_1/xreg_reg[206]  ( .D(\modmult_1/N1235 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[206] ) );
  DFF \modmult_1/xreg_reg[205]  ( .D(\modmult_1/N1234 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[205] ) );
  DFF \modmult_1/xreg_reg[204]  ( .D(\modmult_1/N1233 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[204] ) );
  DFF \modmult_1/xreg_reg[203]  ( .D(\modmult_1/N1232 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[203] ) );
  DFF \modmult_1/xreg_reg[202]  ( .D(\modmult_1/N1231 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[202] ) );
  DFF \modmult_1/xreg_reg[201]  ( .D(\modmult_1/N1230 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[201] ) );
  DFF \modmult_1/xreg_reg[200]  ( .D(\modmult_1/N1229 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[200] ) );
  DFF \modmult_1/xreg_reg[199]  ( .D(\modmult_1/N1228 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[199] ) );
  DFF \modmult_1/xreg_reg[198]  ( .D(\modmult_1/N1227 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[198] ) );
  DFF \modmult_1/xreg_reg[197]  ( .D(\modmult_1/N1226 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[197] ) );
  DFF \modmult_1/xreg_reg[196]  ( .D(\modmult_1/N1225 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[196] ) );
  DFF \modmult_1/xreg_reg[195]  ( .D(\modmult_1/N1224 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[195] ) );
  DFF \modmult_1/xreg_reg[194]  ( .D(\modmult_1/N1223 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[194] ) );
  DFF \modmult_1/xreg_reg[193]  ( .D(\modmult_1/N1222 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[193] ) );
  DFF \modmult_1/xreg_reg[192]  ( .D(\modmult_1/N1221 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[192] ) );
  DFF \modmult_1/xreg_reg[191]  ( .D(\modmult_1/N1220 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[191] ) );
  DFF \modmult_1/xreg_reg[190]  ( .D(\modmult_1/N1219 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[190] ) );
  DFF \modmult_1/xreg_reg[189]  ( .D(\modmult_1/N1218 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[189] ) );
  DFF \modmult_1/xreg_reg[188]  ( .D(\modmult_1/N1217 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[188] ) );
  DFF \modmult_1/xreg_reg[187]  ( .D(\modmult_1/N1216 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[187] ) );
  DFF \modmult_1/xreg_reg[186]  ( .D(\modmult_1/N1215 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[186] ) );
  DFF \modmult_1/xreg_reg[185]  ( .D(\modmult_1/N1214 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[185] ) );
  DFF \modmult_1/xreg_reg[184]  ( .D(\modmult_1/N1213 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[184] ) );
  DFF \modmult_1/xreg_reg[183]  ( .D(\modmult_1/N1212 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[183] ) );
  DFF \modmult_1/xreg_reg[182]  ( .D(\modmult_1/N1211 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[182] ) );
  DFF \modmult_1/xreg_reg[181]  ( .D(\modmult_1/N1210 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[181] ) );
  DFF \modmult_1/xreg_reg[180]  ( .D(\modmult_1/N1209 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[180] ) );
  DFF \modmult_1/xreg_reg[179]  ( .D(\modmult_1/N1208 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[179] ) );
  DFF \modmult_1/xreg_reg[178]  ( .D(\modmult_1/N1207 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[178] ) );
  DFF \modmult_1/xreg_reg[177]  ( .D(\modmult_1/N1206 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[177] ) );
  DFF \modmult_1/xreg_reg[176]  ( .D(\modmult_1/N1205 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[176] ) );
  DFF \modmult_1/xreg_reg[175]  ( .D(\modmult_1/N1204 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[175] ) );
  DFF \modmult_1/xreg_reg[174]  ( .D(\modmult_1/N1203 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[174] ) );
  DFF \modmult_1/xreg_reg[173]  ( .D(\modmult_1/N1202 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[173] ) );
  DFF \modmult_1/xreg_reg[172]  ( .D(\modmult_1/N1201 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[172] ) );
  DFF \modmult_1/xreg_reg[171]  ( .D(\modmult_1/N1200 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[171] ) );
  DFF \modmult_1/xreg_reg[170]  ( .D(\modmult_1/N1199 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[170] ) );
  DFF \modmult_1/xreg_reg[169]  ( .D(\modmult_1/N1198 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[169] ) );
  DFF \modmult_1/xreg_reg[168]  ( .D(\modmult_1/N1197 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[168] ) );
  DFF \modmult_1/xreg_reg[167]  ( .D(\modmult_1/N1196 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[167] ) );
  DFF \modmult_1/xreg_reg[166]  ( .D(\modmult_1/N1195 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[166] ) );
  DFF \modmult_1/xreg_reg[165]  ( .D(\modmult_1/N1194 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[165] ) );
  DFF \modmult_1/xreg_reg[164]  ( .D(\modmult_1/N1193 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[164] ) );
  DFF \modmult_1/xreg_reg[163]  ( .D(\modmult_1/N1192 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[163] ) );
  DFF \modmult_1/xreg_reg[162]  ( .D(\modmult_1/N1191 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[162] ) );
  DFF \modmult_1/xreg_reg[161]  ( .D(\modmult_1/N1190 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[161] ) );
  DFF \modmult_1/xreg_reg[160]  ( .D(\modmult_1/N1189 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[160] ) );
  DFF \modmult_1/xreg_reg[159]  ( .D(\modmult_1/N1188 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[159] ) );
  DFF \modmult_1/xreg_reg[158]  ( .D(\modmult_1/N1187 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[158] ) );
  DFF \modmult_1/xreg_reg[157]  ( .D(\modmult_1/N1186 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[157] ) );
  DFF \modmult_1/xreg_reg[156]  ( .D(\modmult_1/N1185 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[156] ) );
  DFF \modmult_1/xreg_reg[155]  ( .D(\modmult_1/N1184 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[155] ) );
  DFF \modmult_1/xreg_reg[154]  ( .D(\modmult_1/N1183 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[154] ) );
  DFF \modmult_1/xreg_reg[153]  ( .D(\modmult_1/N1182 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[153] ) );
  DFF \modmult_1/xreg_reg[152]  ( .D(\modmult_1/N1181 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[152] ) );
  DFF \modmult_1/xreg_reg[151]  ( .D(\modmult_1/N1180 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[151] ) );
  DFF \modmult_1/xreg_reg[150]  ( .D(\modmult_1/N1179 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[150] ) );
  DFF \modmult_1/xreg_reg[149]  ( .D(\modmult_1/N1178 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[149] ) );
  DFF \modmult_1/xreg_reg[148]  ( .D(\modmult_1/N1177 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[148] ) );
  DFF \modmult_1/xreg_reg[147]  ( .D(\modmult_1/N1176 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[147] ) );
  DFF \modmult_1/xreg_reg[146]  ( .D(\modmult_1/N1175 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[146] ) );
  DFF \modmult_1/xreg_reg[145]  ( .D(\modmult_1/N1174 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[145] ) );
  DFF \modmult_1/xreg_reg[144]  ( .D(\modmult_1/N1173 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[144] ) );
  DFF \modmult_1/xreg_reg[143]  ( .D(\modmult_1/N1172 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[143] ) );
  DFF \modmult_1/xreg_reg[142]  ( .D(\modmult_1/N1171 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[142] ) );
  DFF \modmult_1/xreg_reg[141]  ( .D(\modmult_1/N1170 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[141] ) );
  DFF \modmult_1/xreg_reg[140]  ( .D(\modmult_1/N1169 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[140] ) );
  DFF \modmult_1/xreg_reg[139]  ( .D(\modmult_1/N1168 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[139] ) );
  DFF \modmult_1/xreg_reg[138]  ( .D(\modmult_1/N1167 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[138] ) );
  DFF \modmult_1/xreg_reg[137]  ( .D(\modmult_1/N1166 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[137] ) );
  DFF \modmult_1/xreg_reg[136]  ( .D(\modmult_1/N1165 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[136] ) );
  DFF \modmult_1/xreg_reg[135]  ( .D(\modmult_1/N1164 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[135] ) );
  DFF \modmult_1/xreg_reg[134]  ( .D(\modmult_1/N1163 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[134] ) );
  DFF \modmult_1/xreg_reg[133]  ( .D(\modmult_1/N1162 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[133] ) );
  DFF \modmult_1/xreg_reg[132]  ( .D(\modmult_1/N1161 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[132] ) );
  DFF \modmult_1/xreg_reg[131]  ( .D(\modmult_1/N1160 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[131] ) );
  DFF \modmult_1/xreg_reg[130]  ( .D(\modmult_1/N1159 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[130] ) );
  DFF \modmult_1/xreg_reg[129]  ( .D(\modmult_1/N1158 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[129] ) );
  DFF \modmult_1/xreg_reg[128]  ( .D(\modmult_1/N1157 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[128] ) );
  DFF \modmult_1/xreg_reg[127]  ( .D(\modmult_1/N1156 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[127] ) );
  DFF \modmult_1/xreg_reg[126]  ( .D(\modmult_1/N1155 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[126] ) );
  DFF \modmult_1/xreg_reg[125]  ( .D(\modmult_1/N1154 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[125] ) );
  DFF \modmult_1/xreg_reg[124]  ( .D(\modmult_1/N1153 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[124] ) );
  DFF \modmult_1/xreg_reg[123]  ( .D(\modmult_1/N1152 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[123] ) );
  DFF \modmult_1/xreg_reg[122]  ( .D(\modmult_1/N1151 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[122] ) );
  DFF \modmult_1/xreg_reg[121]  ( .D(\modmult_1/N1150 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[121] ) );
  DFF \modmult_1/xreg_reg[120]  ( .D(\modmult_1/N1149 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[120] ) );
  DFF \modmult_1/xreg_reg[119]  ( .D(\modmult_1/N1148 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[119] ) );
  DFF \modmult_1/xreg_reg[118]  ( .D(\modmult_1/N1147 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[118] ) );
  DFF \modmult_1/xreg_reg[117]  ( .D(\modmult_1/N1146 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[117] ) );
  DFF \modmult_1/xreg_reg[116]  ( .D(\modmult_1/N1145 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[116] ) );
  DFF \modmult_1/xreg_reg[115]  ( .D(\modmult_1/N1144 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[115] ) );
  DFF \modmult_1/xreg_reg[114]  ( .D(\modmult_1/N1143 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[114] ) );
  DFF \modmult_1/xreg_reg[113]  ( .D(\modmult_1/N1142 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[113] ) );
  DFF \modmult_1/xreg_reg[112]  ( .D(\modmult_1/N1141 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[112] ) );
  DFF \modmult_1/xreg_reg[111]  ( .D(\modmult_1/N1140 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[111] ) );
  DFF \modmult_1/xreg_reg[110]  ( .D(\modmult_1/N1139 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[110] ) );
  DFF \modmult_1/xreg_reg[109]  ( .D(\modmult_1/N1138 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[109] ) );
  DFF \modmult_1/xreg_reg[108]  ( .D(\modmult_1/N1137 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[108] ) );
  DFF \modmult_1/xreg_reg[107]  ( .D(\modmult_1/N1136 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[107] ) );
  DFF \modmult_1/xreg_reg[106]  ( .D(\modmult_1/N1135 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[106] ) );
  DFF \modmult_1/xreg_reg[105]  ( .D(\modmult_1/N1134 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[105] ) );
  DFF \modmult_1/xreg_reg[104]  ( .D(\modmult_1/N1133 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[104] ) );
  DFF \modmult_1/xreg_reg[103]  ( .D(\modmult_1/N1132 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[103] ) );
  DFF \modmult_1/xreg_reg[102]  ( .D(\modmult_1/N1131 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[102] ) );
  DFF \modmult_1/xreg_reg[101]  ( .D(\modmult_1/N1130 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[101] ) );
  DFF \modmult_1/xreg_reg[100]  ( .D(\modmult_1/N1129 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[100] ) );
  DFF \modmult_1/xreg_reg[99]  ( .D(\modmult_1/N1128 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[99] ) );
  DFF \modmult_1/xreg_reg[98]  ( .D(\modmult_1/N1127 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[98] ) );
  DFF \modmult_1/xreg_reg[97]  ( .D(\modmult_1/N1126 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[97] ) );
  DFF \modmult_1/xreg_reg[96]  ( .D(\modmult_1/N1125 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[96] ) );
  DFF \modmult_1/xreg_reg[95]  ( .D(\modmult_1/N1124 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[95] ) );
  DFF \modmult_1/xreg_reg[94]  ( .D(\modmult_1/N1123 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[94] ) );
  DFF \modmult_1/xreg_reg[93]  ( .D(\modmult_1/N1122 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[93] ) );
  DFF \modmult_1/xreg_reg[92]  ( .D(\modmult_1/N1121 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[92] ) );
  DFF \modmult_1/xreg_reg[91]  ( .D(\modmult_1/N1120 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[91] ) );
  DFF \modmult_1/xreg_reg[90]  ( .D(\modmult_1/N1119 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[90] ) );
  DFF \modmult_1/xreg_reg[89]  ( .D(\modmult_1/N1118 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[89] ) );
  DFF \modmult_1/xreg_reg[88]  ( .D(\modmult_1/N1117 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[88] ) );
  DFF \modmult_1/xreg_reg[87]  ( .D(\modmult_1/N1116 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[87] ) );
  DFF \modmult_1/xreg_reg[86]  ( .D(\modmult_1/N1115 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[86] ) );
  DFF \modmult_1/xreg_reg[85]  ( .D(\modmult_1/N1114 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[85] ) );
  DFF \modmult_1/xreg_reg[84]  ( .D(\modmult_1/N1113 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[84] ) );
  DFF \modmult_1/xreg_reg[83]  ( .D(\modmult_1/N1112 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[83] ) );
  DFF \modmult_1/xreg_reg[82]  ( .D(\modmult_1/N1111 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[82] ) );
  DFF \modmult_1/xreg_reg[81]  ( .D(\modmult_1/N1110 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[81] ) );
  DFF \modmult_1/xreg_reg[80]  ( .D(\modmult_1/N1109 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[80] ) );
  DFF \modmult_1/xreg_reg[79]  ( .D(\modmult_1/N1108 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[79] ) );
  DFF \modmult_1/xreg_reg[78]  ( .D(\modmult_1/N1107 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[78] ) );
  DFF \modmult_1/xreg_reg[77]  ( .D(\modmult_1/N1106 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[77] ) );
  DFF \modmult_1/xreg_reg[76]  ( .D(\modmult_1/N1105 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[76] ) );
  DFF \modmult_1/xreg_reg[75]  ( .D(\modmult_1/N1104 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[75] ) );
  DFF \modmult_1/xreg_reg[74]  ( .D(\modmult_1/N1103 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[74] ) );
  DFF \modmult_1/xreg_reg[73]  ( .D(\modmult_1/N1102 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[73] ) );
  DFF \modmult_1/xreg_reg[72]  ( .D(\modmult_1/N1101 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[72] ) );
  DFF \modmult_1/xreg_reg[71]  ( .D(\modmult_1/N1100 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[71] ) );
  DFF \modmult_1/xreg_reg[70]  ( .D(\modmult_1/N1099 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[70] ) );
  DFF \modmult_1/xreg_reg[69]  ( .D(\modmult_1/N1098 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[69] ) );
  DFF \modmult_1/xreg_reg[68]  ( .D(\modmult_1/N1097 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[68] ) );
  DFF \modmult_1/xreg_reg[67]  ( .D(\modmult_1/N1096 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[67] ) );
  DFF \modmult_1/xreg_reg[66]  ( .D(\modmult_1/N1095 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[66] ) );
  DFF \modmult_1/xreg_reg[65]  ( .D(\modmult_1/N1094 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[65] ) );
  DFF \modmult_1/xreg_reg[64]  ( .D(\modmult_1/N1093 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[64] ) );
  DFF \modmult_1/xreg_reg[63]  ( .D(\modmult_1/N1092 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[63] ) );
  DFF \modmult_1/xreg_reg[62]  ( .D(\modmult_1/N1091 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[62] ) );
  DFF \modmult_1/xreg_reg[61]  ( .D(\modmult_1/N1090 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[61] ) );
  DFF \modmult_1/xreg_reg[60]  ( .D(\modmult_1/N1089 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[60] ) );
  DFF \modmult_1/xreg_reg[59]  ( .D(\modmult_1/N1088 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[59] ) );
  DFF \modmult_1/xreg_reg[58]  ( .D(\modmult_1/N1087 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[58] ) );
  DFF \modmult_1/xreg_reg[57]  ( .D(\modmult_1/N1086 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[57] ) );
  DFF \modmult_1/xreg_reg[56]  ( .D(\modmult_1/N1085 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[56] ) );
  DFF \modmult_1/xreg_reg[55]  ( .D(\modmult_1/N1084 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[55] ) );
  DFF \modmult_1/xreg_reg[54]  ( .D(\modmult_1/N1083 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[54] ) );
  DFF \modmult_1/xreg_reg[53]  ( .D(\modmult_1/N1082 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[53] ) );
  DFF \modmult_1/xreg_reg[52]  ( .D(\modmult_1/N1081 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[52] ) );
  DFF \modmult_1/xreg_reg[51]  ( .D(\modmult_1/N1080 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[51] ) );
  DFF \modmult_1/xreg_reg[50]  ( .D(\modmult_1/N1079 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[50] ) );
  DFF \modmult_1/xreg_reg[49]  ( .D(\modmult_1/N1078 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[49] ) );
  DFF \modmult_1/xreg_reg[48]  ( .D(\modmult_1/N1077 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[48] ) );
  DFF \modmult_1/xreg_reg[47]  ( .D(\modmult_1/N1076 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[47] ) );
  DFF \modmult_1/xreg_reg[46]  ( .D(\modmult_1/N1075 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[46] ) );
  DFF \modmult_1/xreg_reg[45]  ( .D(\modmult_1/N1074 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[45] ) );
  DFF \modmult_1/xreg_reg[44]  ( .D(\modmult_1/N1073 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[44] ) );
  DFF \modmult_1/xreg_reg[43]  ( .D(\modmult_1/N1072 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[43] ) );
  DFF \modmult_1/xreg_reg[42]  ( .D(\modmult_1/N1071 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[42] ) );
  DFF \modmult_1/xreg_reg[41]  ( .D(\modmult_1/N1070 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[41] ) );
  DFF \modmult_1/xreg_reg[40]  ( .D(\modmult_1/N1069 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[40] ) );
  DFF \modmult_1/xreg_reg[39]  ( .D(\modmult_1/N1068 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[39] ) );
  DFF \modmult_1/xreg_reg[38]  ( .D(\modmult_1/N1067 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[38] ) );
  DFF \modmult_1/xreg_reg[37]  ( .D(\modmult_1/N1066 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[37] ) );
  DFF \modmult_1/xreg_reg[36]  ( .D(\modmult_1/N1065 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[36] ) );
  DFF \modmult_1/xreg_reg[35]  ( .D(\modmult_1/N1064 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[35] ) );
  DFF \modmult_1/xreg_reg[34]  ( .D(\modmult_1/N1063 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[34] ) );
  DFF \modmult_1/xreg_reg[33]  ( .D(\modmult_1/N1062 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[33] ) );
  DFF \modmult_1/xreg_reg[32]  ( .D(\modmult_1/N1061 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[32] ) );
  DFF \modmult_1/xreg_reg[31]  ( .D(\modmult_1/N1060 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[31] ) );
  DFF \modmult_1/xreg_reg[30]  ( .D(\modmult_1/N1059 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[30] ) );
  DFF \modmult_1/xreg_reg[29]  ( .D(\modmult_1/N1058 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[29] ) );
  DFF \modmult_1/xreg_reg[28]  ( .D(\modmult_1/N1057 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[28] ) );
  DFF \modmult_1/xreg_reg[27]  ( .D(\modmult_1/N1056 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[27] ) );
  DFF \modmult_1/xreg_reg[26]  ( .D(\modmult_1/N1055 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[26] ) );
  DFF \modmult_1/xreg_reg[25]  ( .D(\modmult_1/N1054 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[25] ) );
  DFF \modmult_1/xreg_reg[24]  ( .D(\modmult_1/N1053 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[24] ) );
  DFF \modmult_1/xreg_reg[23]  ( .D(\modmult_1/N1052 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[23] ) );
  DFF \modmult_1/xreg_reg[22]  ( .D(\modmult_1/N1051 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[22] ) );
  DFF \modmult_1/xreg_reg[21]  ( .D(\modmult_1/N1050 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[21] ) );
  DFF \modmult_1/xreg_reg[20]  ( .D(\modmult_1/N1049 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[20] ) );
  DFF \modmult_1/xreg_reg[19]  ( .D(\modmult_1/N1048 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[19] ) );
  DFF \modmult_1/xreg_reg[18]  ( .D(\modmult_1/N1047 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[18] ) );
  DFF \modmult_1/xreg_reg[17]  ( .D(\modmult_1/N1046 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[17] ) );
  DFF \modmult_1/xreg_reg[16]  ( .D(\modmult_1/N1045 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[16] ) );
  DFF \modmult_1/xreg_reg[15]  ( .D(\modmult_1/N1044 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[15] ) );
  DFF \modmult_1/xreg_reg[14]  ( .D(\modmult_1/N1043 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[14] ) );
  DFF \modmult_1/xreg_reg[13]  ( .D(\modmult_1/N1042 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[13] ) );
  DFF \modmult_1/xreg_reg[12]  ( .D(\modmult_1/N1041 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[12] ) );
  DFF \modmult_1/xreg_reg[11]  ( .D(\modmult_1/N1040 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[11] ) );
  DFF \modmult_1/xreg_reg[10]  ( .D(\modmult_1/N1039 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[10] ) );
  DFF \modmult_1/xreg_reg[9]  ( .D(\modmult_1/N1038 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[9] ) );
  DFF \modmult_1/xreg_reg[8]  ( .D(\modmult_1/N1037 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[8] ) );
  DFF \modmult_1/xreg_reg[7]  ( .D(\modmult_1/N1036 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[7] ) );
  DFF \modmult_1/xreg_reg[6]  ( .D(\modmult_1/N1035 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[6] ) );
  DFF \modmult_1/xreg_reg[5]  ( .D(\modmult_1/N1034 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[5] ) );
  DFF \modmult_1/xreg_reg[4]  ( .D(\modmult_1/N1033 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[4] ) );
  DFF \modmult_1/xreg_reg[3]  ( .D(\modmult_1/N1032 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[3] ) );
  DFF \modmult_1/xreg_reg[2]  ( .D(\modmult_1/N1031 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[2] ) );
  DFF \modmult_1/xreg_reg[1]  ( .D(\modmult_1/N1030 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[1] ) );
  DFF \modmult_1/xreg_reg[0]  ( .D(\modmult_1/N1029 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\modmult_1/xin[0] ) );
  XNOR U1037 ( .A(n1033), .B(n1034), .Z(o[9]) );
  AND U1038 ( .A(n1035), .B(n1036), .Z(n1033) );
  XNOR U1039 ( .A(creg[9]), .B(n1034), .Z(n1036) );
  XNOR U1040 ( .A(n1037), .B(n1038), .Z(o[99]) );
  AND U1041 ( .A(n1035), .B(n1039), .Z(n1037) );
  XNOR U1042 ( .A(creg[99]), .B(n1038), .Z(n1039) );
  XNOR U1043 ( .A(n1040), .B(n1041), .Z(o[999]) );
  AND U1044 ( .A(n1035), .B(n1042), .Z(n1040) );
  XNOR U1045 ( .A(creg[999]), .B(n1041), .Z(n1042) );
  XNOR U1046 ( .A(n1043), .B(n1044), .Z(o[998]) );
  AND U1047 ( .A(n1035), .B(n1045), .Z(n1043) );
  XNOR U1048 ( .A(creg[998]), .B(n1044), .Z(n1045) );
  XNOR U1049 ( .A(n1046), .B(n1047), .Z(o[997]) );
  AND U1050 ( .A(n1035), .B(n1048), .Z(n1046) );
  XNOR U1051 ( .A(creg[997]), .B(n1047), .Z(n1048) );
  XNOR U1052 ( .A(n1049), .B(n1050), .Z(o[996]) );
  AND U1053 ( .A(n1035), .B(n1051), .Z(n1049) );
  XNOR U1054 ( .A(creg[996]), .B(n1050), .Z(n1051) );
  XNOR U1055 ( .A(n1052), .B(n1053), .Z(o[995]) );
  AND U1056 ( .A(n1035), .B(n1054), .Z(n1052) );
  XNOR U1057 ( .A(creg[995]), .B(n1053), .Z(n1054) );
  XNOR U1058 ( .A(n1055), .B(n1056), .Z(o[994]) );
  AND U1059 ( .A(n1035), .B(n1057), .Z(n1055) );
  XNOR U1060 ( .A(creg[994]), .B(n1056), .Z(n1057) );
  XNOR U1061 ( .A(n1058), .B(n1059), .Z(o[993]) );
  AND U1062 ( .A(n1035), .B(n1060), .Z(n1058) );
  XNOR U1063 ( .A(creg[993]), .B(n1059), .Z(n1060) );
  XNOR U1064 ( .A(n1061), .B(n1062), .Z(o[992]) );
  AND U1065 ( .A(n1035), .B(n1063), .Z(n1061) );
  XNOR U1066 ( .A(creg[992]), .B(n1062), .Z(n1063) );
  XNOR U1067 ( .A(n1064), .B(n1065), .Z(o[991]) );
  AND U1068 ( .A(n1035), .B(n1066), .Z(n1064) );
  XNOR U1069 ( .A(creg[991]), .B(n1065), .Z(n1066) );
  XNOR U1070 ( .A(n1067), .B(n1068), .Z(o[990]) );
  AND U1071 ( .A(n1035), .B(n1069), .Z(n1067) );
  XNOR U1072 ( .A(creg[990]), .B(n1068), .Z(n1069) );
  XNOR U1073 ( .A(n1070), .B(n1071), .Z(o[98]) );
  AND U1074 ( .A(n1035), .B(n1072), .Z(n1070) );
  XNOR U1075 ( .A(creg[98]), .B(n1071), .Z(n1072) );
  XNOR U1076 ( .A(n1073), .B(n1074), .Z(o[989]) );
  AND U1077 ( .A(n1035), .B(n1075), .Z(n1073) );
  XNOR U1078 ( .A(creg[989]), .B(n1074), .Z(n1075) );
  XNOR U1079 ( .A(n1076), .B(n1077), .Z(o[988]) );
  AND U1080 ( .A(n1035), .B(n1078), .Z(n1076) );
  XNOR U1081 ( .A(creg[988]), .B(n1077), .Z(n1078) );
  XNOR U1082 ( .A(n1079), .B(n1080), .Z(o[987]) );
  AND U1083 ( .A(n1035), .B(n1081), .Z(n1079) );
  XNOR U1084 ( .A(creg[987]), .B(n1080), .Z(n1081) );
  XNOR U1085 ( .A(n1082), .B(n1083), .Z(o[986]) );
  AND U1086 ( .A(n1035), .B(n1084), .Z(n1082) );
  XNOR U1087 ( .A(creg[986]), .B(n1083), .Z(n1084) );
  XNOR U1088 ( .A(n1085), .B(n1086), .Z(o[985]) );
  AND U1089 ( .A(n1035), .B(n1087), .Z(n1085) );
  XNOR U1090 ( .A(creg[985]), .B(n1086), .Z(n1087) );
  XNOR U1091 ( .A(n1088), .B(n1089), .Z(o[984]) );
  AND U1092 ( .A(n1035), .B(n1090), .Z(n1088) );
  XNOR U1093 ( .A(creg[984]), .B(n1089), .Z(n1090) );
  XNOR U1094 ( .A(n1091), .B(n1092), .Z(o[983]) );
  AND U1095 ( .A(n1035), .B(n1093), .Z(n1091) );
  XNOR U1096 ( .A(creg[983]), .B(n1092), .Z(n1093) );
  XNOR U1097 ( .A(n1094), .B(n1095), .Z(o[982]) );
  AND U1098 ( .A(n1035), .B(n1096), .Z(n1094) );
  XNOR U1099 ( .A(creg[982]), .B(n1095), .Z(n1096) );
  XNOR U1100 ( .A(n1097), .B(n1098), .Z(o[981]) );
  AND U1101 ( .A(n1035), .B(n1099), .Z(n1097) );
  XNOR U1102 ( .A(creg[981]), .B(n1098), .Z(n1099) );
  XNOR U1103 ( .A(n1100), .B(n1101), .Z(o[980]) );
  AND U1104 ( .A(n1035), .B(n1102), .Z(n1100) );
  XNOR U1105 ( .A(creg[980]), .B(n1101), .Z(n1102) );
  XNOR U1106 ( .A(n1103), .B(n1104), .Z(o[97]) );
  AND U1107 ( .A(n1035), .B(n1105), .Z(n1103) );
  XNOR U1108 ( .A(creg[97]), .B(n1104), .Z(n1105) );
  XNOR U1109 ( .A(n1106), .B(n1107), .Z(o[979]) );
  AND U1110 ( .A(n1035), .B(n1108), .Z(n1106) );
  XNOR U1111 ( .A(creg[979]), .B(n1107), .Z(n1108) );
  XNOR U1112 ( .A(n1109), .B(n1110), .Z(o[978]) );
  AND U1113 ( .A(n1035), .B(n1111), .Z(n1109) );
  XNOR U1114 ( .A(creg[978]), .B(n1110), .Z(n1111) );
  XNOR U1115 ( .A(n1112), .B(n1113), .Z(o[977]) );
  AND U1116 ( .A(n1035), .B(n1114), .Z(n1112) );
  XNOR U1117 ( .A(creg[977]), .B(n1113), .Z(n1114) );
  XNOR U1118 ( .A(n1115), .B(n1116), .Z(o[976]) );
  AND U1119 ( .A(n1035), .B(n1117), .Z(n1115) );
  XNOR U1120 ( .A(creg[976]), .B(n1116), .Z(n1117) );
  XNOR U1121 ( .A(n1118), .B(n1119), .Z(o[975]) );
  AND U1122 ( .A(n1035), .B(n1120), .Z(n1118) );
  XNOR U1123 ( .A(creg[975]), .B(n1119), .Z(n1120) );
  XNOR U1124 ( .A(n1121), .B(n1122), .Z(o[974]) );
  AND U1125 ( .A(n1035), .B(n1123), .Z(n1121) );
  XNOR U1126 ( .A(creg[974]), .B(n1122), .Z(n1123) );
  XNOR U1127 ( .A(n1124), .B(n1125), .Z(o[973]) );
  AND U1128 ( .A(n1035), .B(n1126), .Z(n1124) );
  XNOR U1129 ( .A(creg[973]), .B(n1125), .Z(n1126) );
  XNOR U1130 ( .A(n1127), .B(n1128), .Z(o[972]) );
  AND U1131 ( .A(n1035), .B(n1129), .Z(n1127) );
  XNOR U1132 ( .A(creg[972]), .B(n1128), .Z(n1129) );
  XNOR U1133 ( .A(n1130), .B(n1131), .Z(o[971]) );
  AND U1134 ( .A(n1035), .B(n1132), .Z(n1130) );
  XNOR U1135 ( .A(creg[971]), .B(n1131), .Z(n1132) );
  XNOR U1136 ( .A(n1133), .B(n1134), .Z(o[970]) );
  AND U1137 ( .A(n1035), .B(n1135), .Z(n1133) );
  XNOR U1138 ( .A(creg[970]), .B(n1134), .Z(n1135) );
  XNOR U1139 ( .A(n1136), .B(n1137), .Z(o[96]) );
  AND U1140 ( .A(n1035), .B(n1138), .Z(n1136) );
  XNOR U1141 ( .A(creg[96]), .B(n1137), .Z(n1138) );
  XNOR U1142 ( .A(n1139), .B(n1140), .Z(o[969]) );
  AND U1143 ( .A(n1035), .B(n1141), .Z(n1139) );
  XNOR U1144 ( .A(creg[969]), .B(n1140), .Z(n1141) );
  XNOR U1145 ( .A(n1142), .B(n1143), .Z(o[968]) );
  AND U1146 ( .A(n1035), .B(n1144), .Z(n1142) );
  XNOR U1147 ( .A(creg[968]), .B(n1143), .Z(n1144) );
  XNOR U1148 ( .A(n1145), .B(n1146), .Z(o[967]) );
  AND U1149 ( .A(n1035), .B(n1147), .Z(n1145) );
  XNOR U1150 ( .A(creg[967]), .B(n1146), .Z(n1147) );
  XNOR U1151 ( .A(n1148), .B(n1149), .Z(o[966]) );
  AND U1152 ( .A(n1035), .B(n1150), .Z(n1148) );
  XNOR U1153 ( .A(creg[966]), .B(n1149), .Z(n1150) );
  XNOR U1154 ( .A(n1151), .B(n1152), .Z(o[965]) );
  AND U1155 ( .A(n1035), .B(n1153), .Z(n1151) );
  XNOR U1156 ( .A(creg[965]), .B(n1152), .Z(n1153) );
  XNOR U1157 ( .A(n1154), .B(n1155), .Z(o[964]) );
  AND U1158 ( .A(n1035), .B(n1156), .Z(n1154) );
  XNOR U1159 ( .A(creg[964]), .B(n1155), .Z(n1156) );
  XNOR U1160 ( .A(n1157), .B(n1158), .Z(o[963]) );
  AND U1161 ( .A(n1035), .B(n1159), .Z(n1157) );
  XNOR U1162 ( .A(creg[963]), .B(n1158), .Z(n1159) );
  XNOR U1163 ( .A(n1160), .B(n1161), .Z(o[962]) );
  AND U1164 ( .A(n1035), .B(n1162), .Z(n1160) );
  XNOR U1165 ( .A(creg[962]), .B(n1161), .Z(n1162) );
  XNOR U1166 ( .A(n1163), .B(n1164), .Z(o[961]) );
  AND U1167 ( .A(n1035), .B(n1165), .Z(n1163) );
  XNOR U1168 ( .A(creg[961]), .B(n1164), .Z(n1165) );
  XNOR U1169 ( .A(n1166), .B(n1167), .Z(o[960]) );
  AND U1170 ( .A(n1035), .B(n1168), .Z(n1166) );
  XNOR U1171 ( .A(creg[960]), .B(n1167), .Z(n1168) );
  XNOR U1172 ( .A(n1169), .B(n1170), .Z(o[95]) );
  AND U1173 ( .A(n1035), .B(n1171), .Z(n1169) );
  XNOR U1174 ( .A(creg[95]), .B(n1170), .Z(n1171) );
  XNOR U1175 ( .A(n1172), .B(n1173), .Z(o[959]) );
  AND U1176 ( .A(n1035), .B(n1174), .Z(n1172) );
  XNOR U1177 ( .A(creg[959]), .B(n1173), .Z(n1174) );
  XNOR U1178 ( .A(n1175), .B(n1176), .Z(o[958]) );
  AND U1179 ( .A(n1035), .B(n1177), .Z(n1175) );
  XNOR U1180 ( .A(creg[958]), .B(n1176), .Z(n1177) );
  XNOR U1181 ( .A(n1178), .B(n1179), .Z(o[957]) );
  AND U1182 ( .A(n1035), .B(n1180), .Z(n1178) );
  XNOR U1183 ( .A(creg[957]), .B(n1179), .Z(n1180) );
  XNOR U1184 ( .A(n1181), .B(n1182), .Z(o[956]) );
  AND U1185 ( .A(n1035), .B(n1183), .Z(n1181) );
  XNOR U1186 ( .A(creg[956]), .B(n1182), .Z(n1183) );
  XNOR U1187 ( .A(n1184), .B(n1185), .Z(o[955]) );
  AND U1188 ( .A(n1035), .B(n1186), .Z(n1184) );
  XNOR U1189 ( .A(creg[955]), .B(n1185), .Z(n1186) );
  XNOR U1190 ( .A(n1187), .B(n1188), .Z(o[954]) );
  AND U1191 ( .A(n1035), .B(n1189), .Z(n1187) );
  XNOR U1192 ( .A(creg[954]), .B(n1188), .Z(n1189) );
  XNOR U1193 ( .A(n1190), .B(n1191), .Z(o[953]) );
  AND U1194 ( .A(n1035), .B(n1192), .Z(n1190) );
  XNOR U1195 ( .A(creg[953]), .B(n1191), .Z(n1192) );
  XNOR U1196 ( .A(n1193), .B(n1194), .Z(o[952]) );
  AND U1197 ( .A(n1035), .B(n1195), .Z(n1193) );
  XNOR U1198 ( .A(creg[952]), .B(n1194), .Z(n1195) );
  XNOR U1199 ( .A(n1196), .B(n1197), .Z(o[951]) );
  AND U1200 ( .A(n1035), .B(n1198), .Z(n1196) );
  XNOR U1201 ( .A(creg[951]), .B(n1197), .Z(n1198) );
  XNOR U1202 ( .A(n1199), .B(n1200), .Z(o[950]) );
  AND U1203 ( .A(n1035), .B(n1201), .Z(n1199) );
  XNOR U1204 ( .A(creg[950]), .B(n1200), .Z(n1201) );
  XNOR U1205 ( .A(n1202), .B(n1203), .Z(o[94]) );
  AND U1206 ( .A(n1035), .B(n1204), .Z(n1202) );
  XNOR U1207 ( .A(creg[94]), .B(n1203), .Z(n1204) );
  XNOR U1208 ( .A(n1205), .B(n1206), .Z(o[949]) );
  AND U1209 ( .A(n1035), .B(n1207), .Z(n1205) );
  XNOR U1210 ( .A(creg[949]), .B(n1206), .Z(n1207) );
  XNOR U1211 ( .A(n1208), .B(n1209), .Z(o[948]) );
  AND U1212 ( .A(n1035), .B(n1210), .Z(n1208) );
  XNOR U1213 ( .A(creg[948]), .B(n1209), .Z(n1210) );
  XNOR U1214 ( .A(n1211), .B(n1212), .Z(o[947]) );
  AND U1215 ( .A(n1035), .B(n1213), .Z(n1211) );
  XNOR U1216 ( .A(creg[947]), .B(n1212), .Z(n1213) );
  XNOR U1217 ( .A(n1214), .B(n1215), .Z(o[946]) );
  AND U1218 ( .A(n1035), .B(n1216), .Z(n1214) );
  XNOR U1219 ( .A(creg[946]), .B(n1215), .Z(n1216) );
  XNOR U1220 ( .A(n1217), .B(n1218), .Z(o[945]) );
  AND U1221 ( .A(n1035), .B(n1219), .Z(n1217) );
  XNOR U1222 ( .A(creg[945]), .B(n1218), .Z(n1219) );
  XNOR U1223 ( .A(n1220), .B(n1221), .Z(o[944]) );
  AND U1224 ( .A(n1035), .B(n1222), .Z(n1220) );
  XNOR U1225 ( .A(creg[944]), .B(n1221), .Z(n1222) );
  XNOR U1226 ( .A(n1223), .B(n1224), .Z(o[943]) );
  AND U1227 ( .A(n1035), .B(n1225), .Z(n1223) );
  XNOR U1228 ( .A(creg[943]), .B(n1224), .Z(n1225) );
  XNOR U1229 ( .A(n1226), .B(n1227), .Z(o[942]) );
  AND U1230 ( .A(n1035), .B(n1228), .Z(n1226) );
  XNOR U1231 ( .A(creg[942]), .B(n1227), .Z(n1228) );
  XNOR U1232 ( .A(n1229), .B(n1230), .Z(o[941]) );
  AND U1233 ( .A(n1035), .B(n1231), .Z(n1229) );
  XNOR U1234 ( .A(creg[941]), .B(n1230), .Z(n1231) );
  XNOR U1235 ( .A(n1232), .B(n1233), .Z(o[940]) );
  AND U1236 ( .A(n1035), .B(n1234), .Z(n1232) );
  XNOR U1237 ( .A(creg[940]), .B(n1233), .Z(n1234) );
  XNOR U1238 ( .A(n1235), .B(n1236), .Z(o[93]) );
  AND U1239 ( .A(n1035), .B(n1237), .Z(n1235) );
  XNOR U1240 ( .A(creg[93]), .B(n1236), .Z(n1237) );
  XNOR U1241 ( .A(n1238), .B(n1239), .Z(o[939]) );
  AND U1242 ( .A(n1035), .B(n1240), .Z(n1238) );
  XNOR U1243 ( .A(creg[939]), .B(n1239), .Z(n1240) );
  XNOR U1244 ( .A(n1241), .B(n1242), .Z(o[938]) );
  AND U1245 ( .A(n1035), .B(n1243), .Z(n1241) );
  XNOR U1246 ( .A(creg[938]), .B(n1242), .Z(n1243) );
  XNOR U1247 ( .A(n1244), .B(n1245), .Z(o[937]) );
  AND U1248 ( .A(n1035), .B(n1246), .Z(n1244) );
  XNOR U1249 ( .A(creg[937]), .B(n1245), .Z(n1246) );
  XNOR U1250 ( .A(n1247), .B(n1248), .Z(o[936]) );
  AND U1251 ( .A(n1035), .B(n1249), .Z(n1247) );
  XNOR U1252 ( .A(creg[936]), .B(n1248), .Z(n1249) );
  XNOR U1253 ( .A(n1250), .B(n1251), .Z(o[935]) );
  AND U1254 ( .A(n1035), .B(n1252), .Z(n1250) );
  XNOR U1255 ( .A(creg[935]), .B(n1251), .Z(n1252) );
  XNOR U1256 ( .A(n1253), .B(n1254), .Z(o[934]) );
  AND U1257 ( .A(n1035), .B(n1255), .Z(n1253) );
  XNOR U1258 ( .A(creg[934]), .B(n1254), .Z(n1255) );
  XNOR U1259 ( .A(n1256), .B(n1257), .Z(o[933]) );
  AND U1260 ( .A(n1035), .B(n1258), .Z(n1256) );
  XNOR U1261 ( .A(creg[933]), .B(n1257), .Z(n1258) );
  XNOR U1262 ( .A(n1259), .B(n1260), .Z(o[932]) );
  AND U1263 ( .A(n1035), .B(n1261), .Z(n1259) );
  XNOR U1264 ( .A(creg[932]), .B(n1260), .Z(n1261) );
  XNOR U1265 ( .A(n1262), .B(n1263), .Z(o[931]) );
  AND U1266 ( .A(n1035), .B(n1264), .Z(n1262) );
  XNOR U1267 ( .A(creg[931]), .B(n1263), .Z(n1264) );
  XNOR U1268 ( .A(n1265), .B(n1266), .Z(o[930]) );
  AND U1269 ( .A(n1035), .B(n1267), .Z(n1265) );
  XNOR U1270 ( .A(creg[930]), .B(n1266), .Z(n1267) );
  XNOR U1271 ( .A(n1268), .B(n1269), .Z(o[92]) );
  AND U1272 ( .A(n1035), .B(n1270), .Z(n1268) );
  XNOR U1273 ( .A(creg[92]), .B(n1269), .Z(n1270) );
  XNOR U1274 ( .A(n1271), .B(n1272), .Z(o[929]) );
  AND U1275 ( .A(n1035), .B(n1273), .Z(n1271) );
  XNOR U1276 ( .A(creg[929]), .B(n1272), .Z(n1273) );
  XNOR U1277 ( .A(n1274), .B(n1275), .Z(o[928]) );
  AND U1278 ( .A(n1035), .B(n1276), .Z(n1274) );
  XNOR U1279 ( .A(creg[928]), .B(n1275), .Z(n1276) );
  XNOR U1280 ( .A(n1277), .B(n1278), .Z(o[927]) );
  AND U1281 ( .A(n1035), .B(n1279), .Z(n1277) );
  XNOR U1282 ( .A(creg[927]), .B(n1278), .Z(n1279) );
  XNOR U1283 ( .A(n1280), .B(n1281), .Z(o[926]) );
  AND U1284 ( .A(n1035), .B(n1282), .Z(n1280) );
  XNOR U1285 ( .A(creg[926]), .B(n1281), .Z(n1282) );
  XNOR U1286 ( .A(n1283), .B(n1284), .Z(o[925]) );
  AND U1287 ( .A(n1035), .B(n1285), .Z(n1283) );
  XNOR U1288 ( .A(creg[925]), .B(n1284), .Z(n1285) );
  XNOR U1289 ( .A(n1286), .B(n1287), .Z(o[924]) );
  AND U1290 ( .A(n1035), .B(n1288), .Z(n1286) );
  XNOR U1291 ( .A(creg[924]), .B(n1287), .Z(n1288) );
  XNOR U1292 ( .A(n1289), .B(n1290), .Z(o[923]) );
  AND U1293 ( .A(n1035), .B(n1291), .Z(n1289) );
  XNOR U1294 ( .A(creg[923]), .B(n1290), .Z(n1291) );
  XNOR U1295 ( .A(n1292), .B(n1293), .Z(o[922]) );
  AND U1296 ( .A(n1035), .B(n1294), .Z(n1292) );
  XNOR U1297 ( .A(creg[922]), .B(n1293), .Z(n1294) );
  XNOR U1298 ( .A(n1295), .B(n1296), .Z(o[921]) );
  AND U1299 ( .A(n1035), .B(n1297), .Z(n1295) );
  XNOR U1300 ( .A(creg[921]), .B(n1296), .Z(n1297) );
  XNOR U1301 ( .A(n1298), .B(n1299), .Z(o[920]) );
  AND U1302 ( .A(n1035), .B(n1300), .Z(n1298) );
  XNOR U1303 ( .A(creg[920]), .B(n1299), .Z(n1300) );
  XNOR U1304 ( .A(n1301), .B(n1302), .Z(o[91]) );
  AND U1305 ( .A(n1035), .B(n1303), .Z(n1301) );
  XNOR U1306 ( .A(creg[91]), .B(n1302), .Z(n1303) );
  XNOR U1307 ( .A(n1304), .B(n1305), .Z(o[919]) );
  AND U1308 ( .A(n1035), .B(n1306), .Z(n1304) );
  XNOR U1309 ( .A(creg[919]), .B(n1305), .Z(n1306) );
  XNOR U1310 ( .A(n1307), .B(n1308), .Z(o[918]) );
  AND U1311 ( .A(n1035), .B(n1309), .Z(n1307) );
  XNOR U1312 ( .A(creg[918]), .B(n1308), .Z(n1309) );
  XNOR U1313 ( .A(n1310), .B(n1311), .Z(o[917]) );
  AND U1314 ( .A(n1035), .B(n1312), .Z(n1310) );
  XNOR U1315 ( .A(creg[917]), .B(n1311), .Z(n1312) );
  XNOR U1316 ( .A(n1313), .B(n1314), .Z(o[916]) );
  AND U1317 ( .A(n1035), .B(n1315), .Z(n1313) );
  XNOR U1318 ( .A(creg[916]), .B(n1314), .Z(n1315) );
  XNOR U1319 ( .A(n1316), .B(n1317), .Z(o[915]) );
  AND U1320 ( .A(n1035), .B(n1318), .Z(n1316) );
  XNOR U1321 ( .A(creg[915]), .B(n1317), .Z(n1318) );
  XNOR U1322 ( .A(n1319), .B(n1320), .Z(o[914]) );
  AND U1323 ( .A(n1035), .B(n1321), .Z(n1319) );
  XNOR U1324 ( .A(creg[914]), .B(n1320), .Z(n1321) );
  XNOR U1325 ( .A(n1322), .B(n1323), .Z(o[913]) );
  AND U1326 ( .A(n1035), .B(n1324), .Z(n1322) );
  XNOR U1327 ( .A(creg[913]), .B(n1323), .Z(n1324) );
  XNOR U1328 ( .A(n1325), .B(n1326), .Z(o[912]) );
  AND U1329 ( .A(n1035), .B(n1327), .Z(n1325) );
  XNOR U1330 ( .A(creg[912]), .B(n1326), .Z(n1327) );
  XNOR U1331 ( .A(n1328), .B(n1329), .Z(o[911]) );
  AND U1332 ( .A(n1035), .B(n1330), .Z(n1328) );
  XNOR U1333 ( .A(creg[911]), .B(n1329), .Z(n1330) );
  XNOR U1334 ( .A(n1331), .B(n1332), .Z(o[910]) );
  AND U1335 ( .A(n1035), .B(n1333), .Z(n1331) );
  XNOR U1336 ( .A(creg[910]), .B(n1332), .Z(n1333) );
  XNOR U1337 ( .A(n1334), .B(n1335), .Z(o[90]) );
  AND U1338 ( .A(n1035), .B(n1336), .Z(n1334) );
  XNOR U1339 ( .A(creg[90]), .B(n1335), .Z(n1336) );
  XNOR U1340 ( .A(n1337), .B(n1338), .Z(o[909]) );
  AND U1341 ( .A(n1035), .B(n1339), .Z(n1337) );
  XNOR U1342 ( .A(creg[909]), .B(n1338), .Z(n1339) );
  XNOR U1343 ( .A(n1340), .B(n1341), .Z(o[908]) );
  AND U1344 ( .A(n1035), .B(n1342), .Z(n1340) );
  XNOR U1345 ( .A(creg[908]), .B(n1341), .Z(n1342) );
  XNOR U1346 ( .A(n1343), .B(n1344), .Z(o[907]) );
  AND U1347 ( .A(n1035), .B(n1345), .Z(n1343) );
  XNOR U1348 ( .A(creg[907]), .B(n1344), .Z(n1345) );
  XNOR U1349 ( .A(n1346), .B(n1347), .Z(o[906]) );
  AND U1350 ( .A(n1035), .B(n1348), .Z(n1346) );
  XNOR U1351 ( .A(creg[906]), .B(n1347), .Z(n1348) );
  XNOR U1352 ( .A(n1349), .B(n1350), .Z(o[905]) );
  AND U1353 ( .A(n1035), .B(n1351), .Z(n1349) );
  XNOR U1354 ( .A(creg[905]), .B(n1350), .Z(n1351) );
  XNOR U1355 ( .A(n1352), .B(n1353), .Z(o[904]) );
  AND U1356 ( .A(n1035), .B(n1354), .Z(n1352) );
  XNOR U1357 ( .A(creg[904]), .B(n1353), .Z(n1354) );
  XNOR U1358 ( .A(n1355), .B(n1356), .Z(o[903]) );
  AND U1359 ( .A(n1035), .B(n1357), .Z(n1355) );
  XNOR U1360 ( .A(creg[903]), .B(n1356), .Z(n1357) );
  XNOR U1361 ( .A(n1358), .B(n1359), .Z(o[902]) );
  AND U1362 ( .A(n1035), .B(n1360), .Z(n1358) );
  XNOR U1363 ( .A(creg[902]), .B(n1359), .Z(n1360) );
  XNOR U1364 ( .A(n1361), .B(n1362), .Z(o[901]) );
  AND U1365 ( .A(n1035), .B(n1363), .Z(n1361) );
  XNOR U1366 ( .A(creg[901]), .B(n1362), .Z(n1363) );
  XNOR U1367 ( .A(n1364), .B(n1365), .Z(o[900]) );
  AND U1368 ( .A(n1035), .B(n1366), .Z(n1364) );
  XNOR U1369 ( .A(creg[900]), .B(n1365), .Z(n1366) );
  XNOR U1370 ( .A(n1367), .B(n1368), .Z(o[8]) );
  AND U1371 ( .A(n1035), .B(n1369), .Z(n1367) );
  XNOR U1372 ( .A(creg[8]), .B(n1368), .Z(n1369) );
  XNOR U1373 ( .A(n1370), .B(n1371), .Z(o[89]) );
  AND U1374 ( .A(n1035), .B(n1372), .Z(n1370) );
  XNOR U1375 ( .A(creg[89]), .B(n1371), .Z(n1372) );
  XNOR U1376 ( .A(n1373), .B(n1374), .Z(o[899]) );
  AND U1377 ( .A(n1035), .B(n1375), .Z(n1373) );
  XNOR U1378 ( .A(creg[899]), .B(n1374), .Z(n1375) );
  XNOR U1379 ( .A(n1376), .B(n1377), .Z(o[898]) );
  AND U1380 ( .A(n1035), .B(n1378), .Z(n1376) );
  XNOR U1381 ( .A(creg[898]), .B(n1377), .Z(n1378) );
  XNOR U1382 ( .A(n1379), .B(n1380), .Z(o[897]) );
  AND U1383 ( .A(n1035), .B(n1381), .Z(n1379) );
  XNOR U1384 ( .A(creg[897]), .B(n1380), .Z(n1381) );
  XNOR U1385 ( .A(n1382), .B(n1383), .Z(o[896]) );
  AND U1386 ( .A(n1035), .B(n1384), .Z(n1382) );
  XNOR U1387 ( .A(creg[896]), .B(n1383), .Z(n1384) );
  XNOR U1388 ( .A(n1385), .B(n1386), .Z(o[895]) );
  AND U1389 ( .A(n1035), .B(n1387), .Z(n1385) );
  XNOR U1390 ( .A(creg[895]), .B(n1386), .Z(n1387) );
  XNOR U1391 ( .A(n1388), .B(n1389), .Z(o[894]) );
  AND U1392 ( .A(n1035), .B(n1390), .Z(n1388) );
  XNOR U1393 ( .A(creg[894]), .B(n1389), .Z(n1390) );
  XNOR U1394 ( .A(n1391), .B(n1392), .Z(o[893]) );
  AND U1395 ( .A(n1035), .B(n1393), .Z(n1391) );
  XNOR U1396 ( .A(creg[893]), .B(n1392), .Z(n1393) );
  XNOR U1397 ( .A(n1394), .B(n1395), .Z(o[892]) );
  AND U1398 ( .A(n1035), .B(n1396), .Z(n1394) );
  XNOR U1399 ( .A(creg[892]), .B(n1395), .Z(n1396) );
  XNOR U1400 ( .A(n1397), .B(n1398), .Z(o[891]) );
  AND U1401 ( .A(n1035), .B(n1399), .Z(n1397) );
  XNOR U1402 ( .A(creg[891]), .B(n1398), .Z(n1399) );
  XNOR U1403 ( .A(n1400), .B(n1401), .Z(o[890]) );
  AND U1404 ( .A(n1035), .B(n1402), .Z(n1400) );
  XNOR U1405 ( .A(creg[890]), .B(n1401), .Z(n1402) );
  XNOR U1406 ( .A(n1403), .B(n1404), .Z(o[88]) );
  AND U1407 ( .A(n1035), .B(n1405), .Z(n1403) );
  XNOR U1408 ( .A(creg[88]), .B(n1404), .Z(n1405) );
  XNOR U1409 ( .A(n1406), .B(n1407), .Z(o[889]) );
  AND U1410 ( .A(n1035), .B(n1408), .Z(n1406) );
  XNOR U1411 ( .A(creg[889]), .B(n1407), .Z(n1408) );
  XNOR U1412 ( .A(n1409), .B(n1410), .Z(o[888]) );
  AND U1413 ( .A(n1035), .B(n1411), .Z(n1409) );
  XNOR U1414 ( .A(creg[888]), .B(n1410), .Z(n1411) );
  XNOR U1415 ( .A(n1412), .B(n1413), .Z(o[887]) );
  AND U1416 ( .A(n1035), .B(n1414), .Z(n1412) );
  XNOR U1417 ( .A(creg[887]), .B(n1413), .Z(n1414) );
  XNOR U1418 ( .A(n1415), .B(n1416), .Z(o[886]) );
  AND U1419 ( .A(n1035), .B(n1417), .Z(n1415) );
  XNOR U1420 ( .A(creg[886]), .B(n1416), .Z(n1417) );
  XNOR U1421 ( .A(n1418), .B(n1419), .Z(o[885]) );
  AND U1422 ( .A(n1035), .B(n1420), .Z(n1418) );
  XNOR U1423 ( .A(creg[885]), .B(n1419), .Z(n1420) );
  XNOR U1424 ( .A(n1421), .B(n1422), .Z(o[884]) );
  AND U1425 ( .A(n1035), .B(n1423), .Z(n1421) );
  XNOR U1426 ( .A(creg[884]), .B(n1422), .Z(n1423) );
  XNOR U1427 ( .A(n1424), .B(n1425), .Z(o[883]) );
  AND U1428 ( .A(n1035), .B(n1426), .Z(n1424) );
  XNOR U1429 ( .A(creg[883]), .B(n1425), .Z(n1426) );
  XNOR U1430 ( .A(n1427), .B(n1428), .Z(o[882]) );
  AND U1431 ( .A(n1035), .B(n1429), .Z(n1427) );
  XNOR U1432 ( .A(creg[882]), .B(n1428), .Z(n1429) );
  XNOR U1433 ( .A(n1430), .B(n1431), .Z(o[881]) );
  AND U1434 ( .A(n1035), .B(n1432), .Z(n1430) );
  XNOR U1435 ( .A(creg[881]), .B(n1431), .Z(n1432) );
  XNOR U1436 ( .A(n1433), .B(n1434), .Z(o[880]) );
  AND U1437 ( .A(n1035), .B(n1435), .Z(n1433) );
  XNOR U1438 ( .A(creg[880]), .B(n1434), .Z(n1435) );
  XNOR U1439 ( .A(n1436), .B(n1437), .Z(o[87]) );
  AND U1440 ( .A(n1035), .B(n1438), .Z(n1436) );
  XNOR U1441 ( .A(creg[87]), .B(n1437), .Z(n1438) );
  XNOR U1442 ( .A(n1439), .B(n1440), .Z(o[879]) );
  AND U1443 ( .A(n1035), .B(n1441), .Z(n1439) );
  XNOR U1444 ( .A(creg[879]), .B(n1440), .Z(n1441) );
  XNOR U1445 ( .A(n1442), .B(n1443), .Z(o[878]) );
  AND U1446 ( .A(n1035), .B(n1444), .Z(n1442) );
  XNOR U1447 ( .A(creg[878]), .B(n1443), .Z(n1444) );
  XNOR U1448 ( .A(n1445), .B(n1446), .Z(o[877]) );
  AND U1449 ( .A(n1035), .B(n1447), .Z(n1445) );
  XNOR U1450 ( .A(creg[877]), .B(n1446), .Z(n1447) );
  XNOR U1451 ( .A(n1448), .B(n1449), .Z(o[876]) );
  AND U1452 ( .A(n1035), .B(n1450), .Z(n1448) );
  XNOR U1453 ( .A(creg[876]), .B(n1449), .Z(n1450) );
  XNOR U1454 ( .A(n1451), .B(n1452), .Z(o[875]) );
  AND U1455 ( .A(n1035), .B(n1453), .Z(n1451) );
  XNOR U1456 ( .A(creg[875]), .B(n1452), .Z(n1453) );
  XNOR U1457 ( .A(n1454), .B(n1455), .Z(o[874]) );
  AND U1458 ( .A(n1035), .B(n1456), .Z(n1454) );
  XNOR U1459 ( .A(creg[874]), .B(n1455), .Z(n1456) );
  XNOR U1460 ( .A(n1457), .B(n1458), .Z(o[873]) );
  AND U1461 ( .A(n1035), .B(n1459), .Z(n1457) );
  XNOR U1462 ( .A(creg[873]), .B(n1458), .Z(n1459) );
  XNOR U1463 ( .A(n1460), .B(n1461), .Z(o[872]) );
  AND U1464 ( .A(n1035), .B(n1462), .Z(n1460) );
  XNOR U1465 ( .A(creg[872]), .B(n1461), .Z(n1462) );
  XNOR U1466 ( .A(n1463), .B(n1464), .Z(o[871]) );
  AND U1467 ( .A(n1035), .B(n1465), .Z(n1463) );
  XNOR U1468 ( .A(creg[871]), .B(n1464), .Z(n1465) );
  XNOR U1469 ( .A(n1466), .B(n1467), .Z(o[870]) );
  AND U1470 ( .A(n1035), .B(n1468), .Z(n1466) );
  XNOR U1471 ( .A(creg[870]), .B(n1467), .Z(n1468) );
  XNOR U1472 ( .A(n1469), .B(n1470), .Z(o[86]) );
  AND U1473 ( .A(n1035), .B(n1471), .Z(n1469) );
  XNOR U1474 ( .A(creg[86]), .B(n1470), .Z(n1471) );
  XNOR U1475 ( .A(n1472), .B(n1473), .Z(o[869]) );
  AND U1476 ( .A(n1035), .B(n1474), .Z(n1472) );
  XNOR U1477 ( .A(creg[869]), .B(n1473), .Z(n1474) );
  XNOR U1478 ( .A(n1475), .B(n1476), .Z(o[868]) );
  AND U1479 ( .A(n1035), .B(n1477), .Z(n1475) );
  XNOR U1480 ( .A(creg[868]), .B(n1476), .Z(n1477) );
  XNOR U1481 ( .A(n1478), .B(n1479), .Z(o[867]) );
  AND U1482 ( .A(n1035), .B(n1480), .Z(n1478) );
  XNOR U1483 ( .A(creg[867]), .B(n1479), .Z(n1480) );
  XNOR U1484 ( .A(n1481), .B(n1482), .Z(o[866]) );
  AND U1485 ( .A(n1035), .B(n1483), .Z(n1481) );
  XNOR U1486 ( .A(creg[866]), .B(n1482), .Z(n1483) );
  XNOR U1487 ( .A(n1484), .B(n1485), .Z(o[865]) );
  AND U1488 ( .A(n1035), .B(n1486), .Z(n1484) );
  XNOR U1489 ( .A(creg[865]), .B(n1485), .Z(n1486) );
  XNOR U1490 ( .A(n1487), .B(n1488), .Z(o[864]) );
  AND U1491 ( .A(n1035), .B(n1489), .Z(n1487) );
  XNOR U1492 ( .A(creg[864]), .B(n1488), .Z(n1489) );
  XNOR U1493 ( .A(n1490), .B(n1491), .Z(o[863]) );
  AND U1494 ( .A(n1035), .B(n1492), .Z(n1490) );
  XNOR U1495 ( .A(creg[863]), .B(n1491), .Z(n1492) );
  XNOR U1496 ( .A(n1493), .B(n1494), .Z(o[862]) );
  AND U1497 ( .A(n1035), .B(n1495), .Z(n1493) );
  XNOR U1498 ( .A(creg[862]), .B(n1494), .Z(n1495) );
  XNOR U1499 ( .A(n1496), .B(n1497), .Z(o[861]) );
  AND U1500 ( .A(n1035), .B(n1498), .Z(n1496) );
  XNOR U1501 ( .A(creg[861]), .B(n1497), .Z(n1498) );
  XNOR U1502 ( .A(n1499), .B(n1500), .Z(o[860]) );
  AND U1503 ( .A(n1035), .B(n1501), .Z(n1499) );
  XNOR U1504 ( .A(creg[860]), .B(n1500), .Z(n1501) );
  XNOR U1505 ( .A(n1502), .B(n1503), .Z(o[85]) );
  AND U1506 ( .A(n1035), .B(n1504), .Z(n1502) );
  XNOR U1507 ( .A(creg[85]), .B(n1503), .Z(n1504) );
  XNOR U1508 ( .A(n1505), .B(n1506), .Z(o[859]) );
  AND U1509 ( .A(n1035), .B(n1507), .Z(n1505) );
  XNOR U1510 ( .A(creg[859]), .B(n1506), .Z(n1507) );
  XNOR U1511 ( .A(n1508), .B(n1509), .Z(o[858]) );
  AND U1512 ( .A(n1035), .B(n1510), .Z(n1508) );
  XNOR U1513 ( .A(creg[858]), .B(n1509), .Z(n1510) );
  XNOR U1514 ( .A(n1511), .B(n1512), .Z(o[857]) );
  AND U1515 ( .A(n1035), .B(n1513), .Z(n1511) );
  XNOR U1516 ( .A(creg[857]), .B(n1512), .Z(n1513) );
  XNOR U1517 ( .A(n1514), .B(n1515), .Z(o[856]) );
  AND U1518 ( .A(n1035), .B(n1516), .Z(n1514) );
  XNOR U1519 ( .A(creg[856]), .B(n1515), .Z(n1516) );
  XNOR U1520 ( .A(n1517), .B(n1518), .Z(o[855]) );
  AND U1521 ( .A(n1035), .B(n1519), .Z(n1517) );
  XNOR U1522 ( .A(creg[855]), .B(n1518), .Z(n1519) );
  XNOR U1523 ( .A(n1520), .B(n1521), .Z(o[854]) );
  AND U1524 ( .A(n1035), .B(n1522), .Z(n1520) );
  XNOR U1525 ( .A(creg[854]), .B(n1521), .Z(n1522) );
  XNOR U1526 ( .A(n1523), .B(n1524), .Z(o[853]) );
  AND U1527 ( .A(n1035), .B(n1525), .Z(n1523) );
  XNOR U1528 ( .A(creg[853]), .B(n1524), .Z(n1525) );
  XNOR U1529 ( .A(n1526), .B(n1527), .Z(o[852]) );
  AND U1530 ( .A(n1035), .B(n1528), .Z(n1526) );
  XNOR U1531 ( .A(creg[852]), .B(n1527), .Z(n1528) );
  XNOR U1532 ( .A(n1529), .B(n1530), .Z(o[851]) );
  AND U1533 ( .A(n1035), .B(n1531), .Z(n1529) );
  XNOR U1534 ( .A(creg[851]), .B(n1530), .Z(n1531) );
  XNOR U1535 ( .A(n1532), .B(n1533), .Z(o[850]) );
  AND U1536 ( .A(n1035), .B(n1534), .Z(n1532) );
  XNOR U1537 ( .A(creg[850]), .B(n1533), .Z(n1534) );
  XNOR U1538 ( .A(n1535), .B(n1536), .Z(o[84]) );
  AND U1539 ( .A(n1035), .B(n1537), .Z(n1535) );
  XNOR U1540 ( .A(creg[84]), .B(n1536), .Z(n1537) );
  XNOR U1541 ( .A(n1538), .B(n1539), .Z(o[849]) );
  AND U1542 ( .A(n1035), .B(n1540), .Z(n1538) );
  XNOR U1543 ( .A(creg[849]), .B(n1539), .Z(n1540) );
  XNOR U1544 ( .A(n1541), .B(n1542), .Z(o[848]) );
  AND U1545 ( .A(n1035), .B(n1543), .Z(n1541) );
  XNOR U1546 ( .A(creg[848]), .B(n1542), .Z(n1543) );
  XNOR U1547 ( .A(n1544), .B(n1545), .Z(o[847]) );
  AND U1548 ( .A(n1035), .B(n1546), .Z(n1544) );
  XNOR U1549 ( .A(creg[847]), .B(n1545), .Z(n1546) );
  XNOR U1550 ( .A(n1547), .B(n1548), .Z(o[846]) );
  AND U1551 ( .A(n1035), .B(n1549), .Z(n1547) );
  XNOR U1552 ( .A(creg[846]), .B(n1548), .Z(n1549) );
  XNOR U1553 ( .A(n1550), .B(n1551), .Z(o[845]) );
  AND U1554 ( .A(n1035), .B(n1552), .Z(n1550) );
  XNOR U1555 ( .A(creg[845]), .B(n1551), .Z(n1552) );
  XNOR U1556 ( .A(n1553), .B(n1554), .Z(o[844]) );
  AND U1557 ( .A(n1035), .B(n1555), .Z(n1553) );
  XNOR U1558 ( .A(creg[844]), .B(n1554), .Z(n1555) );
  XNOR U1559 ( .A(n1556), .B(n1557), .Z(o[843]) );
  AND U1560 ( .A(n1035), .B(n1558), .Z(n1556) );
  XNOR U1561 ( .A(creg[843]), .B(n1557), .Z(n1558) );
  XNOR U1562 ( .A(n1559), .B(n1560), .Z(o[842]) );
  AND U1563 ( .A(n1035), .B(n1561), .Z(n1559) );
  XNOR U1564 ( .A(creg[842]), .B(n1560), .Z(n1561) );
  XNOR U1565 ( .A(n1562), .B(n1563), .Z(o[841]) );
  AND U1566 ( .A(n1035), .B(n1564), .Z(n1562) );
  XNOR U1567 ( .A(creg[841]), .B(n1563), .Z(n1564) );
  XNOR U1568 ( .A(n1565), .B(n1566), .Z(o[840]) );
  AND U1569 ( .A(n1035), .B(n1567), .Z(n1565) );
  XNOR U1570 ( .A(creg[840]), .B(n1566), .Z(n1567) );
  XNOR U1571 ( .A(n1568), .B(n1569), .Z(o[83]) );
  AND U1572 ( .A(n1035), .B(n1570), .Z(n1568) );
  XNOR U1573 ( .A(creg[83]), .B(n1569), .Z(n1570) );
  XNOR U1574 ( .A(n1571), .B(n1572), .Z(o[839]) );
  AND U1575 ( .A(n1035), .B(n1573), .Z(n1571) );
  XNOR U1576 ( .A(creg[839]), .B(n1572), .Z(n1573) );
  XNOR U1577 ( .A(n1574), .B(n1575), .Z(o[838]) );
  AND U1578 ( .A(n1035), .B(n1576), .Z(n1574) );
  XNOR U1579 ( .A(creg[838]), .B(n1575), .Z(n1576) );
  XNOR U1580 ( .A(n1577), .B(n1578), .Z(o[837]) );
  AND U1581 ( .A(n1035), .B(n1579), .Z(n1577) );
  XNOR U1582 ( .A(creg[837]), .B(n1578), .Z(n1579) );
  XNOR U1583 ( .A(n1580), .B(n1581), .Z(o[836]) );
  AND U1584 ( .A(n1035), .B(n1582), .Z(n1580) );
  XNOR U1585 ( .A(creg[836]), .B(n1581), .Z(n1582) );
  XNOR U1586 ( .A(n1583), .B(n1584), .Z(o[835]) );
  AND U1587 ( .A(n1035), .B(n1585), .Z(n1583) );
  XNOR U1588 ( .A(creg[835]), .B(n1584), .Z(n1585) );
  XNOR U1589 ( .A(n1586), .B(n1587), .Z(o[834]) );
  AND U1590 ( .A(n1035), .B(n1588), .Z(n1586) );
  XNOR U1591 ( .A(creg[834]), .B(n1587), .Z(n1588) );
  XNOR U1592 ( .A(n1589), .B(n1590), .Z(o[833]) );
  AND U1593 ( .A(n1035), .B(n1591), .Z(n1589) );
  XNOR U1594 ( .A(creg[833]), .B(n1590), .Z(n1591) );
  XNOR U1595 ( .A(n1592), .B(n1593), .Z(o[832]) );
  AND U1596 ( .A(n1035), .B(n1594), .Z(n1592) );
  XNOR U1597 ( .A(creg[832]), .B(n1593), .Z(n1594) );
  XNOR U1598 ( .A(n1595), .B(n1596), .Z(o[831]) );
  AND U1599 ( .A(n1035), .B(n1597), .Z(n1595) );
  XNOR U1600 ( .A(creg[831]), .B(n1596), .Z(n1597) );
  XNOR U1601 ( .A(n1598), .B(n1599), .Z(o[830]) );
  AND U1602 ( .A(n1035), .B(n1600), .Z(n1598) );
  XNOR U1603 ( .A(creg[830]), .B(n1599), .Z(n1600) );
  XNOR U1604 ( .A(n1601), .B(n1602), .Z(o[82]) );
  AND U1605 ( .A(n1035), .B(n1603), .Z(n1601) );
  XNOR U1606 ( .A(creg[82]), .B(n1602), .Z(n1603) );
  XNOR U1607 ( .A(n1604), .B(n1605), .Z(o[829]) );
  AND U1608 ( .A(n1035), .B(n1606), .Z(n1604) );
  XNOR U1609 ( .A(creg[829]), .B(n1605), .Z(n1606) );
  XNOR U1610 ( .A(n1607), .B(n1608), .Z(o[828]) );
  AND U1611 ( .A(n1035), .B(n1609), .Z(n1607) );
  XNOR U1612 ( .A(creg[828]), .B(n1608), .Z(n1609) );
  XNOR U1613 ( .A(n1610), .B(n1611), .Z(o[827]) );
  AND U1614 ( .A(n1035), .B(n1612), .Z(n1610) );
  XNOR U1615 ( .A(creg[827]), .B(n1611), .Z(n1612) );
  XNOR U1616 ( .A(n1613), .B(n1614), .Z(o[826]) );
  AND U1617 ( .A(n1035), .B(n1615), .Z(n1613) );
  XNOR U1618 ( .A(creg[826]), .B(n1614), .Z(n1615) );
  XNOR U1619 ( .A(n1616), .B(n1617), .Z(o[825]) );
  AND U1620 ( .A(n1035), .B(n1618), .Z(n1616) );
  XNOR U1621 ( .A(creg[825]), .B(n1617), .Z(n1618) );
  XNOR U1622 ( .A(n1619), .B(n1620), .Z(o[824]) );
  AND U1623 ( .A(n1035), .B(n1621), .Z(n1619) );
  XNOR U1624 ( .A(creg[824]), .B(n1620), .Z(n1621) );
  XNOR U1625 ( .A(n1622), .B(n1623), .Z(o[823]) );
  AND U1626 ( .A(n1035), .B(n1624), .Z(n1622) );
  XNOR U1627 ( .A(creg[823]), .B(n1623), .Z(n1624) );
  XNOR U1628 ( .A(n1625), .B(n1626), .Z(o[822]) );
  AND U1629 ( .A(n1035), .B(n1627), .Z(n1625) );
  XNOR U1630 ( .A(creg[822]), .B(n1626), .Z(n1627) );
  XNOR U1631 ( .A(n1628), .B(n1629), .Z(o[821]) );
  AND U1632 ( .A(n1035), .B(n1630), .Z(n1628) );
  XNOR U1633 ( .A(creg[821]), .B(n1629), .Z(n1630) );
  XNOR U1634 ( .A(n1631), .B(n1632), .Z(o[820]) );
  AND U1635 ( .A(n1035), .B(n1633), .Z(n1631) );
  XNOR U1636 ( .A(creg[820]), .B(n1632), .Z(n1633) );
  XNOR U1637 ( .A(n1634), .B(n1635), .Z(o[81]) );
  AND U1638 ( .A(n1035), .B(n1636), .Z(n1634) );
  XNOR U1639 ( .A(creg[81]), .B(n1635), .Z(n1636) );
  XNOR U1640 ( .A(n1637), .B(n1638), .Z(o[819]) );
  AND U1641 ( .A(n1035), .B(n1639), .Z(n1637) );
  XNOR U1642 ( .A(creg[819]), .B(n1638), .Z(n1639) );
  XNOR U1643 ( .A(n1640), .B(n1641), .Z(o[818]) );
  AND U1644 ( .A(n1035), .B(n1642), .Z(n1640) );
  XNOR U1645 ( .A(creg[818]), .B(n1641), .Z(n1642) );
  XNOR U1646 ( .A(n1643), .B(n1644), .Z(o[817]) );
  AND U1647 ( .A(n1035), .B(n1645), .Z(n1643) );
  XNOR U1648 ( .A(creg[817]), .B(n1644), .Z(n1645) );
  XNOR U1649 ( .A(n1646), .B(n1647), .Z(o[816]) );
  AND U1650 ( .A(n1035), .B(n1648), .Z(n1646) );
  XNOR U1651 ( .A(creg[816]), .B(n1647), .Z(n1648) );
  XNOR U1652 ( .A(n1649), .B(n1650), .Z(o[815]) );
  AND U1653 ( .A(n1035), .B(n1651), .Z(n1649) );
  XNOR U1654 ( .A(creg[815]), .B(n1650), .Z(n1651) );
  XNOR U1655 ( .A(n1652), .B(n1653), .Z(o[814]) );
  AND U1656 ( .A(n1035), .B(n1654), .Z(n1652) );
  XNOR U1657 ( .A(creg[814]), .B(n1653), .Z(n1654) );
  XNOR U1658 ( .A(n1655), .B(n1656), .Z(o[813]) );
  AND U1659 ( .A(n1035), .B(n1657), .Z(n1655) );
  XNOR U1660 ( .A(creg[813]), .B(n1656), .Z(n1657) );
  XNOR U1661 ( .A(n1658), .B(n1659), .Z(o[812]) );
  AND U1662 ( .A(n1035), .B(n1660), .Z(n1658) );
  XNOR U1663 ( .A(creg[812]), .B(n1659), .Z(n1660) );
  XNOR U1664 ( .A(n1661), .B(n1662), .Z(o[811]) );
  AND U1665 ( .A(n1035), .B(n1663), .Z(n1661) );
  XNOR U1666 ( .A(creg[811]), .B(n1662), .Z(n1663) );
  XNOR U1667 ( .A(n1664), .B(n1665), .Z(o[810]) );
  AND U1668 ( .A(n1035), .B(n1666), .Z(n1664) );
  XNOR U1669 ( .A(creg[810]), .B(n1665), .Z(n1666) );
  XNOR U1670 ( .A(n1667), .B(n1668), .Z(o[80]) );
  AND U1671 ( .A(n1035), .B(n1669), .Z(n1667) );
  XNOR U1672 ( .A(creg[80]), .B(n1668), .Z(n1669) );
  XNOR U1673 ( .A(n1670), .B(n1671), .Z(o[809]) );
  AND U1674 ( .A(n1035), .B(n1672), .Z(n1670) );
  XNOR U1675 ( .A(creg[809]), .B(n1671), .Z(n1672) );
  XNOR U1676 ( .A(n1673), .B(n1674), .Z(o[808]) );
  AND U1677 ( .A(n1035), .B(n1675), .Z(n1673) );
  XNOR U1678 ( .A(creg[808]), .B(n1674), .Z(n1675) );
  XNOR U1679 ( .A(n1676), .B(n1677), .Z(o[807]) );
  AND U1680 ( .A(n1035), .B(n1678), .Z(n1676) );
  XNOR U1681 ( .A(creg[807]), .B(n1677), .Z(n1678) );
  XNOR U1682 ( .A(n1679), .B(n1680), .Z(o[806]) );
  AND U1683 ( .A(n1035), .B(n1681), .Z(n1679) );
  XNOR U1684 ( .A(creg[806]), .B(n1680), .Z(n1681) );
  XNOR U1685 ( .A(n1682), .B(n1683), .Z(o[805]) );
  AND U1686 ( .A(n1035), .B(n1684), .Z(n1682) );
  XNOR U1687 ( .A(creg[805]), .B(n1683), .Z(n1684) );
  XNOR U1688 ( .A(n1685), .B(n1686), .Z(o[804]) );
  AND U1689 ( .A(n1035), .B(n1687), .Z(n1685) );
  XNOR U1690 ( .A(creg[804]), .B(n1686), .Z(n1687) );
  XNOR U1691 ( .A(n1688), .B(n1689), .Z(o[803]) );
  AND U1692 ( .A(n1035), .B(n1690), .Z(n1688) );
  XNOR U1693 ( .A(creg[803]), .B(n1689), .Z(n1690) );
  XNOR U1694 ( .A(n1691), .B(n1692), .Z(o[802]) );
  AND U1695 ( .A(n1035), .B(n1693), .Z(n1691) );
  XNOR U1696 ( .A(creg[802]), .B(n1692), .Z(n1693) );
  XNOR U1697 ( .A(n1694), .B(n1695), .Z(o[801]) );
  AND U1698 ( .A(n1035), .B(n1696), .Z(n1694) );
  XNOR U1699 ( .A(creg[801]), .B(n1695), .Z(n1696) );
  XNOR U1700 ( .A(n1697), .B(n1698), .Z(o[800]) );
  AND U1701 ( .A(n1035), .B(n1699), .Z(n1697) );
  XNOR U1702 ( .A(creg[800]), .B(n1698), .Z(n1699) );
  XNOR U1703 ( .A(n1700), .B(n1701), .Z(o[7]) );
  AND U1704 ( .A(n1035), .B(n1702), .Z(n1700) );
  XNOR U1705 ( .A(creg[7]), .B(n1701), .Z(n1702) );
  XNOR U1706 ( .A(n1703), .B(n1704), .Z(o[79]) );
  AND U1707 ( .A(n1035), .B(n1705), .Z(n1703) );
  XNOR U1708 ( .A(creg[79]), .B(n1704), .Z(n1705) );
  XNOR U1709 ( .A(n1706), .B(n1707), .Z(o[799]) );
  AND U1710 ( .A(n1035), .B(n1708), .Z(n1706) );
  XNOR U1711 ( .A(creg[799]), .B(n1707), .Z(n1708) );
  XNOR U1712 ( .A(n1709), .B(n1710), .Z(o[798]) );
  AND U1713 ( .A(n1035), .B(n1711), .Z(n1709) );
  XNOR U1714 ( .A(creg[798]), .B(n1710), .Z(n1711) );
  XNOR U1715 ( .A(n1712), .B(n1713), .Z(o[797]) );
  AND U1716 ( .A(n1035), .B(n1714), .Z(n1712) );
  XNOR U1717 ( .A(creg[797]), .B(n1713), .Z(n1714) );
  XNOR U1718 ( .A(n1715), .B(n1716), .Z(o[796]) );
  AND U1719 ( .A(n1035), .B(n1717), .Z(n1715) );
  XNOR U1720 ( .A(creg[796]), .B(n1716), .Z(n1717) );
  XNOR U1721 ( .A(n1718), .B(n1719), .Z(o[795]) );
  AND U1722 ( .A(n1035), .B(n1720), .Z(n1718) );
  XNOR U1723 ( .A(creg[795]), .B(n1719), .Z(n1720) );
  XNOR U1724 ( .A(n1721), .B(n1722), .Z(o[794]) );
  AND U1725 ( .A(n1035), .B(n1723), .Z(n1721) );
  XNOR U1726 ( .A(creg[794]), .B(n1722), .Z(n1723) );
  XNOR U1727 ( .A(n1724), .B(n1725), .Z(o[793]) );
  AND U1728 ( .A(n1035), .B(n1726), .Z(n1724) );
  XNOR U1729 ( .A(creg[793]), .B(n1725), .Z(n1726) );
  XNOR U1730 ( .A(n1727), .B(n1728), .Z(o[792]) );
  AND U1731 ( .A(n1035), .B(n1729), .Z(n1727) );
  XNOR U1732 ( .A(creg[792]), .B(n1728), .Z(n1729) );
  XNOR U1733 ( .A(n1730), .B(n1731), .Z(o[791]) );
  AND U1734 ( .A(n1035), .B(n1732), .Z(n1730) );
  XNOR U1735 ( .A(creg[791]), .B(n1731), .Z(n1732) );
  XNOR U1736 ( .A(n1733), .B(n1734), .Z(o[790]) );
  AND U1737 ( .A(n1035), .B(n1735), .Z(n1733) );
  XNOR U1738 ( .A(creg[790]), .B(n1734), .Z(n1735) );
  XNOR U1739 ( .A(n1736), .B(n1737), .Z(o[78]) );
  AND U1740 ( .A(n1035), .B(n1738), .Z(n1736) );
  XNOR U1741 ( .A(creg[78]), .B(n1737), .Z(n1738) );
  XNOR U1742 ( .A(n1739), .B(n1740), .Z(o[789]) );
  AND U1743 ( .A(n1035), .B(n1741), .Z(n1739) );
  XNOR U1744 ( .A(creg[789]), .B(n1740), .Z(n1741) );
  XNOR U1745 ( .A(n1742), .B(n1743), .Z(o[788]) );
  AND U1746 ( .A(n1035), .B(n1744), .Z(n1742) );
  XNOR U1747 ( .A(creg[788]), .B(n1743), .Z(n1744) );
  XNOR U1748 ( .A(n1745), .B(n1746), .Z(o[787]) );
  AND U1749 ( .A(n1035), .B(n1747), .Z(n1745) );
  XNOR U1750 ( .A(creg[787]), .B(n1746), .Z(n1747) );
  XNOR U1751 ( .A(n1748), .B(n1749), .Z(o[786]) );
  AND U1752 ( .A(n1035), .B(n1750), .Z(n1748) );
  XNOR U1753 ( .A(creg[786]), .B(n1749), .Z(n1750) );
  XNOR U1754 ( .A(n1751), .B(n1752), .Z(o[785]) );
  AND U1755 ( .A(n1035), .B(n1753), .Z(n1751) );
  XNOR U1756 ( .A(creg[785]), .B(n1752), .Z(n1753) );
  XNOR U1757 ( .A(n1754), .B(n1755), .Z(o[784]) );
  AND U1758 ( .A(n1035), .B(n1756), .Z(n1754) );
  XNOR U1759 ( .A(creg[784]), .B(n1755), .Z(n1756) );
  XNOR U1760 ( .A(n1757), .B(n1758), .Z(o[783]) );
  AND U1761 ( .A(n1035), .B(n1759), .Z(n1757) );
  XNOR U1762 ( .A(creg[783]), .B(n1758), .Z(n1759) );
  XNOR U1763 ( .A(n1760), .B(n1761), .Z(o[782]) );
  AND U1764 ( .A(n1035), .B(n1762), .Z(n1760) );
  XNOR U1765 ( .A(creg[782]), .B(n1761), .Z(n1762) );
  XNOR U1766 ( .A(n1763), .B(n1764), .Z(o[781]) );
  AND U1767 ( .A(n1035), .B(n1765), .Z(n1763) );
  XNOR U1768 ( .A(creg[781]), .B(n1764), .Z(n1765) );
  XNOR U1769 ( .A(n1766), .B(n1767), .Z(o[780]) );
  AND U1770 ( .A(n1035), .B(n1768), .Z(n1766) );
  XNOR U1771 ( .A(creg[780]), .B(n1767), .Z(n1768) );
  XNOR U1772 ( .A(n1769), .B(n1770), .Z(o[77]) );
  AND U1773 ( .A(n1035), .B(n1771), .Z(n1769) );
  XNOR U1774 ( .A(creg[77]), .B(n1770), .Z(n1771) );
  XNOR U1775 ( .A(n1772), .B(n1773), .Z(o[779]) );
  AND U1776 ( .A(n1035), .B(n1774), .Z(n1772) );
  XNOR U1777 ( .A(creg[779]), .B(n1773), .Z(n1774) );
  XNOR U1778 ( .A(n1775), .B(n1776), .Z(o[778]) );
  AND U1779 ( .A(n1035), .B(n1777), .Z(n1775) );
  XNOR U1780 ( .A(creg[778]), .B(n1776), .Z(n1777) );
  XNOR U1781 ( .A(n1778), .B(n1779), .Z(o[777]) );
  AND U1782 ( .A(n1035), .B(n1780), .Z(n1778) );
  XNOR U1783 ( .A(creg[777]), .B(n1779), .Z(n1780) );
  XNOR U1784 ( .A(n1781), .B(n1782), .Z(o[776]) );
  AND U1785 ( .A(n1035), .B(n1783), .Z(n1781) );
  XNOR U1786 ( .A(creg[776]), .B(n1782), .Z(n1783) );
  XNOR U1787 ( .A(n1784), .B(n1785), .Z(o[775]) );
  AND U1788 ( .A(n1035), .B(n1786), .Z(n1784) );
  XNOR U1789 ( .A(creg[775]), .B(n1785), .Z(n1786) );
  XNOR U1790 ( .A(n1787), .B(n1788), .Z(o[774]) );
  AND U1791 ( .A(n1035), .B(n1789), .Z(n1787) );
  XNOR U1792 ( .A(creg[774]), .B(n1788), .Z(n1789) );
  XNOR U1793 ( .A(n1790), .B(n1791), .Z(o[773]) );
  AND U1794 ( .A(n1035), .B(n1792), .Z(n1790) );
  XNOR U1795 ( .A(creg[773]), .B(n1791), .Z(n1792) );
  XNOR U1796 ( .A(n1793), .B(n1794), .Z(o[772]) );
  AND U1797 ( .A(n1035), .B(n1795), .Z(n1793) );
  XNOR U1798 ( .A(creg[772]), .B(n1794), .Z(n1795) );
  XNOR U1799 ( .A(n1796), .B(n1797), .Z(o[771]) );
  AND U1800 ( .A(n1035), .B(n1798), .Z(n1796) );
  XNOR U1801 ( .A(creg[771]), .B(n1797), .Z(n1798) );
  XNOR U1802 ( .A(n1799), .B(n1800), .Z(o[770]) );
  AND U1803 ( .A(n1035), .B(n1801), .Z(n1799) );
  XNOR U1804 ( .A(creg[770]), .B(n1800), .Z(n1801) );
  XNOR U1805 ( .A(n1802), .B(n1803), .Z(o[76]) );
  AND U1806 ( .A(n1035), .B(n1804), .Z(n1802) );
  XNOR U1807 ( .A(creg[76]), .B(n1803), .Z(n1804) );
  XNOR U1808 ( .A(n1805), .B(n1806), .Z(o[769]) );
  AND U1809 ( .A(n1035), .B(n1807), .Z(n1805) );
  XNOR U1810 ( .A(creg[769]), .B(n1806), .Z(n1807) );
  XNOR U1811 ( .A(n1808), .B(n1809), .Z(o[768]) );
  AND U1812 ( .A(n1035), .B(n1810), .Z(n1808) );
  XNOR U1813 ( .A(creg[768]), .B(n1809), .Z(n1810) );
  XNOR U1814 ( .A(n1811), .B(n1812), .Z(o[767]) );
  AND U1815 ( .A(n1035), .B(n1813), .Z(n1811) );
  XNOR U1816 ( .A(creg[767]), .B(n1812), .Z(n1813) );
  XNOR U1817 ( .A(n1814), .B(n1815), .Z(o[766]) );
  AND U1818 ( .A(n1035), .B(n1816), .Z(n1814) );
  XNOR U1819 ( .A(creg[766]), .B(n1815), .Z(n1816) );
  XNOR U1820 ( .A(n1817), .B(n1818), .Z(o[765]) );
  AND U1821 ( .A(n1035), .B(n1819), .Z(n1817) );
  XNOR U1822 ( .A(creg[765]), .B(n1818), .Z(n1819) );
  XNOR U1823 ( .A(n1820), .B(n1821), .Z(o[764]) );
  AND U1824 ( .A(n1035), .B(n1822), .Z(n1820) );
  XNOR U1825 ( .A(creg[764]), .B(n1821), .Z(n1822) );
  XNOR U1826 ( .A(n1823), .B(n1824), .Z(o[763]) );
  AND U1827 ( .A(n1035), .B(n1825), .Z(n1823) );
  XNOR U1828 ( .A(creg[763]), .B(n1824), .Z(n1825) );
  XNOR U1829 ( .A(n1826), .B(n1827), .Z(o[762]) );
  AND U1830 ( .A(n1035), .B(n1828), .Z(n1826) );
  XNOR U1831 ( .A(creg[762]), .B(n1827), .Z(n1828) );
  XNOR U1832 ( .A(n1829), .B(n1830), .Z(o[761]) );
  AND U1833 ( .A(n1035), .B(n1831), .Z(n1829) );
  XNOR U1834 ( .A(creg[761]), .B(n1830), .Z(n1831) );
  XNOR U1835 ( .A(n1832), .B(n1833), .Z(o[760]) );
  AND U1836 ( .A(n1035), .B(n1834), .Z(n1832) );
  XNOR U1837 ( .A(creg[760]), .B(n1833), .Z(n1834) );
  XNOR U1838 ( .A(n1835), .B(n1836), .Z(o[75]) );
  AND U1839 ( .A(n1035), .B(n1837), .Z(n1835) );
  XNOR U1840 ( .A(creg[75]), .B(n1836), .Z(n1837) );
  XNOR U1841 ( .A(n1838), .B(n1839), .Z(o[759]) );
  AND U1842 ( .A(n1035), .B(n1840), .Z(n1838) );
  XNOR U1843 ( .A(creg[759]), .B(n1839), .Z(n1840) );
  XNOR U1844 ( .A(n1841), .B(n1842), .Z(o[758]) );
  AND U1845 ( .A(n1035), .B(n1843), .Z(n1841) );
  XNOR U1846 ( .A(creg[758]), .B(n1842), .Z(n1843) );
  XNOR U1847 ( .A(n1844), .B(n1845), .Z(o[757]) );
  AND U1848 ( .A(n1035), .B(n1846), .Z(n1844) );
  XNOR U1849 ( .A(creg[757]), .B(n1845), .Z(n1846) );
  XNOR U1850 ( .A(n1847), .B(n1848), .Z(o[756]) );
  AND U1851 ( .A(n1035), .B(n1849), .Z(n1847) );
  XNOR U1852 ( .A(creg[756]), .B(n1848), .Z(n1849) );
  XNOR U1853 ( .A(n1850), .B(n1851), .Z(o[755]) );
  AND U1854 ( .A(n1035), .B(n1852), .Z(n1850) );
  XNOR U1855 ( .A(creg[755]), .B(n1851), .Z(n1852) );
  XNOR U1856 ( .A(n1853), .B(n1854), .Z(o[754]) );
  AND U1857 ( .A(n1035), .B(n1855), .Z(n1853) );
  XNOR U1858 ( .A(creg[754]), .B(n1854), .Z(n1855) );
  XNOR U1859 ( .A(n1856), .B(n1857), .Z(o[753]) );
  AND U1860 ( .A(n1035), .B(n1858), .Z(n1856) );
  XNOR U1861 ( .A(creg[753]), .B(n1857), .Z(n1858) );
  XNOR U1862 ( .A(n1859), .B(n1860), .Z(o[752]) );
  AND U1863 ( .A(n1035), .B(n1861), .Z(n1859) );
  XNOR U1864 ( .A(creg[752]), .B(n1860), .Z(n1861) );
  XNOR U1865 ( .A(n1862), .B(n1863), .Z(o[751]) );
  AND U1866 ( .A(n1035), .B(n1864), .Z(n1862) );
  XNOR U1867 ( .A(creg[751]), .B(n1863), .Z(n1864) );
  XNOR U1868 ( .A(n1865), .B(n1866), .Z(o[750]) );
  AND U1869 ( .A(n1035), .B(n1867), .Z(n1865) );
  XNOR U1870 ( .A(creg[750]), .B(n1866), .Z(n1867) );
  XNOR U1871 ( .A(n1868), .B(n1869), .Z(o[74]) );
  AND U1872 ( .A(n1035), .B(n1870), .Z(n1868) );
  XNOR U1873 ( .A(creg[74]), .B(n1869), .Z(n1870) );
  XNOR U1874 ( .A(n1871), .B(n1872), .Z(o[749]) );
  AND U1875 ( .A(n1035), .B(n1873), .Z(n1871) );
  XNOR U1876 ( .A(creg[749]), .B(n1872), .Z(n1873) );
  XNOR U1877 ( .A(n1874), .B(n1875), .Z(o[748]) );
  AND U1878 ( .A(n1035), .B(n1876), .Z(n1874) );
  XNOR U1879 ( .A(creg[748]), .B(n1875), .Z(n1876) );
  XNOR U1880 ( .A(n1877), .B(n1878), .Z(o[747]) );
  AND U1881 ( .A(n1035), .B(n1879), .Z(n1877) );
  XNOR U1882 ( .A(creg[747]), .B(n1878), .Z(n1879) );
  XNOR U1883 ( .A(n1880), .B(n1881), .Z(o[746]) );
  AND U1884 ( .A(n1035), .B(n1882), .Z(n1880) );
  XNOR U1885 ( .A(creg[746]), .B(n1881), .Z(n1882) );
  XNOR U1886 ( .A(n1883), .B(n1884), .Z(o[745]) );
  AND U1887 ( .A(n1035), .B(n1885), .Z(n1883) );
  XNOR U1888 ( .A(creg[745]), .B(n1884), .Z(n1885) );
  XNOR U1889 ( .A(n1886), .B(n1887), .Z(o[744]) );
  AND U1890 ( .A(n1035), .B(n1888), .Z(n1886) );
  XNOR U1891 ( .A(creg[744]), .B(n1887), .Z(n1888) );
  XNOR U1892 ( .A(n1889), .B(n1890), .Z(o[743]) );
  AND U1893 ( .A(n1035), .B(n1891), .Z(n1889) );
  XNOR U1894 ( .A(creg[743]), .B(n1890), .Z(n1891) );
  XNOR U1895 ( .A(n1892), .B(n1893), .Z(o[742]) );
  AND U1896 ( .A(n1035), .B(n1894), .Z(n1892) );
  XNOR U1897 ( .A(creg[742]), .B(n1893), .Z(n1894) );
  XNOR U1898 ( .A(n1895), .B(n1896), .Z(o[741]) );
  AND U1899 ( .A(n1035), .B(n1897), .Z(n1895) );
  XNOR U1900 ( .A(creg[741]), .B(n1896), .Z(n1897) );
  XNOR U1901 ( .A(n1898), .B(n1899), .Z(o[740]) );
  AND U1902 ( .A(n1035), .B(n1900), .Z(n1898) );
  XNOR U1903 ( .A(creg[740]), .B(n1899), .Z(n1900) );
  XNOR U1904 ( .A(n1901), .B(n1902), .Z(o[73]) );
  AND U1905 ( .A(n1035), .B(n1903), .Z(n1901) );
  XNOR U1906 ( .A(creg[73]), .B(n1902), .Z(n1903) );
  XNOR U1907 ( .A(n1904), .B(n1905), .Z(o[739]) );
  AND U1908 ( .A(n1035), .B(n1906), .Z(n1904) );
  XNOR U1909 ( .A(creg[739]), .B(n1905), .Z(n1906) );
  XNOR U1910 ( .A(n1907), .B(n1908), .Z(o[738]) );
  AND U1911 ( .A(n1035), .B(n1909), .Z(n1907) );
  XNOR U1912 ( .A(creg[738]), .B(n1908), .Z(n1909) );
  XNOR U1913 ( .A(n1910), .B(n1911), .Z(o[737]) );
  AND U1914 ( .A(n1035), .B(n1912), .Z(n1910) );
  XNOR U1915 ( .A(creg[737]), .B(n1911), .Z(n1912) );
  XNOR U1916 ( .A(n1913), .B(n1914), .Z(o[736]) );
  AND U1917 ( .A(n1035), .B(n1915), .Z(n1913) );
  XNOR U1918 ( .A(creg[736]), .B(n1914), .Z(n1915) );
  XNOR U1919 ( .A(n1916), .B(n1917), .Z(o[735]) );
  AND U1920 ( .A(n1035), .B(n1918), .Z(n1916) );
  XNOR U1921 ( .A(creg[735]), .B(n1917), .Z(n1918) );
  XNOR U1922 ( .A(n1919), .B(n1920), .Z(o[734]) );
  AND U1923 ( .A(n1035), .B(n1921), .Z(n1919) );
  XNOR U1924 ( .A(creg[734]), .B(n1920), .Z(n1921) );
  XNOR U1925 ( .A(n1922), .B(n1923), .Z(o[733]) );
  AND U1926 ( .A(n1035), .B(n1924), .Z(n1922) );
  XNOR U1927 ( .A(creg[733]), .B(n1923), .Z(n1924) );
  XNOR U1928 ( .A(n1925), .B(n1926), .Z(o[732]) );
  AND U1929 ( .A(n1035), .B(n1927), .Z(n1925) );
  XNOR U1930 ( .A(creg[732]), .B(n1926), .Z(n1927) );
  XNOR U1931 ( .A(n1928), .B(n1929), .Z(o[731]) );
  AND U1932 ( .A(n1035), .B(n1930), .Z(n1928) );
  XNOR U1933 ( .A(creg[731]), .B(n1929), .Z(n1930) );
  XNOR U1934 ( .A(n1931), .B(n1932), .Z(o[730]) );
  AND U1935 ( .A(n1035), .B(n1933), .Z(n1931) );
  XNOR U1936 ( .A(creg[730]), .B(n1932), .Z(n1933) );
  XNOR U1937 ( .A(n1934), .B(n1935), .Z(o[72]) );
  AND U1938 ( .A(n1035), .B(n1936), .Z(n1934) );
  XNOR U1939 ( .A(creg[72]), .B(n1935), .Z(n1936) );
  XNOR U1940 ( .A(n1937), .B(n1938), .Z(o[729]) );
  AND U1941 ( .A(n1035), .B(n1939), .Z(n1937) );
  XNOR U1942 ( .A(creg[729]), .B(n1938), .Z(n1939) );
  XNOR U1943 ( .A(n1940), .B(n1941), .Z(o[728]) );
  AND U1944 ( .A(n1035), .B(n1942), .Z(n1940) );
  XNOR U1945 ( .A(creg[728]), .B(n1941), .Z(n1942) );
  XNOR U1946 ( .A(n1943), .B(n1944), .Z(o[727]) );
  AND U1947 ( .A(n1035), .B(n1945), .Z(n1943) );
  XNOR U1948 ( .A(creg[727]), .B(n1944), .Z(n1945) );
  XNOR U1949 ( .A(n1946), .B(n1947), .Z(o[726]) );
  AND U1950 ( .A(n1035), .B(n1948), .Z(n1946) );
  XNOR U1951 ( .A(creg[726]), .B(n1947), .Z(n1948) );
  XNOR U1952 ( .A(n1949), .B(n1950), .Z(o[725]) );
  AND U1953 ( .A(n1035), .B(n1951), .Z(n1949) );
  XNOR U1954 ( .A(creg[725]), .B(n1950), .Z(n1951) );
  XNOR U1955 ( .A(n1952), .B(n1953), .Z(o[724]) );
  AND U1956 ( .A(n1035), .B(n1954), .Z(n1952) );
  XNOR U1957 ( .A(creg[724]), .B(n1953), .Z(n1954) );
  XNOR U1958 ( .A(n1955), .B(n1956), .Z(o[723]) );
  AND U1959 ( .A(n1035), .B(n1957), .Z(n1955) );
  XNOR U1960 ( .A(creg[723]), .B(n1956), .Z(n1957) );
  XNOR U1961 ( .A(n1958), .B(n1959), .Z(o[722]) );
  AND U1962 ( .A(n1035), .B(n1960), .Z(n1958) );
  XNOR U1963 ( .A(creg[722]), .B(n1959), .Z(n1960) );
  XNOR U1964 ( .A(n1961), .B(n1962), .Z(o[721]) );
  AND U1965 ( .A(n1035), .B(n1963), .Z(n1961) );
  XNOR U1966 ( .A(creg[721]), .B(n1962), .Z(n1963) );
  XNOR U1967 ( .A(n1964), .B(n1965), .Z(o[720]) );
  AND U1968 ( .A(n1035), .B(n1966), .Z(n1964) );
  XNOR U1969 ( .A(creg[720]), .B(n1965), .Z(n1966) );
  XNOR U1970 ( .A(n1967), .B(n1968), .Z(o[71]) );
  AND U1971 ( .A(n1035), .B(n1969), .Z(n1967) );
  XNOR U1972 ( .A(creg[71]), .B(n1968), .Z(n1969) );
  XNOR U1973 ( .A(n1970), .B(n1971), .Z(o[719]) );
  AND U1974 ( .A(n1035), .B(n1972), .Z(n1970) );
  XNOR U1975 ( .A(creg[719]), .B(n1971), .Z(n1972) );
  XNOR U1976 ( .A(n1973), .B(n1974), .Z(o[718]) );
  AND U1977 ( .A(n1035), .B(n1975), .Z(n1973) );
  XNOR U1978 ( .A(creg[718]), .B(n1974), .Z(n1975) );
  XNOR U1979 ( .A(n1976), .B(n1977), .Z(o[717]) );
  AND U1980 ( .A(n1035), .B(n1978), .Z(n1976) );
  XNOR U1981 ( .A(creg[717]), .B(n1977), .Z(n1978) );
  XNOR U1982 ( .A(n1979), .B(n1980), .Z(o[716]) );
  AND U1983 ( .A(n1035), .B(n1981), .Z(n1979) );
  XNOR U1984 ( .A(creg[716]), .B(n1980), .Z(n1981) );
  XNOR U1985 ( .A(n1982), .B(n1983), .Z(o[715]) );
  AND U1986 ( .A(n1035), .B(n1984), .Z(n1982) );
  XNOR U1987 ( .A(creg[715]), .B(n1983), .Z(n1984) );
  XNOR U1988 ( .A(n1985), .B(n1986), .Z(o[714]) );
  AND U1989 ( .A(n1035), .B(n1987), .Z(n1985) );
  XNOR U1990 ( .A(creg[714]), .B(n1986), .Z(n1987) );
  XNOR U1991 ( .A(n1988), .B(n1989), .Z(o[713]) );
  AND U1992 ( .A(n1035), .B(n1990), .Z(n1988) );
  XNOR U1993 ( .A(creg[713]), .B(n1989), .Z(n1990) );
  XNOR U1994 ( .A(n1991), .B(n1992), .Z(o[712]) );
  AND U1995 ( .A(n1035), .B(n1993), .Z(n1991) );
  XNOR U1996 ( .A(creg[712]), .B(n1992), .Z(n1993) );
  XNOR U1997 ( .A(n1994), .B(n1995), .Z(o[711]) );
  AND U1998 ( .A(n1035), .B(n1996), .Z(n1994) );
  XNOR U1999 ( .A(creg[711]), .B(n1995), .Z(n1996) );
  XNOR U2000 ( .A(n1997), .B(n1998), .Z(o[710]) );
  AND U2001 ( .A(n1035), .B(n1999), .Z(n1997) );
  XNOR U2002 ( .A(creg[710]), .B(n1998), .Z(n1999) );
  XNOR U2003 ( .A(n2000), .B(n2001), .Z(o[70]) );
  AND U2004 ( .A(n1035), .B(n2002), .Z(n2000) );
  XNOR U2005 ( .A(creg[70]), .B(n2001), .Z(n2002) );
  XNOR U2006 ( .A(n2003), .B(n2004), .Z(o[709]) );
  AND U2007 ( .A(n1035), .B(n2005), .Z(n2003) );
  XNOR U2008 ( .A(creg[709]), .B(n2004), .Z(n2005) );
  XNOR U2009 ( .A(n2006), .B(n2007), .Z(o[708]) );
  AND U2010 ( .A(n1035), .B(n2008), .Z(n2006) );
  XNOR U2011 ( .A(creg[708]), .B(n2007), .Z(n2008) );
  XNOR U2012 ( .A(n2009), .B(n2010), .Z(o[707]) );
  AND U2013 ( .A(n1035), .B(n2011), .Z(n2009) );
  XNOR U2014 ( .A(creg[707]), .B(n2010), .Z(n2011) );
  XNOR U2015 ( .A(n2012), .B(n2013), .Z(o[706]) );
  AND U2016 ( .A(n1035), .B(n2014), .Z(n2012) );
  XNOR U2017 ( .A(creg[706]), .B(n2013), .Z(n2014) );
  XNOR U2018 ( .A(n2015), .B(n2016), .Z(o[705]) );
  AND U2019 ( .A(n1035), .B(n2017), .Z(n2015) );
  XNOR U2020 ( .A(creg[705]), .B(n2016), .Z(n2017) );
  XNOR U2021 ( .A(n2018), .B(n2019), .Z(o[704]) );
  AND U2022 ( .A(n1035), .B(n2020), .Z(n2018) );
  XNOR U2023 ( .A(creg[704]), .B(n2019), .Z(n2020) );
  XNOR U2024 ( .A(n2021), .B(n2022), .Z(o[703]) );
  AND U2025 ( .A(n1035), .B(n2023), .Z(n2021) );
  XNOR U2026 ( .A(creg[703]), .B(n2022), .Z(n2023) );
  XNOR U2027 ( .A(n2024), .B(n2025), .Z(o[702]) );
  AND U2028 ( .A(n1035), .B(n2026), .Z(n2024) );
  XNOR U2029 ( .A(creg[702]), .B(n2025), .Z(n2026) );
  XNOR U2030 ( .A(n2027), .B(n2028), .Z(o[701]) );
  AND U2031 ( .A(n1035), .B(n2029), .Z(n2027) );
  XNOR U2032 ( .A(creg[701]), .B(n2028), .Z(n2029) );
  XNOR U2033 ( .A(n2030), .B(n2031), .Z(o[700]) );
  AND U2034 ( .A(n1035), .B(n2032), .Z(n2030) );
  XNOR U2035 ( .A(creg[700]), .B(n2031), .Z(n2032) );
  XNOR U2036 ( .A(n2033), .B(n2034), .Z(o[6]) );
  AND U2037 ( .A(n1035), .B(n2035), .Z(n2033) );
  XNOR U2038 ( .A(creg[6]), .B(n2034), .Z(n2035) );
  XNOR U2039 ( .A(n2036), .B(n2037), .Z(o[69]) );
  AND U2040 ( .A(n1035), .B(n2038), .Z(n2036) );
  XNOR U2041 ( .A(creg[69]), .B(n2037), .Z(n2038) );
  XNOR U2042 ( .A(n2039), .B(n2040), .Z(o[699]) );
  AND U2043 ( .A(n1035), .B(n2041), .Z(n2039) );
  XNOR U2044 ( .A(creg[699]), .B(n2040), .Z(n2041) );
  XNOR U2045 ( .A(n2042), .B(n2043), .Z(o[698]) );
  AND U2046 ( .A(n1035), .B(n2044), .Z(n2042) );
  XNOR U2047 ( .A(creg[698]), .B(n2043), .Z(n2044) );
  XNOR U2048 ( .A(n2045), .B(n2046), .Z(o[697]) );
  AND U2049 ( .A(n1035), .B(n2047), .Z(n2045) );
  XNOR U2050 ( .A(creg[697]), .B(n2046), .Z(n2047) );
  XNOR U2051 ( .A(n2048), .B(n2049), .Z(o[696]) );
  AND U2052 ( .A(n1035), .B(n2050), .Z(n2048) );
  XNOR U2053 ( .A(creg[696]), .B(n2049), .Z(n2050) );
  XNOR U2054 ( .A(n2051), .B(n2052), .Z(o[695]) );
  AND U2055 ( .A(n1035), .B(n2053), .Z(n2051) );
  XNOR U2056 ( .A(creg[695]), .B(n2052), .Z(n2053) );
  XNOR U2057 ( .A(n2054), .B(n2055), .Z(o[694]) );
  AND U2058 ( .A(n1035), .B(n2056), .Z(n2054) );
  XNOR U2059 ( .A(creg[694]), .B(n2055), .Z(n2056) );
  XNOR U2060 ( .A(n2057), .B(n2058), .Z(o[693]) );
  AND U2061 ( .A(n1035), .B(n2059), .Z(n2057) );
  XNOR U2062 ( .A(creg[693]), .B(n2058), .Z(n2059) );
  XNOR U2063 ( .A(n2060), .B(n2061), .Z(o[692]) );
  AND U2064 ( .A(n1035), .B(n2062), .Z(n2060) );
  XNOR U2065 ( .A(creg[692]), .B(n2061), .Z(n2062) );
  XNOR U2066 ( .A(n2063), .B(n2064), .Z(o[691]) );
  AND U2067 ( .A(n1035), .B(n2065), .Z(n2063) );
  XNOR U2068 ( .A(creg[691]), .B(n2064), .Z(n2065) );
  XNOR U2069 ( .A(n2066), .B(n2067), .Z(o[690]) );
  AND U2070 ( .A(n1035), .B(n2068), .Z(n2066) );
  XNOR U2071 ( .A(creg[690]), .B(n2067), .Z(n2068) );
  XNOR U2072 ( .A(n2069), .B(n2070), .Z(o[68]) );
  AND U2073 ( .A(n1035), .B(n2071), .Z(n2069) );
  XNOR U2074 ( .A(creg[68]), .B(n2070), .Z(n2071) );
  XNOR U2075 ( .A(n2072), .B(n2073), .Z(o[689]) );
  AND U2076 ( .A(n1035), .B(n2074), .Z(n2072) );
  XNOR U2077 ( .A(creg[689]), .B(n2073), .Z(n2074) );
  XNOR U2078 ( .A(n2075), .B(n2076), .Z(o[688]) );
  AND U2079 ( .A(n1035), .B(n2077), .Z(n2075) );
  XNOR U2080 ( .A(creg[688]), .B(n2076), .Z(n2077) );
  XNOR U2081 ( .A(n2078), .B(n2079), .Z(o[687]) );
  AND U2082 ( .A(n1035), .B(n2080), .Z(n2078) );
  XNOR U2083 ( .A(creg[687]), .B(n2079), .Z(n2080) );
  XNOR U2084 ( .A(n2081), .B(n2082), .Z(o[686]) );
  AND U2085 ( .A(n1035), .B(n2083), .Z(n2081) );
  XNOR U2086 ( .A(creg[686]), .B(n2082), .Z(n2083) );
  XNOR U2087 ( .A(n2084), .B(n2085), .Z(o[685]) );
  AND U2088 ( .A(n1035), .B(n2086), .Z(n2084) );
  XNOR U2089 ( .A(creg[685]), .B(n2085), .Z(n2086) );
  XNOR U2090 ( .A(n2087), .B(n2088), .Z(o[684]) );
  AND U2091 ( .A(n1035), .B(n2089), .Z(n2087) );
  XNOR U2092 ( .A(creg[684]), .B(n2088), .Z(n2089) );
  XNOR U2093 ( .A(n2090), .B(n2091), .Z(o[683]) );
  AND U2094 ( .A(n1035), .B(n2092), .Z(n2090) );
  XNOR U2095 ( .A(creg[683]), .B(n2091), .Z(n2092) );
  XNOR U2096 ( .A(n2093), .B(n2094), .Z(o[682]) );
  AND U2097 ( .A(n1035), .B(n2095), .Z(n2093) );
  XNOR U2098 ( .A(creg[682]), .B(n2094), .Z(n2095) );
  XNOR U2099 ( .A(n2096), .B(n2097), .Z(o[681]) );
  AND U2100 ( .A(n1035), .B(n2098), .Z(n2096) );
  XNOR U2101 ( .A(creg[681]), .B(n2097), .Z(n2098) );
  XNOR U2102 ( .A(n2099), .B(n2100), .Z(o[680]) );
  AND U2103 ( .A(n1035), .B(n2101), .Z(n2099) );
  XNOR U2104 ( .A(creg[680]), .B(n2100), .Z(n2101) );
  XNOR U2105 ( .A(n2102), .B(n2103), .Z(o[67]) );
  AND U2106 ( .A(n1035), .B(n2104), .Z(n2102) );
  XNOR U2107 ( .A(creg[67]), .B(n2103), .Z(n2104) );
  XNOR U2108 ( .A(n2105), .B(n2106), .Z(o[679]) );
  AND U2109 ( .A(n1035), .B(n2107), .Z(n2105) );
  XNOR U2110 ( .A(creg[679]), .B(n2106), .Z(n2107) );
  XNOR U2111 ( .A(n2108), .B(n2109), .Z(o[678]) );
  AND U2112 ( .A(n1035), .B(n2110), .Z(n2108) );
  XNOR U2113 ( .A(creg[678]), .B(n2109), .Z(n2110) );
  XNOR U2114 ( .A(n2111), .B(n2112), .Z(o[677]) );
  AND U2115 ( .A(n1035), .B(n2113), .Z(n2111) );
  XNOR U2116 ( .A(creg[677]), .B(n2112), .Z(n2113) );
  XNOR U2117 ( .A(n2114), .B(n2115), .Z(o[676]) );
  AND U2118 ( .A(n1035), .B(n2116), .Z(n2114) );
  XNOR U2119 ( .A(creg[676]), .B(n2115), .Z(n2116) );
  XNOR U2120 ( .A(n2117), .B(n2118), .Z(o[675]) );
  AND U2121 ( .A(n1035), .B(n2119), .Z(n2117) );
  XNOR U2122 ( .A(creg[675]), .B(n2118), .Z(n2119) );
  XNOR U2123 ( .A(n2120), .B(n2121), .Z(o[674]) );
  AND U2124 ( .A(n1035), .B(n2122), .Z(n2120) );
  XNOR U2125 ( .A(creg[674]), .B(n2121), .Z(n2122) );
  XNOR U2126 ( .A(n2123), .B(n2124), .Z(o[673]) );
  AND U2127 ( .A(n1035), .B(n2125), .Z(n2123) );
  XNOR U2128 ( .A(creg[673]), .B(n2124), .Z(n2125) );
  XNOR U2129 ( .A(n2126), .B(n2127), .Z(o[672]) );
  AND U2130 ( .A(n1035), .B(n2128), .Z(n2126) );
  XNOR U2131 ( .A(creg[672]), .B(n2127), .Z(n2128) );
  XNOR U2132 ( .A(n2129), .B(n2130), .Z(o[671]) );
  AND U2133 ( .A(n1035), .B(n2131), .Z(n2129) );
  XNOR U2134 ( .A(creg[671]), .B(n2130), .Z(n2131) );
  XNOR U2135 ( .A(n2132), .B(n2133), .Z(o[670]) );
  AND U2136 ( .A(n1035), .B(n2134), .Z(n2132) );
  XNOR U2137 ( .A(creg[670]), .B(n2133), .Z(n2134) );
  XNOR U2138 ( .A(n2135), .B(n2136), .Z(o[66]) );
  AND U2139 ( .A(n1035), .B(n2137), .Z(n2135) );
  XNOR U2140 ( .A(creg[66]), .B(n2136), .Z(n2137) );
  XNOR U2141 ( .A(n2138), .B(n2139), .Z(o[669]) );
  AND U2142 ( .A(n1035), .B(n2140), .Z(n2138) );
  XNOR U2143 ( .A(creg[669]), .B(n2139), .Z(n2140) );
  XNOR U2144 ( .A(n2141), .B(n2142), .Z(o[668]) );
  AND U2145 ( .A(n1035), .B(n2143), .Z(n2141) );
  XNOR U2146 ( .A(creg[668]), .B(n2142), .Z(n2143) );
  XNOR U2147 ( .A(n2144), .B(n2145), .Z(o[667]) );
  AND U2148 ( .A(n1035), .B(n2146), .Z(n2144) );
  XNOR U2149 ( .A(creg[667]), .B(n2145), .Z(n2146) );
  XNOR U2150 ( .A(n2147), .B(n2148), .Z(o[666]) );
  AND U2151 ( .A(n1035), .B(n2149), .Z(n2147) );
  XNOR U2152 ( .A(creg[666]), .B(n2148), .Z(n2149) );
  XNOR U2153 ( .A(n2150), .B(n2151), .Z(o[665]) );
  AND U2154 ( .A(n1035), .B(n2152), .Z(n2150) );
  XNOR U2155 ( .A(creg[665]), .B(n2151), .Z(n2152) );
  XNOR U2156 ( .A(n2153), .B(n2154), .Z(o[664]) );
  AND U2157 ( .A(n1035), .B(n2155), .Z(n2153) );
  XNOR U2158 ( .A(creg[664]), .B(n2154), .Z(n2155) );
  XNOR U2159 ( .A(n2156), .B(n2157), .Z(o[663]) );
  AND U2160 ( .A(n1035), .B(n2158), .Z(n2156) );
  XNOR U2161 ( .A(creg[663]), .B(n2157), .Z(n2158) );
  XNOR U2162 ( .A(n2159), .B(n2160), .Z(o[662]) );
  AND U2163 ( .A(n1035), .B(n2161), .Z(n2159) );
  XNOR U2164 ( .A(creg[662]), .B(n2160), .Z(n2161) );
  XNOR U2165 ( .A(n2162), .B(n2163), .Z(o[661]) );
  AND U2166 ( .A(n1035), .B(n2164), .Z(n2162) );
  XNOR U2167 ( .A(creg[661]), .B(n2163), .Z(n2164) );
  XNOR U2168 ( .A(n2165), .B(n2166), .Z(o[660]) );
  AND U2169 ( .A(n1035), .B(n2167), .Z(n2165) );
  XNOR U2170 ( .A(creg[660]), .B(n2166), .Z(n2167) );
  XNOR U2171 ( .A(n2168), .B(n2169), .Z(o[65]) );
  AND U2172 ( .A(n1035), .B(n2170), .Z(n2168) );
  XNOR U2173 ( .A(creg[65]), .B(n2169), .Z(n2170) );
  XNOR U2174 ( .A(n2171), .B(n2172), .Z(o[659]) );
  AND U2175 ( .A(n1035), .B(n2173), .Z(n2171) );
  XNOR U2176 ( .A(creg[659]), .B(n2172), .Z(n2173) );
  XNOR U2177 ( .A(n2174), .B(n2175), .Z(o[658]) );
  AND U2178 ( .A(n1035), .B(n2176), .Z(n2174) );
  XNOR U2179 ( .A(creg[658]), .B(n2175), .Z(n2176) );
  XNOR U2180 ( .A(n2177), .B(n2178), .Z(o[657]) );
  AND U2181 ( .A(n1035), .B(n2179), .Z(n2177) );
  XNOR U2182 ( .A(creg[657]), .B(n2178), .Z(n2179) );
  XNOR U2183 ( .A(n2180), .B(n2181), .Z(o[656]) );
  AND U2184 ( .A(n1035), .B(n2182), .Z(n2180) );
  XNOR U2185 ( .A(creg[656]), .B(n2181), .Z(n2182) );
  XNOR U2186 ( .A(n2183), .B(n2184), .Z(o[655]) );
  AND U2187 ( .A(n1035), .B(n2185), .Z(n2183) );
  XNOR U2188 ( .A(creg[655]), .B(n2184), .Z(n2185) );
  XNOR U2189 ( .A(n2186), .B(n2187), .Z(o[654]) );
  AND U2190 ( .A(n1035), .B(n2188), .Z(n2186) );
  XNOR U2191 ( .A(creg[654]), .B(n2187), .Z(n2188) );
  XNOR U2192 ( .A(n2189), .B(n2190), .Z(o[653]) );
  AND U2193 ( .A(n1035), .B(n2191), .Z(n2189) );
  XNOR U2194 ( .A(creg[653]), .B(n2190), .Z(n2191) );
  XNOR U2195 ( .A(n2192), .B(n2193), .Z(o[652]) );
  AND U2196 ( .A(n1035), .B(n2194), .Z(n2192) );
  XNOR U2197 ( .A(creg[652]), .B(n2193), .Z(n2194) );
  XNOR U2198 ( .A(n2195), .B(n2196), .Z(o[651]) );
  AND U2199 ( .A(n1035), .B(n2197), .Z(n2195) );
  XNOR U2200 ( .A(creg[651]), .B(n2196), .Z(n2197) );
  XNOR U2201 ( .A(n2198), .B(n2199), .Z(o[650]) );
  AND U2202 ( .A(n1035), .B(n2200), .Z(n2198) );
  XNOR U2203 ( .A(creg[650]), .B(n2199), .Z(n2200) );
  XNOR U2204 ( .A(n2201), .B(n2202), .Z(o[64]) );
  AND U2205 ( .A(n1035), .B(n2203), .Z(n2201) );
  XNOR U2206 ( .A(creg[64]), .B(n2202), .Z(n2203) );
  XNOR U2207 ( .A(n2204), .B(n2205), .Z(o[649]) );
  AND U2208 ( .A(n1035), .B(n2206), .Z(n2204) );
  XNOR U2209 ( .A(creg[649]), .B(n2205), .Z(n2206) );
  XNOR U2210 ( .A(n2207), .B(n2208), .Z(o[648]) );
  AND U2211 ( .A(n1035), .B(n2209), .Z(n2207) );
  XNOR U2212 ( .A(creg[648]), .B(n2208), .Z(n2209) );
  XNOR U2213 ( .A(n2210), .B(n2211), .Z(o[647]) );
  AND U2214 ( .A(n1035), .B(n2212), .Z(n2210) );
  XNOR U2215 ( .A(creg[647]), .B(n2211), .Z(n2212) );
  XNOR U2216 ( .A(n2213), .B(n2214), .Z(o[646]) );
  AND U2217 ( .A(n1035), .B(n2215), .Z(n2213) );
  XNOR U2218 ( .A(creg[646]), .B(n2214), .Z(n2215) );
  XNOR U2219 ( .A(n2216), .B(n2217), .Z(o[645]) );
  AND U2220 ( .A(n1035), .B(n2218), .Z(n2216) );
  XNOR U2221 ( .A(creg[645]), .B(n2217), .Z(n2218) );
  XNOR U2222 ( .A(n2219), .B(n2220), .Z(o[644]) );
  AND U2223 ( .A(n1035), .B(n2221), .Z(n2219) );
  XNOR U2224 ( .A(creg[644]), .B(n2220), .Z(n2221) );
  XNOR U2225 ( .A(n2222), .B(n2223), .Z(o[643]) );
  AND U2226 ( .A(n1035), .B(n2224), .Z(n2222) );
  XNOR U2227 ( .A(creg[643]), .B(n2223), .Z(n2224) );
  XNOR U2228 ( .A(n2225), .B(n2226), .Z(o[642]) );
  AND U2229 ( .A(n1035), .B(n2227), .Z(n2225) );
  XNOR U2230 ( .A(creg[642]), .B(n2226), .Z(n2227) );
  XNOR U2231 ( .A(n2228), .B(n2229), .Z(o[641]) );
  AND U2232 ( .A(n1035), .B(n2230), .Z(n2228) );
  XNOR U2233 ( .A(creg[641]), .B(n2229), .Z(n2230) );
  XNOR U2234 ( .A(n2231), .B(n2232), .Z(o[640]) );
  AND U2235 ( .A(n1035), .B(n2233), .Z(n2231) );
  XNOR U2236 ( .A(creg[640]), .B(n2232), .Z(n2233) );
  XNOR U2237 ( .A(n2234), .B(n2235), .Z(o[63]) );
  AND U2238 ( .A(n1035), .B(n2236), .Z(n2234) );
  XNOR U2239 ( .A(creg[63]), .B(n2235), .Z(n2236) );
  XNOR U2240 ( .A(n2237), .B(n2238), .Z(o[639]) );
  AND U2241 ( .A(n1035), .B(n2239), .Z(n2237) );
  XNOR U2242 ( .A(creg[639]), .B(n2238), .Z(n2239) );
  XNOR U2243 ( .A(n2240), .B(n2241), .Z(o[638]) );
  AND U2244 ( .A(n1035), .B(n2242), .Z(n2240) );
  XNOR U2245 ( .A(creg[638]), .B(n2241), .Z(n2242) );
  XNOR U2246 ( .A(n2243), .B(n2244), .Z(o[637]) );
  AND U2247 ( .A(n1035), .B(n2245), .Z(n2243) );
  XNOR U2248 ( .A(creg[637]), .B(n2244), .Z(n2245) );
  XNOR U2249 ( .A(n2246), .B(n2247), .Z(o[636]) );
  AND U2250 ( .A(n1035), .B(n2248), .Z(n2246) );
  XNOR U2251 ( .A(creg[636]), .B(n2247), .Z(n2248) );
  XNOR U2252 ( .A(n2249), .B(n2250), .Z(o[635]) );
  AND U2253 ( .A(n1035), .B(n2251), .Z(n2249) );
  XNOR U2254 ( .A(creg[635]), .B(n2250), .Z(n2251) );
  XNOR U2255 ( .A(n2252), .B(n2253), .Z(o[634]) );
  AND U2256 ( .A(n1035), .B(n2254), .Z(n2252) );
  XNOR U2257 ( .A(creg[634]), .B(n2253), .Z(n2254) );
  XNOR U2258 ( .A(n2255), .B(n2256), .Z(o[633]) );
  AND U2259 ( .A(n1035), .B(n2257), .Z(n2255) );
  XNOR U2260 ( .A(creg[633]), .B(n2256), .Z(n2257) );
  XNOR U2261 ( .A(n2258), .B(n2259), .Z(o[632]) );
  AND U2262 ( .A(n1035), .B(n2260), .Z(n2258) );
  XNOR U2263 ( .A(creg[632]), .B(n2259), .Z(n2260) );
  XNOR U2264 ( .A(n2261), .B(n2262), .Z(o[631]) );
  AND U2265 ( .A(n1035), .B(n2263), .Z(n2261) );
  XNOR U2266 ( .A(creg[631]), .B(n2262), .Z(n2263) );
  XNOR U2267 ( .A(n2264), .B(n2265), .Z(o[630]) );
  AND U2268 ( .A(n1035), .B(n2266), .Z(n2264) );
  XNOR U2269 ( .A(creg[630]), .B(n2265), .Z(n2266) );
  XNOR U2270 ( .A(n2267), .B(n2268), .Z(o[62]) );
  AND U2271 ( .A(n1035), .B(n2269), .Z(n2267) );
  XNOR U2272 ( .A(creg[62]), .B(n2268), .Z(n2269) );
  XNOR U2273 ( .A(n2270), .B(n2271), .Z(o[629]) );
  AND U2274 ( .A(n1035), .B(n2272), .Z(n2270) );
  XNOR U2275 ( .A(creg[629]), .B(n2271), .Z(n2272) );
  XNOR U2276 ( .A(n2273), .B(n2274), .Z(o[628]) );
  AND U2277 ( .A(n1035), .B(n2275), .Z(n2273) );
  XNOR U2278 ( .A(creg[628]), .B(n2274), .Z(n2275) );
  XNOR U2279 ( .A(n2276), .B(n2277), .Z(o[627]) );
  AND U2280 ( .A(n1035), .B(n2278), .Z(n2276) );
  XNOR U2281 ( .A(creg[627]), .B(n2277), .Z(n2278) );
  XNOR U2282 ( .A(n2279), .B(n2280), .Z(o[626]) );
  AND U2283 ( .A(n1035), .B(n2281), .Z(n2279) );
  XNOR U2284 ( .A(creg[626]), .B(n2280), .Z(n2281) );
  XNOR U2285 ( .A(n2282), .B(n2283), .Z(o[625]) );
  AND U2286 ( .A(n1035), .B(n2284), .Z(n2282) );
  XNOR U2287 ( .A(creg[625]), .B(n2283), .Z(n2284) );
  XNOR U2288 ( .A(n2285), .B(n2286), .Z(o[624]) );
  AND U2289 ( .A(n1035), .B(n2287), .Z(n2285) );
  XNOR U2290 ( .A(creg[624]), .B(n2286), .Z(n2287) );
  XNOR U2291 ( .A(n2288), .B(n2289), .Z(o[623]) );
  AND U2292 ( .A(n1035), .B(n2290), .Z(n2288) );
  XNOR U2293 ( .A(creg[623]), .B(n2289), .Z(n2290) );
  XNOR U2294 ( .A(n2291), .B(n2292), .Z(o[622]) );
  AND U2295 ( .A(n1035), .B(n2293), .Z(n2291) );
  XNOR U2296 ( .A(creg[622]), .B(n2292), .Z(n2293) );
  XNOR U2297 ( .A(n2294), .B(n2295), .Z(o[621]) );
  AND U2298 ( .A(n1035), .B(n2296), .Z(n2294) );
  XNOR U2299 ( .A(creg[621]), .B(n2295), .Z(n2296) );
  XNOR U2300 ( .A(n2297), .B(n2298), .Z(o[620]) );
  AND U2301 ( .A(n1035), .B(n2299), .Z(n2297) );
  XNOR U2302 ( .A(creg[620]), .B(n2298), .Z(n2299) );
  XNOR U2303 ( .A(n2300), .B(n2301), .Z(o[61]) );
  AND U2304 ( .A(n1035), .B(n2302), .Z(n2300) );
  XNOR U2305 ( .A(creg[61]), .B(n2301), .Z(n2302) );
  XNOR U2306 ( .A(n2303), .B(n2304), .Z(o[619]) );
  AND U2307 ( .A(n1035), .B(n2305), .Z(n2303) );
  XNOR U2308 ( .A(creg[619]), .B(n2304), .Z(n2305) );
  XNOR U2309 ( .A(n2306), .B(n2307), .Z(o[618]) );
  AND U2310 ( .A(n1035), .B(n2308), .Z(n2306) );
  XNOR U2311 ( .A(creg[618]), .B(n2307), .Z(n2308) );
  XNOR U2312 ( .A(n2309), .B(n2310), .Z(o[617]) );
  AND U2313 ( .A(n1035), .B(n2311), .Z(n2309) );
  XNOR U2314 ( .A(creg[617]), .B(n2310), .Z(n2311) );
  XNOR U2315 ( .A(n2312), .B(n2313), .Z(o[616]) );
  AND U2316 ( .A(n1035), .B(n2314), .Z(n2312) );
  XNOR U2317 ( .A(creg[616]), .B(n2313), .Z(n2314) );
  XNOR U2318 ( .A(n2315), .B(n2316), .Z(o[615]) );
  AND U2319 ( .A(n1035), .B(n2317), .Z(n2315) );
  XNOR U2320 ( .A(creg[615]), .B(n2316), .Z(n2317) );
  XNOR U2321 ( .A(n2318), .B(n2319), .Z(o[614]) );
  AND U2322 ( .A(n1035), .B(n2320), .Z(n2318) );
  XNOR U2323 ( .A(creg[614]), .B(n2319), .Z(n2320) );
  XNOR U2324 ( .A(n2321), .B(n2322), .Z(o[613]) );
  AND U2325 ( .A(n1035), .B(n2323), .Z(n2321) );
  XNOR U2326 ( .A(creg[613]), .B(n2322), .Z(n2323) );
  XNOR U2327 ( .A(n2324), .B(n2325), .Z(o[612]) );
  AND U2328 ( .A(n1035), .B(n2326), .Z(n2324) );
  XNOR U2329 ( .A(creg[612]), .B(n2325), .Z(n2326) );
  XNOR U2330 ( .A(n2327), .B(n2328), .Z(o[611]) );
  AND U2331 ( .A(n1035), .B(n2329), .Z(n2327) );
  XNOR U2332 ( .A(creg[611]), .B(n2328), .Z(n2329) );
  XNOR U2333 ( .A(n2330), .B(n2331), .Z(o[610]) );
  AND U2334 ( .A(n1035), .B(n2332), .Z(n2330) );
  XNOR U2335 ( .A(creg[610]), .B(n2331), .Z(n2332) );
  XNOR U2336 ( .A(n2333), .B(n2334), .Z(o[60]) );
  AND U2337 ( .A(n1035), .B(n2335), .Z(n2333) );
  XNOR U2338 ( .A(creg[60]), .B(n2334), .Z(n2335) );
  XNOR U2339 ( .A(n2336), .B(n2337), .Z(o[609]) );
  AND U2340 ( .A(n1035), .B(n2338), .Z(n2336) );
  XNOR U2341 ( .A(creg[609]), .B(n2337), .Z(n2338) );
  XNOR U2342 ( .A(n2339), .B(n2340), .Z(o[608]) );
  AND U2343 ( .A(n1035), .B(n2341), .Z(n2339) );
  XNOR U2344 ( .A(creg[608]), .B(n2340), .Z(n2341) );
  XNOR U2345 ( .A(n2342), .B(n2343), .Z(o[607]) );
  AND U2346 ( .A(n1035), .B(n2344), .Z(n2342) );
  XNOR U2347 ( .A(creg[607]), .B(n2343), .Z(n2344) );
  XNOR U2348 ( .A(n2345), .B(n2346), .Z(o[606]) );
  AND U2349 ( .A(n1035), .B(n2347), .Z(n2345) );
  XNOR U2350 ( .A(creg[606]), .B(n2346), .Z(n2347) );
  XNOR U2351 ( .A(n2348), .B(n2349), .Z(o[605]) );
  AND U2352 ( .A(n1035), .B(n2350), .Z(n2348) );
  XNOR U2353 ( .A(creg[605]), .B(n2349), .Z(n2350) );
  XNOR U2354 ( .A(n2351), .B(n2352), .Z(o[604]) );
  AND U2355 ( .A(n1035), .B(n2353), .Z(n2351) );
  XNOR U2356 ( .A(creg[604]), .B(n2352), .Z(n2353) );
  XNOR U2357 ( .A(n2354), .B(n2355), .Z(o[603]) );
  AND U2358 ( .A(n1035), .B(n2356), .Z(n2354) );
  XNOR U2359 ( .A(creg[603]), .B(n2355), .Z(n2356) );
  XNOR U2360 ( .A(n2357), .B(n2358), .Z(o[602]) );
  AND U2361 ( .A(n1035), .B(n2359), .Z(n2357) );
  XNOR U2362 ( .A(creg[602]), .B(n2358), .Z(n2359) );
  XNOR U2363 ( .A(n2360), .B(n2361), .Z(o[601]) );
  AND U2364 ( .A(n1035), .B(n2362), .Z(n2360) );
  XNOR U2365 ( .A(creg[601]), .B(n2361), .Z(n2362) );
  XNOR U2366 ( .A(n2363), .B(n2364), .Z(o[600]) );
  AND U2367 ( .A(n1035), .B(n2365), .Z(n2363) );
  XNOR U2368 ( .A(creg[600]), .B(n2364), .Z(n2365) );
  XNOR U2369 ( .A(n2366), .B(n2367), .Z(o[5]) );
  AND U2370 ( .A(n1035), .B(n2368), .Z(n2366) );
  XNOR U2371 ( .A(creg[5]), .B(n2367), .Z(n2368) );
  XNOR U2372 ( .A(n2369), .B(n2370), .Z(o[59]) );
  AND U2373 ( .A(n1035), .B(n2371), .Z(n2369) );
  XNOR U2374 ( .A(creg[59]), .B(n2370), .Z(n2371) );
  XNOR U2375 ( .A(n2372), .B(n2373), .Z(o[599]) );
  AND U2376 ( .A(n1035), .B(n2374), .Z(n2372) );
  XNOR U2377 ( .A(creg[599]), .B(n2373), .Z(n2374) );
  XNOR U2378 ( .A(n2375), .B(n2376), .Z(o[598]) );
  AND U2379 ( .A(n1035), .B(n2377), .Z(n2375) );
  XNOR U2380 ( .A(creg[598]), .B(n2376), .Z(n2377) );
  XNOR U2381 ( .A(n2378), .B(n2379), .Z(o[597]) );
  AND U2382 ( .A(n1035), .B(n2380), .Z(n2378) );
  XNOR U2383 ( .A(creg[597]), .B(n2379), .Z(n2380) );
  XNOR U2384 ( .A(n2381), .B(n2382), .Z(o[596]) );
  AND U2385 ( .A(n1035), .B(n2383), .Z(n2381) );
  XNOR U2386 ( .A(creg[596]), .B(n2382), .Z(n2383) );
  XNOR U2387 ( .A(n2384), .B(n2385), .Z(o[595]) );
  AND U2388 ( .A(n1035), .B(n2386), .Z(n2384) );
  XNOR U2389 ( .A(creg[595]), .B(n2385), .Z(n2386) );
  XNOR U2390 ( .A(n2387), .B(n2388), .Z(o[594]) );
  AND U2391 ( .A(n1035), .B(n2389), .Z(n2387) );
  XNOR U2392 ( .A(creg[594]), .B(n2388), .Z(n2389) );
  XNOR U2393 ( .A(n2390), .B(n2391), .Z(o[593]) );
  AND U2394 ( .A(n1035), .B(n2392), .Z(n2390) );
  XNOR U2395 ( .A(creg[593]), .B(n2391), .Z(n2392) );
  XNOR U2396 ( .A(n2393), .B(n2394), .Z(o[592]) );
  AND U2397 ( .A(n1035), .B(n2395), .Z(n2393) );
  XNOR U2398 ( .A(creg[592]), .B(n2394), .Z(n2395) );
  XNOR U2399 ( .A(n2396), .B(n2397), .Z(o[591]) );
  AND U2400 ( .A(n1035), .B(n2398), .Z(n2396) );
  XNOR U2401 ( .A(creg[591]), .B(n2397), .Z(n2398) );
  XNOR U2402 ( .A(n2399), .B(n2400), .Z(o[590]) );
  AND U2403 ( .A(n1035), .B(n2401), .Z(n2399) );
  XNOR U2404 ( .A(creg[590]), .B(n2400), .Z(n2401) );
  XNOR U2405 ( .A(n2402), .B(n2403), .Z(o[58]) );
  AND U2406 ( .A(n1035), .B(n2404), .Z(n2402) );
  XNOR U2407 ( .A(creg[58]), .B(n2403), .Z(n2404) );
  XNOR U2408 ( .A(n2405), .B(n2406), .Z(o[589]) );
  AND U2409 ( .A(n1035), .B(n2407), .Z(n2405) );
  XNOR U2410 ( .A(creg[589]), .B(n2406), .Z(n2407) );
  XNOR U2411 ( .A(n2408), .B(n2409), .Z(o[588]) );
  AND U2412 ( .A(n1035), .B(n2410), .Z(n2408) );
  XNOR U2413 ( .A(creg[588]), .B(n2409), .Z(n2410) );
  XNOR U2414 ( .A(n2411), .B(n2412), .Z(o[587]) );
  AND U2415 ( .A(n1035), .B(n2413), .Z(n2411) );
  XNOR U2416 ( .A(creg[587]), .B(n2412), .Z(n2413) );
  XNOR U2417 ( .A(n2414), .B(n2415), .Z(o[586]) );
  AND U2418 ( .A(n1035), .B(n2416), .Z(n2414) );
  XNOR U2419 ( .A(creg[586]), .B(n2415), .Z(n2416) );
  XNOR U2420 ( .A(n2417), .B(n2418), .Z(o[585]) );
  AND U2421 ( .A(n1035), .B(n2419), .Z(n2417) );
  XNOR U2422 ( .A(creg[585]), .B(n2418), .Z(n2419) );
  XNOR U2423 ( .A(n2420), .B(n2421), .Z(o[584]) );
  AND U2424 ( .A(n1035), .B(n2422), .Z(n2420) );
  XNOR U2425 ( .A(creg[584]), .B(n2421), .Z(n2422) );
  XNOR U2426 ( .A(n2423), .B(n2424), .Z(o[583]) );
  AND U2427 ( .A(n1035), .B(n2425), .Z(n2423) );
  XNOR U2428 ( .A(creg[583]), .B(n2424), .Z(n2425) );
  XNOR U2429 ( .A(n2426), .B(n2427), .Z(o[582]) );
  AND U2430 ( .A(n1035), .B(n2428), .Z(n2426) );
  XNOR U2431 ( .A(creg[582]), .B(n2427), .Z(n2428) );
  XNOR U2432 ( .A(n2429), .B(n2430), .Z(o[581]) );
  AND U2433 ( .A(n1035), .B(n2431), .Z(n2429) );
  XNOR U2434 ( .A(creg[581]), .B(n2430), .Z(n2431) );
  XNOR U2435 ( .A(n2432), .B(n2433), .Z(o[580]) );
  AND U2436 ( .A(n1035), .B(n2434), .Z(n2432) );
  XNOR U2437 ( .A(creg[580]), .B(n2433), .Z(n2434) );
  XNOR U2438 ( .A(n2435), .B(n2436), .Z(o[57]) );
  AND U2439 ( .A(n1035), .B(n2437), .Z(n2435) );
  XNOR U2440 ( .A(creg[57]), .B(n2436), .Z(n2437) );
  XNOR U2441 ( .A(n2438), .B(n2439), .Z(o[579]) );
  AND U2442 ( .A(n1035), .B(n2440), .Z(n2438) );
  XNOR U2443 ( .A(creg[579]), .B(n2439), .Z(n2440) );
  XNOR U2444 ( .A(n2441), .B(n2442), .Z(o[578]) );
  AND U2445 ( .A(n1035), .B(n2443), .Z(n2441) );
  XNOR U2446 ( .A(creg[578]), .B(n2442), .Z(n2443) );
  XNOR U2447 ( .A(n2444), .B(n2445), .Z(o[577]) );
  AND U2448 ( .A(n1035), .B(n2446), .Z(n2444) );
  XNOR U2449 ( .A(creg[577]), .B(n2445), .Z(n2446) );
  XNOR U2450 ( .A(n2447), .B(n2448), .Z(o[576]) );
  AND U2451 ( .A(n1035), .B(n2449), .Z(n2447) );
  XNOR U2452 ( .A(creg[576]), .B(n2448), .Z(n2449) );
  XNOR U2453 ( .A(n2450), .B(n2451), .Z(o[575]) );
  AND U2454 ( .A(n1035), .B(n2452), .Z(n2450) );
  XNOR U2455 ( .A(creg[575]), .B(n2451), .Z(n2452) );
  XNOR U2456 ( .A(n2453), .B(n2454), .Z(o[574]) );
  AND U2457 ( .A(n1035), .B(n2455), .Z(n2453) );
  XNOR U2458 ( .A(creg[574]), .B(n2454), .Z(n2455) );
  XNOR U2459 ( .A(n2456), .B(n2457), .Z(o[573]) );
  AND U2460 ( .A(n1035), .B(n2458), .Z(n2456) );
  XNOR U2461 ( .A(creg[573]), .B(n2457), .Z(n2458) );
  XNOR U2462 ( .A(n2459), .B(n2460), .Z(o[572]) );
  AND U2463 ( .A(n1035), .B(n2461), .Z(n2459) );
  XNOR U2464 ( .A(creg[572]), .B(n2460), .Z(n2461) );
  XNOR U2465 ( .A(n2462), .B(n2463), .Z(o[571]) );
  AND U2466 ( .A(n1035), .B(n2464), .Z(n2462) );
  XNOR U2467 ( .A(creg[571]), .B(n2463), .Z(n2464) );
  XNOR U2468 ( .A(n2465), .B(n2466), .Z(o[570]) );
  AND U2469 ( .A(n1035), .B(n2467), .Z(n2465) );
  XNOR U2470 ( .A(creg[570]), .B(n2466), .Z(n2467) );
  XNOR U2471 ( .A(n2468), .B(n2469), .Z(o[56]) );
  AND U2472 ( .A(n1035), .B(n2470), .Z(n2468) );
  XNOR U2473 ( .A(creg[56]), .B(n2469), .Z(n2470) );
  XNOR U2474 ( .A(n2471), .B(n2472), .Z(o[569]) );
  AND U2475 ( .A(n1035), .B(n2473), .Z(n2471) );
  XNOR U2476 ( .A(creg[569]), .B(n2472), .Z(n2473) );
  XNOR U2477 ( .A(n2474), .B(n2475), .Z(o[568]) );
  AND U2478 ( .A(n1035), .B(n2476), .Z(n2474) );
  XNOR U2479 ( .A(creg[568]), .B(n2475), .Z(n2476) );
  XNOR U2480 ( .A(n2477), .B(n2478), .Z(o[567]) );
  AND U2481 ( .A(n1035), .B(n2479), .Z(n2477) );
  XNOR U2482 ( .A(creg[567]), .B(n2478), .Z(n2479) );
  XNOR U2483 ( .A(n2480), .B(n2481), .Z(o[566]) );
  AND U2484 ( .A(n1035), .B(n2482), .Z(n2480) );
  XNOR U2485 ( .A(creg[566]), .B(n2481), .Z(n2482) );
  XNOR U2486 ( .A(n2483), .B(n2484), .Z(o[565]) );
  AND U2487 ( .A(n1035), .B(n2485), .Z(n2483) );
  XNOR U2488 ( .A(creg[565]), .B(n2484), .Z(n2485) );
  XNOR U2489 ( .A(n2486), .B(n2487), .Z(o[564]) );
  AND U2490 ( .A(n1035), .B(n2488), .Z(n2486) );
  XNOR U2491 ( .A(creg[564]), .B(n2487), .Z(n2488) );
  XNOR U2492 ( .A(n2489), .B(n2490), .Z(o[563]) );
  AND U2493 ( .A(n1035), .B(n2491), .Z(n2489) );
  XNOR U2494 ( .A(creg[563]), .B(n2490), .Z(n2491) );
  XNOR U2495 ( .A(n2492), .B(n2493), .Z(o[562]) );
  AND U2496 ( .A(n1035), .B(n2494), .Z(n2492) );
  XNOR U2497 ( .A(creg[562]), .B(n2493), .Z(n2494) );
  XNOR U2498 ( .A(n2495), .B(n2496), .Z(o[561]) );
  AND U2499 ( .A(n1035), .B(n2497), .Z(n2495) );
  XNOR U2500 ( .A(creg[561]), .B(n2496), .Z(n2497) );
  XNOR U2501 ( .A(n2498), .B(n2499), .Z(o[560]) );
  AND U2502 ( .A(n1035), .B(n2500), .Z(n2498) );
  XNOR U2503 ( .A(creg[560]), .B(n2499), .Z(n2500) );
  XNOR U2504 ( .A(n2501), .B(n2502), .Z(o[55]) );
  AND U2505 ( .A(n1035), .B(n2503), .Z(n2501) );
  XNOR U2506 ( .A(creg[55]), .B(n2502), .Z(n2503) );
  XNOR U2507 ( .A(n2504), .B(n2505), .Z(o[559]) );
  AND U2508 ( .A(n1035), .B(n2506), .Z(n2504) );
  XNOR U2509 ( .A(creg[559]), .B(n2505), .Z(n2506) );
  XNOR U2510 ( .A(n2507), .B(n2508), .Z(o[558]) );
  AND U2511 ( .A(n1035), .B(n2509), .Z(n2507) );
  XNOR U2512 ( .A(creg[558]), .B(n2508), .Z(n2509) );
  XNOR U2513 ( .A(n2510), .B(n2511), .Z(o[557]) );
  AND U2514 ( .A(n1035), .B(n2512), .Z(n2510) );
  XNOR U2515 ( .A(creg[557]), .B(n2511), .Z(n2512) );
  XNOR U2516 ( .A(n2513), .B(n2514), .Z(o[556]) );
  AND U2517 ( .A(n1035), .B(n2515), .Z(n2513) );
  XNOR U2518 ( .A(creg[556]), .B(n2514), .Z(n2515) );
  XNOR U2519 ( .A(n2516), .B(n2517), .Z(o[555]) );
  AND U2520 ( .A(n1035), .B(n2518), .Z(n2516) );
  XNOR U2521 ( .A(creg[555]), .B(n2517), .Z(n2518) );
  XNOR U2522 ( .A(n2519), .B(n2520), .Z(o[554]) );
  AND U2523 ( .A(n1035), .B(n2521), .Z(n2519) );
  XNOR U2524 ( .A(creg[554]), .B(n2520), .Z(n2521) );
  XNOR U2525 ( .A(n2522), .B(n2523), .Z(o[553]) );
  AND U2526 ( .A(n1035), .B(n2524), .Z(n2522) );
  XNOR U2527 ( .A(creg[553]), .B(n2523), .Z(n2524) );
  XNOR U2528 ( .A(n2525), .B(n2526), .Z(o[552]) );
  AND U2529 ( .A(n1035), .B(n2527), .Z(n2525) );
  XNOR U2530 ( .A(creg[552]), .B(n2526), .Z(n2527) );
  XNOR U2531 ( .A(n2528), .B(n2529), .Z(o[551]) );
  AND U2532 ( .A(n1035), .B(n2530), .Z(n2528) );
  XNOR U2533 ( .A(creg[551]), .B(n2529), .Z(n2530) );
  XNOR U2534 ( .A(n2531), .B(n2532), .Z(o[550]) );
  AND U2535 ( .A(n1035), .B(n2533), .Z(n2531) );
  XNOR U2536 ( .A(creg[550]), .B(n2532), .Z(n2533) );
  XNOR U2537 ( .A(n2534), .B(n2535), .Z(o[54]) );
  AND U2538 ( .A(n1035), .B(n2536), .Z(n2534) );
  XNOR U2539 ( .A(creg[54]), .B(n2535), .Z(n2536) );
  XNOR U2540 ( .A(n2537), .B(n2538), .Z(o[549]) );
  AND U2541 ( .A(n1035), .B(n2539), .Z(n2537) );
  XNOR U2542 ( .A(creg[549]), .B(n2538), .Z(n2539) );
  XNOR U2543 ( .A(n2540), .B(n2541), .Z(o[548]) );
  AND U2544 ( .A(n1035), .B(n2542), .Z(n2540) );
  XNOR U2545 ( .A(creg[548]), .B(n2541), .Z(n2542) );
  XNOR U2546 ( .A(n2543), .B(n2544), .Z(o[547]) );
  AND U2547 ( .A(n1035), .B(n2545), .Z(n2543) );
  XNOR U2548 ( .A(creg[547]), .B(n2544), .Z(n2545) );
  XNOR U2549 ( .A(n2546), .B(n2547), .Z(o[546]) );
  AND U2550 ( .A(n1035), .B(n2548), .Z(n2546) );
  XNOR U2551 ( .A(creg[546]), .B(n2547), .Z(n2548) );
  XNOR U2552 ( .A(n2549), .B(n2550), .Z(o[545]) );
  AND U2553 ( .A(n1035), .B(n2551), .Z(n2549) );
  XNOR U2554 ( .A(creg[545]), .B(n2550), .Z(n2551) );
  XNOR U2555 ( .A(n2552), .B(n2553), .Z(o[544]) );
  AND U2556 ( .A(n1035), .B(n2554), .Z(n2552) );
  XNOR U2557 ( .A(creg[544]), .B(n2553), .Z(n2554) );
  XNOR U2558 ( .A(n2555), .B(n2556), .Z(o[543]) );
  AND U2559 ( .A(n1035), .B(n2557), .Z(n2555) );
  XNOR U2560 ( .A(creg[543]), .B(n2556), .Z(n2557) );
  XNOR U2561 ( .A(n2558), .B(n2559), .Z(o[542]) );
  AND U2562 ( .A(n1035), .B(n2560), .Z(n2558) );
  XNOR U2563 ( .A(creg[542]), .B(n2559), .Z(n2560) );
  XNOR U2564 ( .A(n2561), .B(n2562), .Z(o[541]) );
  AND U2565 ( .A(n1035), .B(n2563), .Z(n2561) );
  XNOR U2566 ( .A(creg[541]), .B(n2562), .Z(n2563) );
  XNOR U2567 ( .A(n2564), .B(n2565), .Z(o[540]) );
  AND U2568 ( .A(n1035), .B(n2566), .Z(n2564) );
  XNOR U2569 ( .A(creg[540]), .B(n2565), .Z(n2566) );
  XNOR U2570 ( .A(n2567), .B(n2568), .Z(o[53]) );
  AND U2571 ( .A(n1035), .B(n2569), .Z(n2567) );
  XNOR U2572 ( .A(creg[53]), .B(n2568), .Z(n2569) );
  XNOR U2573 ( .A(n2570), .B(n2571), .Z(o[539]) );
  AND U2574 ( .A(n1035), .B(n2572), .Z(n2570) );
  XNOR U2575 ( .A(creg[539]), .B(n2571), .Z(n2572) );
  XNOR U2576 ( .A(n2573), .B(n2574), .Z(o[538]) );
  AND U2577 ( .A(n1035), .B(n2575), .Z(n2573) );
  XNOR U2578 ( .A(creg[538]), .B(n2574), .Z(n2575) );
  XNOR U2579 ( .A(n2576), .B(n2577), .Z(o[537]) );
  AND U2580 ( .A(n1035), .B(n2578), .Z(n2576) );
  XNOR U2581 ( .A(creg[537]), .B(n2577), .Z(n2578) );
  XNOR U2582 ( .A(n2579), .B(n2580), .Z(o[536]) );
  AND U2583 ( .A(n1035), .B(n2581), .Z(n2579) );
  XNOR U2584 ( .A(creg[536]), .B(n2580), .Z(n2581) );
  XNOR U2585 ( .A(n2582), .B(n2583), .Z(o[535]) );
  AND U2586 ( .A(n1035), .B(n2584), .Z(n2582) );
  XNOR U2587 ( .A(creg[535]), .B(n2583), .Z(n2584) );
  XNOR U2588 ( .A(n2585), .B(n2586), .Z(o[534]) );
  AND U2589 ( .A(n1035), .B(n2587), .Z(n2585) );
  XNOR U2590 ( .A(creg[534]), .B(n2586), .Z(n2587) );
  XNOR U2591 ( .A(n2588), .B(n2589), .Z(o[533]) );
  AND U2592 ( .A(n1035), .B(n2590), .Z(n2588) );
  XNOR U2593 ( .A(creg[533]), .B(n2589), .Z(n2590) );
  XNOR U2594 ( .A(n2591), .B(n2592), .Z(o[532]) );
  AND U2595 ( .A(n1035), .B(n2593), .Z(n2591) );
  XNOR U2596 ( .A(creg[532]), .B(n2592), .Z(n2593) );
  XNOR U2597 ( .A(n2594), .B(n2595), .Z(o[531]) );
  AND U2598 ( .A(n1035), .B(n2596), .Z(n2594) );
  XNOR U2599 ( .A(creg[531]), .B(n2595), .Z(n2596) );
  XNOR U2600 ( .A(n2597), .B(n2598), .Z(o[530]) );
  AND U2601 ( .A(n1035), .B(n2599), .Z(n2597) );
  XNOR U2602 ( .A(creg[530]), .B(n2598), .Z(n2599) );
  XNOR U2603 ( .A(n2600), .B(n2601), .Z(o[52]) );
  AND U2604 ( .A(n1035), .B(n2602), .Z(n2600) );
  XNOR U2605 ( .A(creg[52]), .B(n2601), .Z(n2602) );
  XNOR U2606 ( .A(n2603), .B(n2604), .Z(o[529]) );
  AND U2607 ( .A(n1035), .B(n2605), .Z(n2603) );
  XNOR U2608 ( .A(creg[529]), .B(n2604), .Z(n2605) );
  XNOR U2609 ( .A(n2606), .B(n2607), .Z(o[528]) );
  AND U2610 ( .A(n1035), .B(n2608), .Z(n2606) );
  XNOR U2611 ( .A(creg[528]), .B(n2607), .Z(n2608) );
  XNOR U2612 ( .A(n2609), .B(n2610), .Z(o[527]) );
  AND U2613 ( .A(n1035), .B(n2611), .Z(n2609) );
  XNOR U2614 ( .A(creg[527]), .B(n2610), .Z(n2611) );
  XNOR U2615 ( .A(n2612), .B(n2613), .Z(o[526]) );
  AND U2616 ( .A(n1035), .B(n2614), .Z(n2612) );
  XNOR U2617 ( .A(creg[526]), .B(n2613), .Z(n2614) );
  XNOR U2618 ( .A(n2615), .B(n2616), .Z(o[525]) );
  AND U2619 ( .A(n1035), .B(n2617), .Z(n2615) );
  XNOR U2620 ( .A(creg[525]), .B(n2616), .Z(n2617) );
  XNOR U2621 ( .A(n2618), .B(n2619), .Z(o[524]) );
  AND U2622 ( .A(n1035), .B(n2620), .Z(n2618) );
  XNOR U2623 ( .A(creg[524]), .B(n2619), .Z(n2620) );
  XNOR U2624 ( .A(n2621), .B(n2622), .Z(o[523]) );
  AND U2625 ( .A(n1035), .B(n2623), .Z(n2621) );
  XNOR U2626 ( .A(creg[523]), .B(n2622), .Z(n2623) );
  XNOR U2627 ( .A(n2624), .B(n2625), .Z(o[522]) );
  AND U2628 ( .A(n1035), .B(n2626), .Z(n2624) );
  XNOR U2629 ( .A(creg[522]), .B(n2625), .Z(n2626) );
  XNOR U2630 ( .A(n2627), .B(n2628), .Z(o[521]) );
  AND U2631 ( .A(n1035), .B(n2629), .Z(n2627) );
  XNOR U2632 ( .A(creg[521]), .B(n2628), .Z(n2629) );
  XNOR U2633 ( .A(n2630), .B(n2631), .Z(o[520]) );
  AND U2634 ( .A(n1035), .B(n2632), .Z(n2630) );
  XNOR U2635 ( .A(creg[520]), .B(n2631), .Z(n2632) );
  XNOR U2636 ( .A(n2633), .B(n2634), .Z(o[51]) );
  AND U2637 ( .A(n1035), .B(n2635), .Z(n2633) );
  XNOR U2638 ( .A(creg[51]), .B(n2634), .Z(n2635) );
  XNOR U2639 ( .A(n2636), .B(n2637), .Z(o[519]) );
  AND U2640 ( .A(n1035), .B(n2638), .Z(n2636) );
  XNOR U2641 ( .A(creg[519]), .B(n2637), .Z(n2638) );
  XNOR U2642 ( .A(n2639), .B(n2640), .Z(o[518]) );
  AND U2643 ( .A(n1035), .B(n2641), .Z(n2639) );
  XNOR U2644 ( .A(creg[518]), .B(n2640), .Z(n2641) );
  XNOR U2645 ( .A(n2642), .B(n2643), .Z(o[517]) );
  AND U2646 ( .A(n1035), .B(n2644), .Z(n2642) );
  XNOR U2647 ( .A(creg[517]), .B(n2643), .Z(n2644) );
  XNOR U2648 ( .A(n2645), .B(n2646), .Z(o[516]) );
  AND U2649 ( .A(n1035), .B(n2647), .Z(n2645) );
  XNOR U2650 ( .A(creg[516]), .B(n2646), .Z(n2647) );
  XNOR U2651 ( .A(n2648), .B(n2649), .Z(o[515]) );
  AND U2652 ( .A(n1035), .B(n2650), .Z(n2648) );
  XNOR U2653 ( .A(creg[515]), .B(n2649), .Z(n2650) );
  XNOR U2654 ( .A(n2651), .B(n2652), .Z(o[514]) );
  AND U2655 ( .A(n1035), .B(n2653), .Z(n2651) );
  XNOR U2656 ( .A(creg[514]), .B(n2652), .Z(n2653) );
  XNOR U2657 ( .A(n2654), .B(n2655), .Z(o[513]) );
  AND U2658 ( .A(n1035), .B(n2656), .Z(n2654) );
  XNOR U2659 ( .A(creg[513]), .B(n2655), .Z(n2656) );
  XNOR U2660 ( .A(n2657), .B(n2658), .Z(o[512]) );
  AND U2661 ( .A(n1035), .B(n2659), .Z(n2657) );
  XNOR U2662 ( .A(creg[512]), .B(n2658), .Z(n2659) );
  XNOR U2663 ( .A(n2660), .B(n2661), .Z(o[511]) );
  AND U2664 ( .A(n1035), .B(n2662), .Z(n2660) );
  XNOR U2665 ( .A(creg[511]), .B(n2661), .Z(n2662) );
  XNOR U2666 ( .A(n2663), .B(n2664), .Z(o[510]) );
  AND U2667 ( .A(n1035), .B(n2665), .Z(n2663) );
  XNOR U2668 ( .A(creg[510]), .B(n2664), .Z(n2665) );
  XNOR U2669 ( .A(n2666), .B(n2667), .Z(o[50]) );
  AND U2670 ( .A(n1035), .B(n2668), .Z(n2666) );
  XNOR U2671 ( .A(creg[50]), .B(n2667), .Z(n2668) );
  XNOR U2672 ( .A(n2669), .B(n2670), .Z(o[509]) );
  AND U2673 ( .A(n1035), .B(n2671), .Z(n2669) );
  XNOR U2674 ( .A(creg[509]), .B(n2670), .Z(n2671) );
  XNOR U2675 ( .A(n2672), .B(n2673), .Z(o[508]) );
  AND U2676 ( .A(n1035), .B(n2674), .Z(n2672) );
  XNOR U2677 ( .A(creg[508]), .B(n2673), .Z(n2674) );
  XNOR U2678 ( .A(n2675), .B(n2676), .Z(o[507]) );
  AND U2679 ( .A(n1035), .B(n2677), .Z(n2675) );
  XNOR U2680 ( .A(creg[507]), .B(n2676), .Z(n2677) );
  XNOR U2681 ( .A(n2678), .B(n2679), .Z(o[506]) );
  AND U2682 ( .A(n1035), .B(n2680), .Z(n2678) );
  XNOR U2683 ( .A(creg[506]), .B(n2679), .Z(n2680) );
  XNOR U2684 ( .A(n2681), .B(n2682), .Z(o[505]) );
  AND U2685 ( .A(n1035), .B(n2683), .Z(n2681) );
  XNOR U2686 ( .A(creg[505]), .B(n2682), .Z(n2683) );
  XNOR U2687 ( .A(n2684), .B(n2685), .Z(o[504]) );
  AND U2688 ( .A(n1035), .B(n2686), .Z(n2684) );
  XNOR U2689 ( .A(creg[504]), .B(n2685), .Z(n2686) );
  XNOR U2690 ( .A(n2687), .B(n2688), .Z(o[503]) );
  AND U2691 ( .A(n1035), .B(n2689), .Z(n2687) );
  XNOR U2692 ( .A(creg[503]), .B(n2688), .Z(n2689) );
  XNOR U2693 ( .A(n2690), .B(n2691), .Z(o[502]) );
  AND U2694 ( .A(n1035), .B(n2692), .Z(n2690) );
  XNOR U2695 ( .A(creg[502]), .B(n2691), .Z(n2692) );
  XNOR U2696 ( .A(n2693), .B(n2694), .Z(o[501]) );
  AND U2697 ( .A(n1035), .B(n2695), .Z(n2693) );
  XNOR U2698 ( .A(creg[501]), .B(n2694), .Z(n2695) );
  XNOR U2699 ( .A(n2696), .B(n2697), .Z(o[500]) );
  AND U2700 ( .A(n1035), .B(n2698), .Z(n2696) );
  XNOR U2701 ( .A(creg[500]), .B(n2697), .Z(n2698) );
  XNOR U2702 ( .A(n2699), .B(n2700), .Z(o[4]) );
  AND U2703 ( .A(n1035), .B(n2701), .Z(n2699) );
  XNOR U2704 ( .A(creg[4]), .B(n2700), .Z(n2701) );
  XNOR U2705 ( .A(n2702), .B(n2703), .Z(o[49]) );
  AND U2706 ( .A(n1035), .B(n2704), .Z(n2702) );
  XNOR U2707 ( .A(creg[49]), .B(n2703), .Z(n2704) );
  XNOR U2708 ( .A(n2705), .B(n2706), .Z(o[499]) );
  AND U2709 ( .A(n1035), .B(n2707), .Z(n2705) );
  XNOR U2710 ( .A(creg[499]), .B(n2706), .Z(n2707) );
  XNOR U2711 ( .A(n2708), .B(n2709), .Z(o[498]) );
  AND U2712 ( .A(n1035), .B(n2710), .Z(n2708) );
  XNOR U2713 ( .A(creg[498]), .B(n2709), .Z(n2710) );
  XNOR U2714 ( .A(n2711), .B(n2712), .Z(o[497]) );
  AND U2715 ( .A(n1035), .B(n2713), .Z(n2711) );
  XNOR U2716 ( .A(creg[497]), .B(n2712), .Z(n2713) );
  XNOR U2717 ( .A(n2714), .B(n2715), .Z(o[496]) );
  AND U2718 ( .A(n1035), .B(n2716), .Z(n2714) );
  XNOR U2719 ( .A(creg[496]), .B(n2715), .Z(n2716) );
  XNOR U2720 ( .A(n2717), .B(n2718), .Z(o[495]) );
  AND U2721 ( .A(n1035), .B(n2719), .Z(n2717) );
  XNOR U2722 ( .A(creg[495]), .B(n2718), .Z(n2719) );
  XNOR U2723 ( .A(n2720), .B(n2721), .Z(o[494]) );
  AND U2724 ( .A(n1035), .B(n2722), .Z(n2720) );
  XNOR U2725 ( .A(creg[494]), .B(n2721), .Z(n2722) );
  XNOR U2726 ( .A(n2723), .B(n2724), .Z(o[493]) );
  AND U2727 ( .A(n1035), .B(n2725), .Z(n2723) );
  XNOR U2728 ( .A(creg[493]), .B(n2724), .Z(n2725) );
  XNOR U2729 ( .A(n2726), .B(n2727), .Z(o[492]) );
  AND U2730 ( .A(n1035), .B(n2728), .Z(n2726) );
  XNOR U2731 ( .A(creg[492]), .B(n2727), .Z(n2728) );
  XNOR U2732 ( .A(n2729), .B(n2730), .Z(o[491]) );
  AND U2733 ( .A(n1035), .B(n2731), .Z(n2729) );
  XNOR U2734 ( .A(creg[491]), .B(n2730), .Z(n2731) );
  XNOR U2735 ( .A(n2732), .B(n2733), .Z(o[490]) );
  AND U2736 ( .A(n1035), .B(n2734), .Z(n2732) );
  XNOR U2737 ( .A(creg[490]), .B(n2733), .Z(n2734) );
  XNOR U2738 ( .A(n2735), .B(n2736), .Z(o[48]) );
  AND U2739 ( .A(n1035), .B(n2737), .Z(n2735) );
  XNOR U2740 ( .A(creg[48]), .B(n2736), .Z(n2737) );
  XNOR U2741 ( .A(n2738), .B(n2739), .Z(o[489]) );
  AND U2742 ( .A(n1035), .B(n2740), .Z(n2738) );
  XNOR U2743 ( .A(creg[489]), .B(n2739), .Z(n2740) );
  XNOR U2744 ( .A(n2741), .B(n2742), .Z(o[488]) );
  AND U2745 ( .A(n1035), .B(n2743), .Z(n2741) );
  XNOR U2746 ( .A(creg[488]), .B(n2742), .Z(n2743) );
  XNOR U2747 ( .A(n2744), .B(n2745), .Z(o[487]) );
  AND U2748 ( .A(n1035), .B(n2746), .Z(n2744) );
  XNOR U2749 ( .A(creg[487]), .B(n2745), .Z(n2746) );
  XNOR U2750 ( .A(n2747), .B(n2748), .Z(o[486]) );
  AND U2751 ( .A(n1035), .B(n2749), .Z(n2747) );
  XNOR U2752 ( .A(creg[486]), .B(n2748), .Z(n2749) );
  XNOR U2753 ( .A(n2750), .B(n2751), .Z(o[485]) );
  AND U2754 ( .A(n1035), .B(n2752), .Z(n2750) );
  XNOR U2755 ( .A(creg[485]), .B(n2751), .Z(n2752) );
  XNOR U2756 ( .A(n2753), .B(n2754), .Z(o[484]) );
  AND U2757 ( .A(n1035), .B(n2755), .Z(n2753) );
  XNOR U2758 ( .A(creg[484]), .B(n2754), .Z(n2755) );
  XNOR U2759 ( .A(n2756), .B(n2757), .Z(o[483]) );
  AND U2760 ( .A(n1035), .B(n2758), .Z(n2756) );
  XNOR U2761 ( .A(creg[483]), .B(n2757), .Z(n2758) );
  XNOR U2762 ( .A(n2759), .B(n2760), .Z(o[482]) );
  AND U2763 ( .A(n1035), .B(n2761), .Z(n2759) );
  XNOR U2764 ( .A(creg[482]), .B(n2760), .Z(n2761) );
  XNOR U2765 ( .A(n2762), .B(n2763), .Z(o[481]) );
  AND U2766 ( .A(n1035), .B(n2764), .Z(n2762) );
  XNOR U2767 ( .A(creg[481]), .B(n2763), .Z(n2764) );
  XNOR U2768 ( .A(n2765), .B(n2766), .Z(o[480]) );
  AND U2769 ( .A(n1035), .B(n2767), .Z(n2765) );
  XNOR U2770 ( .A(creg[480]), .B(n2766), .Z(n2767) );
  XNOR U2771 ( .A(n2768), .B(n2769), .Z(o[47]) );
  AND U2772 ( .A(n1035), .B(n2770), .Z(n2768) );
  XNOR U2773 ( .A(creg[47]), .B(n2769), .Z(n2770) );
  XNOR U2774 ( .A(n2771), .B(n2772), .Z(o[479]) );
  AND U2775 ( .A(n1035), .B(n2773), .Z(n2771) );
  XNOR U2776 ( .A(creg[479]), .B(n2772), .Z(n2773) );
  XNOR U2777 ( .A(n2774), .B(n2775), .Z(o[478]) );
  AND U2778 ( .A(n1035), .B(n2776), .Z(n2774) );
  XNOR U2779 ( .A(creg[478]), .B(n2775), .Z(n2776) );
  XNOR U2780 ( .A(n2777), .B(n2778), .Z(o[477]) );
  AND U2781 ( .A(n1035), .B(n2779), .Z(n2777) );
  XNOR U2782 ( .A(creg[477]), .B(n2778), .Z(n2779) );
  XNOR U2783 ( .A(n2780), .B(n2781), .Z(o[476]) );
  AND U2784 ( .A(n1035), .B(n2782), .Z(n2780) );
  XNOR U2785 ( .A(creg[476]), .B(n2781), .Z(n2782) );
  XNOR U2786 ( .A(n2783), .B(n2784), .Z(o[475]) );
  AND U2787 ( .A(n1035), .B(n2785), .Z(n2783) );
  XNOR U2788 ( .A(creg[475]), .B(n2784), .Z(n2785) );
  XNOR U2789 ( .A(n2786), .B(n2787), .Z(o[474]) );
  AND U2790 ( .A(n1035), .B(n2788), .Z(n2786) );
  XNOR U2791 ( .A(creg[474]), .B(n2787), .Z(n2788) );
  XNOR U2792 ( .A(n2789), .B(n2790), .Z(o[473]) );
  AND U2793 ( .A(n1035), .B(n2791), .Z(n2789) );
  XNOR U2794 ( .A(creg[473]), .B(n2790), .Z(n2791) );
  XNOR U2795 ( .A(n2792), .B(n2793), .Z(o[472]) );
  AND U2796 ( .A(n1035), .B(n2794), .Z(n2792) );
  XNOR U2797 ( .A(creg[472]), .B(n2793), .Z(n2794) );
  XNOR U2798 ( .A(n2795), .B(n2796), .Z(o[471]) );
  AND U2799 ( .A(n1035), .B(n2797), .Z(n2795) );
  XNOR U2800 ( .A(creg[471]), .B(n2796), .Z(n2797) );
  XNOR U2801 ( .A(n2798), .B(n2799), .Z(o[470]) );
  AND U2802 ( .A(n1035), .B(n2800), .Z(n2798) );
  XNOR U2803 ( .A(creg[470]), .B(n2799), .Z(n2800) );
  XNOR U2804 ( .A(n2801), .B(n2802), .Z(o[46]) );
  AND U2805 ( .A(n1035), .B(n2803), .Z(n2801) );
  XNOR U2806 ( .A(creg[46]), .B(n2802), .Z(n2803) );
  XNOR U2807 ( .A(n2804), .B(n2805), .Z(o[469]) );
  AND U2808 ( .A(n1035), .B(n2806), .Z(n2804) );
  XNOR U2809 ( .A(creg[469]), .B(n2805), .Z(n2806) );
  XNOR U2810 ( .A(n2807), .B(n2808), .Z(o[468]) );
  AND U2811 ( .A(n1035), .B(n2809), .Z(n2807) );
  XNOR U2812 ( .A(creg[468]), .B(n2808), .Z(n2809) );
  XNOR U2813 ( .A(n2810), .B(n2811), .Z(o[467]) );
  AND U2814 ( .A(n1035), .B(n2812), .Z(n2810) );
  XNOR U2815 ( .A(creg[467]), .B(n2811), .Z(n2812) );
  XNOR U2816 ( .A(n2813), .B(n2814), .Z(o[466]) );
  AND U2817 ( .A(n1035), .B(n2815), .Z(n2813) );
  XNOR U2818 ( .A(creg[466]), .B(n2814), .Z(n2815) );
  XNOR U2819 ( .A(n2816), .B(n2817), .Z(o[465]) );
  AND U2820 ( .A(n1035), .B(n2818), .Z(n2816) );
  XNOR U2821 ( .A(creg[465]), .B(n2817), .Z(n2818) );
  XNOR U2822 ( .A(n2819), .B(n2820), .Z(o[464]) );
  AND U2823 ( .A(n1035), .B(n2821), .Z(n2819) );
  XNOR U2824 ( .A(creg[464]), .B(n2820), .Z(n2821) );
  XNOR U2825 ( .A(n2822), .B(n2823), .Z(o[463]) );
  AND U2826 ( .A(n1035), .B(n2824), .Z(n2822) );
  XNOR U2827 ( .A(creg[463]), .B(n2823), .Z(n2824) );
  XNOR U2828 ( .A(n2825), .B(n2826), .Z(o[462]) );
  AND U2829 ( .A(n1035), .B(n2827), .Z(n2825) );
  XNOR U2830 ( .A(creg[462]), .B(n2826), .Z(n2827) );
  XNOR U2831 ( .A(n2828), .B(n2829), .Z(o[461]) );
  AND U2832 ( .A(n1035), .B(n2830), .Z(n2828) );
  XNOR U2833 ( .A(creg[461]), .B(n2829), .Z(n2830) );
  XNOR U2834 ( .A(n2831), .B(n2832), .Z(o[460]) );
  AND U2835 ( .A(n1035), .B(n2833), .Z(n2831) );
  XNOR U2836 ( .A(creg[460]), .B(n2832), .Z(n2833) );
  XNOR U2837 ( .A(n2834), .B(n2835), .Z(o[45]) );
  AND U2838 ( .A(n1035), .B(n2836), .Z(n2834) );
  XNOR U2839 ( .A(creg[45]), .B(n2835), .Z(n2836) );
  XNOR U2840 ( .A(n2837), .B(n2838), .Z(o[459]) );
  AND U2841 ( .A(n1035), .B(n2839), .Z(n2837) );
  XNOR U2842 ( .A(creg[459]), .B(n2838), .Z(n2839) );
  XNOR U2843 ( .A(n2840), .B(n2841), .Z(o[458]) );
  AND U2844 ( .A(n1035), .B(n2842), .Z(n2840) );
  XNOR U2845 ( .A(creg[458]), .B(n2841), .Z(n2842) );
  XNOR U2846 ( .A(n2843), .B(n2844), .Z(o[457]) );
  AND U2847 ( .A(n1035), .B(n2845), .Z(n2843) );
  XNOR U2848 ( .A(creg[457]), .B(n2844), .Z(n2845) );
  XNOR U2849 ( .A(n2846), .B(n2847), .Z(o[456]) );
  AND U2850 ( .A(n1035), .B(n2848), .Z(n2846) );
  XNOR U2851 ( .A(creg[456]), .B(n2847), .Z(n2848) );
  XNOR U2852 ( .A(n2849), .B(n2850), .Z(o[455]) );
  AND U2853 ( .A(n1035), .B(n2851), .Z(n2849) );
  XNOR U2854 ( .A(creg[455]), .B(n2850), .Z(n2851) );
  XNOR U2855 ( .A(n2852), .B(n2853), .Z(o[454]) );
  AND U2856 ( .A(n1035), .B(n2854), .Z(n2852) );
  XNOR U2857 ( .A(creg[454]), .B(n2853), .Z(n2854) );
  XNOR U2858 ( .A(n2855), .B(n2856), .Z(o[453]) );
  AND U2859 ( .A(n1035), .B(n2857), .Z(n2855) );
  XNOR U2860 ( .A(creg[453]), .B(n2856), .Z(n2857) );
  XNOR U2861 ( .A(n2858), .B(n2859), .Z(o[452]) );
  AND U2862 ( .A(n1035), .B(n2860), .Z(n2858) );
  XNOR U2863 ( .A(creg[452]), .B(n2859), .Z(n2860) );
  XNOR U2864 ( .A(n2861), .B(n2862), .Z(o[451]) );
  AND U2865 ( .A(n1035), .B(n2863), .Z(n2861) );
  XNOR U2866 ( .A(creg[451]), .B(n2862), .Z(n2863) );
  XNOR U2867 ( .A(n2864), .B(n2865), .Z(o[450]) );
  AND U2868 ( .A(n1035), .B(n2866), .Z(n2864) );
  XNOR U2869 ( .A(creg[450]), .B(n2865), .Z(n2866) );
  XNOR U2870 ( .A(n2867), .B(n2868), .Z(o[44]) );
  AND U2871 ( .A(n1035), .B(n2869), .Z(n2867) );
  XNOR U2872 ( .A(creg[44]), .B(n2868), .Z(n2869) );
  XNOR U2873 ( .A(n2870), .B(n2871), .Z(o[449]) );
  AND U2874 ( .A(n1035), .B(n2872), .Z(n2870) );
  XNOR U2875 ( .A(creg[449]), .B(n2871), .Z(n2872) );
  XNOR U2876 ( .A(n2873), .B(n2874), .Z(o[448]) );
  AND U2877 ( .A(n1035), .B(n2875), .Z(n2873) );
  XNOR U2878 ( .A(creg[448]), .B(n2874), .Z(n2875) );
  XNOR U2879 ( .A(n2876), .B(n2877), .Z(o[447]) );
  AND U2880 ( .A(n1035), .B(n2878), .Z(n2876) );
  XNOR U2881 ( .A(creg[447]), .B(n2877), .Z(n2878) );
  XNOR U2882 ( .A(n2879), .B(n2880), .Z(o[446]) );
  AND U2883 ( .A(n1035), .B(n2881), .Z(n2879) );
  XNOR U2884 ( .A(creg[446]), .B(n2880), .Z(n2881) );
  XNOR U2885 ( .A(n2882), .B(n2883), .Z(o[445]) );
  AND U2886 ( .A(n1035), .B(n2884), .Z(n2882) );
  XNOR U2887 ( .A(creg[445]), .B(n2883), .Z(n2884) );
  XNOR U2888 ( .A(n2885), .B(n2886), .Z(o[444]) );
  AND U2889 ( .A(n1035), .B(n2887), .Z(n2885) );
  XNOR U2890 ( .A(creg[444]), .B(n2886), .Z(n2887) );
  XNOR U2891 ( .A(n2888), .B(n2889), .Z(o[443]) );
  AND U2892 ( .A(n1035), .B(n2890), .Z(n2888) );
  XNOR U2893 ( .A(creg[443]), .B(n2889), .Z(n2890) );
  XNOR U2894 ( .A(n2891), .B(n2892), .Z(o[442]) );
  AND U2895 ( .A(n1035), .B(n2893), .Z(n2891) );
  XNOR U2896 ( .A(creg[442]), .B(n2892), .Z(n2893) );
  XNOR U2897 ( .A(n2894), .B(n2895), .Z(o[441]) );
  AND U2898 ( .A(n1035), .B(n2896), .Z(n2894) );
  XNOR U2899 ( .A(creg[441]), .B(n2895), .Z(n2896) );
  XNOR U2900 ( .A(n2897), .B(n2898), .Z(o[440]) );
  AND U2901 ( .A(n1035), .B(n2899), .Z(n2897) );
  XNOR U2902 ( .A(creg[440]), .B(n2898), .Z(n2899) );
  XNOR U2903 ( .A(n2900), .B(n2901), .Z(o[43]) );
  AND U2904 ( .A(n1035), .B(n2902), .Z(n2900) );
  XNOR U2905 ( .A(creg[43]), .B(n2901), .Z(n2902) );
  XNOR U2906 ( .A(n2903), .B(n2904), .Z(o[439]) );
  AND U2907 ( .A(n1035), .B(n2905), .Z(n2903) );
  XNOR U2908 ( .A(creg[439]), .B(n2904), .Z(n2905) );
  XNOR U2909 ( .A(n2906), .B(n2907), .Z(o[438]) );
  AND U2910 ( .A(n1035), .B(n2908), .Z(n2906) );
  XNOR U2911 ( .A(creg[438]), .B(n2907), .Z(n2908) );
  XNOR U2912 ( .A(n2909), .B(n2910), .Z(o[437]) );
  AND U2913 ( .A(n1035), .B(n2911), .Z(n2909) );
  XNOR U2914 ( .A(creg[437]), .B(n2910), .Z(n2911) );
  XNOR U2915 ( .A(n2912), .B(n2913), .Z(o[436]) );
  AND U2916 ( .A(n1035), .B(n2914), .Z(n2912) );
  XNOR U2917 ( .A(creg[436]), .B(n2913), .Z(n2914) );
  XNOR U2918 ( .A(n2915), .B(n2916), .Z(o[435]) );
  AND U2919 ( .A(n1035), .B(n2917), .Z(n2915) );
  XNOR U2920 ( .A(creg[435]), .B(n2916), .Z(n2917) );
  XNOR U2921 ( .A(n2918), .B(n2919), .Z(o[434]) );
  AND U2922 ( .A(n1035), .B(n2920), .Z(n2918) );
  XNOR U2923 ( .A(creg[434]), .B(n2919), .Z(n2920) );
  XNOR U2924 ( .A(n2921), .B(n2922), .Z(o[433]) );
  AND U2925 ( .A(n1035), .B(n2923), .Z(n2921) );
  XNOR U2926 ( .A(creg[433]), .B(n2922), .Z(n2923) );
  XNOR U2927 ( .A(n2924), .B(n2925), .Z(o[432]) );
  AND U2928 ( .A(n1035), .B(n2926), .Z(n2924) );
  XNOR U2929 ( .A(creg[432]), .B(n2925), .Z(n2926) );
  XNOR U2930 ( .A(n2927), .B(n2928), .Z(o[431]) );
  AND U2931 ( .A(n1035), .B(n2929), .Z(n2927) );
  XNOR U2932 ( .A(creg[431]), .B(n2928), .Z(n2929) );
  XNOR U2933 ( .A(n2930), .B(n2931), .Z(o[430]) );
  AND U2934 ( .A(n1035), .B(n2932), .Z(n2930) );
  XNOR U2935 ( .A(creg[430]), .B(n2931), .Z(n2932) );
  XNOR U2936 ( .A(n2933), .B(n2934), .Z(o[42]) );
  AND U2937 ( .A(n1035), .B(n2935), .Z(n2933) );
  XNOR U2938 ( .A(creg[42]), .B(n2934), .Z(n2935) );
  XNOR U2939 ( .A(n2936), .B(n2937), .Z(o[429]) );
  AND U2940 ( .A(n1035), .B(n2938), .Z(n2936) );
  XNOR U2941 ( .A(creg[429]), .B(n2937), .Z(n2938) );
  XNOR U2942 ( .A(n2939), .B(n2940), .Z(o[428]) );
  AND U2943 ( .A(n1035), .B(n2941), .Z(n2939) );
  XNOR U2944 ( .A(creg[428]), .B(n2940), .Z(n2941) );
  XNOR U2945 ( .A(n2942), .B(n2943), .Z(o[427]) );
  AND U2946 ( .A(n1035), .B(n2944), .Z(n2942) );
  XNOR U2947 ( .A(creg[427]), .B(n2943), .Z(n2944) );
  XNOR U2948 ( .A(n2945), .B(n2946), .Z(o[426]) );
  AND U2949 ( .A(n1035), .B(n2947), .Z(n2945) );
  XNOR U2950 ( .A(creg[426]), .B(n2946), .Z(n2947) );
  XNOR U2951 ( .A(n2948), .B(n2949), .Z(o[425]) );
  AND U2952 ( .A(n1035), .B(n2950), .Z(n2948) );
  XNOR U2953 ( .A(creg[425]), .B(n2949), .Z(n2950) );
  XNOR U2954 ( .A(n2951), .B(n2952), .Z(o[424]) );
  AND U2955 ( .A(n1035), .B(n2953), .Z(n2951) );
  XNOR U2956 ( .A(creg[424]), .B(n2952), .Z(n2953) );
  XNOR U2957 ( .A(n2954), .B(n2955), .Z(o[423]) );
  AND U2958 ( .A(n1035), .B(n2956), .Z(n2954) );
  XNOR U2959 ( .A(creg[423]), .B(n2955), .Z(n2956) );
  XNOR U2960 ( .A(n2957), .B(n2958), .Z(o[422]) );
  AND U2961 ( .A(n1035), .B(n2959), .Z(n2957) );
  XNOR U2962 ( .A(creg[422]), .B(n2958), .Z(n2959) );
  XNOR U2963 ( .A(n2960), .B(n2961), .Z(o[421]) );
  AND U2964 ( .A(n1035), .B(n2962), .Z(n2960) );
  XNOR U2965 ( .A(creg[421]), .B(n2961), .Z(n2962) );
  XNOR U2966 ( .A(n2963), .B(n2964), .Z(o[420]) );
  AND U2967 ( .A(n1035), .B(n2965), .Z(n2963) );
  XNOR U2968 ( .A(creg[420]), .B(n2964), .Z(n2965) );
  XNOR U2969 ( .A(n2966), .B(n2967), .Z(o[41]) );
  AND U2970 ( .A(n1035), .B(n2968), .Z(n2966) );
  XNOR U2971 ( .A(creg[41]), .B(n2967), .Z(n2968) );
  XNOR U2972 ( .A(n2969), .B(n2970), .Z(o[419]) );
  AND U2973 ( .A(n1035), .B(n2971), .Z(n2969) );
  XNOR U2974 ( .A(creg[419]), .B(n2970), .Z(n2971) );
  XNOR U2975 ( .A(n2972), .B(n2973), .Z(o[418]) );
  AND U2976 ( .A(n1035), .B(n2974), .Z(n2972) );
  XNOR U2977 ( .A(creg[418]), .B(n2973), .Z(n2974) );
  XNOR U2978 ( .A(n2975), .B(n2976), .Z(o[417]) );
  AND U2979 ( .A(n1035), .B(n2977), .Z(n2975) );
  XNOR U2980 ( .A(creg[417]), .B(n2976), .Z(n2977) );
  XNOR U2981 ( .A(n2978), .B(n2979), .Z(o[416]) );
  AND U2982 ( .A(n1035), .B(n2980), .Z(n2978) );
  XNOR U2983 ( .A(creg[416]), .B(n2979), .Z(n2980) );
  XNOR U2984 ( .A(n2981), .B(n2982), .Z(o[415]) );
  AND U2985 ( .A(n1035), .B(n2983), .Z(n2981) );
  XNOR U2986 ( .A(creg[415]), .B(n2982), .Z(n2983) );
  XNOR U2987 ( .A(n2984), .B(n2985), .Z(o[414]) );
  AND U2988 ( .A(n1035), .B(n2986), .Z(n2984) );
  XNOR U2989 ( .A(creg[414]), .B(n2985), .Z(n2986) );
  XNOR U2990 ( .A(n2987), .B(n2988), .Z(o[413]) );
  AND U2991 ( .A(n1035), .B(n2989), .Z(n2987) );
  XNOR U2992 ( .A(creg[413]), .B(n2988), .Z(n2989) );
  XNOR U2993 ( .A(n2990), .B(n2991), .Z(o[412]) );
  AND U2994 ( .A(n1035), .B(n2992), .Z(n2990) );
  XNOR U2995 ( .A(creg[412]), .B(n2991), .Z(n2992) );
  XNOR U2996 ( .A(n2993), .B(n2994), .Z(o[411]) );
  AND U2997 ( .A(n1035), .B(n2995), .Z(n2993) );
  XNOR U2998 ( .A(creg[411]), .B(n2994), .Z(n2995) );
  XNOR U2999 ( .A(n2996), .B(n2997), .Z(o[410]) );
  AND U3000 ( .A(n1035), .B(n2998), .Z(n2996) );
  XNOR U3001 ( .A(creg[410]), .B(n2997), .Z(n2998) );
  XNOR U3002 ( .A(n2999), .B(n3000), .Z(o[40]) );
  AND U3003 ( .A(n1035), .B(n3001), .Z(n2999) );
  XNOR U3004 ( .A(creg[40]), .B(n3000), .Z(n3001) );
  XNOR U3005 ( .A(n3002), .B(n3003), .Z(o[409]) );
  AND U3006 ( .A(n1035), .B(n3004), .Z(n3002) );
  XNOR U3007 ( .A(creg[409]), .B(n3003), .Z(n3004) );
  XNOR U3008 ( .A(n3005), .B(n3006), .Z(o[408]) );
  AND U3009 ( .A(n1035), .B(n3007), .Z(n3005) );
  XNOR U3010 ( .A(creg[408]), .B(n3006), .Z(n3007) );
  XNOR U3011 ( .A(n3008), .B(n3009), .Z(o[407]) );
  AND U3012 ( .A(n1035), .B(n3010), .Z(n3008) );
  XNOR U3013 ( .A(creg[407]), .B(n3009), .Z(n3010) );
  XNOR U3014 ( .A(n3011), .B(n3012), .Z(o[406]) );
  AND U3015 ( .A(n1035), .B(n3013), .Z(n3011) );
  XNOR U3016 ( .A(creg[406]), .B(n3012), .Z(n3013) );
  XNOR U3017 ( .A(n3014), .B(n3015), .Z(o[405]) );
  AND U3018 ( .A(n1035), .B(n3016), .Z(n3014) );
  XNOR U3019 ( .A(creg[405]), .B(n3015), .Z(n3016) );
  XNOR U3020 ( .A(n3017), .B(n3018), .Z(o[404]) );
  AND U3021 ( .A(n1035), .B(n3019), .Z(n3017) );
  XNOR U3022 ( .A(creg[404]), .B(n3018), .Z(n3019) );
  XNOR U3023 ( .A(n3020), .B(n3021), .Z(o[403]) );
  AND U3024 ( .A(n1035), .B(n3022), .Z(n3020) );
  XNOR U3025 ( .A(creg[403]), .B(n3021), .Z(n3022) );
  XNOR U3026 ( .A(n3023), .B(n3024), .Z(o[402]) );
  AND U3027 ( .A(n1035), .B(n3025), .Z(n3023) );
  XNOR U3028 ( .A(creg[402]), .B(n3024), .Z(n3025) );
  XNOR U3029 ( .A(n3026), .B(n3027), .Z(o[401]) );
  AND U3030 ( .A(n1035), .B(n3028), .Z(n3026) );
  XNOR U3031 ( .A(creg[401]), .B(n3027), .Z(n3028) );
  XNOR U3032 ( .A(n3029), .B(n3030), .Z(o[400]) );
  AND U3033 ( .A(n1035), .B(n3031), .Z(n3029) );
  XNOR U3034 ( .A(creg[400]), .B(n3030), .Z(n3031) );
  XNOR U3035 ( .A(n3032), .B(n3033), .Z(o[3]) );
  AND U3036 ( .A(n1035), .B(n3034), .Z(n3032) );
  XNOR U3037 ( .A(creg[3]), .B(n3033), .Z(n3034) );
  XNOR U3038 ( .A(n3035), .B(n3036), .Z(o[39]) );
  AND U3039 ( .A(n1035), .B(n3037), .Z(n3035) );
  XNOR U3040 ( .A(creg[39]), .B(n3036), .Z(n3037) );
  XNOR U3041 ( .A(n3038), .B(n3039), .Z(o[399]) );
  AND U3042 ( .A(n1035), .B(n3040), .Z(n3038) );
  XNOR U3043 ( .A(creg[399]), .B(n3039), .Z(n3040) );
  XNOR U3044 ( .A(n3041), .B(n3042), .Z(o[398]) );
  AND U3045 ( .A(n1035), .B(n3043), .Z(n3041) );
  XNOR U3046 ( .A(creg[398]), .B(n3042), .Z(n3043) );
  XNOR U3047 ( .A(n3044), .B(n3045), .Z(o[397]) );
  AND U3048 ( .A(n1035), .B(n3046), .Z(n3044) );
  XNOR U3049 ( .A(creg[397]), .B(n3045), .Z(n3046) );
  XNOR U3050 ( .A(n3047), .B(n3048), .Z(o[396]) );
  AND U3051 ( .A(n1035), .B(n3049), .Z(n3047) );
  XNOR U3052 ( .A(creg[396]), .B(n3048), .Z(n3049) );
  XNOR U3053 ( .A(n3050), .B(n3051), .Z(o[395]) );
  AND U3054 ( .A(n1035), .B(n3052), .Z(n3050) );
  XNOR U3055 ( .A(creg[395]), .B(n3051), .Z(n3052) );
  XNOR U3056 ( .A(n3053), .B(n3054), .Z(o[394]) );
  AND U3057 ( .A(n1035), .B(n3055), .Z(n3053) );
  XNOR U3058 ( .A(creg[394]), .B(n3054), .Z(n3055) );
  XNOR U3059 ( .A(n3056), .B(n3057), .Z(o[393]) );
  AND U3060 ( .A(n1035), .B(n3058), .Z(n3056) );
  XNOR U3061 ( .A(creg[393]), .B(n3057), .Z(n3058) );
  XNOR U3062 ( .A(n3059), .B(n3060), .Z(o[392]) );
  AND U3063 ( .A(n1035), .B(n3061), .Z(n3059) );
  XNOR U3064 ( .A(creg[392]), .B(n3060), .Z(n3061) );
  XNOR U3065 ( .A(n3062), .B(n3063), .Z(o[391]) );
  AND U3066 ( .A(n1035), .B(n3064), .Z(n3062) );
  XNOR U3067 ( .A(creg[391]), .B(n3063), .Z(n3064) );
  XNOR U3068 ( .A(n3065), .B(n3066), .Z(o[390]) );
  AND U3069 ( .A(n1035), .B(n3067), .Z(n3065) );
  XNOR U3070 ( .A(creg[390]), .B(n3066), .Z(n3067) );
  XNOR U3071 ( .A(n3068), .B(n3069), .Z(o[38]) );
  AND U3072 ( .A(n1035), .B(n3070), .Z(n3068) );
  XNOR U3073 ( .A(creg[38]), .B(n3069), .Z(n3070) );
  XNOR U3074 ( .A(n3071), .B(n3072), .Z(o[389]) );
  AND U3075 ( .A(n1035), .B(n3073), .Z(n3071) );
  XNOR U3076 ( .A(creg[389]), .B(n3072), .Z(n3073) );
  XNOR U3077 ( .A(n3074), .B(n3075), .Z(o[388]) );
  AND U3078 ( .A(n1035), .B(n3076), .Z(n3074) );
  XNOR U3079 ( .A(creg[388]), .B(n3075), .Z(n3076) );
  XNOR U3080 ( .A(n3077), .B(n3078), .Z(o[387]) );
  AND U3081 ( .A(n1035), .B(n3079), .Z(n3077) );
  XNOR U3082 ( .A(creg[387]), .B(n3078), .Z(n3079) );
  XNOR U3083 ( .A(n3080), .B(n3081), .Z(o[386]) );
  AND U3084 ( .A(n1035), .B(n3082), .Z(n3080) );
  XNOR U3085 ( .A(creg[386]), .B(n3081), .Z(n3082) );
  XNOR U3086 ( .A(n3083), .B(n3084), .Z(o[385]) );
  AND U3087 ( .A(n1035), .B(n3085), .Z(n3083) );
  XNOR U3088 ( .A(creg[385]), .B(n3084), .Z(n3085) );
  XNOR U3089 ( .A(n3086), .B(n3087), .Z(o[384]) );
  AND U3090 ( .A(n1035), .B(n3088), .Z(n3086) );
  XNOR U3091 ( .A(creg[384]), .B(n3087), .Z(n3088) );
  XNOR U3092 ( .A(n3089), .B(n3090), .Z(o[383]) );
  AND U3093 ( .A(n1035), .B(n3091), .Z(n3089) );
  XNOR U3094 ( .A(creg[383]), .B(n3090), .Z(n3091) );
  XNOR U3095 ( .A(n3092), .B(n3093), .Z(o[382]) );
  AND U3096 ( .A(n1035), .B(n3094), .Z(n3092) );
  XNOR U3097 ( .A(creg[382]), .B(n3093), .Z(n3094) );
  XNOR U3098 ( .A(n3095), .B(n3096), .Z(o[381]) );
  AND U3099 ( .A(n1035), .B(n3097), .Z(n3095) );
  XNOR U3100 ( .A(creg[381]), .B(n3096), .Z(n3097) );
  XNOR U3101 ( .A(n3098), .B(n3099), .Z(o[380]) );
  AND U3102 ( .A(n1035), .B(n3100), .Z(n3098) );
  XNOR U3103 ( .A(creg[380]), .B(n3099), .Z(n3100) );
  XNOR U3104 ( .A(n3101), .B(n3102), .Z(o[37]) );
  AND U3105 ( .A(n1035), .B(n3103), .Z(n3101) );
  XNOR U3106 ( .A(creg[37]), .B(n3102), .Z(n3103) );
  XNOR U3107 ( .A(n3104), .B(n3105), .Z(o[379]) );
  AND U3108 ( .A(n1035), .B(n3106), .Z(n3104) );
  XNOR U3109 ( .A(creg[379]), .B(n3105), .Z(n3106) );
  XNOR U3110 ( .A(n3107), .B(n3108), .Z(o[378]) );
  AND U3111 ( .A(n1035), .B(n3109), .Z(n3107) );
  XNOR U3112 ( .A(creg[378]), .B(n3108), .Z(n3109) );
  XNOR U3113 ( .A(n3110), .B(n3111), .Z(o[377]) );
  AND U3114 ( .A(n1035), .B(n3112), .Z(n3110) );
  XNOR U3115 ( .A(creg[377]), .B(n3111), .Z(n3112) );
  XNOR U3116 ( .A(n3113), .B(n3114), .Z(o[376]) );
  AND U3117 ( .A(n1035), .B(n3115), .Z(n3113) );
  XNOR U3118 ( .A(creg[376]), .B(n3114), .Z(n3115) );
  XNOR U3119 ( .A(n3116), .B(n3117), .Z(o[375]) );
  AND U3120 ( .A(n1035), .B(n3118), .Z(n3116) );
  XNOR U3121 ( .A(creg[375]), .B(n3117), .Z(n3118) );
  XNOR U3122 ( .A(n3119), .B(n3120), .Z(o[374]) );
  AND U3123 ( .A(n1035), .B(n3121), .Z(n3119) );
  XNOR U3124 ( .A(creg[374]), .B(n3120), .Z(n3121) );
  XNOR U3125 ( .A(n3122), .B(n3123), .Z(o[373]) );
  AND U3126 ( .A(n1035), .B(n3124), .Z(n3122) );
  XNOR U3127 ( .A(creg[373]), .B(n3123), .Z(n3124) );
  XNOR U3128 ( .A(n3125), .B(n3126), .Z(o[372]) );
  AND U3129 ( .A(n1035), .B(n3127), .Z(n3125) );
  XNOR U3130 ( .A(creg[372]), .B(n3126), .Z(n3127) );
  XNOR U3131 ( .A(n3128), .B(n3129), .Z(o[371]) );
  AND U3132 ( .A(n1035), .B(n3130), .Z(n3128) );
  XNOR U3133 ( .A(creg[371]), .B(n3129), .Z(n3130) );
  XNOR U3134 ( .A(n3131), .B(n3132), .Z(o[370]) );
  AND U3135 ( .A(n1035), .B(n3133), .Z(n3131) );
  XNOR U3136 ( .A(creg[370]), .B(n3132), .Z(n3133) );
  XNOR U3137 ( .A(n3134), .B(n3135), .Z(o[36]) );
  AND U3138 ( .A(n1035), .B(n3136), .Z(n3134) );
  XNOR U3139 ( .A(creg[36]), .B(n3135), .Z(n3136) );
  XNOR U3140 ( .A(n3137), .B(n3138), .Z(o[369]) );
  AND U3141 ( .A(n1035), .B(n3139), .Z(n3137) );
  XNOR U3142 ( .A(creg[369]), .B(n3138), .Z(n3139) );
  XNOR U3143 ( .A(n3140), .B(n3141), .Z(o[368]) );
  AND U3144 ( .A(n1035), .B(n3142), .Z(n3140) );
  XNOR U3145 ( .A(creg[368]), .B(n3141), .Z(n3142) );
  XNOR U3146 ( .A(n3143), .B(n3144), .Z(o[367]) );
  AND U3147 ( .A(n1035), .B(n3145), .Z(n3143) );
  XNOR U3148 ( .A(creg[367]), .B(n3144), .Z(n3145) );
  XNOR U3149 ( .A(n3146), .B(n3147), .Z(o[366]) );
  AND U3150 ( .A(n1035), .B(n3148), .Z(n3146) );
  XNOR U3151 ( .A(creg[366]), .B(n3147), .Z(n3148) );
  XNOR U3152 ( .A(n3149), .B(n3150), .Z(o[365]) );
  AND U3153 ( .A(n1035), .B(n3151), .Z(n3149) );
  XNOR U3154 ( .A(creg[365]), .B(n3150), .Z(n3151) );
  XNOR U3155 ( .A(n3152), .B(n3153), .Z(o[364]) );
  AND U3156 ( .A(n1035), .B(n3154), .Z(n3152) );
  XNOR U3157 ( .A(creg[364]), .B(n3153), .Z(n3154) );
  XNOR U3158 ( .A(n3155), .B(n3156), .Z(o[363]) );
  AND U3159 ( .A(n1035), .B(n3157), .Z(n3155) );
  XNOR U3160 ( .A(creg[363]), .B(n3156), .Z(n3157) );
  XNOR U3161 ( .A(n3158), .B(n3159), .Z(o[362]) );
  AND U3162 ( .A(n1035), .B(n3160), .Z(n3158) );
  XNOR U3163 ( .A(creg[362]), .B(n3159), .Z(n3160) );
  XNOR U3164 ( .A(n3161), .B(n3162), .Z(o[361]) );
  AND U3165 ( .A(n1035), .B(n3163), .Z(n3161) );
  XNOR U3166 ( .A(creg[361]), .B(n3162), .Z(n3163) );
  XNOR U3167 ( .A(n3164), .B(n3165), .Z(o[360]) );
  AND U3168 ( .A(n1035), .B(n3166), .Z(n3164) );
  XNOR U3169 ( .A(creg[360]), .B(n3165), .Z(n3166) );
  XNOR U3170 ( .A(n3167), .B(n3168), .Z(o[35]) );
  AND U3171 ( .A(n1035), .B(n3169), .Z(n3167) );
  XNOR U3172 ( .A(creg[35]), .B(n3168), .Z(n3169) );
  XNOR U3173 ( .A(n3170), .B(n3171), .Z(o[359]) );
  AND U3174 ( .A(n1035), .B(n3172), .Z(n3170) );
  XNOR U3175 ( .A(creg[359]), .B(n3171), .Z(n3172) );
  XNOR U3176 ( .A(n3173), .B(n3174), .Z(o[358]) );
  AND U3177 ( .A(n1035), .B(n3175), .Z(n3173) );
  XNOR U3178 ( .A(creg[358]), .B(n3174), .Z(n3175) );
  XNOR U3179 ( .A(n3176), .B(n3177), .Z(o[357]) );
  AND U3180 ( .A(n1035), .B(n3178), .Z(n3176) );
  XNOR U3181 ( .A(creg[357]), .B(n3177), .Z(n3178) );
  XNOR U3182 ( .A(n3179), .B(n3180), .Z(o[356]) );
  AND U3183 ( .A(n1035), .B(n3181), .Z(n3179) );
  XNOR U3184 ( .A(creg[356]), .B(n3180), .Z(n3181) );
  XNOR U3185 ( .A(n3182), .B(n3183), .Z(o[355]) );
  AND U3186 ( .A(n1035), .B(n3184), .Z(n3182) );
  XNOR U3187 ( .A(creg[355]), .B(n3183), .Z(n3184) );
  XNOR U3188 ( .A(n3185), .B(n3186), .Z(o[354]) );
  AND U3189 ( .A(n1035), .B(n3187), .Z(n3185) );
  XNOR U3190 ( .A(creg[354]), .B(n3186), .Z(n3187) );
  XNOR U3191 ( .A(n3188), .B(n3189), .Z(o[353]) );
  AND U3192 ( .A(n1035), .B(n3190), .Z(n3188) );
  XNOR U3193 ( .A(creg[353]), .B(n3189), .Z(n3190) );
  XNOR U3194 ( .A(n3191), .B(n3192), .Z(o[352]) );
  AND U3195 ( .A(n1035), .B(n3193), .Z(n3191) );
  XNOR U3196 ( .A(creg[352]), .B(n3192), .Z(n3193) );
  XNOR U3197 ( .A(n3194), .B(n3195), .Z(o[351]) );
  AND U3198 ( .A(n1035), .B(n3196), .Z(n3194) );
  XNOR U3199 ( .A(creg[351]), .B(n3195), .Z(n3196) );
  XNOR U3200 ( .A(n3197), .B(n3198), .Z(o[350]) );
  AND U3201 ( .A(n1035), .B(n3199), .Z(n3197) );
  XNOR U3202 ( .A(creg[350]), .B(n3198), .Z(n3199) );
  XNOR U3203 ( .A(n3200), .B(n3201), .Z(o[34]) );
  AND U3204 ( .A(n1035), .B(n3202), .Z(n3200) );
  XNOR U3205 ( .A(creg[34]), .B(n3201), .Z(n3202) );
  XNOR U3206 ( .A(n3203), .B(n3204), .Z(o[349]) );
  AND U3207 ( .A(n1035), .B(n3205), .Z(n3203) );
  XNOR U3208 ( .A(creg[349]), .B(n3204), .Z(n3205) );
  XNOR U3209 ( .A(n3206), .B(n3207), .Z(o[348]) );
  AND U3210 ( .A(n1035), .B(n3208), .Z(n3206) );
  XNOR U3211 ( .A(creg[348]), .B(n3207), .Z(n3208) );
  XNOR U3212 ( .A(n3209), .B(n3210), .Z(o[347]) );
  AND U3213 ( .A(n1035), .B(n3211), .Z(n3209) );
  XNOR U3214 ( .A(creg[347]), .B(n3210), .Z(n3211) );
  XNOR U3215 ( .A(n3212), .B(n3213), .Z(o[346]) );
  AND U3216 ( .A(n1035), .B(n3214), .Z(n3212) );
  XNOR U3217 ( .A(creg[346]), .B(n3213), .Z(n3214) );
  XNOR U3218 ( .A(n3215), .B(n3216), .Z(o[345]) );
  AND U3219 ( .A(n1035), .B(n3217), .Z(n3215) );
  XNOR U3220 ( .A(creg[345]), .B(n3216), .Z(n3217) );
  XNOR U3221 ( .A(n3218), .B(n3219), .Z(o[344]) );
  AND U3222 ( .A(n1035), .B(n3220), .Z(n3218) );
  XNOR U3223 ( .A(creg[344]), .B(n3219), .Z(n3220) );
  XNOR U3224 ( .A(n3221), .B(n3222), .Z(o[343]) );
  AND U3225 ( .A(n1035), .B(n3223), .Z(n3221) );
  XNOR U3226 ( .A(creg[343]), .B(n3222), .Z(n3223) );
  XNOR U3227 ( .A(n3224), .B(n3225), .Z(o[342]) );
  AND U3228 ( .A(n1035), .B(n3226), .Z(n3224) );
  XNOR U3229 ( .A(creg[342]), .B(n3225), .Z(n3226) );
  XNOR U3230 ( .A(n3227), .B(n3228), .Z(o[341]) );
  AND U3231 ( .A(n1035), .B(n3229), .Z(n3227) );
  XNOR U3232 ( .A(creg[341]), .B(n3228), .Z(n3229) );
  XNOR U3233 ( .A(n3230), .B(n3231), .Z(o[340]) );
  AND U3234 ( .A(n1035), .B(n3232), .Z(n3230) );
  XNOR U3235 ( .A(creg[340]), .B(n3231), .Z(n3232) );
  XNOR U3236 ( .A(n3233), .B(n3234), .Z(o[33]) );
  AND U3237 ( .A(n1035), .B(n3235), .Z(n3233) );
  XNOR U3238 ( .A(creg[33]), .B(n3234), .Z(n3235) );
  XNOR U3239 ( .A(n3236), .B(n3237), .Z(o[339]) );
  AND U3240 ( .A(n1035), .B(n3238), .Z(n3236) );
  XNOR U3241 ( .A(creg[339]), .B(n3237), .Z(n3238) );
  XNOR U3242 ( .A(n3239), .B(n3240), .Z(o[338]) );
  AND U3243 ( .A(n1035), .B(n3241), .Z(n3239) );
  XNOR U3244 ( .A(creg[338]), .B(n3240), .Z(n3241) );
  XNOR U3245 ( .A(n3242), .B(n3243), .Z(o[337]) );
  AND U3246 ( .A(n1035), .B(n3244), .Z(n3242) );
  XNOR U3247 ( .A(creg[337]), .B(n3243), .Z(n3244) );
  XNOR U3248 ( .A(n3245), .B(n3246), .Z(o[336]) );
  AND U3249 ( .A(n1035), .B(n3247), .Z(n3245) );
  XNOR U3250 ( .A(creg[336]), .B(n3246), .Z(n3247) );
  XNOR U3251 ( .A(n3248), .B(n3249), .Z(o[335]) );
  AND U3252 ( .A(n1035), .B(n3250), .Z(n3248) );
  XNOR U3253 ( .A(creg[335]), .B(n3249), .Z(n3250) );
  XNOR U3254 ( .A(n3251), .B(n3252), .Z(o[334]) );
  AND U3255 ( .A(n1035), .B(n3253), .Z(n3251) );
  XNOR U3256 ( .A(creg[334]), .B(n3252), .Z(n3253) );
  XNOR U3257 ( .A(n3254), .B(n3255), .Z(o[333]) );
  AND U3258 ( .A(n1035), .B(n3256), .Z(n3254) );
  XNOR U3259 ( .A(creg[333]), .B(n3255), .Z(n3256) );
  XNOR U3260 ( .A(n3257), .B(n3258), .Z(o[332]) );
  AND U3261 ( .A(n1035), .B(n3259), .Z(n3257) );
  XNOR U3262 ( .A(creg[332]), .B(n3258), .Z(n3259) );
  XNOR U3263 ( .A(n3260), .B(n3261), .Z(o[331]) );
  AND U3264 ( .A(n1035), .B(n3262), .Z(n3260) );
  XNOR U3265 ( .A(creg[331]), .B(n3261), .Z(n3262) );
  XNOR U3266 ( .A(n3263), .B(n3264), .Z(o[330]) );
  AND U3267 ( .A(n1035), .B(n3265), .Z(n3263) );
  XNOR U3268 ( .A(creg[330]), .B(n3264), .Z(n3265) );
  XNOR U3269 ( .A(n3266), .B(n3267), .Z(o[32]) );
  AND U3270 ( .A(n1035), .B(n3268), .Z(n3266) );
  XNOR U3271 ( .A(creg[32]), .B(n3267), .Z(n3268) );
  XNOR U3272 ( .A(n3269), .B(n3270), .Z(o[329]) );
  AND U3273 ( .A(n1035), .B(n3271), .Z(n3269) );
  XNOR U3274 ( .A(creg[329]), .B(n3270), .Z(n3271) );
  XNOR U3275 ( .A(n3272), .B(n3273), .Z(o[328]) );
  AND U3276 ( .A(n1035), .B(n3274), .Z(n3272) );
  XNOR U3277 ( .A(creg[328]), .B(n3273), .Z(n3274) );
  XNOR U3278 ( .A(n3275), .B(n3276), .Z(o[327]) );
  AND U3279 ( .A(n1035), .B(n3277), .Z(n3275) );
  XNOR U3280 ( .A(creg[327]), .B(n3276), .Z(n3277) );
  XNOR U3281 ( .A(n3278), .B(n3279), .Z(o[326]) );
  AND U3282 ( .A(n1035), .B(n3280), .Z(n3278) );
  XNOR U3283 ( .A(creg[326]), .B(n3279), .Z(n3280) );
  XNOR U3284 ( .A(n3281), .B(n3282), .Z(o[325]) );
  AND U3285 ( .A(n1035), .B(n3283), .Z(n3281) );
  XNOR U3286 ( .A(creg[325]), .B(n3282), .Z(n3283) );
  XNOR U3287 ( .A(n3284), .B(n3285), .Z(o[324]) );
  AND U3288 ( .A(n1035), .B(n3286), .Z(n3284) );
  XNOR U3289 ( .A(creg[324]), .B(n3285), .Z(n3286) );
  XNOR U3290 ( .A(n3287), .B(n3288), .Z(o[323]) );
  AND U3291 ( .A(n1035), .B(n3289), .Z(n3287) );
  XNOR U3292 ( .A(creg[323]), .B(n3288), .Z(n3289) );
  XNOR U3293 ( .A(n3290), .B(n3291), .Z(o[322]) );
  AND U3294 ( .A(n1035), .B(n3292), .Z(n3290) );
  XNOR U3295 ( .A(creg[322]), .B(n3291), .Z(n3292) );
  XNOR U3296 ( .A(n3293), .B(n3294), .Z(o[321]) );
  AND U3297 ( .A(n1035), .B(n3295), .Z(n3293) );
  XNOR U3298 ( .A(creg[321]), .B(n3294), .Z(n3295) );
  XNOR U3299 ( .A(n3296), .B(n3297), .Z(o[320]) );
  AND U3300 ( .A(n1035), .B(n3298), .Z(n3296) );
  XNOR U3301 ( .A(creg[320]), .B(n3297), .Z(n3298) );
  XNOR U3302 ( .A(n3299), .B(n3300), .Z(o[31]) );
  AND U3303 ( .A(n1035), .B(n3301), .Z(n3299) );
  XNOR U3304 ( .A(creg[31]), .B(n3300), .Z(n3301) );
  XNOR U3305 ( .A(n3302), .B(n3303), .Z(o[319]) );
  AND U3306 ( .A(n1035), .B(n3304), .Z(n3302) );
  XNOR U3307 ( .A(creg[319]), .B(n3303), .Z(n3304) );
  XNOR U3308 ( .A(n3305), .B(n3306), .Z(o[318]) );
  AND U3309 ( .A(n1035), .B(n3307), .Z(n3305) );
  XNOR U3310 ( .A(creg[318]), .B(n3306), .Z(n3307) );
  XNOR U3311 ( .A(n3308), .B(n3309), .Z(o[317]) );
  AND U3312 ( .A(n1035), .B(n3310), .Z(n3308) );
  XNOR U3313 ( .A(creg[317]), .B(n3309), .Z(n3310) );
  XNOR U3314 ( .A(n3311), .B(n3312), .Z(o[316]) );
  AND U3315 ( .A(n1035), .B(n3313), .Z(n3311) );
  XNOR U3316 ( .A(creg[316]), .B(n3312), .Z(n3313) );
  XNOR U3317 ( .A(n3314), .B(n3315), .Z(o[315]) );
  AND U3318 ( .A(n1035), .B(n3316), .Z(n3314) );
  XNOR U3319 ( .A(creg[315]), .B(n3315), .Z(n3316) );
  XNOR U3320 ( .A(n3317), .B(n3318), .Z(o[314]) );
  AND U3321 ( .A(n1035), .B(n3319), .Z(n3317) );
  XNOR U3322 ( .A(creg[314]), .B(n3318), .Z(n3319) );
  XNOR U3323 ( .A(n3320), .B(n3321), .Z(o[313]) );
  AND U3324 ( .A(n1035), .B(n3322), .Z(n3320) );
  XNOR U3325 ( .A(creg[313]), .B(n3321), .Z(n3322) );
  XNOR U3326 ( .A(n3323), .B(n3324), .Z(o[312]) );
  AND U3327 ( .A(n1035), .B(n3325), .Z(n3323) );
  XNOR U3328 ( .A(creg[312]), .B(n3324), .Z(n3325) );
  XNOR U3329 ( .A(n3326), .B(n3327), .Z(o[311]) );
  AND U3330 ( .A(n1035), .B(n3328), .Z(n3326) );
  XNOR U3331 ( .A(creg[311]), .B(n3327), .Z(n3328) );
  XNOR U3332 ( .A(n3329), .B(n3330), .Z(o[310]) );
  AND U3333 ( .A(n1035), .B(n3331), .Z(n3329) );
  XNOR U3334 ( .A(creg[310]), .B(n3330), .Z(n3331) );
  XNOR U3335 ( .A(n3332), .B(n3333), .Z(o[30]) );
  AND U3336 ( .A(n1035), .B(n3334), .Z(n3332) );
  XNOR U3337 ( .A(creg[30]), .B(n3333), .Z(n3334) );
  XNOR U3338 ( .A(n3335), .B(n3336), .Z(o[309]) );
  AND U3339 ( .A(n1035), .B(n3337), .Z(n3335) );
  XNOR U3340 ( .A(creg[309]), .B(n3336), .Z(n3337) );
  XNOR U3341 ( .A(n3338), .B(n3339), .Z(o[308]) );
  AND U3342 ( .A(n1035), .B(n3340), .Z(n3338) );
  XNOR U3343 ( .A(creg[308]), .B(n3339), .Z(n3340) );
  XNOR U3344 ( .A(n3341), .B(n3342), .Z(o[307]) );
  AND U3345 ( .A(n1035), .B(n3343), .Z(n3341) );
  XNOR U3346 ( .A(creg[307]), .B(n3342), .Z(n3343) );
  XNOR U3347 ( .A(n3344), .B(n3345), .Z(o[306]) );
  AND U3348 ( .A(n1035), .B(n3346), .Z(n3344) );
  XNOR U3349 ( .A(creg[306]), .B(n3345), .Z(n3346) );
  XNOR U3350 ( .A(n3347), .B(n3348), .Z(o[305]) );
  AND U3351 ( .A(n1035), .B(n3349), .Z(n3347) );
  XNOR U3352 ( .A(creg[305]), .B(n3348), .Z(n3349) );
  XNOR U3353 ( .A(n3350), .B(n3351), .Z(o[304]) );
  AND U3354 ( .A(n1035), .B(n3352), .Z(n3350) );
  XNOR U3355 ( .A(creg[304]), .B(n3351), .Z(n3352) );
  XNOR U3356 ( .A(n3353), .B(n3354), .Z(o[303]) );
  AND U3357 ( .A(n1035), .B(n3355), .Z(n3353) );
  XNOR U3358 ( .A(creg[303]), .B(n3354), .Z(n3355) );
  XNOR U3359 ( .A(n3356), .B(n3357), .Z(o[302]) );
  AND U3360 ( .A(n1035), .B(n3358), .Z(n3356) );
  XNOR U3361 ( .A(creg[302]), .B(n3357), .Z(n3358) );
  XNOR U3362 ( .A(n3359), .B(n3360), .Z(o[301]) );
  AND U3363 ( .A(n1035), .B(n3361), .Z(n3359) );
  XNOR U3364 ( .A(creg[301]), .B(n3360), .Z(n3361) );
  XNOR U3365 ( .A(n3362), .B(n3363), .Z(o[300]) );
  AND U3366 ( .A(n1035), .B(n3364), .Z(n3362) );
  XNOR U3367 ( .A(creg[300]), .B(n3363), .Z(n3364) );
  XNOR U3368 ( .A(n3365), .B(n3366), .Z(o[2]) );
  AND U3369 ( .A(n1035), .B(n3367), .Z(n3365) );
  XNOR U3370 ( .A(creg[2]), .B(n3366), .Z(n3367) );
  XNOR U3371 ( .A(n3368), .B(n3369), .Z(o[29]) );
  AND U3372 ( .A(n1035), .B(n3370), .Z(n3368) );
  XNOR U3373 ( .A(creg[29]), .B(n3369), .Z(n3370) );
  XNOR U3374 ( .A(n3371), .B(n3372), .Z(o[299]) );
  AND U3375 ( .A(n1035), .B(n3373), .Z(n3371) );
  XNOR U3376 ( .A(creg[299]), .B(n3372), .Z(n3373) );
  XNOR U3377 ( .A(n3374), .B(n3375), .Z(o[298]) );
  AND U3378 ( .A(n1035), .B(n3376), .Z(n3374) );
  XNOR U3379 ( .A(creg[298]), .B(n3375), .Z(n3376) );
  XNOR U3380 ( .A(n3377), .B(n3378), .Z(o[297]) );
  AND U3381 ( .A(n1035), .B(n3379), .Z(n3377) );
  XNOR U3382 ( .A(creg[297]), .B(n3378), .Z(n3379) );
  XNOR U3383 ( .A(n3380), .B(n3381), .Z(o[296]) );
  AND U3384 ( .A(n1035), .B(n3382), .Z(n3380) );
  XNOR U3385 ( .A(creg[296]), .B(n3381), .Z(n3382) );
  XNOR U3386 ( .A(n3383), .B(n3384), .Z(o[295]) );
  AND U3387 ( .A(n1035), .B(n3385), .Z(n3383) );
  XNOR U3388 ( .A(creg[295]), .B(n3384), .Z(n3385) );
  XNOR U3389 ( .A(n3386), .B(n3387), .Z(o[294]) );
  AND U3390 ( .A(n1035), .B(n3388), .Z(n3386) );
  XNOR U3391 ( .A(creg[294]), .B(n3387), .Z(n3388) );
  XNOR U3392 ( .A(n3389), .B(n3390), .Z(o[293]) );
  AND U3393 ( .A(n1035), .B(n3391), .Z(n3389) );
  XNOR U3394 ( .A(creg[293]), .B(n3390), .Z(n3391) );
  XNOR U3395 ( .A(n3392), .B(n3393), .Z(o[292]) );
  AND U3396 ( .A(n1035), .B(n3394), .Z(n3392) );
  XNOR U3397 ( .A(creg[292]), .B(n3393), .Z(n3394) );
  XNOR U3398 ( .A(n3395), .B(n3396), .Z(o[291]) );
  AND U3399 ( .A(n1035), .B(n3397), .Z(n3395) );
  XNOR U3400 ( .A(creg[291]), .B(n3396), .Z(n3397) );
  XNOR U3401 ( .A(n3398), .B(n3399), .Z(o[290]) );
  AND U3402 ( .A(n1035), .B(n3400), .Z(n3398) );
  XNOR U3403 ( .A(creg[290]), .B(n3399), .Z(n3400) );
  XNOR U3404 ( .A(n3401), .B(n3402), .Z(o[28]) );
  AND U3405 ( .A(n1035), .B(n3403), .Z(n3401) );
  XNOR U3406 ( .A(creg[28]), .B(n3402), .Z(n3403) );
  XNOR U3407 ( .A(n3404), .B(n3405), .Z(o[289]) );
  AND U3408 ( .A(n1035), .B(n3406), .Z(n3404) );
  XNOR U3409 ( .A(creg[289]), .B(n3405), .Z(n3406) );
  XNOR U3410 ( .A(n3407), .B(n3408), .Z(o[288]) );
  AND U3411 ( .A(n1035), .B(n3409), .Z(n3407) );
  XNOR U3412 ( .A(creg[288]), .B(n3408), .Z(n3409) );
  XNOR U3413 ( .A(n3410), .B(n3411), .Z(o[287]) );
  AND U3414 ( .A(n1035), .B(n3412), .Z(n3410) );
  XNOR U3415 ( .A(creg[287]), .B(n3411), .Z(n3412) );
  XNOR U3416 ( .A(n3413), .B(n3414), .Z(o[286]) );
  AND U3417 ( .A(n1035), .B(n3415), .Z(n3413) );
  XNOR U3418 ( .A(creg[286]), .B(n3414), .Z(n3415) );
  XNOR U3419 ( .A(n3416), .B(n3417), .Z(o[285]) );
  AND U3420 ( .A(n1035), .B(n3418), .Z(n3416) );
  XNOR U3421 ( .A(creg[285]), .B(n3417), .Z(n3418) );
  XNOR U3422 ( .A(n3419), .B(n3420), .Z(o[284]) );
  AND U3423 ( .A(n1035), .B(n3421), .Z(n3419) );
  XNOR U3424 ( .A(creg[284]), .B(n3420), .Z(n3421) );
  XNOR U3425 ( .A(n3422), .B(n3423), .Z(o[283]) );
  AND U3426 ( .A(n1035), .B(n3424), .Z(n3422) );
  XNOR U3427 ( .A(creg[283]), .B(n3423), .Z(n3424) );
  XNOR U3428 ( .A(n3425), .B(n3426), .Z(o[282]) );
  AND U3429 ( .A(n1035), .B(n3427), .Z(n3425) );
  XNOR U3430 ( .A(creg[282]), .B(n3426), .Z(n3427) );
  XNOR U3431 ( .A(n3428), .B(n3429), .Z(o[281]) );
  AND U3432 ( .A(n1035), .B(n3430), .Z(n3428) );
  XNOR U3433 ( .A(creg[281]), .B(n3429), .Z(n3430) );
  XNOR U3434 ( .A(n3431), .B(n3432), .Z(o[280]) );
  AND U3435 ( .A(n1035), .B(n3433), .Z(n3431) );
  XNOR U3436 ( .A(creg[280]), .B(n3432), .Z(n3433) );
  XNOR U3437 ( .A(n3434), .B(n3435), .Z(o[27]) );
  AND U3438 ( .A(n1035), .B(n3436), .Z(n3434) );
  XNOR U3439 ( .A(creg[27]), .B(n3435), .Z(n3436) );
  XNOR U3440 ( .A(n3437), .B(n3438), .Z(o[279]) );
  AND U3441 ( .A(n1035), .B(n3439), .Z(n3437) );
  XNOR U3442 ( .A(creg[279]), .B(n3438), .Z(n3439) );
  XNOR U3443 ( .A(n3440), .B(n3441), .Z(o[278]) );
  AND U3444 ( .A(n1035), .B(n3442), .Z(n3440) );
  XNOR U3445 ( .A(creg[278]), .B(n3441), .Z(n3442) );
  XNOR U3446 ( .A(n3443), .B(n3444), .Z(o[277]) );
  AND U3447 ( .A(n1035), .B(n3445), .Z(n3443) );
  XNOR U3448 ( .A(creg[277]), .B(n3444), .Z(n3445) );
  XNOR U3449 ( .A(n3446), .B(n3447), .Z(o[276]) );
  AND U3450 ( .A(n1035), .B(n3448), .Z(n3446) );
  XNOR U3451 ( .A(creg[276]), .B(n3447), .Z(n3448) );
  XNOR U3452 ( .A(n3449), .B(n3450), .Z(o[275]) );
  AND U3453 ( .A(n1035), .B(n3451), .Z(n3449) );
  XNOR U3454 ( .A(creg[275]), .B(n3450), .Z(n3451) );
  XNOR U3455 ( .A(n3452), .B(n3453), .Z(o[274]) );
  AND U3456 ( .A(n1035), .B(n3454), .Z(n3452) );
  XNOR U3457 ( .A(creg[274]), .B(n3453), .Z(n3454) );
  XNOR U3458 ( .A(n3455), .B(n3456), .Z(o[273]) );
  AND U3459 ( .A(n1035), .B(n3457), .Z(n3455) );
  XNOR U3460 ( .A(creg[273]), .B(n3456), .Z(n3457) );
  XNOR U3461 ( .A(n3458), .B(n3459), .Z(o[272]) );
  AND U3462 ( .A(n1035), .B(n3460), .Z(n3458) );
  XNOR U3463 ( .A(creg[272]), .B(n3459), .Z(n3460) );
  XNOR U3464 ( .A(n3461), .B(n3462), .Z(o[271]) );
  AND U3465 ( .A(n1035), .B(n3463), .Z(n3461) );
  XNOR U3466 ( .A(creg[271]), .B(n3462), .Z(n3463) );
  XNOR U3467 ( .A(n3464), .B(n3465), .Z(o[270]) );
  AND U3468 ( .A(n1035), .B(n3466), .Z(n3464) );
  XNOR U3469 ( .A(creg[270]), .B(n3465), .Z(n3466) );
  XNOR U3470 ( .A(n3467), .B(n3468), .Z(o[26]) );
  AND U3471 ( .A(n1035), .B(n3469), .Z(n3467) );
  XNOR U3472 ( .A(creg[26]), .B(n3468), .Z(n3469) );
  XNOR U3473 ( .A(n3470), .B(n3471), .Z(o[269]) );
  AND U3474 ( .A(n1035), .B(n3472), .Z(n3470) );
  XNOR U3475 ( .A(creg[269]), .B(n3471), .Z(n3472) );
  XNOR U3476 ( .A(n3473), .B(n3474), .Z(o[268]) );
  AND U3477 ( .A(n1035), .B(n3475), .Z(n3473) );
  XNOR U3478 ( .A(creg[268]), .B(n3474), .Z(n3475) );
  XNOR U3479 ( .A(n3476), .B(n3477), .Z(o[267]) );
  AND U3480 ( .A(n1035), .B(n3478), .Z(n3476) );
  XNOR U3481 ( .A(creg[267]), .B(n3477), .Z(n3478) );
  XNOR U3482 ( .A(n3479), .B(n3480), .Z(o[266]) );
  AND U3483 ( .A(n1035), .B(n3481), .Z(n3479) );
  XNOR U3484 ( .A(creg[266]), .B(n3480), .Z(n3481) );
  XNOR U3485 ( .A(n3482), .B(n3483), .Z(o[265]) );
  AND U3486 ( .A(n1035), .B(n3484), .Z(n3482) );
  XNOR U3487 ( .A(creg[265]), .B(n3483), .Z(n3484) );
  XNOR U3488 ( .A(n3485), .B(n3486), .Z(o[264]) );
  AND U3489 ( .A(n1035), .B(n3487), .Z(n3485) );
  XNOR U3490 ( .A(creg[264]), .B(n3486), .Z(n3487) );
  XNOR U3491 ( .A(n3488), .B(n3489), .Z(o[263]) );
  AND U3492 ( .A(n1035), .B(n3490), .Z(n3488) );
  XNOR U3493 ( .A(creg[263]), .B(n3489), .Z(n3490) );
  XNOR U3494 ( .A(n3491), .B(n3492), .Z(o[262]) );
  AND U3495 ( .A(n1035), .B(n3493), .Z(n3491) );
  XNOR U3496 ( .A(creg[262]), .B(n3492), .Z(n3493) );
  XNOR U3497 ( .A(n3494), .B(n3495), .Z(o[261]) );
  AND U3498 ( .A(n1035), .B(n3496), .Z(n3494) );
  XNOR U3499 ( .A(creg[261]), .B(n3495), .Z(n3496) );
  XNOR U3500 ( .A(n3497), .B(n3498), .Z(o[260]) );
  AND U3501 ( .A(n1035), .B(n3499), .Z(n3497) );
  XNOR U3502 ( .A(creg[260]), .B(n3498), .Z(n3499) );
  XNOR U3503 ( .A(n3500), .B(n3501), .Z(o[25]) );
  AND U3504 ( .A(n1035), .B(n3502), .Z(n3500) );
  XNOR U3505 ( .A(creg[25]), .B(n3501), .Z(n3502) );
  XNOR U3506 ( .A(n3503), .B(n3504), .Z(o[259]) );
  AND U3507 ( .A(n1035), .B(n3505), .Z(n3503) );
  XNOR U3508 ( .A(creg[259]), .B(n3504), .Z(n3505) );
  XNOR U3509 ( .A(n3506), .B(n3507), .Z(o[258]) );
  AND U3510 ( .A(n1035), .B(n3508), .Z(n3506) );
  XNOR U3511 ( .A(creg[258]), .B(n3507), .Z(n3508) );
  XNOR U3512 ( .A(n3509), .B(n3510), .Z(o[257]) );
  AND U3513 ( .A(n1035), .B(n3511), .Z(n3509) );
  XNOR U3514 ( .A(creg[257]), .B(n3510), .Z(n3511) );
  XNOR U3515 ( .A(n3512), .B(n3513), .Z(o[256]) );
  AND U3516 ( .A(n1035), .B(n3514), .Z(n3512) );
  XNOR U3517 ( .A(creg[256]), .B(n3513), .Z(n3514) );
  XNOR U3518 ( .A(n3515), .B(n3516), .Z(o[255]) );
  AND U3519 ( .A(n1035), .B(n3517), .Z(n3515) );
  XNOR U3520 ( .A(creg[255]), .B(n3516), .Z(n3517) );
  XNOR U3521 ( .A(n3518), .B(n3519), .Z(o[254]) );
  AND U3522 ( .A(n1035), .B(n3520), .Z(n3518) );
  XNOR U3523 ( .A(creg[254]), .B(n3519), .Z(n3520) );
  XNOR U3524 ( .A(n3521), .B(n3522), .Z(o[253]) );
  AND U3525 ( .A(n1035), .B(n3523), .Z(n3521) );
  XNOR U3526 ( .A(creg[253]), .B(n3522), .Z(n3523) );
  XNOR U3527 ( .A(n3524), .B(n3525), .Z(o[252]) );
  AND U3528 ( .A(n1035), .B(n3526), .Z(n3524) );
  XNOR U3529 ( .A(creg[252]), .B(n3525), .Z(n3526) );
  XNOR U3530 ( .A(n3527), .B(n3528), .Z(o[251]) );
  AND U3531 ( .A(n1035), .B(n3529), .Z(n3527) );
  XNOR U3532 ( .A(creg[251]), .B(n3528), .Z(n3529) );
  XNOR U3533 ( .A(n3530), .B(n3531), .Z(o[250]) );
  AND U3534 ( .A(n1035), .B(n3532), .Z(n3530) );
  XNOR U3535 ( .A(creg[250]), .B(n3531), .Z(n3532) );
  XNOR U3536 ( .A(n3533), .B(n3534), .Z(o[24]) );
  AND U3537 ( .A(n1035), .B(n3535), .Z(n3533) );
  XNOR U3538 ( .A(creg[24]), .B(n3534), .Z(n3535) );
  XNOR U3539 ( .A(n3536), .B(n3537), .Z(o[249]) );
  AND U3540 ( .A(n1035), .B(n3538), .Z(n3536) );
  XNOR U3541 ( .A(creg[249]), .B(n3537), .Z(n3538) );
  XNOR U3542 ( .A(n3539), .B(n3540), .Z(o[248]) );
  AND U3543 ( .A(n1035), .B(n3541), .Z(n3539) );
  XNOR U3544 ( .A(creg[248]), .B(n3540), .Z(n3541) );
  XNOR U3545 ( .A(n3542), .B(n3543), .Z(o[247]) );
  AND U3546 ( .A(n1035), .B(n3544), .Z(n3542) );
  XNOR U3547 ( .A(creg[247]), .B(n3543), .Z(n3544) );
  XNOR U3548 ( .A(n3545), .B(n3546), .Z(o[246]) );
  AND U3549 ( .A(n1035), .B(n3547), .Z(n3545) );
  XNOR U3550 ( .A(creg[246]), .B(n3546), .Z(n3547) );
  XNOR U3551 ( .A(n3548), .B(n3549), .Z(o[245]) );
  AND U3552 ( .A(n1035), .B(n3550), .Z(n3548) );
  XNOR U3553 ( .A(creg[245]), .B(n3549), .Z(n3550) );
  XNOR U3554 ( .A(n3551), .B(n3552), .Z(o[244]) );
  AND U3555 ( .A(n1035), .B(n3553), .Z(n3551) );
  XNOR U3556 ( .A(creg[244]), .B(n3552), .Z(n3553) );
  XNOR U3557 ( .A(n3554), .B(n3555), .Z(o[243]) );
  AND U3558 ( .A(n1035), .B(n3556), .Z(n3554) );
  XNOR U3559 ( .A(creg[243]), .B(n3555), .Z(n3556) );
  XNOR U3560 ( .A(n3557), .B(n3558), .Z(o[242]) );
  AND U3561 ( .A(n1035), .B(n3559), .Z(n3557) );
  XNOR U3562 ( .A(creg[242]), .B(n3558), .Z(n3559) );
  XNOR U3563 ( .A(n3560), .B(n3561), .Z(o[241]) );
  AND U3564 ( .A(n1035), .B(n3562), .Z(n3560) );
  XNOR U3565 ( .A(creg[241]), .B(n3561), .Z(n3562) );
  XNOR U3566 ( .A(n3563), .B(n3564), .Z(o[240]) );
  AND U3567 ( .A(n1035), .B(n3565), .Z(n3563) );
  XNOR U3568 ( .A(creg[240]), .B(n3564), .Z(n3565) );
  XNOR U3569 ( .A(n3566), .B(n3567), .Z(o[23]) );
  AND U3570 ( .A(n1035), .B(n3568), .Z(n3566) );
  XNOR U3571 ( .A(creg[23]), .B(n3567), .Z(n3568) );
  XNOR U3572 ( .A(n3569), .B(n3570), .Z(o[239]) );
  AND U3573 ( .A(n1035), .B(n3571), .Z(n3569) );
  XNOR U3574 ( .A(creg[239]), .B(n3570), .Z(n3571) );
  XNOR U3575 ( .A(n3572), .B(n3573), .Z(o[238]) );
  AND U3576 ( .A(n1035), .B(n3574), .Z(n3572) );
  XNOR U3577 ( .A(creg[238]), .B(n3573), .Z(n3574) );
  XNOR U3578 ( .A(n3575), .B(n3576), .Z(o[237]) );
  AND U3579 ( .A(n1035), .B(n3577), .Z(n3575) );
  XNOR U3580 ( .A(creg[237]), .B(n3576), .Z(n3577) );
  XNOR U3581 ( .A(n3578), .B(n3579), .Z(o[236]) );
  AND U3582 ( .A(n1035), .B(n3580), .Z(n3578) );
  XNOR U3583 ( .A(creg[236]), .B(n3579), .Z(n3580) );
  XNOR U3584 ( .A(n3581), .B(n3582), .Z(o[235]) );
  AND U3585 ( .A(n1035), .B(n3583), .Z(n3581) );
  XNOR U3586 ( .A(creg[235]), .B(n3582), .Z(n3583) );
  XNOR U3587 ( .A(n3584), .B(n3585), .Z(o[234]) );
  AND U3588 ( .A(n1035), .B(n3586), .Z(n3584) );
  XNOR U3589 ( .A(creg[234]), .B(n3585), .Z(n3586) );
  XNOR U3590 ( .A(n3587), .B(n3588), .Z(o[233]) );
  AND U3591 ( .A(n1035), .B(n3589), .Z(n3587) );
  XNOR U3592 ( .A(creg[233]), .B(n3588), .Z(n3589) );
  XNOR U3593 ( .A(n3590), .B(n3591), .Z(o[232]) );
  AND U3594 ( .A(n1035), .B(n3592), .Z(n3590) );
  XNOR U3595 ( .A(creg[232]), .B(n3591), .Z(n3592) );
  XNOR U3596 ( .A(n3593), .B(n3594), .Z(o[231]) );
  AND U3597 ( .A(n1035), .B(n3595), .Z(n3593) );
  XNOR U3598 ( .A(creg[231]), .B(n3594), .Z(n3595) );
  XNOR U3599 ( .A(n3596), .B(n3597), .Z(o[230]) );
  AND U3600 ( .A(n1035), .B(n3598), .Z(n3596) );
  XNOR U3601 ( .A(creg[230]), .B(n3597), .Z(n3598) );
  XNOR U3602 ( .A(n3599), .B(n3600), .Z(o[22]) );
  AND U3603 ( .A(n1035), .B(n3601), .Z(n3599) );
  XNOR U3604 ( .A(creg[22]), .B(n3600), .Z(n3601) );
  XNOR U3605 ( .A(n3602), .B(n3603), .Z(o[229]) );
  AND U3606 ( .A(n1035), .B(n3604), .Z(n3602) );
  XNOR U3607 ( .A(creg[229]), .B(n3603), .Z(n3604) );
  XNOR U3608 ( .A(n3605), .B(n3606), .Z(o[228]) );
  AND U3609 ( .A(n1035), .B(n3607), .Z(n3605) );
  XNOR U3610 ( .A(creg[228]), .B(n3606), .Z(n3607) );
  XNOR U3611 ( .A(n3608), .B(n3609), .Z(o[227]) );
  AND U3612 ( .A(n1035), .B(n3610), .Z(n3608) );
  XNOR U3613 ( .A(creg[227]), .B(n3609), .Z(n3610) );
  XNOR U3614 ( .A(n3611), .B(n3612), .Z(o[226]) );
  AND U3615 ( .A(n1035), .B(n3613), .Z(n3611) );
  XNOR U3616 ( .A(creg[226]), .B(n3612), .Z(n3613) );
  XNOR U3617 ( .A(n3614), .B(n3615), .Z(o[225]) );
  AND U3618 ( .A(n1035), .B(n3616), .Z(n3614) );
  XNOR U3619 ( .A(creg[225]), .B(n3615), .Z(n3616) );
  XNOR U3620 ( .A(n3617), .B(n3618), .Z(o[224]) );
  AND U3621 ( .A(n1035), .B(n3619), .Z(n3617) );
  XNOR U3622 ( .A(creg[224]), .B(n3618), .Z(n3619) );
  XNOR U3623 ( .A(n3620), .B(n3621), .Z(o[223]) );
  AND U3624 ( .A(n1035), .B(n3622), .Z(n3620) );
  XNOR U3625 ( .A(creg[223]), .B(n3621), .Z(n3622) );
  XNOR U3626 ( .A(n3623), .B(n3624), .Z(o[222]) );
  AND U3627 ( .A(n1035), .B(n3625), .Z(n3623) );
  XNOR U3628 ( .A(creg[222]), .B(n3624), .Z(n3625) );
  XNOR U3629 ( .A(n3626), .B(n3627), .Z(o[221]) );
  AND U3630 ( .A(n1035), .B(n3628), .Z(n3626) );
  XNOR U3631 ( .A(creg[221]), .B(n3627), .Z(n3628) );
  XNOR U3632 ( .A(n3629), .B(n3630), .Z(o[220]) );
  AND U3633 ( .A(n1035), .B(n3631), .Z(n3629) );
  XNOR U3634 ( .A(creg[220]), .B(n3630), .Z(n3631) );
  XNOR U3635 ( .A(n3632), .B(n3633), .Z(o[21]) );
  AND U3636 ( .A(n1035), .B(n3634), .Z(n3632) );
  XNOR U3637 ( .A(creg[21]), .B(n3633), .Z(n3634) );
  XNOR U3638 ( .A(n3635), .B(n3636), .Z(o[219]) );
  AND U3639 ( .A(n1035), .B(n3637), .Z(n3635) );
  XNOR U3640 ( .A(creg[219]), .B(n3636), .Z(n3637) );
  XNOR U3641 ( .A(n3638), .B(n3639), .Z(o[218]) );
  AND U3642 ( .A(n1035), .B(n3640), .Z(n3638) );
  XNOR U3643 ( .A(creg[218]), .B(n3639), .Z(n3640) );
  XNOR U3644 ( .A(n3641), .B(n3642), .Z(o[217]) );
  AND U3645 ( .A(n1035), .B(n3643), .Z(n3641) );
  XNOR U3646 ( .A(creg[217]), .B(n3642), .Z(n3643) );
  XNOR U3647 ( .A(n3644), .B(n3645), .Z(o[216]) );
  AND U3648 ( .A(n1035), .B(n3646), .Z(n3644) );
  XNOR U3649 ( .A(creg[216]), .B(n3645), .Z(n3646) );
  XNOR U3650 ( .A(n3647), .B(n3648), .Z(o[215]) );
  AND U3651 ( .A(n1035), .B(n3649), .Z(n3647) );
  XNOR U3652 ( .A(creg[215]), .B(n3648), .Z(n3649) );
  XNOR U3653 ( .A(n3650), .B(n3651), .Z(o[214]) );
  AND U3654 ( .A(n1035), .B(n3652), .Z(n3650) );
  XNOR U3655 ( .A(creg[214]), .B(n3651), .Z(n3652) );
  XNOR U3656 ( .A(n3653), .B(n3654), .Z(o[213]) );
  AND U3657 ( .A(n1035), .B(n3655), .Z(n3653) );
  XNOR U3658 ( .A(creg[213]), .B(n3654), .Z(n3655) );
  XNOR U3659 ( .A(n3656), .B(n3657), .Z(o[212]) );
  AND U3660 ( .A(n1035), .B(n3658), .Z(n3656) );
  XNOR U3661 ( .A(creg[212]), .B(n3657), .Z(n3658) );
  XNOR U3662 ( .A(n3659), .B(n3660), .Z(o[211]) );
  AND U3663 ( .A(n1035), .B(n3661), .Z(n3659) );
  XNOR U3664 ( .A(creg[211]), .B(n3660), .Z(n3661) );
  XNOR U3665 ( .A(n3662), .B(n3663), .Z(o[210]) );
  AND U3666 ( .A(n1035), .B(n3664), .Z(n3662) );
  XNOR U3667 ( .A(creg[210]), .B(n3663), .Z(n3664) );
  XNOR U3668 ( .A(n3665), .B(n3666), .Z(o[20]) );
  AND U3669 ( .A(n1035), .B(n3667), .Z(n3665) );
  XNOR U3670 ( .A(creg[20]), .B(n3666), .Z(n3667) );
  XNOR U3671 ( .A(n3668), .B(n3669), .Z(o[209]) );
  AND U3672 ( .A(n1035), .B(n3670), .Z(n3668) );
  XNOR U3673 ( .A(creg[209]), .B(n3669), .Z(n3670) );
  XNOR U3674 ( .A(n3671), .B(n3672), .Z(o[208]) );
  AND U3675 ( .A(n1035), .B(n3673), .Z(n3671) );
  XNOR U3676 ( .A(creg[208]), .B(n3672), .Z(n3673) );
  XNOR U3677 ( .A(n3674), .B(n3675), .Z(o[207]) );
  AND U3678 ( .A(n1035), .B(n3676), .Z(n3674) );
  XNOR U3679 ( .A(creg[207]), .B(n3675), .Z(n3676) );
  XNOR U3680 ( .A(n3677), .B(n3678), .Z(o[206]) );
  AND U3681 ( .A(n1035), .B(n3679), .Z(n3677) );
  XNOR U3682 ( .A(creg[206]), .B(n3678), .Z(n3679) );
  XNOR U3683 ( .A(n3680), .B(n3681), .Z(o[205]) );
  AND U3684 ( .A(n1035), .B(n3682), .Z(n3680) );
  XNOR U3685 ( .A(creg[205]), .B(n3681), .Z(n3682) );
  XNOR U3686 ( .A(n3683), .B(n3684), .Z(o[204]) );
  AND U3687 ( .A(n1035), .B(n3685), .Z(n3683) );
  XNOR U3688 ( .A(creg[204]), .B(n3684), .Z(n3685) );
  XNOR U3689 ( .A(n3686), .B(n3687), .Z(o[203]) );
  AND U3690 ( .A(n1035), .B(n3688), .Z(n3686) );
  XNOR U3691 ( .A(creg[203]), .B(n3687), .Z(n3688) );
  XNOR U3692 ( .A(n3689), .B(n3690), .Z(o[202]) );
  AND U3693 ( .A(n1035), .B(n3691), .Z(n3689) );
  XNOR U3694 ( .A(creg[202]), .B(n3690), .Z(n3691) );
  XNOR U3695 ( .A(n3692), .B(n3693), .Z(o[201]) );
  AND U3696 ( .A(n1035), .B(n3694), .Z(n3692) );
  XNOR U3697 ( .A(creg[201]), .B(n3693), .Z(n3694) );
  XNOR U3698 ( .A(n3695), .B(n3696), .Z(o[200]) );
  AND U3699 ( .A(n1035), .B(n3697), .Z(n3695) );
  XNOR U3700 ( .A(creg[200]), .B(n3696), .Z(n3697) );
  XNOR U3701 ( .A(n3698), .B(n3699), .Z(o[1]) );
  AND U3702 ( .A(n1035), .B(n3700), .Z(n3698) );
  XNOR U3703 ( .A(creg[1]), .B(n3699), .Z(n3700) );
  XNOR U3704 ( .A(n3701), .B(n3702), .Z(o[19]) );
  AND U3705 ( .A(n1035), .B(n3703), .Z(n3701) );
  XNOR U3706 ( .A(creg[19]), .B(n3702), .Z(n3703) );
  XNOR U3707 ( .A(n3704), .B(n3705), .Z(o[199]) );
  AND U3708 ( .A(n1035), .B(n3706), .Z(n3704) );
  XNOR U3709 ( .A(creg[199]), .B(n3705), .Z(n3706) );
  XNOR U3710 ( .A(n3707), .B(n3708), .Z(o[198]) );
  AND U3711 ( .A(n1035), .B(n3709), .Z(n3707) );
  XNOR U3712 ( .A(creg[198]), .B(n3708), .Z(n3709) );
  XNOR U3713 ( .A(n3710), .B(n3711), .Z(o[197]) );
  AND U3714 ( .A(n1035), .B(n3712), .Z(n3710) );
  XNOR U3715 ( .A(creg[197]), .B(n3711), .Z(n3712) );
  XNOR U3716 ( .A(n3713), .B(n3714), .Z(o[196]) );
  AND U3717 ( .A(n1035), .B(n3715), .Z(n3713) );
  XNOR U3718 ( .A(creg[196]), .B(n3714), .Z(n3715) );
  XNOR U3719 ( .A(n3716), .B(n3717), .Z(o[195]) );
  AND U3720 ( .A(n1035), .B(n3718), .Z(n3716) );
  XNOR U3721 ( .A(creg[195]), .B(n3717), .Z(n3718) );
  XNOR U3722 ( .A(n3719), .B(n3720), .Z(o[194]) );
  AND U3723 ( .A(n1035), .B(n3721), .Z(n3719) );
  XNOR U3724 ( .A(creg[194]), .B(n3720), .Z(n3721) );
  XNOR U3725 ( .A(n3722), .B(n3723), .Z(o[193]) );
  AND U3726 ( .A(n1035), .B(n3724), .Z(n3722) );
  XNOR U3727 ( .A(creg[193]), .B(n3723), .Z(n3724) );
  XNOR U3728 ( .A(n3725), .B(n3726), .Z(o[192]) );
  AND U3729 ( .A(n1035), .B(n3727), .Z(n3725) );
  XNOR U3730 ( .A(creg[192]), .B(n3726), .Z(n3727) );
  XNOR U3731 ( .A(n3728), .B(n3729), .Z(o[191]) );
  AND U3732 ( .A(n1035), .B(n3730), .Z(n3728) );
  XNOR U3733 ( .A(creg[191]), .B(n3729), .Z(n3730) );
  XNOR U3734 ( .A(n3731), .B(n3732), .Z(o[190]) );
  AND U3735 ( .A(n1035), .B(n3733), .Z(n3731) );
  XNOR U3736 ( .A(creg[190]), .B(n3732), .Z(n3733) );
  XNOR U3737 ( .A(n3734), .B(n3735), .Z(o[18]) );
  AND U3738 ( .A(n1035), .B(n3736), .Z(n3734) );
  XNOR U3739 ( .A(creg[18]), .B(n3735), .Z(n3736) );
  XNOR U3740 ( .A(n3737), .B(n3738), .Z(o[189]) );
  AND U3741 ( .A(n1035), .B(n3739), .Z(n3737) );
  XNOR U3742 ( .A(creg[189]), .B(n3738), .Z(n3739) );
  XNOR U3743 ( .A(n3740), .B(n3741), .Z(o[188]) );
  AND U3744 ( .A(n1035), .B(n3742), .Z(n3740) );
  XNOR U3745 ( .A(creg[188]), .B(n3741), .Z(n3742) );
  XNOR U3746 ( .A(n3743), .B(n3744), .Z(o[187]) );
  AND U3747 ( .A(n1035), .B(n3745), .Z(n3743) );
  XNOR U3748 ( .A(creg[187]), .B(n3744), .Z(n3745) );
  XNOR U3749 ( .A(n3746), .B(n3747), .Z(o[186]) );
  AND U3750 ( .A(n1035), .B(n3748), .Z(n3746) );
  XNOR U3751 ( .A(creg[186]), .B(n3747), .Z(n3748) );
  XNOR U3752 ( .A(n3749), .B(n3750), .Z(o[185]) );
  AND U3753 ( .A(n1035), .B(n3751), .Z(n3749) );
  XNOR U3754 ( .A(creg[185]), .B(n3750), .Z(n3751) );
  XNOR U3755 ( .A(n3752), .B(n3753), .Z(o[184]) );
  AND U3756 ( .A(n1035), .B(n3754), .Z(n3752) );
  XNOR U3757 ( .A(creg[184]), .B(n3753), .Z(n3754) );
  XNOR U3758 ( .A(n3755), .B(n3756), .Z(o[183]) );
  AND U3759 ( .A(n1035), .B(n3757), .Z(n3755) );
  XNOR U3760 ( .A(creg[183]), .B(n3756), .Z(n3757) );
  XNOR U3761 ( .A(n3758), .B(n3759), .Z(o[182]) );
  AND U3762 ( .A(n1035), .B(n3760), .Z(n3758) );
  XNOR U3763 ( .A(creg[182]), .B(n3759), .Z(n3760) );
  XNOR U3764 ( .A(n3761), .B(n3762), .Z(o[181]) );
  AND U3765 ( .A(n1035), .B(n3763), .Z(n3761) );
  XNOR U3766 ( .A(creg[181]), .B(n3762), .Z(n3763) );
  XNOR U3767 ( .A(n3764), .B(n3765), .Z(o[180]) );
  AND U3768 ( .A(n1035), .B(n3766), .Z(n3764) );
  XNOR U3769 ( .A(creg[180]), .B(n3765), .Z(n3766) );
  XNOR U3770 ( .A(n3767), .B(n3768), .Z(o[17]) );
  AND U3771 ( .A(n1035), .B(n3769), .Z(n3767) );
  XNOR U3772 ( .A(creg[17]), .B(n3768), .Z(n3769) );
  XNOR U3773 ( .A(n3770), .B(n3771), .Z(o[179]) );
  AND U3774 ( .A(n1035), .B(n3772), .Z(n3770) );
  XNOR U3775 ( .A(creg[179]), .B(n3771), .Z(n3772) );
  XNOR U3776 ( .A(n3773), .B(n3774), .Z(o[178]) );
  AND U3777 ( .A(n1035), .B(n3775), .Z(n3773) );
  XNOR U3778 ( .A(creg[178]), .B(n3774), .Z(n3775) );
  XNOR U3779 ( .A(n3776), .B(n3777), .Z(o[177]) );
  AND U3780 ( .A(n1035), .B(n3778), .Z(n3776) );
  XNOR U3781 ( .A(creg[177]), .B(n3777), .Z(n3778) );
  XNOR U3782 ( .A(n3779), .B(n3780), .Z(o[176]) );
  AND U3783 ( .A(n1035), .B(n3781), .Z(n3779) );
  XNOR U3784 ( .A(creg[176]), .B(n3780), .Z(n3781) );
  XNOR U3785 ( .A(n3782), .B(n3783), .Z(o[175]) );
  AND U3786 ( .A(n1035), .B(n3784), .Z(n3782) );
  XNOR U3787 ( .A(creg[175]), .B(n3783), .Z(n3784) );
  XNOR U3788 ( .A(n3785), .B(n3786), .Z(o[174]) );
  AND U3789 ( .A(n1035), .B(n3787), .Z(n3785) );
  XNOR U3790 ( .A(creg[174]), .B(n3786), .Z(n3787) );
  XNOR U3791 ( .A(n3788), .B(n3789), .Z(o[173]) );
  AND U3792 ( .A(n1035), .B(n3790), .Z(n3788) );
  XNOR U3793 ( .A(creg[173]), .B(n3789), .Z(n3790) );
  XNOR U3794 ( .A(n3791), .B(n3792), .Z(o[172]) );
  AND U3795 ( .A(n1035), .B(n3793), .Z(n3791) );
  XNOR U3796 ( .A(creg[172]), .B(n3792), .Z(n3793) );
  XNOR U3797 ( .A(n3794), .B(n3795), .Z(o[171]) );
  AND U3798 ( .A(n1035), .B(n3796), .Z(n3794) );
  XNOR U3799 ( .A(creg[171]), .B(n3795), .Z(n3796) );
  XNOR U3800 ( .A(n3797), .B(n3798), .Z(o[170]) );
  AND U3801 ( .A(n1035), .B(n3799), .Z(n3797) );
  XNOR U3802 ( .A(creg[170]), .B(n3798), .Z(n3799) );
  XNOR U3803 ( .A(n3800), .B(n3801), .Z(o[16]) );
  AND U3804 ( .A(n1035), .B(n3802), .Z(n3800) );
  XNOR U3805 ( .A(creg[16]), .B(n3801), .Z(n3802) );
  XNOR U3806 ( .A(n3803), .B(n3804), .Z(o[169]) );
  AND U3807 ( .A(n1035), .B(n3805), .Z(n3803) );
  XNOR U3808 ( .A(creg[169]), .B(n3804), .Z(n3805) );
  XNOR U3809 ( .A(n3806), .B(n3807), .Z(o[168]) );
  AND U3810 ( .A(n1035), .B(n3808), .Z(n3806) );
  XNOR U3811 ( .A(creg[168]), .B(n3807), .Z(n3808) );
  XNOR U3812 ( .A(n3809), .B(n3810), .Z(o[167]) );
  AND U3813 ( .A(n1035), .B(n3811), .Z(n3809) );
  XNOR U3814 ( .A(creg[167]), .B(n3810), .Z(n3811) );
  XNOR U3815 ( .A(n3812), .B(n3813), .Z(o[166]) );
  AND U3816 ( .A(n1035), .B(n3814), .Z(n3812) );
  XNOR U3817 ( .A(creg[166]), .B(n3813), .Z(n3814) );
  XNOR U3818 ( .A(n3815), .B(n3816), .Z(o[165]) );
  AND U3819 ( .A(n1035), .B(n3817), .Z(n3815) );
  XNOR U3820 ( .A(creg[165]), .B(n3816), .Z(n3817) );
  XNOR U3821 ( .A(n3818), .B(n3819), .Z(o[164]) );
  AND U3822 ( .A(n1035), .B(n3820), .Z(n3818) );
  XNOR U3823 ( .A(creg[164]), .B(n3819), .Z(n3820) );
  XNOR U3824 ( .A(n3821), .B(n3822), .Z(o[163]) );
  AND U3825 ( .A(n1035), .B(n3823), .Z(n3821) );
  XNOR U3826 ( .A(creg[163]), .B(n3822), .Z(n3823) );
  XNOR U3827 ( .A(n3824), .B(n3825), .Z(o[162]) );
  AND U3828 ( .A(n1035), .B(n3826), .Z(n3824) );
  XNOR U3829 ( .A(creg[162]), .B(n3825), .Z(n3826) );
  XNOR U3830 ( .A(n3827), .B(n3828), .Z(o[161]) );
  AND U3831 ( .A(n1035), .B(n3829), .Z(n3827) );
  XNOR U3832 ( .A(creg[161]), .B(n3828), .Z(n3829) );
  XNOR U3833 ( .A(n3830), .B(n3831), .Z(o[160]) );
  AND U3834 ( .A(n1035), .B(n3832), .Z(n3830) );
  XNOR U3835 ( .A(creg[160]), .B(n3831), .Z(n3832) );
  XNOR U3836 ( .A(n3833), .B(n3834), .Z(o[15]) );
  AND U3837 ( .A(n1035), .B(n3835), .Z(n3833) );
  XNOR U3838 ( .A(creg[15]), .B(n3834), .Z(n3835) );
  XNOR U3839 ( .A(n3836), .B(n3837), .Z(o[159]) );
  AND U3840 ( .A(n1035), .B(n3838), .Z(n3836) );
  XNOR U3841 ( .A(creg[159]), .B(n3837), .Z(n3838) );
  XNOR U3842 ( .A(n3839), .B(n3840), .Z(o[158]) );
  AND U3843 ( .A(n1035), .B(n3841), .Z(n3839) );
  XNOR U3844 ( .A(creg[158]), .B(n3840), .Z(n3841) );
  XNOR U3845 ( .A(n3842), .B(n3843), .Z(o[157]) );
  AND U3846 ( .A(n1035), .B(n3844), .Z(n3842) );
  XNOR U3847 ( .A(creg[157]), .B(n3843), .Z(n3844) );
  XNOR U3848 ( .A(n3845), .B(n3846), .Z(o[156]) );
  AND U3849 ( .A(n1035), .B(n3847), .Z(n3845) );
  XNOR U3850 ( .A(creg[156]), .B(n3846), .Z(n3847) );
  XNOR U3851 ( .A(n3848), .B(n3849), .Z(o[155]) );
  AND U3852 ( .A(n1035), .B(n3850), .Z(n3848) );
  XNOR U3853 ( .A(creg[155]), .B(n3849), .Z(n3850) );
  XNOR U3854 ( .A(n3851), .B(n3852), .Z(o[154]) );
  AND U3855 ( .A(n1035), .B(n3853), .Z(n3851) );
  XNOR U3856 ( .A(creg[154]), .B(n3852), .Z(n3853) );
  XNOR U3857 ( .A(n3854), .B(n3855), .Z(o[153]) );
  AND U3858 ( .A(n1035), .B(n3856), .Z(n3854) );
  XNOR U3859 ( .A(creg[153]), .B(n3855), .Z(n3856) );
  XNOR U3860 ( .A(n3857), .B(n3858), .Z(o[152]) );
  AND U3861 ( .A(n1035), .B(n3859), .Z(n3857) );
  XNOR U3862 ( .A(creg[152]), .B(n3858), .Z(n3859) );
  XNOR U3863 ( .A(n3860), .B(n3861), .Z(o[151]) );
  AND U3864 ( .A(n1035), .B(n3862), .Z(n3860) );
  XNOR U3865 ( .A(creg[151]), .B(n3861), .Z(n3862) );
  XNOR U3866 ( .A(n3863), .B(n3864), .Z(o[150]) );
  AND U3867 ( .A(n1035), .B(n3865), .Z(n3863) );
  XNOR U3868 ( .A(creg[150]), .B(n3864), .Z(n3865) );
  XNOR U3869 ( .A(n3866), .B(n3867), .Z(o[14]) );
  AND U3870 ( .A(n1035), .B(n3868), .Z(n3866) );
  XNOR U3871 ( .A(creg[14]), .B(n3867), .Z(n3868) );
  XNOR U3872 ( .A(n3869), .B(n3870), .Z(o[149]) );
  AND U3873 ( .A(n1035), .B(n3871), .Z(n3869) );
  XNOR U3874 ( .A(creg[149]), .B(n3870), .Z(n3871) );
  XNOR U3875 ( .A(n3872), .B(n3873), .Z(o[148]) );
  AND U3876 ( .A(n1035), .B(n3874), .Z(n3872) );
  XNOR U3877 ( .A(creg[148]), .B(n3873), .Z(n3874) );
  XNOR U3878 ( .A(n3875), .B(n3876), .Z(o[147]) );
  AND U3879 ( .A(n1035), .B(n3877), .Z(n3875) );
  XNOR U3880 ( .A(creg[147]), .B(n3876), .Z(n3877) );
  XNOR U3881 ( .A(n3878), .B(n3879), .Z(o[146]) );
  AND U3882 ( .A(n1035), .B(n3880), .Z(n3878) );
  XNOR U3883 ( .A(creg[146]), .B(n3879), .Z(n3880) );
  XNOR U3884 ( .A(n3881), .B(n3882), .Z(o[145]) );
  AND U3885 ( .A(n1035), .B(n3883), .Z(n3881) );
  XNOR U3886 ( .A(creg[145]), .B(n3882), .Z(n3883) );
  XNOR U3887 ( .A(n3884), .B(n3885), .Z(o[144]) );
  AND U3888 ( .A(n1035), .B(n3886), .Z(n3884) );
  XNOR U3889 ( .A(creg[144]), .B(n3885), .Z(n3886) );
  XNOR U3890 ( .A(n3887), .B(n3888), .Z(o[143]) );
  AND U3891 ( .A(n1035), .B(n3889), .Z(n3887) );
  XNOR U3892 ( .A(creg[143]), .B(n3888), .Z(n3889) );
  XNOR U3893 ( .A(n3890), .B(n3891), .Z(o[142]) );
  AND U3894 ( .A(n1035), .B(n3892), .Z(n3890) );
  XNOR U3895 ( .A(creg[142]), .B(n3891), .Z(n3892) );
  XNOR U3896 ( .A(n3893), .B(n3894), .Z(o[141]) );
  AND U3897 ( .A(n1035), .B(n3895), .Z(n3893) );
  XNOR U3898 ( .A(creg[141]), .B(n3894), .Z(n3895) );
  XNOR U3899 ( .A(n3896), .B(n3897), .Z(o[140]) );
  AND U3900 ( .A(n1035), .B(n3898), .Z(n3896) );
  XNOR U3901 ( .A(creg[140]), .B(n3897), .Z(n3898) );
  XNOR U3902 ( .A(n3899), .B(n3900), .Z(o[13]) );
  AND U3903 ( .A(n1035), .B(n3901), .Z(n3899) );
  XNOR U3904 ( .A(creg[13]), .B(n3900), .Z(n3901) );
  XNOR U3905 ( .A(n3902), .B(n3903), .Z(o[139]) );
  AND U3906 ( .A(n1035), .B(n3904), .Z(n3902) );
  XNOR U3907 ( .A(creg[139]), .B(n3903), .Z(n3904) );
  XNOR U3908 ( .A(n3905), .B(n3906), .Z(o[138]) );
  AND U3909 ( .A(n1035), .B(n3907), .Z(n3905) );
  XNOR U3910 ( .A(creg[138]), .B(n3906), .Z(n3907) );
  XNOR U3911 ( .A(n3908), .B(n3909), .Z(o[137]) );
  AND U3912 ( .A(n1035), .B(n3910), .Z(n3908) );
  XNOR U3913 ( .A(creg[137]), .B(n3909), .Z(n3910) );
  XNOR U3914 ( .A(n3911), .B(n3912), .Z(o[136]) );
  AND U3915 ( .A(n1035), .B(n3913), .Z(n3911) );
  XNOR U3916 ( .A(creg[136]), .B(n3912), .Z(n3913) );
  XNOR U3917 ( .A(n3914), .B(n3915), .Z(o[135]) );
  AND U3918 ( .A(n1035), .B(n3916), .Z(n3914) );
  XNOR U3919 ( .A(creg[135]), .B(n3915), .Z(n3916) );
  XNOR U3920 ( .A(n3917), .B(n3918), .Z(o[134]) );
  AND U3921 ( .A(n1035), .B(n3919), .Z(n3917) );
  XNOR U3922 ( .A(creg[134]), .B(n3918), .Z(n3919) );
  XNOR U3923 ( .A(n3920), .B(n3921), .Z(o[133]) );
  AND U3924 ( .A(n1035), .B(n3922), .Z(n3920) );
  XNOR U3925 ( .A(creg[133]), .B(n3921), .Z(n3922) );
  XNOR U3926 ( .A(n3923), .B(n3924), .Z(o[132]) );
  AND U3927 ( .A(n1035), .B(n3925), .Z(n3923) );
  XNOR U3928 ( .A(creg[132]), .B(n3924), .Z(n3925) );
  XNOR U3929 ( .A(n3926), .B(n3927), .Z(o[131]) );
  AND U3930 ( .A(n1035), .B(n3928), .Z(n3926) );
  XNOR U3931 ( .A(creg[131]), .B(n3927), .Z(n3928) );
  XNOR U3932 ( .A(n3929), .B(n3930), .Z(o[130]) );
  AND U3933 ( .A(n1035), .B(n3931), .Z(n3929) );
  XNOR U3934 ( .A(creg[130]), .B(n3930), .Z(n3931) );
  XNOR U3935 ( .A(n3932), .B(n3933), .Z(o[12]) );
  AND U3936 ( .A(n1035), .B(n3934), .Z(n3932) );
  XNOR U3937 ( .A(creg[12]), .B(n3933), .Z(n3934) );
  XNOR U3938 ( .A(n3935), .B(n3936), .Z(o[129]) );
  AND U3939 ( .A(n1035), .B(n3937), .Z(n3935) );
  XNOR U3940 ( .A(creg[129]), .B(n3936), .Z(n3937) );
  XNOR U3941 ( .A(n3938), .B(n3939), .Z(o[128]) );
  AND U3942 ( .A(n1035), .B(n3940), .Z(n3938) );
  XNOR U3943 ( .A(creg[128]), .B(n3939), .Z(n3940) );
  XNOR U3944 ( .A(n3941), .B(n3942), .Z(o[127]) );
  AND U3945 ( .A(n1035), .B(n3943), .Z(n3941) );
  XNOR U3946 ( .A(creg[127]), .B(n3942), .Z(n3943) );
  XNOR U3947 ( .A(n3944), .B(n3945), .Z(o[126]) );
  AND U3948 ( .A(n1035), .B(n3946), .Z(n3944) );
  XNOR U3949 ( .A(creg[126]), .B(n3945), .Z(n3946) );
  XNOR U3950 ( .A(n3947), .B(n3948), .Z(o[125]) );
  AND U3951 ( .A(n1035), .B(n3949), .Z(n3947) );
  XNOR U3952 ( .A(creg[125]), .B(n3948), .Z(n3949) );
  XNOR U3953 ( .A(n3950), .B(n3951), .Z(o[124]) );
  AND U3954 ( .A(n1035), .B(n3952), .Z(n3950) );
  XNOR U3955 ( .A(creg[124]), .B(n3951), .Z(n3952) );
  XNOR U3956 ( .A(n3953), .B(n3954), .Z(o[123]) );
  AND U3957 ( .A(n1035), .B(n3955), .Z(n3953) );
  XNOR U3958 ( .A(creg[123]), .B(n3954), .Z(n3955) );
  XNOR U3959 ( .A(n3956), .B(n3957), .Z(o[122]) );
  AND U3960 ( .A(n1035), .B(n3958), .Z(n3956) );
  XNOR U3961 ( .A(creg[122]), .B(n3957), .Z(n3958) );
  XNOR U3962 ( .A(n3959), .B(n3960), .Z(o[121]) );
  AND U3963 ( .A(n1035), .B(n3961), .Z(n3959) );
  XNOR U3964 ( .A(creg[121]), .B(n3960), .Z(n3961) );
  XNOR U3965 ( .A(n3962), .B(n3963), .Z(o[120]) );
  AND U3966 ( .A(n1035), .B(n3964), .Z(n3962) );
  XNOR U3967 ( .A(creg[120]), .B(n3963), .Z(n3964) );
  XNOR U3968 ( .A(n3965), .B(n3966), .Z(o[11]) );
  AND U3969 ( .A(n1035), .B(n3967), .Z(n3965) );
  XNOR U3970 ( .A(creg[11]), .B(n3966), .Z(n3967) );
  XNOR U3971 ( .A(n3968), .B(n3969), .Z(o[119]) );
  AND U3972 ( .A(n1035), .B(n3970), .Z(n3968) );
  XNOR U3973 ( .A(creg[119]), .B(n3969), .Z(n3970) );
  XNOR U3974 ( .A(n3971), .B(n3972), .Z(o[118]) );
  AND U3975 ( .A(n1035), .B(n3973), .Z(n3971) );
  XNOR U3976 ( .A(creg[118]), .B(n3972), .Z(n3973) );
  XNOR U3977 ( .A(n3974), .B(n3975), .Z(o[117]) );
  AND U3978 ( .A(n1035), .B(n3976), .Z(n3974) );
  XNOR U3979 ( .A(creg[117]), .B(n3975), .Z(n3976) );
  XNOR U3980 ( .A(n3977), .B(n3978), .Z(o[116]) );
  AND U3981 ( .A(n1035), .B(n3979), .Z(n3977) );
  XNOR U3982 ( .A(creg[116]), .B(n3978), .Z(n3979) );
  XNOR U3983 ( .A(n3980), .B(n3981), .Z(o[115]) );
  AND U3984 ( .A(n1035), .B(n3982), .Z(n3980) );
  XNOR U3985 ( .A(creg[115]), .B(n3981), .Z(n3982) );
  XNOR U3986 ( .A(n3983), .B(n3984), .Z(o[114]) );
  AND U3987 ( .A(n1035), .B(n3985), .Z(n3983) );
  XNOR U3988 ( .A(creg[114]), .B(n3984), .Z(n3985) );
  XNOR U3989 ( .A(n3986), .B(n3987), .Z(o[113]) );
  AND U3990 ( .A(n1035), .B(n3988), .Z(n3986) );
  XNOR U3991 ( .A(creg[113]), .B(n3987), .Z(n3988) );
  XNOR U3992 ( .A(n3989), .B(n3990), .Z(o[112]) );
  AND U3993 ( .A(n1035), .B(n3991), .Z(n3989) );
  XNOR U3994 ( .A(creg[112]), .B(n3990), .Z(n3991) );
  XNOR U3995 ( .A(n3992), .B(n3993), .Z(o[111]) );
  AND U3996 ( .A(n1035), .B(n3994), .Z(n3992) );
  XNOR U3997 ( .A(creg[111]), .B(n3993), .Z(n3994) );
  XNOR U3998 ( .A(n3995), .B(n3996), .Z(o[110]) );
  AND U3999 ( .A(n1035), .B(n3997), .Z(n3995) );
  XNOR U4000 ( .A(creg[110]), .B(n3996), .Z(n3997) );
  XNOR U4001 ( .A(n3998), .B(n3999), .Z(o[10]) );
  AND U4002 ( .A(n1035), .B(n4000), .Z(n3998) );
  XNOR U4003 ( .A(creg[10]), .B(n3999), .Z(n4000) );
  XNOR U4004 ( .A(n4001), .B(n4002), .Z(o[109]) );
  AND U4005 ( .A(n1035), .B(n4003), .Z(n4001) );
  XNOR U4006 ( .A(creg[109]), .B(n4002), .Z(n4003) );
  XNOR U4007 ( .A(n4004), .B(n4005), .Z(o[108]) );
  AND U4008 ( .A(n1035), .B(n4006), .Z(n4004) );
  XNOR U4009 ( .A(creg[108]), .B(n4005), .Z(n4006) );
  XNOR U4010 ( .A(n4007), .B(n4008), .Z(o[107]) );
  AND U4011 ( .A(n1035), .B(n4009), .Z(n4007) );
  XNOR U4012 ( .A(creg[107]), .B(n4008), .Z(n4009) );
  XNOR U4013 ( .A(n4010), .B(n4011), .Z(o[106]) );
  AND U4014 ( .A(n1035), .B(n4012), .Z(n4010) );
  XNOR U4015 ( .A(creg[106]), .B(n4011), .Z(n4012) );
  XNOR U4016 ( .A(n4013), .B(n4014), .Z(o[105]) );
  AND U4017 ( .A(n1035), .B(n4015), .Z(n4013) );
  XNOR U4018 ( .A(creg[105]), .B(n4014), .Z(n4015) );
  XNOR U4019 ( .A(n4016), .B(n4017), .Z(o[104]) );
  AND U4020 ( .A(n1035), .B(n4018), .Z(n4016) );
  XNOR U4021 ( .A(creg[104]), .B(n4017), .Z(n4018) );
  XNOR U4022 ( .A(n4019), .B(n4020), .Z(o[103]) );
  AND U4023 ( .A(n1035), .B(n4021), .Z(n4019) );
  XNOR U4024 ( .A(creg[103]), .B(n4020), .Z(n4021) );
  XNOR U4025 ( .A(n4022), .B(n4023), .Z(o[102]) );
  AND U4026 ( .A(n1035), .B(n4024), .Z(n4022) );
  XNOR U4027 ( .A(creg[102]), .B(n4023), .Z(n4024) );
  XNOR U4028 ( .A(n4025), .B(n4026), .Z(o[1023]) );
  AND U4029 ( .A(n1035), .B(n4027), .Z(n4025) );
  XNOR U4030 ( .A(creg[1023]), .B(n4026), .Z(n4027) );
  XNOR U4031 ( .A(n4028), .B(n4029), .Z(o[1022]) );
  AND U4032 ( .A(n1035), .B(n4030), .Z(n4028) );
  XNOR U4033 ( .A(creg[1022]), .B(n4029), .Z(n4030) );
  XNOR U4034 ( .A(n4031), .B(n4032), .Z(o[1021]) );
  AND U4035 ( .A(n1035), .B(n4033), .Z(n4031) );
  XNOR U4036 ( .A(creg[1021]), .B(n4032), .Z(n4033) );
  XNOR U4037 ( .A(n4034), .B(n4035), .Z(o[1020]) );
  AND U4038 ( .A(n1035), .B(n4036), .Z(n4034) );
  XNOR U4039 ( .A(creg[1020]), .B(n4035), .Z(n4036) );
  XNOR U4040 ( .A(n4037), .B(n4038), .Z(o[101]) );
  AND U4041 ( .A(n1035), .B(n4039), .Z(n4037) );
  XNOR U4042 ( .A(creg[101]), .B(n4038), .Z(n4039) );
  XNOR U4043 ( .A(n4040), .B(n4041), .Z(o[1019]) );
  AND U4044 ( .A(n1035), .B(n4042), .Z(n4040) );
  XNOR U4045 ( .A(creg[1019]), .B(n4041), .Z(n4042) );
  XNOR U4046 ( .A(n4043), .B(n4044), .Z(o[1018]) );
  AND U4047 ( .A(n1035), .B(n4045), .Z(n4043) );
  XNOR U4048 ( .A(creg[1018]), .B(n4044), .Z(n4045) );
  XNOR U4049 ( .A(n4046), .B(n4047), .Z(o[1017]) );
  AND U4050 ( .A(n1035), .B(n4048), .Z(n4046) );
  XNOR U4051 ( .A(creg[1017]), .B(n4047), .Z(n4048) );
  XNOR U4052 ( .A(n4049), .B(n4050), .Z(o[1016]) );
  AND U4053 ( .A(n1035), .B(n4051), .Z(n4049) );
  XNOR U4054 ( .A(creg[1016]), .B(n4050), .Z(n4051) );
  XNOR U4055 ( .A(n4052), .B(n4053), .Z(o[1015]) );
  AND U4056 ( .A(n1035), .B(n4054), .Z(n4052) );
  XNOR U4057 ( .A(creg[1015]), .B(n4053), .Z(n4054) );
  XNOR U4058 ( .A(n4055), .B(n4056), .Z(o[1014]) );
  AND U4059 ( .A(n1035), .B(n4057), .Z(n4055) );
  XNOR U4060 ( .A(creg[1014]), .B(n4056), .Z(n4057) );
  XNOR U4061 ( .A(n4058), .B(n4059), .Z(o[1013]) );
  AND U4062 ( .A(n1035), .B(n4060), .Z(n4058) );
  XNOR U4063 ( .A(creg[1013]), .B(n4059), .Z(n4060) );
  XNOR U4064 ( .A(n4061), .B(n4062), .Z(o[1012]) );
  AND U4065 ( .A(n1035), .B(n4063), .Z(n4061) );
  XNOR U4066 ( .A(creg[1012]), .B(n4062), .Z(n4063) );
  XNOR U4067 ( .A(n4064), .B(n4065), .Z(o[1011]) );
  AND U4068 ( .A(n1035), .B(n4066), .Z(n4064) );
  XNOR U4069 ( .A(creg[1011]), .B(n4065), .Z(n4066) );
  XNOR U4070 ( .A(n4067), .B(n4068), .Z(o[1010]) );
  AND U4071 ( .A(n1035), .B(n4069), .Z(n4067) );
  XNOR U4072 ( .A(creg[1010]), .B(n4068), .Z(n4069) );
  XNOR U4073 ( .A(n4070), .B(n4071), .Z(o[100]) );
  AND U4074 ( .A(n1035), .B(n4072), .Z(n4070) );
  XNOR U4075 ( .A(creg[100]), .B(n4071), .Z(n4072) );
  XNOR U4076 ( .A(n4073), .B(n4074), .Z(o[1009]) );
  AND U4077 ( .A(n1035), .B(n4075), .Z(n4073) );
  XNOR U4078 ( .A(creg[1009]), .B(n4074), .Z(n4075) );
  XNOR U4079 ( .A(n4076), .B(n4077), .Z(o[1008]) );
  AND U4080 ( .A(n1035), .B(n4078), .Z(n4076) );
  XNOR U4081 ( .A(creg[1008]), .B(n4077), .Z(n4078) );
  XNOR U4082 ( .A(n4079), .B(n4080), .Z(o[1007]) );
  AND U4083 ( .A(n1035), .B(n4081), .Z(n4079) );
  XNOR U4084 ( .A(creg[1007]), .B(n4080), .Z(n4081) );
  XNOR U4085 ( .A(n4082), .B(n4083), .Z(o[1006]) );
  AND U4086 ( .A(n1035), .B(n4084), .Z(n4082) );
  XNOR U4087 ( .A(creg[1006]), .B(n4083), .Z(n4084) );
  XNOR U4088 ( .A(n4085), .B(n4086), .Z(o[1005]) );
  AND U4089 ( .A(n1035), .B(n4087), .Z(n4085) );
  XNOR U4090 ( .A(creg[1005]), .B(n4086), .Z(n4087) );
  XNOR U4091 ( .A(n4088), .B(n4089), .Z(o[1004]) );
  AND U4092 ( .A(n1035), .B(n4090), .Z(n4088) );
  XNOR U4093 ( .A(creg[1004]), .B(n4089), .Z(n4090) );
  XNOR U4094 ( .A(n4091), .B(n4092), .Z(o[1003]) );
  AND U4095 ( .A(n1035), .B(n4093), .Z(n4091) );
  XNOR U4096 ( .A(creg[1003]), .B(n4092), .Z(n4093) );
  XNOR U4097 ( .A(n4094), .B(n4095), .Z(o[1002]) );
  AND U4098 ( .A(n1035), .B(n4096), .Z(n4094) );
  XNOR U4099 ( .A(creg[1002]), .B(n4095), .Z(n4096) );
  XNOR U4100 ( .A(n4097), .B(n4098), .Z(o[1001]) );
  AND U4101 ( .A(n1035), .B(n4099), .Z(n4097) );
  XNOR U4102 ( .A(creg[1001]), .B(n4098), .Z(n4099) );
  XNOR U4103 ( .A(n4100), .B(n4101), .Z(o[1000]) );
  AND U4104 ( .A(n1035), .B(n4102), .Z(n4100) );
  XNOR U4105 ( .A(creg[1000]), .B(n4101), .Z(n4102) );
  XOR U4106 ( .A(n4103), .B(n4104), .Z(o[0]) );
  AND U4107 ( .A(n1035), .B(n4105), .Z(n4103) );
  XOR U4108 ( .A(creg[0]), .B(n4104), .Z(n4105) );
  NAND U4109 ( .A(n4106), .B(n4107), .Z(n1035) );
  NANDN U4110 ( .B(mul_pow), .A(first_one), .Z(n4107) );
  NAND U4111 ( .A(first_one), .B(ein[1023]), .Z(n4106) );
  XOR U4112 ( .A(start_in[1023]), .B(mul_pow), .Z(n8) );
  NANDN U4113 ( .B(first_one), .A(n4108), .Z(n6) );
  NAND U4114 ( .A(n4109), .B(start_in[1023]), .Z(n4108) );
  AND U4115 ( .A(ein[1023]), .B(mul_pow), .Z(n4109) );
  ANDN U4116 ( .A(n4110), .B(n1050), .Z(\modmult_1/N999 ) );
  XOR U4117 ( .A(n4111), .B(n4112), .Z(n1050) );
  ANDN U4118 ( .A(n4110), .B(n1053), .Z(\modmult_1/N998 ) );
  XOR U4119 ( .A(n4113), .B(n4114), .Z(n1053) );
  ANDN U4120 ( .A(n4110), .B(n1056), .Z(\modmult_1/N997 ) );
  XOR U4121 ( .A(n4115), .B(n4116), .Z(n1056) );
  ANDN U4122 ( .A(n4110), .B(n1059), .Z(\modmult_1/N996 ) );
  XOR U4123 ( .A(n4117), .B(n4118), .Z(n1059) );
  ANDN U4124 ( .A(n4110), .B(n1062), .Z(\modmult_1/N995 ) );
  XOR U4125 ( .A(n4119), .B(n4120), .Z(n1062) );
  ANDN U4126 ( .A(n4110), .B(n1065), .Z(\modmult_1/N994 ) );
  XOR U4127 ( .A(n4121), .B(n4122), .Z(n1065) );
  ANDN U4128 ( .A(n4110), .B(n1068), .Z(\modmult_1/N993 ) );
  XOR U4129 ( .A(n4123), .B(n4124), .Z(n1068) );
  ANDN U4130 ( .A(n4110), .B(n1074), .Z(\modmult_1/N992 ) );
  XOR U4131 ( .A(n4125), .B(n4126), .Z(n1074) );
  ANDN U4132 ( .A(n4110), .B(n1077), .Z(\modmult_1/N991 ) );
  XOR U4133 ( .A(n4127), .B(n4128), .Z(n1077) );
  ANDN U4134 ( .A(n4110), .B(n1080), .Z(\modmult_1/N990 ) );
  XOR U4135 ( .A(n4129), .B(n4130), .Z(n1080) );
  ANDN U4136 ( .A(n4110), .B(n1137), .Z(\modmult_1/N99 ) );
  XOR U4137 ( .A(n4131), .B(n4132), .Z(n1137) );
  ANDN U4138 ( .A(n4110), .B(n1083), .Z(\modmult_1/N989 ) );
  XOR U4139 ( .A(n4133), .B(n4134), .Z(n1083) );
  ANDN U4140 ( .A(n4110), .B(n1086), .Z(\modmult_1/N988 ) );
  XOR U4141 ( .A(n4135), .B(n4136), .Z(n1086) );
  ANDN U4142 ( .A(n4110), .B(n1089), .Z(\modmult_1/N987 ) );
  XOR U4143 ( .A(n4137), .B(n4138), .Z(n1089) );
  ANDN U4144 ( .A(n4110), .B(n1092), .Z(\modmult_1/N986 ) );
  XOR U4145 ( .A(n4139), .B(n4140), .Z(n1092) );
  ANDN U4146 ( .A(n4110), .B(n1095), .Z(\modmult_1/N985 ) );
  XOR U4147 ( .A(n4141), .B(n4142), .Z(n1095) );
  ANDN U4148 ( .A(n4110), .B(n1098), .Z(\modmult_1/N984 ) );
  XOR U4149 ( .A(n4143), .B(n4144), .Z(n1098) );
  ANDN U4150 ( .A(n4110), .B(n1101), .Z(\modmult_1/N983 ) );
  XOR U4151 ( .A(n4145), .B(n4146), .Z(n1101) );
  ANDN U4152 ( .A(n4110), .B(n1107), .Z(\modmult_1/N982 ) );
  XOR U4153 ( .A(n4147), .B(n4148), .Z(n1107) );
  ANDN U4154 ( .A(n4110), .B(n1110), .Z(\modmult_1/N981 ) );
  XOR U4155 ( .A(n4149), .B(n4150), .Z(n1110) );
  ANDN U4156 ( .A(n4110), .B(n1113), .Z(\modmult_1/N980 ) );
  XOR U4157 ( .A(n4151), .B(n4152), .Z(n1113) );
  ANDN U4158 ( .A(n4110), .B(n1170), .Z(\modmult_1/N98 ) );
  XOR U4159 ( .A(n4153), .B(n4154), .Z(n1170) );
  ANDN U4160 ( .A(n4110), .B(n1116), .Z(\modmult_1/N979 ) );
  XOR U4161 ( .A(n4155), .B(n4156), .Z(n1116) );
  ANDN U4162 ( .A(n4110), .B(n1119), .Z(\modmult_1/N978 ) );
  XOR U4163 ( .A(n4157), .B(n4158), .Z(n1119) );
  ANDN U4164 ( .A(n4110), .B(n1122), .Z(\modmult_1/N977 ) );
  XOR U4165 ( .A(n4159), .B(n4160), .Z(n1122) );
  ANDN U4166 ( .A(n4110), .B(n1125), .Z(\modmult_1/N976 ) );
  XOR U4167 ( .A(n4161), .B(n4162), .Z(n1125) );
  ANDN U4168 ( .A(n4110), .B(n1128), .Z(\modmult_1/N975 ) );
  XOR U4169 ( .A(n4163), .B(n4164), .Z(n1128) );
  ANDN U4170 ( .A(n4110), .B(n1131), .Z(\modmult_1/N974 ) );
  XOR U4171 ( .A(n4165), .B(n4166), .Z(n1131) );
  ANDN U4172 ( .A(n4110), .B(n1134), .Z(\modmult_1/N973 ) );
  XOR U4173 ( .A(n4167), .B(n4168), .Z(n1134) );
  ANDN U4174 ( .A(n4110), .B(n1140), .Z(\modmult_1/N972 ) );
  XOR U4175 ( .A(n4169), .B(n4170), .Z(n1140) );
  ANDN U4176 ( .A(n4110), .B(n1143), .Z(\modmult_1/N971 ) );
  XOR U4177 ( .A(n4171), .B(n4172), .Z(n1143) );
  ANDN U4178 ( .A(n4110), .B(n1146), .Z(\modmult_1/N970 ) );
  XOR U4179 ( .A(n4173), .B(n4174), .Z(n1146) );
  ANDN U4180 ( .A(n4110), .B(n1203), .Z(\modmult_1/N97 ) );
  XOR U4181 ( .A(n4175), .B(n4176), .Z(n1203) );
  ANDN U4182 ( .A(n4110), .B(n1149), .Z(\modmult_1/N969 ) );
  XOR U4183 ( .A(n4177), .B(n4178), .Z(n1149) );
  ANDN U4184 ( .A(n4110), .B(n1152), .Z(\modmult_1/N968 ) );
  XOR U4185 ( .A(n4179), .B(n4180), .Z(n1152) );
  ANDN U4186 ( .A(n4110), .B(n1155), .Z(\modmult_1/N967 ) );
  XOR U4187 ( .A(n4181), .B(n4182), .Z(n1155) );
  ANDN U4188 ( .A(n4110), .B(n1158), .Z(\modmult_1/N966 ) );
  XOR U4189 ( .A(n4183), .B(n4184), .Z(n1158) );
  ANDN U4190 ( .A(n4110), .B(n1161), .Z(\modmult_1/N965 ) );
  XOR U4191 ( .A(n4185), .B(n4186), .Z(n1161) );
  ANDN U4192 ( .A(n4110), .B(n1164), .Z(\modmult_1/N964 ) );
  XOR U4193 ( .A(n4187), .B(n4188), .Z(n1164) );
  ANDN U4194 ( .A(n4110), .B(n1167), .Z(\modmult_1/N963 ) );
  XOR U4195 ( .A(n4189), .B(n4190), .Z(n1167) );
  ANDN U4196 ( .A(n4110), .B(n1173), .Z(\modmult_1/N962 ) );
  XOR U4197 ( .A(n4191), .B(n4192), .Z(n1173) );
  ANDN U4198 ( .A(n4110), .B(n1176), .Z(\modmult_1/N961 ) );
  XOR U4199 ( .A(n4193), .B(n4194), .Z(n1176) );
  ANDN U4200 ( .A(n4110), .B(n1179), .Z(\modmult_1/N960 ) );
  XOR U4201 ( .A(n4195), .B(n4196), .Z(n1179) );
  ANDN U4202 ( .A(n4110), .B(n1236), .Z(\modmult_1/N96 ) );
  XOR U4203 ( .A(n4197), .B(n4198), .Z(n1236) );
  ANDN U4204 ( .A(n4110), .B(n1182), .Z(\modmult_1/N959 ) );
  XOR U4205 ( .A(n4199), .B(n4200), .Z(n1182) );
  ANDN U4206 ( .A(n4110), .B(n1185), .Z(\modmult_1/N958 ) );
  XOR U4207 ( .A(n4201), .B(n4202), .Z(n1185) );
  ANDN U4208 ( .A(n4110), .B(n1188), .Z(\modmult_1/N957 ) );
  XOR U4209 ( .A(n4203), .B(n4204), .Z(n1188) );
  ANDN U4210 ( .A(n4110), .B(n1191), .Z(\modmult_1/N956 ) );
  XOR U4211 ( .A(n4205), .B(n4206), .Z(n1191) );
  ANDN U4212 ( .A(n4110), .B(n1194), .Z(\modmult_1/N955 ) );
  XOR U4213 ( .A(n4207), .B(n4208), .Z(n1194) );
  ANDN U4214 ( .A(n4110), .B(n1197), .Z(\modmult_1/N954 ) );
  XOR U4215 ( .A(n4209), .B(n4210), .Z(n1197) );
  ANDN U4216 ( .A(n4110), .B(n1200), .Z(\modmult_1/N953 ) );
  XOR U4217 ( .A(n4211), .B(n4212), .Z(n1200) );
  ANDN U4218 ( .A(n4110), .B(n1206), .Z(\modmult_1/N952 ) );
  XOR U4219 ( .A(n4213), .B(n4214), .Z(n1206) );
  ANDN U4220 ( .A(n4110), .B(n1209), .Z(\modmult_1/N951 ) );
  XOR U4221 ( .A(n4215), .B(n4216), .Z(n1209) );
  ANDN U4222 ( .A(n4110), .B(n1212), .Z(\modmult_1/N950 ) );
  XOR U4223 ( .A(n4217), .B(n4218), .Z(n1212) );
  ANDN U4224 ( .A(n4110), .B(n1269), .Z(\modmult_1/N95 ) );
  XOR U4225 ( .A(n4219), .B(n4220), .Z(n1269) );
  ANDN U4226 ( .A(n4110), .B(n1215), .Z(\modmult_1/N949 ) );
  XOR U4227 ( .A(n4221), .B(n4222), .Z(n1215) );
  ANDN U4228 ( .A(n4110), .B(n1218), .Z(\modmult_1/N948 ) );
  XOR U4229 ( .A(n4223), .B(n4224), .Z(n1218) );
  ANDN U4230 ( .A(n4110), .B(n1221), .Z(\modmult_1/N947 ) );
  XOR U4231 ( .A(n4225), .B(n4226), .Z(n1221) );
  ANDN U4232 ( .A(n4110), .B(n1224), .Z(\modmult_1/N946 ) );
  XOR U4233 ( .A(n4227), .B(n4228), .Z(n1224) );
  ANDN U4234 ( .A(n4110), .B(n1227), .Z(\modmult_1/N945 ) );
  XOR U4235 ( .A(n4229), .B(n4230), .Z(n1227) );
  ANDN U4236 ( .A(n4110), .B(n1230), .Z(\modmult_1/N944 ) );
  XOR U4237 ( .A(n4231), .B(n4232), .Z(n1230) );
  ANDN U4238 ( .A(n4110), .B(n1233), .Z(\modmult_1/N943 ) );
  XOR U4239 ( .A(n4233), .B(n4234), .Z(n1233) );
  ANDN U4240 ( .A(n4110), .B(n1239), .Z(\modmult_1/N942 ) );
  XOR U4241 ( .A(n4235), .B(n4236), .Z(n1239) );
  ANDN U4242 ( .A(n4110), .B(n1242), .Z(\modmult_1/N941 ) );
  XOR U4243 ( .A(n4237), .B(n4238), .Z(n1242) );
  ANDN U4244 ( .A(n4110), .B(n1245), .Z(\modmult_1/N940 ) );
  XOR U4245 ( .A(n4239), .B(n4240), .Z(n1245) );
  ANDN U4246 ( .A(n4110), .B(n1302), .Z(\modmult_1/N94 ) );
  XOR U4247 ( .A(n4241), .B(n4242), .Z(n1302) );
  ANDN U4248 ( .A(n4110), .B(n1248), .Z(\modmult_1/N939 ) );
  XOR U4249 ( .A(n4243), .B(n4244), .Z(n1248) );
  ANDN U4250 ( .A(n4110), .B(n1251), .Z(\modmult_1/N938 ) );
  XOR U4251 ( .A(n4245), .B(n4246), .Z(n1251) );
  ANDN U4252 ( .A(n4110), .B(n1254), .Z(\modmult_1/N937 ) );
  XOR U4253 ( .A(n4247), .B(n4248), .Z(n1254) );
  ANDN U4254 ( .A(n4110), .B(n1257), .Z(\modmult_1/N936 ) );
  XOR U4255 ( .A(n4249), .B(n4250), .Z(n1257) );
  ANDN U4256 ( .A(n4110), .B(n1260), .Z(\modmult_1/N935 ) );
  XOR U4257 ( .A(n4251), .B(n4252), .Z(n1260) );
  ANDN U4258 ( .A(n4110), .B(n1263), .Z(\modmult_1/N934 ) );
  XOR U4259 ( .A(n4253), .B(n4254), .Z(n1263) );
  ANDN U4260 ( .A(n4110), .B(n1266), .Z(\modmult_1/N933 ) );
  XOR U4261 ( .A(n4255), .B(n4256), .Z(n1266) );
  ANDN U4262 ( .A(n4110), .B(n1272), .Z(\modmult_1/N932 ) );
  XOR U4263 ( .A(n4257), .B(n4258), .Z(n1272) );
  ANDN U4264 ( .A(n4110), .B(n1275), .Z(\modmult_1/N931 ) );
  XOR U4265 ( .A(n4259), .B(n4260), .Z(n1275) );
  ANDN U4266 ( .A(n4110), .B(n1278), .Z(\modmult_1/N930 ) );
  XOR U4267 ( .A(n4261), .B(n4262), .Z(n1278) );
  ANDN U4268 ( .A(n4110), .B(n1335), .Z(\modmult_1/N93 ) );
  XOR U4269 ( .A(n4263), .B(n4264), .Z(n1335) );
  ANDN U4270 ( .A(n4110), .B(n1281), .Z(\modmult_1/N929 ) );
  XOR U4271 ( .A(n4265), .B(n4266), .Z(n1281) );
  ANDN U4272 ( .A(n4110), .B(n1284), .Z(\modmult_1/N928 ) );
  XOR U4273 ( .A(n4267), .B(n4268), .Z(n1284) );
  ANDN U4274 ( .A(n4110), .B(n1287), .Z(\modmult_1/N927 ) );
  XOR U4275 ( .A(n4269), .B(n4270), .Z(n1287) );
  ANDN U4276 ( .A(n4110), .B(n1290), .Z(\modmult_1/N926 ) );
  XOR U4277 ( .A(n4271), .B(n4272), .Z(n1290) );
  ANDN U4278 ( .A(n4110), .B(n1293), .Z(\modmult_1/N925 ) );
  XOR U4279 ( .A(n4273), .B(n4274), .Z(n1293) );
  ANDN U4280 ( .A(n4110), .B(n1296), .Z(\modmult_1/N924 ) );
  XOR U4281 ( .A(n4275), .B(n4276), .Z(n1296) );
  ANDN U4282 ( .A(n4110), .B(n1299), .Z(\modmult_1/N923 ) );
  XOR U4283 ( .A(n4277), .B(n4278), .Z(n1299) );
  ANDN U4284 ( .A(n4110), .B(n1305), .Z(\modmult_1/N922 ) );
  XOR U4285 ( .A(n4279), .B(n4280), .Z(n1305) );
  ANDN U4286 ( .A(n4110), .B(n1308), .Z(\modmult_1/N921 ) );
  XOR U4287 ( .A(n4281), .B(n4282), .Z(n1308) );
  ANDN U4288 ( .A(n4110), .B(n1311), .Z(\modmult_1/N920 ) );
  XOR U4289 ( .A(n4283), .B(n4284), .Z(n1311) );
  ANDN U4290 ( .A(n4110), .B(n1371), .Z(\modmult_1/N92 ) );
  XOR U4291 ( .A(n4285), .B(n4286), .Z(n1371) );
  ANDN U4292 ( .A(n4110), .B(n1314), .Z(\modmult_1/N919 ) );
  XOR U4293 ( .A(n4287), .B(n4288), .Z(n1314) );
  ANDN U4294 ( .A(n4110), .B(n1317), .Z(\modmult_1/N918 ) );
  XOR U4295 ( .A(n4289), .B(n4290), .Z(n1317) );
  ANDN U4296 ( .A(n4110), .B(n1320), .Z(\modmult_1/N917 ) );
  XOR U4297 ( .A(n4291), .B(n4292), .Z(n1320) );
  ANDN U4298 ( .A(n4110), .B(n1323), .Z(\modmult_1/N916 ) );
  XOR U4299 ( .A(n4293), .B(n4294), .Z(n1323) );
  ANDN U4300 ( .A(n4110), .B(n1326), .Z(\modmult_1/N915 ) );
  XOR U4301 ( .A(n4295), .B(n4296), .Z(n1326) );
  ANDN U4302 ( .A(n4110), .B(n1329), .Z(\modmult_1/N914 ) );
  XOR U4303 ( .A(n4297), .B(n4298), .Z(n1329) );
  ANDN U4304 ( .A(n4110), .B(n1332), .Z(\modmult_1/N913 ) );
  XOR U4305 ( .A(n4299), .B(n4300), .Z(n1332) );
  ANDN U4306 ( .A(n4110), .B(n1338), .Z(\modmult_1/N912 ) );
  XOR U4307 ( .A(n4301), .B(n4302), .Z(n1338) );
  ANDN U4308 ( .A(n4110), .B(n1341), .Z(\modmult_1/N911 ) );
  XOR U4309 ( .A(n4303), .B(n4304), .Z(n1341) );
  ANDN U4310 ( .A(n4110), .B(n1344), .Z(\modmult_1/N910 ) );
  XOR U4311 ( .A(n4305), .B(n4306), .Z(n1344) );
  ANDN U4312 ( .A(n4110), .B(n1404), .Z(\modmult_1/N91 ) );
  XOR U4313 ( .A(n4307), .B(n4308), .Z(n1404) );
  ANDN U4314 ( .A(n4110), .B(n1347), .Z(\modmult_1/N909 ) );
  XOR U4315 ( .A(n4309), .B(n4310), .Z(n1347) );
  ANDN U4316 ( .A(n4110), .B(n1350), .Z(\modmult_1/N908 ) );
  XOR U4317 ( .A(n4311), .B(n4312), .Z(n1350) );
  ANDN U4318 ( .A(n4110), .B(n1353), .Z(\modmult_1/N907 ) );
  XOR U4319 ( .A(n4313), .B(n4314), .Z(n1353) );
  ANDN U4320 ( .A(n4110), .B(n1356), .Z(\modmult_1/N906 ) );
  XOR U4321 ( .A(n4315), .B(n4316), .Z(n1356) );
  ANDN U4322 ( .A(n4110), .B(n1359), .Z(\modmult_1/N905 ) );
  XOR U4323 ( .A(n4317), .B(n4318), .Z(n1359) );
  ANDN U4324 ( .A(n4110), .B(n1362), .Z(\modmult_1/N904 ) );
  XOR U4325 ( .A(n4319), .B(n4320), .Z(n1362) );
  ANDN U4326 ( .A(n4110), .B(n1365), .Z(\modmult_1/N903 ) );
  XOR U4327 ( .A(n4321), .B(n4322), .Z(n1365) );
  ANDN U4328 ( .A(n4110), .B(n1374), .Z(\modmult_1/N902 ) );
  XOR U4329 ( .A(n4323), .B(n4324), .Z(n1374) );
  ANDN U4330 ( .A(n4110), .B(n1377), .Z(\modmult_1/N901 ) );
  XOR U4331 ( .A(n4325), .B(n4326), .Z(n1377) );
  ANDN U4332 ( .A(n4110), .B(n1380), .Z(\modmult_1/N900 ) );
  XOR U4333 ( .A(n4327), .B(n4328), .Z(n1380) );
  ANDN U4334 ( .A(n4110), .B(n1437), .Z(\modmult_1/N90 ) );
  XOR U4335 ( .A(n4329), .B(n4330), .Z(n1437) );
  ANDN U4336 ( .A(n4110), .B(n2034), .Z(\modmult_1/N9 ) );
  XOR U4337 ( .A(n4331), .B(n4332), .Z(n2034) );
  ANDN U4338 ( .A(n4110), .B(n1383), .Z(\modmult_1/N899 ) );
  XOR U4339 ( .A(n4333), .B(n4334), .Z(n1383) );
  ANDN U4340 ( .A(n4110), .B(n1386), .Z(\modmult_1/N898 ) );
  XOR U4341 ( .A(n4335), .B(n4336), .Z(n1386) );
  ANDN U4342 ( .A(n4110), .B(n1389), .Z(\modmult_1/N897 ) );
  XOR U4343 ( .A(n4337), .B(n4338), .Z(n1389) );
  ANDN U4344 ( .A(n4110), .B(n1392), .Z(\modmult_1/N896 ) );
  XOR U4345 ( .A(n4339), .B(n4340), .Z(n1392) );
  ANDN U4346 ( .A(n4110), .B(n1395), .Z(\modmult_1/N895 ) );
  XOR U4347 ( .A(n4341), .B(n4342), .Z(n1395) );
  ANDN U4348 ( .A(n4110), .B(n1398), .Z(\modmult_1/N894 ) );
  XOR U4349 ( .A(n4343), .B(n4344), .Z(n1398) );
  ANDN U4350 ( .A(n4110), .B(n1401), .Z(\modmult_1/N893 ) );
  XOR U4351 ( .A(n4345), .B(n4346), .Z(n1401) );
  ANDN U4352 ( .A(n4110), .B(n1407), .Z(\modmult_1/N892 ) );
  XOR U4353 ( .A(n4347), .B(n4348), .Z(n1407) );
  ANDN U4354 ( .A(n4110), .B(n1410), .Z(\modmult_1/N891 ) );
  XOR U4355 ( .A(n4349), .B(n4350), .Z(n1410) );
  ANDN U4356 ( .A(n4110), .B(n1413), .Z(\modmult_1/N890 ) );
  XOR U4357 ( .A(n4351), .B(n4352), .Z(n1413) );
  ANDN U4358 ( .A(n4110), .B(n1470), .Z(\modmult_1/N89 ) );
  XOR U4359 ( .A(n4353), .B(n4354), .Z(n1470) );
  ANDN U4360 ( .A(n4110), .B(n1416), .Z(\modmult_1/N889 ) );
  XOR U4361 ( .A(n4355), .B(n4356), .Z(n1416) );
  ANDN U4362 ( .A(n4110), .B(n1419), .Z(\modmult_1/N888 ) );
  XOR U4363 ( .A(n4357), .B(n4358), .Z(n1419) );
  ANDN U4364 ( .A(n4110), .B(n1422), .Z(\modmult_1/N887 ) );
  XOR U4365 ( .A(n4359), .B(n4360), .Z(n1422) );
  ANDN U4366 ( .A(n4110), .B(n1425), .Z(\modmult_1/N886 ) );
  XOR U4367 ( .A(n4361), .B(n4362), .Z(n1425) );
  ANDN U4368 ( .A(n4110), .B(n1428), .Z(\modmult_1/N885 ) );
  XOR U4369 ( .A(n4363), .B(n4364), .Z(n1428) );
  ANDN U4370 ( .A(n4110), .B(n1431), .Z(\modmult_1/N884 ) );
  XOR U4371 ( .A(n4365), .B(n4366), .Z(n1431) );
  ANDN U4372 ( .A(n4110), .B(n1434), .Z(\modmult_1/N883 ) );
  XOR U4373 ( .A(n4367), .B(n4368), .Z(n1434) );
  ANDN U4374 ( .A(n4110), .B(n1440), .Z(\modmult_1/N882 ) );
  XOR U4375 ( .A(n4369), .B(n4370), .Z(n1440) );
  ANDN U4376 ( .A(n4110), .B(n1443), .Z(\modmult_1/N881 ) );
  XOR U4377 ( .A(n4371), .B(n4372), .Z(n1443) );
  ANDN U4378 ( .A(n4110), .B(n1446), .Z(\modmult_1/N880 ) );
  XOR U4379 ( .A(n4373), .B(n4374), .Z(n1446) );
  ANDN U4380 ( .A(n4110), .B(n1503), .Z(\modmult_1/N88 ) );
  XOR U4381 ( .A(n4375), .B(n4376), .Z(n1503) );
  ANDN U4382 ( .A(n4110), .B(n1449), .Z(\modmult_1/N879 ) );
  XOR U4383 ( .A(n4377), .B(n4378), .Z(n1449) );
  ANDN U4384 ( .A(n4110), .B(n1452), .Z(\modmult_1/N878 ) );
  XOR U4385 ( .A(n4379), .B(n4380), .Z(n1452) );
  ANDN U4386 ( .A(n4110), .B(n1455), .Z(\modmult_1/N877 ) );
  XOR U4387 ( .A(n4381), .B(n4382), .Z(n1455) );
  ANDN U4388 ( .A(n4110), .B(n1458), .Z(\modmult_1/N876 ) );
  XOR U4389 ( .A(n4383), .B(n4384), .Z(n1458) );
  ANDN U4390 ( .A(n4110), .B(n1461), .Z(\modmult_1/N875 ) );
  XOR U4391 ( .A(n4385), .B(n4386), .Z(n1461) );
  ANDN U4392 ( .A(n4110), .B(n1464), .Z(\modmult_1/N874 ) );
  XOR U4393 ( .A(n4387), .B(n4388), .Z(n1464) );
  ANDN U4394 ( .A(n4110), .B(n1467), .Z(\modmult_1/N873 ) );
  XOR U4395 ( .A(n4389), .B(n4390), .Z(n1467) );
  ANDN U4396 ( .A(n4110), .B(n1473), .Z(\modmult_1/N872 ) );
  XOR U4397 ( .A(n4391), .B(n4392), .Z(n1473) );
  ANDN U4398 ( .A(n4110), .B(n1476), .Z(\modmult_1/N871 ) );
  XOR U4399 ( .A(n4393), .B(n4394), .Z(n1476) );
  ANDN U4400 ( .A(n4110), .B(n1479), .Z(\modmult_1/N870 ) );
  XOR U4401 ( .A(n4395), .B(n4396), .Z(n1479) );
  ANDN U4402 ( .A(n4110), .B(n1536), .Z(\modmult_1/N87 ) );
  XOR U4403 ( .A(n4397), .B(n4398), .Z(n1536) );
  ANDN U4404 ( .A(n4110), .B(n1482), .Z(\modmult_1/N869 ) );
  XOR U4405 ( .A(n4399), .B(n4400), .Z(n1482) );
  ANDN U4406 ( .A(n4110), .B(n1485), .Z(\modmult_1/N868 ) );
  XOR U4407 ( .A(n4401), .B(n4402), .Z(n1485) );
  ANDN U4408 ( .A(n4110), .B(n1488), .Z(\modmult_1/N867 ) );
  XOR U4409 ( .A(n4403), .B(n4404), .Z(n1488) );
  ANDN U4410 ( .A(n4110), .B(n1491), .Z(\modmult_1/N866 ) );
  XOR U4411 ( .A(n4405), .B(n4406), .Z(n1491) );
  ANDN U4412 ( .A(n4110), .B(n1494), .Z(\modmult_1/N865 ) );
  XOR U4413 ( .A(n4407), .B(n4408), .Z(n1494) );
  ANDN U4414 ( .A(n4110), .B(n1497), .Z(\modmult_1/N864 ) );
  XOR U4415 ( .A(n4409), .B(n4410), .Z(n1497) );
  ANDN U4416 ( .A(n4110), .B(n1500), .Z(\modmult_1/N863 ) );
  XOR U4417 ( .A(n4411), .B(n4412), .Z(n1500) );
  ANDN U4418 ( .A(n4110), .B(n1506), .Z(\modmult_1/N862 ) );
  XOR U4419 ( .A(n4413), .B(n4414), .Z(n1506) );
  ANDN U4420 ( .A(n4110), .B(n1509), .Z(\modmult_1/N861 ) );
  XOR U4421 ( .A(n4415), .B(n4416), .Z(n1509) );
  ANDN U4422 ( .A(n4110), .B(n1512), .Z(\modmult_1/N860 ) );
  XOR U4423 ( .A(n4417), .B(n4418), .Z(n1512) );
  ANDN U4424 ( .A(n4110), .B(n1569), .Z(\modmult_1/N86 ) );
  XOR U4425 ( .A(n4419), .B(n4420), .Z(n1569) );
  ANDN U4426 ( .A(n4110), .B(n1515), .Z(\modmult_1/N859 ) );
  XOR U4427 ( .A(n4421), .B(n4422), .Z(n1515) );
  ANDN U4428 ( .A(n4110), .B(n1518), .Z(\modmult_1/N858 ) );
  XOR U4429 ( .A(n4423), .B(n4424), .Z(n1518) );
  ANDN U4430 ( .A(n4110), .B(n1521), .Z(\modmult_1/N857 ) );
  XOR U4431 ( .A(n4425), .B(n4426), .Z(n1521) );
  ANDN U4432 ( .A(n4110), .B(n1524), .Z(\modmult_1/N856 ) );
  XOR U4433 ( .A(n4427), .B(n4428), .Z(n1524) );
  ANDN U4434 ( .A(n4110), .B(n1527), .Z(\modmult_1/N855 ) );
  XOR U4435 ( .A(n4429), .B(n4430), .Z(n1527) );
  ANDN U4436 ( .A(n4110), .B(n1530), .Z(\modmult_1/N854 ) );
  XOR U4437 ( .A(n4431), .B(n4432), .Z(n1530) );
  ANDN U4438 ( .A(n4110), .B(n1533), .Z(\modmult_1/N853 ) );
  XOR U4439 ( .A(n4433), .B(n4434), .Z(n1533) );
  ANDN U4440 ( .A(n4110), .B(n1539), .Z(\modmult_1/N852 ) );
  XOR U4441 ( .A(n4435), .B(n4436), .Z(n1539) );
  ANDN U4442 ( .A(n4110), .B(n1542), .Z(\modmult_1/N851 ) );
  XOR U4443 ( .A(n4437), .B(n4438), .Z(n1542) );
  ANDN U4444 ( .A(n4110), .B(n1545), .Z(\modmult_1/N850 ) );
  XOR U4445 ( .A(n4439), .B(n4440), .Z(n1545) );
  ANDN U4446 ( .A(n4110), .B(n1602), .Z(\modmult_1/N85 ) );
  XOR U4447 ( .A(n4441), .B(n4442), .Z(n1602) );
  ANDN U4448 ( .A(n4110), .B(n1548), .Z(\modmult_1/N849 ) );
  XOR U4449 ( .A(n4443), .B(n4444), .Z(n1548) );
  ANDN U4450 ( .A(n4110), .B(n1551), .Z(\modmult_1/N848 ) );
  XOR U4451 ( .A(n4445), .B(n4446), .Z(n1551) );
  ANDN U4452 ( .A(n4110), .B(n1554), .Z(\modmult_1/N847 ) );
  XOR U4453 ( .A(n4447), .B(n4448), .Z(n1554) );
  ANDN U4454 ( .A(n4110), .B(n1557), .Z(\modmult_1/N846 ) );
  XOR U4455 ( .A(n4449), .B(n4450), .Z(n1557) );
  ANDN U4456 ( .A(n4110), .B(n1560), .Z(\modmult_1/N845 ) );
  XOR U4457 ( .A(n4451), .B(n4452), .Z(n1560) );
  ANDN U4458 ( .A(n4110), .B(n1563), .Z(\modmult_1/N844 ) );
  XOR U4459 ( .A(n4453), .B(n4454), .Z(n1563) );
  ANDN U4460 ( .A(n4110), .B(n1566), .Z(\modmult_1/N843 ) );
  XOR U4461 ( .A(n4455), .B(n4456), .Z(n1566) );
  ANDN U4462 ( .A(n4110), .B(n1572), .Z(\modmult_1/N842 ) );
  XOR U4463 ( .A(n4457), .B(n4458), .Z(n1572) );
  ANDN U4464 ( .A(n4110), .B(n1575), .Z(\modmult_1/N841 ) );
  XOR U4465 ( .A(n4459), .B(n4460), .Z(n1575) );
  ANDN U4466 ( .A(n4110), .B(n1578), .Z(\modmult_1/N840 ) );
  XOR U4467 ( .A(n4461), .B(n4462), .Z(n1578) );
  ANDN U4468 ( .A(n4110), .B(n1635), .Z(\modmult_1/N84 ) );
  XOR U4469 ( .A(n4463), .B(n4464), .Z(n1635) );
  ANDN U4470 ( .A(n4110), .B(n1581), .Z(\modmult_1/N839 ) );
  XOR U4471 ( .A(n4465), .B(n4466), .Z(n1581) );
  ANDN U4472 ( .A(n4110), .B(n1584), .Z(\modmult_1/N838 ) );
  XOR U4473 ( .A(n4467), .B(n4468), .Z(n1584) );
  ANDN U4474 ( .A(n4110), .B(n1587), .Z(\modmult_1/N837 ) );
  XOR U4475 ( .A(n4469), .B(n4470), .Z(n1587) );
  ANDN U4476 ( .A(n4110), .B(n1590), .Z(\modmult_1/N836 ) );
  XOR U4477 ( .A(n4471), .B(n4472), .Z(n1590) );
  ANDN U4478 ( .A(n4110), .B(n1593), .Z(\modmult_1/N835 ) );
  XOR U4479 ( .A(n4473), .B(n4474), .Z(n1593) );
  ANDN U4480 ( .A(n4110), .B(n1596), .Z(\modmult_1/N834 ) );
  XOR U4481 ( .A(n4475), .B(n4476), .Z(n1596) );
  ANDN U4482 ( .A(n4110), .B(n1599), .Z(\modmult_1/N833 ) );
  XOR U4483 ( .A(n4477), .B(n4478), .Z(n1599) );
  ANDN U4484 ( .A(n4110), .B(n1605), .Z(\modmult_1/N832 ) );
  XOR U4485 ( .A(n4479), .B(n4480), .Z(n1605) );
  ANDN U4486 ( .A(n4110), .B(n1608), .Z(\modmult_1/N831 ) );
  XOR U4487 ( .A(n4481), .B(n4482), .Z(n1608) );
  ANDN U4488 ( .A(n4110), .B(n1611), .Z(\modmult_1/N830 ) );
  XOR U4489 ( .A(n4483), .B(n4484), .Z(n1611) );
  ANDN U4490 ( .A(n4110), .B(n1668), .Z(\modmult_1/N83 ) );
  XOR U4491 ( .A(n4485), .B(n4486), .Z(n1668) );
  ANDN U4492 ( .A(n4110), .B(n1614), .Z(\modmult_1/N829 ) );
  XOR U4493 ( .A(n4487), .B(n4488), .Z(n1614) );
  ANDN U4494 ( .A(n4110), .B(n1617), .Z(\modmult_1/N828 ) );
  XOR U4495 ( .A(n4489), .B(n4490), .Z(n1617) );
  ANDN U4496 ( .A(n4110), .B(n1620), .Z(\modmult_1/N827 ) );
  XOR U4497 ( .A(n4491), .B(n4492), .Z(n1620) );
  ANDN U4498 ( .A(n4110), .B(n1623), .Z(\modmult_1/N826 ) );
  XOR U4499 ( .A(n4493), .B(n4494), .Z(n1623) );
  ANDN U4500 ( .A(n4110), .B(n1626), .Z(\modmult_1/N825 ) );
  XOR U4501 ( .A(n4495), .B(n4496), .Z(n1626) );
  ANDN U4502 ( .A(n4110), .B(n1629), .Z(\modmult_1/N824 ) );
  XOR U4503 ( .A(n4497), .B(n4498), .Z(n1629) );
  ANDN U4504 ( .A(n4110), .B(n1632), .Z(\modmult_1/N823 ) );
  XOR U4505 ( .A(n4499), .B(n4500), .Z(n1632) );
  ANDN U4506 ( .A(n4110), .B(n1638), .Z(\modmult_1/N822 ) );
  XOR U4507 ( .A(n4501), .B(n4502), .Z(n1638) );
  ANDN U4508 ( .A(n4110), .B(n1641), .Z(\modmult_1/N821 ) );
  XOR U4509 ( .A(n4503), .B(n4504), .Z(n1641) );
  ANDN U4510 ( .A(n4110), .B(n1644), .Z(\modmult_1/N820 ) );
  XOR U4511 ( .A(n4505), .B(n4506), .Z(n1644) );
  ANDN U4512 ( .A(n4110), .B(n1704), .Z(\modmult_1/N82 ) );
  XOR U4513 ( .A(n4507), .B(n4508), .Z(n1704) );
  ANDN U4514 ( .A(n4110), .B(n1647), .Z(\modmult_1/N819 ) );
  XOR U4515 ( .A(n4509), .B(n4510), .Z(n1647) );
  ANDN U4516 ( .A(n4110), .B(n1650), .Z(\modmult_1/N818 ) );
  XOR U4517 ( .A(n4511), .B(n4512), .Z(n1650) );
  ANDN U4518 ( .A(n4110), .B(n1653), .Z(\modmult_1/N817 ) );
  XOR U4519 ( .A(n4513), .B(n4514), .Z(n1653) );
  ANDN U4520 ( .A(n4110), .B(n1656), .Z(\modmult_1/N816 ) );
  XOR U4521 ( .A(n4515), .B(n4516), .Z(n1656) );
  ANDN U4522 ( .A(n4110), .B(n1659), .Z(\modmult_1/N815 ) );
  XOR U4523 ( .A(n4517), .B(n4518), .Z(n1659) );
  ANDN U4524 ( .A(n4110), .B(n1662), .Z(\modmult_1/N814 ) );
  XOR U4525 ( .A(n4519), .B(n4520), .Z(n1662) );
  ANDN U4526 ( .A(n4110), .B(n1665), .Z(\modmult_1/N813 ) );
  XOR U4527 ( .A(n4521), .B(n4522), .Z(n1665) );
  ANDN U4528 ( .A(n4110), .B(n1671), .Z(\modmult_1/N812 ) );
  XOR U4529 ( .A(n4523), .B(n4524), .Z(n1671) );
  ANDN U4530 ( .A(n4110), .B(n1674), .Z(\modmult_1/N811 ) );
  XOR U4531 ( .A(n4525), .B(n4526), .Z(n1674) );
  ANDN U4532 ( .A(n4110), .B(n1677), .Z(\modmult_1/N810 ) );
  XOR U4533 ( .A(n4527), .B(n4528), .Z(n1677) );
  ANDN U4534 ( .A(n4110), .B(n1737), .Z(\modmult_1/N81 ) );
  XOR U4535 ( .A(n4529), .B(n4530), .Z(n1737) );
  ANDN U4536 ( .A(n4110), .B(n1680), .Z(\modmult_1/N809 ) );
  XOR U4537 ( .A(n4531), .B(n4532), .Z(n1680) );
  ANDN U4538 ( .A(n4110), .B(n1683), .Z(\modmult_1/N808 ) );
  XOR U4539 ( .A(n4533), .B(n4534), .Z(n1683) );
  ANDN U4540 ( .A(n4110), .B(n1686), .Z(\modmult_1/N807 ) );
  XOR U4541 ( .A(n4535), .B(n4536), .Z(n1686) );
  ANDN U4542 ( .A(n4110), .B(n1689), .Z(\modmult_1/N806 ) );
  XOR U4543 ( .A(n4537), .B(n4538), .Z(n1689) );
  ANDN U4544 ( .A(n4110), .B(n1692), .Z(\modmult_1/N805 ) );
  XOR U4545 ( .A(n4539), .B(n4540), .Z(n1692) );
  ANDN U4546 ( .A(n4110), .B(n1695), .Z(\modmult_1/N804 ) );
  XOR U4547 ( .A(n4541), .B(n4542), .Z(n1695) );
  ANDN U4548 ( .A(n4110), .B(n1698), .Z(\modmult_1/N803 ) );
  XOR U4549 ( .A(n4543), .B(n4544), .Z(n1698) );
  ANDN U4550 ( .A(n4110), .B(n1707), .Z(\modmult_1/N802 ) );
  XOR U4551 ( .A(n4545), .B(n4546), .Z(n1707) );
  ANDN U4552 ( .A(n4110), .B(n1710), .Z(\modmult_1/N801 ) );
  XOR U4553 ( .A(n4547), .B(n4548), .Z(n1710) );
  ANDN U4554 ( .A(n4110), .B(n1713), .Z(\modmult_1/N800 ) );
  XOR U4555 ( .A(n4549), .B(n4550), .Z(n1713) );
  ANDN U4556 ( .A(n4110), .B(n1770), .Z(\modmult_1/N80 ) );
  XOR U4557 ( .A(n4551), .B(n4552), .Z(n1770) );
  ANDN U4558 ( .A(n4110), .B(n2367), .Z(\modmult_1/N8 ) );
  XOR U4559 ( .A(n4553), .B(n4554), .Z(n2367) );
  ANDN U4560 ( .A(n4110), .B(n1716), .Z(\modmult_1/N799 ) );
  XOR U4561 ( .A(n4555), .B(n4556), .Z(n1716) );
  ANDN U4562 ( .A(n4110), .B(n1719), .Z(\modmult_1/N798 ) );
  XOR U4563 ( .A(n4557), .B(n4558), .Z(n1719) );
  ANDN U4564 ( .A(n4110), .B(n1722), .Z(\modmult_1/N797 ) );
  XOR U4565 ( .A(n4559), .B(n4560), .Z(n1722) );
  ANDN U4566 ( .A(n4110), .B(n1725), .Z(\modmult_1/N796 ) );
  XOR U4567 ( .A(n4561), .B(n4562), .Z(n1725) );
  ANDN U4568 ( .A(n4110), .B(n1728), .Z(\modmult_1/N795 ) );
  XOR U4569 ( .A(n4563), .B(n4564), .Z(n1728) );
  ANDN U4570 ( .A(n4110), .B(n1731), .Z(\modmult_1/N794 ) );
  XOR U4571 ( .A(n4565), .B(n4566), .Z(n1731) );
  ANDN U4572 ( .A(n4110), .B(n1734), .Z(\modmult_1/N793 ) );
  XOR U4573 ( .A(n4567), .B(n4568), .Z(n1734) );
  ANDN U4574 ( .A(n4110), .B(n1740), .Z(\modmult_1/N792 ) );
  XOR U4575 ( .A(n4569), .B(n4570), .Z(n1740) );
  ANDN U4576 ( .A(n4110), .B(n1743), .Z(\modmult_1/N791 ) );
  XOR U4577 ( .A(n4571), .B(n4572), .Z(n1743) );
  ANDN U4578 ( .A(n4110), .B(n1746), .Z(\modmult_1/N790 ) );
  XOR U4579 ( .A(n4573), .B(n4574), .Z(n1746) );
  ANDN U4580 ( .A(n4110), .B(n1803), .Z(\modmult_1/N79 ) );
  XOR U4581 ( .A(n4575), .B(n4576), .Z(n1803) );
  ANDN U4582 ( .A(n4110), .B(n1749), .Z(\modmult_1/N789 ) );
  XOR U4583 ( .A(n4577), .B(n4578), .Z(n1749) );
  ANDN U4584 ( .A(n4110), .B(n1752), .Z(\modmult_1/N788 ) );
  XOR U4585 ( .A(n4579), .B(n4580), .Z(n1752) );
  ANDN U4586 ( .A(n4110), .B(n1755), .Z(\modmult_1/N787 ) );
  XOR U4587 ( .A(n4581), .B(n4582), .Z(n1755) );
  ANDN U4588 ( .A(n4110), .B(n1758), .Z(\modmult_1/N786 ) );
  XOR U4589 ( .A(n4583), .B(n4584), .Z(n1758) );
  ANDN U4590 ( .A(n4110), .B(n1761), .Z(\modmult_1/N785 ) );
  XOR U4591 ( .A(n4585), .B(n4586), .Z(n1761) );
  ANDN U4592 ( .A(n4110), .B(n1764), .Z(\modmult_1/N784 ) );
  XOR U4593 ( .A(n4587), .B(n4588), .Z(n1764) );
  ANDN U4594 ( .A(n4110), .B(n1767), .Z(\modmult_1/N783 ) );
  XOR U4595 ( .A(n4589), .B(n4590), .Z(n1767) );
  ANDN U4596 ( .A(n4110), .B(n1773), .Z(\modmult_1/N782 ) );
  XOR U4597 ( .A(n4591), .B(n4592), .Z(n1773) );
  ANDN U4598 ( .A(n4110), .B(n1776), .Z(\modmult_1/N781 ) );
  XOR U4599 ( .A(n4593), .B(n4594), .Z(n1776) );
  ANDN U4600 ( .A(n4110), .B(n1779), .Z(\modmult_1/N780 ) );
  XOR U4601 ( .A(n4595), .B(n4596), .Z(n1779) );
  ANDN U4602 ( .A(n4110), .B(n1836), .Z(\modmult_1/N78 ) );
  XOR U4603 ( .A(n4597), .B(n4598), .Z(n1836) );
  ANDN U4604 ( .A(n4110), .B(n1782), .Z(\modmult_1/N779 ) );
  XOR U4605 ( .A(n4599), .B(n4600), .Z(n1782) );
  ANDN U4606 ( .A(n4110), .B(n1785), .Z(\modmult_1/N778 ) );
  XOR U4607 ( .A(n4601), .B(n4602), .Z(n1785) );
  ANDN U4608 ( .A(n4110), .B(n1788), .Z(\modmult_1/N777 ) );
  XOR U4609 ( .A(n4603), .B(n4604), .Z(n1788) );
  ANDN U4610 ( .A(n4110), .B(n1791), .Z(\modmult_1/N776 ) );
  XOR U4611 ( .A(n4605), .B(n4606), .Z(n1791) );
  ANDN U4612 ( .A(n4110), .B(n1794), .Z(\modmult_1/N775 ) );
  XOR U4613 ( .A(n4607), .B(n4608), .Z(n1794) );
  ANDN U4614 ( .A(n4110), .B(n1797), .Z(\modmult_1/N774 ) );
  XOR U4615 ( .A(n4609), .B(n4610), .Z(n1797) );
  ANDN U4616 ( .A(n4110), .B(n1800), .Z(\modmult_1/N773 ) );
  XOR U4617 ( .A(n4611), .B(n4612), .Z(n1800) );
  ANDN U4618 ( .A(n4110), .B(n1806), .Z(\modmult_1/N772 ) );
  XOR U4619 ( .A(n4613), .B(n4614), .Z(n1806) );
  ANDN U4620 ( .A(n4110), .B(n1809), .Z(\modmult_1/N771 ) );
  XOR U4621 ( .A(n4615), .B(n4616), .Z(n1809) );
  ANDN U4622 ( .A(n4110), .B(n1812), .Z(\modmult_1/N770 ) );
  XOR U4623 ( .A(n4617), .B(n4618), .Z(n1812) );
  ANDN U4624 ( .A(n4110), .B(n1869), .Z(\modmult_1/N77 ) );
  XOR U4625 ( .A(n4619), .B(n4620), .Z(n1869) );
  ANDN U4626 ( .A(n4110), .B(n1815), .Z(\modmult_1/N769 ) );
  XOR U4627 ( .A(n4621), .B(n4622), .Z(n1815) );
  ANDN U4628 ( .A(n4110), .B(n1818), .Z(\modmult_1/N768 ) );
  XOR U4629 ( .A(n4623), .B(n4624), .Z(n1818) );
  ANDN U4630 ( .A(n4110), .B(n1821), .Z(\modmult_1/N767 ) );
  XOR U4631 ( .A(n4625), .B(n4626), .Z(n1821) );
  ANDN U4632 ( .A(n4110), .B(n1824), .Z(\modmult_1/N766 ) );
  XOR U4633 ( .A(n4627), .B(n4628), .Z(n1824) );
  ANDN U4634 ( .A(n4110), .B(n1827), .Z(\modmult_1/N765 ) );
  XOR U4635 ( .A(n4629), .B(n4630), .Z(n1827) );
  ANDN U4636 ( .A(n4110), .B(n1830), .Z(\modmult_1/N764 ) );
  XOR U4637 ( .A(n4631), .B(n4632), .Z(n1830) );
  ANDN U4638 ( .A(n4110), .B(n1833), .Z(\modmult_1/N763 ) );
  XOR U4639 ( .A(n4633), .B(n4634), .Z(n1833) );
  ANDN U4640 ( .A(n4110), .B(n1839), .Z(\modmult_1/N762 ) );
  XOR U4641 ( .A(n4635), .B(n4636), .Z(n1839) );
  ANDN U4642 ( .A(n4110), .B(n1842), .Z(\modmult_1/N761 ) );
  XOR U4643 ( .A(n4637), .B(n4638), .Z(n1842) );
  ANDN U4644 ( .A(n4110), .B(n1845), .Z(\modmult_1/N760 ) );
  XOR U4645 ( .A(n4639), .B(n4640), .Z(n1845) );
  ANDN U4646 ( .A(n4110), .B(n1902), .Z(\modmult_1/N76 ) );
  XOR U4647 ( .A(n4641), .B(n4642), .Z(n1902) );
  ANDN U4648 ( .A(n4110), .B(n1848), .Z(\modmult_1/N759 ) );
  XOR U4649 ( .A(n4643), .B(n4644), .Z(n1848) );
  ANDN U4650 ( .A(n4110), .B(n1851), .Z(\modmult_1/N758 ) );
  XOR U4651 ( .A(n4645), .B(n4646), .Z(n1851) );
  ANDN U4652 ( .A(n4110), .B(n1854), .Z(\modmult_1/N757 ) );
  XOR U4653 ( .A(n4647), .B(n4648), .Z(n1854) );
  ANDN U4654 ( .A(n4110), .B(n1857), .Z(\modmult_1/N756 ) );
  XOR U4655 ( .A(n4649), .B(n4650), .Z(n1857) );
  ANDN U4656 ( .A(n4110), .B(n1860), .Z(\modmult_1/N755 ) );
  XOR U4657 ( .A(n4651), .B(n4652), .Z(n1860) );
  ANDN U4658 ( .A(n4110), .B(n1863), .Z(\modmult_1/N754 ) );
  XOR U4659 ( .A(n4653), .B(n4654), .Z(n1863) );
  ANDN U4660 ( .A(n4110), .B(n1866), .Z(\modmult_1/N753 ) );
  XOR U4661 ( .A(n4655), .B(n4656), .Z(n1866) );
  ANDN U4662 ( .A(n4110), .B(n1872), .Z(\modmult_1/N752 ) );
  XOR U4663 ( .A(n4657), .B(n4658), .Z(n1872) );
  ANDN U4664 ( .A(n4110), .B(n1875), .Z(\modmult_1/N751 ) );
  XOR U4665 ( .A(n4659), .B(n4660), .Z(n1875) );
  ANDN U4666 ( .A(n4110), .B(n1878), .Z(\modmult_1/N750 ) );
  XOR U4667 ( .A(n4661), .B(n4662), .Z(n1878) );
  ANDN U4668 ( .A(n4110), .B(n1935), .Z(\modmult_1/N75 ) );
  XOR U4669 ( .A(n4663), .B(n4664), .Z(n1935) );
  ANDN U4670 ( .A(n4110), .B(n1881), .Z(\modmult_1/N749 ) );
  XOR U4671 ( .A(n4665), .B(n4666), .Z(n1881) );
  ANDN U4672 ( .A(n4110), .B(n1884), .Z(\modmult_1/N748 ) );
  XOR U4673 ( .A(n4667), .B(n4668), .Z(n1884) );
  ANDN U4674 ( .A(n4110), .B(n1887), .Z(\modmult_1/N747 ) );
  XOR U4675 ( .A(n4669), .B(n4670), .Z(n1887) );
  ANDN U4676 ( .A(n4110), .B(n1890), .Z(\modmult_1/N746 ) );
  XOR U4677 ( .A(n4671), .B(n4672), .Z(n1890) );
  ANDN U4678 ( .A(n4110), .B(n1893), .Z(\modmult_1/N745 ) );
  XOR U4679 ( .A(n4673), .B(n4674), .Z(n1893) );
  ANDN U4680 ( .A(n4110), .B(n1896), .Z(\modmult_1/N744 ) );
  XOR U4681 ( .A(n4675), .B(n4676), .Z(n1896) );
  ANDN U4682 ( .A(n4110), .B(n1899), .Z(\modmult_1/N743 ) );
  XOR U4683 ( .A(n4677), .B(n4678), .Z(n1899) );
  ANDN U4684 ( .A(n4110), .B(n1905), .Z(\modmult_1/N742 ) );
  XOR U4685 ( .A(n4679), .B(n4680), .Z(n1905) );
  ANDN U4686 ( .A(n4110), .B(n1908), .Z(\modmult_1/N741 ) );
  XOR U4687 ( .A(n4681), .B(n4682), .Z(n1908) );
  ANDN U4688 ( .A(n4110), .B(n1911), .Z(\modmult_1/N740 ) );
  XOR U4689 ( .A(n4683), .B(n4684), .Z(n1911) );
  ANDN U4690 ( .A(n4110), .B(n1968), .Z(\modmult_1/N74 ) );
  XOR U4691 ( .A(n4685), .B(n4686), .Z(n1968) );
  ANDN U4692 ( .A(n4110), .B(n1914), .Z(\modmult_1/N739 ) );
  XOR U4693 ( .A(n4687), .B(n4688), .Z(n1914) );
  ANDN U4694 ( .A(n4110), .B(n1917), .Z(\modmult_1/N738 ) );
  XOR U4695 ( .A(n4689), .B(n4690), .Z(n1917) );
  ANDN U4696 ( .A(n4110), .B(n1920), .Z(\modmult_1/N737 ) );
  XOR U4697 ( .A(n4691), .B(n4692), .Z(n1920) );
  ANDN U4698 ( .A(n4110), .B(n1923), .Z(\modmult_1/N736 ) );
  XOR U4699 ( .A(n4693), .B(n4694), .Z(n1923) );
  ANDN U4700 ( .A(n4110), .B(n1926), .Z(\modmult_1/N735 ) );
  XOR U4701 ( .A(n4695), .B(n4696), .Z(n1926) );
  ANDN U4702 ( .A(n4110), .B(n1929), .Z(\modmult_1/N734 ) );
  XOR U4703 ( .A(n4697), .B(n4698), .Z(n1929) );
  ANDN U4704 ( .A(n4110), .B(n1932), .Z(\modmult_1/N733 ) );
  XOR U4705 ( .A(n4699), .B(n4700), .Z(n1932) );
  ANDN U4706 ( .A(n4110), .B(n1938), .Z(\modmult_1/N732 ) );
  XOR U4707 ( .A(n4701), .B(n4702), .Z(n1938) );
  ANDN U4708 ( .A(n4110), .B(n1941), .Z(\modmult_1/N731 ) );
  XOR U4709 ( .A(n4703), .B(n4704), .Z(n1941) );
  ANDN U4710 ( .A(n4110), .B(n1944), .Z(\modmult_1/N730 ) );
  XOR U4711 ( .A(n4705), .B(n4706), .Z(n1944) );
  ANDN U4712 ( .A(n4110), .B(n2001), .Z(\modmult_1/N73 ) );
  XOR U4713 ( .A(n4707), .B(n4708), .Z(n2001) );
  ANDN U4714 ( .A(n4110), .B(n1947), .Z(\modmult_1/N729 ) );
  XOR U4715 ( .A(n4709), .B(n4710), .Z(n1947) );
  ANDN U4716 ( .A(n4110), .B(n1950), .Z(\modmult_1/N728 ) );
  XOR U4717 ( .A(n4711), .B(n4712), .Z(n1950) );
  ANDN U4718 ( .A(n4110), .B(n1953), .Z(\modmult_1/N727 ) );
  XOR U4719 ( .A(n4713), .B(n4714), .Z(n1953) );
  ANDN U4720 ( .A(n4110), .B(n1956), .Z(\modmult_1/N726 ) );
  XOR U4721 ( .A(n4715), .B(n4716), .Z(n1956) );
  ANDN U4722 ( .A(n4110), .B(n1959), .Z(\modmult_1/N725 ) );
  XOR U4723 ( .A(n4717), .B(n4718), .Z(n1959) );
  ANDN U4724 ( .A(n4110), .B(n1962), .Z(\modmult_1/N724 ) );
  XOR U4725 ( .A(n4719), .B(n4720), .Z(n1962) );
  ANDN U4726 ( .A(n4110), .B(n1965), .Z(\modmult_1/N723 ) );
  XOR U4727 ( .A(n4721), .B(n4722), .Z(n1965) );
  ANDN U4728 ( .A(n4110), .B(n1971), .Z(\modmult_1/N722 ) );
  XOR U4729 ( .A(n4723), .B(n4724), .Z(n1971) );
  ANDN U4730 ( .A(n4110), .B(n1974), .Z(\modmult_1/N721 ) );
  XOR U4731 ( .A(n4725), .B(n4726), .Z(n1974) );
  ANDN U4732 ( .A(n4110), .B(n1977), .Z(\modmult_1/N720 ) );
  XOR U4733 ( .A(n4727), .B(n4728), .Z(n1977) );
  ANDN U4734 ( .A(n4110), .B(n2037), .Z(\modmult_1/N72 ) );
  XOR U4735 ( .A(n4729), .B(n4730), .Z(n2037) );
  ANDN U4736 ( .A(n4110), .B(n1980), .Z(\modmult_1/N719 ) );
  XOR U4737 ( .A(n4731), .B(n4732), .Z(n1980) );
  ANDN U4738 ( .A(n4110), .B(n1983), .Z(\modmult_1/N718 ) );
  XOR U4739 ( .A(n4733), .B(n4734), .Z(n1983) );
  ANDN U4740 ( .A(n4110), .B(n1986), .Z(\modmult_1/N717 ) );
  XOR U4741 ( .A(n4735), .B(n4736), .Z(n1986) );
  ANDN U4742 ( .A(n4110), .B(n1989), .Z(\modmult_1/N716 ) );
  XOR U4743 ( .A(n4737), .B(n4738), .Z(n1989) );
  ANDN U4744 ( .A(n4110), .B(n1992), .Z(\modmult_1/N715 ) );
  XOR U4745 ( .A(n4739), .B(n4740), .Z(n1992) );
  ANDN U4746 ( .A(n4110), .B(n1995), .Z(\modmult_1/N714 ) );
  XOR U4747 ( .A(n4741), .B(n4742), .Z(n1995) );
  ANDN U4748 ( .A(n4110), .B(n1998), .Z(\modmult_1/N713 ) );
  XOR U4749 ( .A(n4743), .B(n4744), .Z(n1998) );
  ANDN U4750 ( .A(n4110), .B(n2004), .Z(\modmult_1/N712 ) );
  XOR U4751 ( .A(n4745), .B(n4746), .Z(n2004) );
  ANDN U4752 ( .A(n4110), .B(n2007), .Z(\modmult_1/N711 ) );
  XOR U4753 ( .A(n4747), .B(n4748), .Z(n2007) );
  ANDN U4754 ( .A(n4110), .B(n2010), .Z(\modmult_1/N710 ) );
  XOR U4755 ( .A(n4749), .B(n4750), .Z(n2010) );
  ANDN U4756 ( .A(n4110), .B(n2070), .Z(\modmult_1/N71 ) );
  XOR U4757 ( .A(n4751), .B(n4752), .Z(n2070) );
  ANDN U4758 ( .A(n4110), .B(n2013), .Z(\modmult_1/N709 ) );
  XOR U4759 ( .A(n4753), .B(n4754), .Z(n2013) );
  ANDN U4760 ( .A(n4110), .B(n2016), .Z(\modmult_1/N708 ) );
  XOR U4761 ( .A(n4755), .B(n4756), .Z(n2016) );
  ANDN U4762 ( .A(n4110), .B(n2019), .Z(\modmult_1/N707 ) );
  XOR U4763 ( .A(n4757), .B(n4758), .Z(n2019) );
  ANDN U4764 ( .A(n4110), .B(n2022), .Z(\modmult_1/N706 ) );
  XOR U4765 ( .A(n4759), .B(n4760), .Z(n2022) );
  ANDN U4766 ( .A(n4110), .B(n2025), .Z(\modmult_1/N705 ) );
  XOR U4767 ( .A(n4761), .B(n4762), .Z(n2025) );
  ANDN U4768 ( .A(n4110), .B(n2028), .Z(\modmult_1/N704 ) );
  XOR U4769 ( .A(n4763), .B(n4764), .Z(n2028) );
  ANDN U4770 ( .A(n4110), .B(n2031), .Z(\modmult_1/N703 ) );
  XOR U4771 ( .A(n4765), .B(n4766), .Z(n2031) );
  ANDN U4772 ( .A(n4110), .B(n2040), .Z(\modmult_1/N702 ) );
  XOR U4773 ( .A(n4767), .B(n4768), .Z(n2040) );
  ANDN U4774 ( .A(n4110), .B(n2043), .Z(\modmult_1/N701 ) );
  XOR U4775 ( .A(n4769), .B(n4770), .Z(n2043) );
  ANDN U4776 ( .A(n4110), .B(n2046), .Z(\modmult_1/N700 ) );
  XOR U4777 ( .A(n4771), .B(n4772), .Z(n2046) );
  ANDN U4778 ( .A(n4110), .B(n2103), .Z(\modmult_1/N70 ) );
  XOR U4779 ( .A(n4773), .B(n4774), .Z(n2103) );
  ANDN U4780 ( .A(n4110), .B(n2700), .Z(\modmult_1/N7 ) );
  XOR U4781 ( .A(n4775), .B(n4776), .Z(n2700) );
  ANDN U4782 ( .A(n4110), .B(n2049), .Z(\modmult_1/N699 ) );
  XOR U4783 ( .A(n4777), .B(n4778), .Z(n2049) );
  ANDN U4784 ( .A(n4110), .B(n2052), .Z(\modmult_1/N698 ) );
  XOR U4785 ( .A(n4779), .B(n4780), .Z(n2052) );
  ANDN U4786 ( .A(n4110), .B(n2055), .Z(\modmult_1/N697 ) );
  XOR U4787 ( .A(n4781), .B(n4782), .Z(n2055) );
  ANDN U4788 ( .A(n4110), .B(n2058), .Z(\modmult_1/N696 ) );
  XOR U4789 ( .A(n4783), .B(n4784), .Z(n2058) );
  ANDN U4790 ( .A(n4110), .B(n2061), .Z(\modmult_1/N695 ) );
  XOR U4791 ( .A(n4785), .B(n4786), .Z(n2061) );
  ANDN U4792 ( .A(n4110), .B(n2064), .Z(\modmult_1/N694 ) );
  XOR U4793 ( .A(n4787), .B(n4788), .Z(n2064) );
  ANDN U4794 ( .A(n4110), .B(n2067), .Z(\modmult_1/N693 ) );
  XOR U4795 ( .A(n4789), .B(n4790), .Z(n2067) );
  ANDN U4796 ( .A(n4110), .B(n2073), .Z(\modmult_1/N692 ) );
  XOR U4797 ( .A(n4791), .B(n4792), .Z(n2073) );
  ANDN U4798 ( .A(n4110), .B(n2076), .Z(\modmult_1/N691 ) );
  XOR U4799 ( .A(n4793), .B(n4794), .Z(n2076) );
  ANDN U4800 ( .A(n4110), .B(n2079), .Z(\modmult_1/N690 ) );
  XOR U4801 ( .A(n4795), .B(n4796), .Z(n2079) );
  ANDN U4802 ( .A(n4110), .B(n2136), .Z(\modmult_1/N69 ) );
  XOR U4803 ( .A(n4797), .B(n4798), .Z(n2136) );
  ANDN U4804 ( .A(n4110), .B(n2082), .Z(\modmult_1/N689 ) );
  XOR U4805 ( .A(n4799), .B(n4800), .Z(n2082) );
  ANDN U4806 ( .A(n4110), .B(n2085), .Z(\modmult_1/N688 ) );
  XOR U4807 ( .A(n4801), .B(n4802), .Z(n2085) );
  ANDN U4808 ( .A(n4110), .B(n2088), .Z(\modmult_1/N687 ) );
  XOR U4809 ( .A(n4803), .B(n4804), .Z(n2088) );
  ANDN U4810 ( .A(n4110), .B(n2091), .Z(\modmult_1/N686 ) );
  XOR U4811 ( .A(n4805), .B(n4806), .Z(n2091) );
  ANDN U4812 ( .A(n4110), .B(n2094), .Z(\modmult_1/N685 ) );
  XOR U4813 ( .A(n4807), .B(n4808), .Z(n2094) );
  ANDN U4814 ( .A(n4110), .B(n2097), .Z(\modmult_1/N684 ) );
  XOR U4815 ( .A(n4809), .B(n4810), .Z(n2097) );
  ANDN U4816 ( .A(n4110), .B(n2100), .Z(\modmult_1/N683 ) );
  XOR U4817 ( .A(n4811), .B(n4812), .Z(n2100) );
  ANDN U4818 ( .A(n4110), .B(n2106), .Z(\modmult_1/N682 ) );
  XOR U4819 ( .A(n4813), .B(n4814), .Z(n2106) );
  ANDN U4820 ( .A(n4110), .B(n2109), .Z(\modmult_1/N681 ) );
  XOR U4821 ( .A(n4815), .B(n4816), .Z(n2109) );
  ANDN U4822 ( .A(n4110), .B(n2112), .Z(\modmult_1/N680 ) );
  XOR U4823 ( .A(n4817), .B(n4818), .Z(n2112) );
  ANDN U4824 ( .A(n4110), .B(n2169), .Z(\modmult_1/N68 ) );
  XOR U4825 ( .A(n4819), .B(n4820), .Z(n2169) );
  ANDN U4826 ( .A(n4110), .B(n2115), .Z(\modmult_1/N679 ) );
  XOR U4827 ( .A(n4821), .B(n4822), .Z(n2115) );
  ANDN U4828 ( .A(n4110), .B(n2118), .Z(\modmult_1/N678 ) );
  XOR U4829 ( .A(n4823), .B(n4824), .Z(n2118) );
  ANDN U4830 ( .A(n4110), .B(n2121), .Z(\modmult_1/N677 ) );
  XOR U4831 ( .A(n4825), .B(n4826), .Z(n2121) );
  ANDN U4832 ( .A(n4110), .B(n2124), .Z(\modmult_1/N676 ) );
  XOR U4833 ( .A(n4827), .B(n4828), .Z(n2124) );
  ANDN U4834 ( .A(n4110), .B(n2127), .Z(\modmult_1/N675 ) );
  XOR U4835 ( .A(n4829), .B(n4830), .Z(n2127) );
  ANDN U4836 ( .A(n4110), .B(n2130), .Z(\modmult_1/N674 ) );
  XOR U4837 ( .A(n4831), .B(n4832), .Z(n2130) );
  ANDN U4838 ( .A(n4110), .B(n2133), .Z(\modmult_1/N673 ) );
  XOR U4839 ( .A(n4833), .B(n4834), .Z(n2133) );
  ANDN U4840 ( .A(n4110), .B(n2139), .Z(\modmult_1/N672 ) );
  XOR U4841 ( .A(n4835), .B(n4836), .Z(n2139) );
  ANDN U4842 ( .A(n4110), .B(n2142), .Z(\modmult_1/N671 ) );
  XOR U4843 ( .A(n4837), .B(n4838), .Z(n2142) );
  ANDN U4844 ( .A(n4110), .B(n2145), .Z(\modmult_1/N670 ) );
  XOR U4845 ( .A(n4839), .B(n4840), .Z(n2145) );
  ANDN U4846 ( .A(n4110), .B(n2202), .Z(\modmult_1/N67 ) );
  XOR U4847 ( .A(n4841), .B(n4842), .Z(n2202) );
  ANDN U4848 ( .A(n4110), .B(n2148), .Z(\modmult_1/N669 ) );
  XOR U4849 ( .A(n4843), .B(n4844), .Z(n2148) );
  ANDN U4850 ( .A(n4110), .B(n2151), .Z(\modmult_1/N668 ) );
  XOR U4851 ( .A(n4845), .B(n4846), .Z(n2151) );
  ANDN U4852 ( .A(n4110), .B(n2154), .Z(\modmult_1/N667 ) );
  XOR U4853 ( .A(n4847), .B(n4848), .Z(n2154) );
  ANDN U4854 ( .A(n4110), .B(n2157), .Z(\modmult_1/N666 ) );
  XOR U4855 ( .A(n4849), .B(n4850), .Z(n2157) );
  ANDN U4856 ( .A(n4110), .B(n2160), .Z(\modmult_1/N665 ) );
  XOR U4857 ( .A(n4851), .B(n4852), .Z(n2160) );
  ANDN U4858 ( .A(n4110), .B(n2163), .Z(\modmult_1/N664 ) );
  XOR U4859 ( .A(n4853), .B(n4854), .Z(n2163) );
  ANDN U4860 ( .A(n4110), .B(n2166), .Z(\modmult_1/N663 ) );
  XOR U4861 ( .A(n4855), .B(n4856), .Z(n2166) );
  ANDN U4862 ( .A(n4110), .B(n2172), .Z(\modmult_1/N662 ) );
  XOR U4863 ( .A(n4857), .B(n4858), .Z(n2172) );
  ANDN U4864 ( .A(n4110), .B(n2175), .Z(\modmult_1/N661 ) );
  XOR U4865 ( .A(n4859), .B(n4860), .Z(n2175) );
  ANDN U4866 ( .A(n4110), .B(n2178), .Z(\modmult_1/N660 ) );
  XOR U4867 ( .A(n4861), .B(n4862), .Z(n2178) );
  ANDN U4868 ( .A(n4110), .B(n2235), .Z(\modmult_1/N66 ) );
  XOR U4869 ( .A(n4863), .B(n4864), .Z(n2235) );
  ANDN U4870 ( .A(n4110), .B(n2181), .Z(\modmult_1/N659 ) );
  XOR U4871 ( .A(n4865), .B(n4866), .Z(n2181) );
  ANDN U4872 ( .A(n4110), .B(n2184), .Z(\modmult_1/N658 ) );
  XOR U4873 ( .A(n4867), .B(n4868), .Z(n2184) );
  ANDN U4874 ( .A(n4110), .B(n2187), .Z(\modmult_1/N657 ) );
  XOR U4875 ( .A(n4869), .B(n4870), .Z(n2187) );
  ANDN U4876 ( .A(n4110), .B(n2190), .Z(\modmult_1/N656 ) );
  XOR U4877 ( .A(n4871), .B(n4872), .Z(n2190) );
  ANDN U4878 ( .A(n4110), .B(n2193), .Z(\modmult_1/N655 ) );
  XOR U4879 ( .A(n4873), .B(n4874), .Z(n2193) );
  ANDN U4880 ( .A(n4110), .B(n2196), .Z(\modmult_1/N654 ) );
  XOR U4881 ( .A(n4875), .B(n4876), .Z(n2196) );
  ANDN U4882 ( .A(n4110), .B(n2199), .Z(\modmult_1/N653 ) );
  XOR U4883 ( .A(n4877), .B(n4878), .Z(n2199) );
  ANDN U4884 ( .A(n4110), .B(n2205), .Z(\modmult_1/N652 ) );
  XOR U4885 ( .A(n4879), .B(n4880), .Z(n2205) );
  ANDN U4886 ( .A(n4110), .B(n2208), .Z(\modmult_1/N651 ) );
  XOR U4887 ( .A(n4881), .B(n4882), .Z(n2208) );
  ANDN U4888 ( .A(n4110), .B(n2211), .Z(\modmult_1/N650 ) );
  XOR U4889 ( .A(n4883), .B(n4884), .Z(n2211) );
  ANDN U4890 ( .A(n4110), .B(n2268), .Z(\modmult_1/N65 ) );
  XOR U4891 ( .A(n4885), .B(n4886), .Z(n2268) );
  ANDN U4892 ( .A(n4110), .B(n2214), .Z(\modmult_1/N649 ) );
  XOR U4893 ( .A(n4887), .B(n4888), .Z(n2214) );
  ANDN U4894 ( .A(n4110), .B(n2217), .Z(\modmult_1/N648 ) );
  XOR U4895 ( .A(n4889), .B(n4890), .Z(n2217) );
  ANDN U4896 ( .A(n4110), .B(n2220), .Z(\modmult_1/N647 ) );
  XOR U4897 ( .A(n4891), .B(n4892), .Z(n2220) );
  ANDN U4898 ( .A(n4110), .B(n2223), .Z(\modmult_1/N646 ) );
  XOR U4899 ( .A(n4893), .B(n4894), .Z(n2223) );
  ANDN U4900 ( .A(n4110), .B(n2226), .Z(\modmult_1/N645 ) );
  XOR U4901 ( .A(n4895), .B(n4896), .Z(n2226) );
  ANDN U4902 ( .A(n4110), .B(n2229), .Z(\modmult_1/N644 ) );
  XOR U4903 ( .A(n4897), .B(n4898), .Z(n2229) );
  ANDN U4904 ( .A(n4110), .B(n2232), .Z(\modmult_1/N643 ) );
  XOR U4905 ( .A(n4899), .B(n4900), .Z(n2232) );
  ANDN U4906 ( .A(n4110), .B(n2238), .Z(\modmult_1/N642 ) );
  XOR U4907 ( .A(n4901), .B(n4902), .Z(n2238) );
  ANDN U4908 ( .A(n4110), .B(n2241), .Z(\modmult_1/N641 ) );
  XOR U4909 ( .A(n4903), .B(n4904), .Z(n2241) );
  ANDN U4910 ( .A(n4110), .B(n2244), .Z(\modmult_1/N640 ) );
  XOR U4911 ( .A(n4905), .B(n4906), .Z(n2244) );
  ANDN U4912 ( .A(n4110), .B(n2301), .Z(\modmult_1/N64 ) );
  XOR U4913 ( .A(n4907), .B(n4908), .Z(n2301) );
  ANDN U4914 ( .A(n4110), .B(n2247), .Z(\modmult_1/N639 ) );
  XOR U4915 ( .A(n4909), .B(n4910), .Z(n2247) );
  ANDN U4916 ( .A(n4110), .B(n2250), .Z(\modmult_1/N638 ) );
  XOR U4917 ( .A(n4911), .B(n4912), .Z(n2250) );
  ANDN U4918 ( .A(n4110), .B(n2253), .Z(\modmult_1/N637 ) );
  XOR U4919 ( .A(n4913), .B(n4914), .Z(n2253) );
  ANDN U4920 ( .A(n4110), .B(n2256), .Z(\modmult_1/N636 ) );
  XOR U4921 ( .A(n4915), .B(n4916), .Z(n2256) );
  ANDN U4922 ( .A(n4110), .B(n2259), .Z(\modmult_1/N635 ) );
  XOR U4923 ( .A(n4917), .B(n4918), .Z(n2259) );
  ANDN U4924 ( .A(n4110), .B(n2262), .Z(\modmult_1/N634 ) );
  XOR U4925 ( .A(n4919), .B(n4920), .Z(n2262) );
  ANDN U4926 ( .A(n4110), .B(n2265), .Z(\modmult_1/N633 ) );
  XOR U4927 ( .A(n4921), .B(n4922), .Z(n2265) );
  ANDN U4928 ( .A(n4110), .B(n2271), .Z(\modmult_1/N632 ) );
  XOR U4929 ( .A(n4923), .B(n4924), .Z(n2271) );
  ANDN U4930 ( .A(n4110), .B(n2274), .Z(\modmult_1/N631 ) );
  XOR U4931 ( .A(n4925), .B(n4926), .Z(n2274) );
  ANDN U4932 ( .A(n4110), .B(n2277), .Z(\modmult_1/N630 ) );
  XOR U4933 ( .A(n4927), .B(n4928), .Z(n2277) );
  ANDN U4934 ( .A(n4110), .B(n2334), .Z(\modmult_1/N63 ) );
  XOR U4935 ( .A(n4929), .B(n4930), .Z(n2334) );
  ANDN U4936 ( .A(n4110), .B(n2280), .Z(\modmult_1/N629 ) );
  XOR U4937 ( .A(n4931), .B(n4932), .Z(n2280) );
  ANDN U4938 ( .A(n4110), .B(n2283), .Z(\modmult_1/N628 ) );
  XOR U4939 ( .A(n4933), .B(n4934), .Z(n2283) );
  ANDN U4940 ( .A(n4110), .B(n2286), .Z(\modmult_1/N627 ) );
  XOR U4941 ( .A(n4935), .B(n4936), .Z(n2286) );
  ANDN U4942 ( .A(n4110), .B(n2289), .Z(\modmult_1/N626 ) );
  XOR U4943 ( .A(n4937), .B(n4938), .Z(n2289) );
  ANDN U4944 ( .A(n4110), .B(n2292), .Z(\modmult_1/N625 ) );
  XOR U4945 ( .A(n4939), .B(n4940), .Z(n2292) );
  ANDN U4946 ( .A(n4110), .B(n2295), .Z(\modmult_1/N624 ) );
  XOR U4947 ( .A(n4941), .B(n4942), .Z(n2295) );
  ANDN U4948 ( .A(n4110), .B(n2298), .Z(\modmult_1/N623 ) );
  XOR U4949 ( .A(n4943), .B(n4944), .Z(n2298) );
  ANDN U4950 ( .A(n4110), .B(n2304), .Z(\modmult_1/N622 ) );
  XOR U4951 ( .A(n4945), .B(n4946), .Z(n2304) );
  ANDN U4952 ( .A(n4110), .B(n2307), .Z(\modmult_1/N621 ) );
  XOR U4953 ( .A(n4947), .B(n4948), .Z(n2307) );
  ANDN U4954 ( .A(n4110), .B(n2310), .Z(\modmult_1/N620 ) );
  XOR U4955 ( .A(n4949), .B(n4950), .Z(n2310) );
  ANDN U4956 ( .A(n4110), .B(n2370), .Z(\modmult_1/N62 ) );
  XOR U4957 ( .A(n4951), .B(n4952), .Z(n2370) );
  ANDN U4958 ( .A(n4110), .B(n2313), .Z(\modmult_1/N619 ) );
  XOR U4959 ( .A(n4953), .B(n4954), .Z(n2313) );
  ANDN U4960 ( .A(n4110), .B(n2316), .Z(\modmult_1/N618 ) );
  XOR U4961 ( .A(n4955), .B(n4956), .Z(n2316) );
  ANDN U4962 ( .A(n4110), .B(n2319), .Z(\modmult_1/N617 ) );
  XOR U4963 ( .A(n4957), .B(n4958), .Z(n2319) );
  ANDN U4964 ( .A(n4110), .B(n2322), .Z(\modmult_1/N616 ) );
  XOR U4965 ( .A(n4959), .B(n4960), .Z(n2322) );
  ANDN U4966 ( .A(n4110), .B(n2325), .Z(\modmult_1/N615 ) );
  XOR U4967 ( .A(n4961), .B(n4962), .Z(n2325) );
  ANDN U4968 ( .A(n4110), .B(n2328), .Z(\modmult_1/N614 ) );
  XOR U4969 ( .A(n4963), .B(n4964), .Z(n2328) );
  ANDN U4970 ( .A(n4110), .B(n2331), .Z(\modmult_1/N613 ) );
  XOR U4971 ( .A(n4965), .B(n4966), .Z(n2331) );
  ANDN U4972 ( .A(n4110), .B(n2337), .Z(\modmult_1/N612 ) );
  XOR U4973 ( .A(n4967), .B(n4968), .Z(n2337) );
  ANDN U4974 ( .A(n4110), .B(n2340), .Z(\modmult_1/N611 ) );
  XOR U4975 ( .A(n4969), .B(n4970), .Z(n2340) );
  ANDN U4976 ( .A(n4110), .B(n2343), .Z(\modmult_1/N610 ) );
  XOR U4977 ( .A(n4971), .B(n4972), .Z(n2343) );
  ANDN U4978 ( .A(n4110), .B(n2403), .Z(\modmult_1/N61 ) );
  XOR U4979 ( .A(n4973), .B(n4974), .Z(n2403) );
  ANDN U4980 ( .A(n4110), .B(n2346), .Z(\modmult_1/N609 ) );
  XOR U4981 ( .A(n4975), .B(n4976), .Z(n2346) );
  ANDN U4982 ( .A(n4110), .B(n2349), .Z(\modmult_1/N608 ) );
  XOR U4983 ( .A(n4977), .B(n4978), .Z(n2349) );
  ANDN U4984 ( .A(n4110), .B(n2352), .Z(\modmult_1/N607 ) );
  XOR U4985 ( .A(n4979), .B(n4980), .Z(n2352) );
  ANDN U4986 ( .A(n4110), .B(n2355), .Z(\modmult_1/N606 ) );
  XOR U4987 ( .A(n4981), .B(n4982), .Z(n2355) );
  ANDN U4988 ( .A(n4110), .B(n2358), .Z(\modmult_1/N605 ) );
  XOR U4989 ( .A(n4983), .B(n4984), .Z(n2358) );
  ANDN U4990 ( .A(n4110), .B(n2361), .Z(\modmult_1/N604 ) );
  XOR U4991 ( .A(n4985), .B(n4986), .Z(n2361) );
  ANDN U4992 ( .A(n4110), .B(n2364), .Z(\modmult_1/N603 ) );
  XOR U4993 ( .A(n4987), .B(n4988), .Z(n2364) );
  ANDN U4994 ( .A(n4110), .B(n2373), .Z(\modmult_1/N602 ) );
  XOR U4995 ( .A(n4989), .B(n4990), .Z(n2373) );
  ANDN U4996 ( .A(n4110), .B(n2376), .Z(\modmult_1/N601 ) );
  XOR U4997 ( .A(n4991), .B(n4992), .Z(n2376) );
  ANDN U4998 ( .A(n4110), .B(n2379), .Z(\modmult_1/N600 ) );
  XOR U4999 ( .A(n4993), .B(n4994), .Z(n2379) );
  ANDN U5000 ( .A(n4110), .B(n2436), .Z(\modmult_1/N60 ) );
  XOR U5001 ( .A(n4995), .B(n4996), .Z(n2436) );
  ANDN U5002 ( .A(n4110), .B(n3033), .Z(\modmult_1/N6 ) );
  XOR U5003 ( .A(n4997), .B(n4998), .Z(n3033) );
  ANDN U5004 ( .A(n4110), .B(n2382), .Z(\modmult_1/N599 ) );
  XOR U5005 ( .A(n4999), .B(n5000), .Z(n2382) );
  ANDN U5006 ( .A(n4110), .B(n2385), .Z(\modmult_1/N598 ) );
  XOR U5007 ( .A(n5001), .B(n5002), .Z(n2385) );
  ANDN U5008 ( .A(n4110), .B(n2388), .Z(\modmult_1/N597 ) );
  XOR U5009 ( .A(n5003), .B(n5004), .Z(n2388) );
  ANDN U5010 ( .A(n4110), .B(n2391), .Z(\modmult_1/N596 ) );
  XOR U5011 ( .A(n5005), .B(n5006), .Z(n2391) );
  ANDN U5012 ( .A(n4110), .B(n2394), .Z(\modmult_1/N595 ) );
  XOR U5013 ( .A(n5007), .B(n5008), .Z(n2394) );
  ANDN U5014 ( .A(n4110), .B(n2397), .Z(\modmult_1/N594 ) );
  XOR U5015 ( .A(n5009), .B(n5010), .Z(n2397) );
  ANDN U5016 ( .A(n4110), .B(n2400), .Z(\modmult_1/N593 ) );
  XOR U5017 ( .A(n5011), .B(n5012), .Z(n2400) );
  ANDN U5018 ( .A(n4110), .B(n2406), .Z(\modmult_1/N592 ) );
  XOR U5019 ( .A(n5013), .B(n5014), .Z(n2406) );
  ANDN U5020 ( .A(n4110), .B(n2409), .Z(\modmult_1/N591 ) );
  XOR U5021 ( .A(n5015), .B(n5016), .Z(n2409) );
  ANDN U5022 ( .A(n4110), .B(n2412), .Z(\modmult_1/N590 ) );
  XOR U5023 ( .A(n5017), .B(n5018), .Z(n2412) );
  ANDN U5024 ( .A(n4110), .B(n2469), .Z(\modmult_1/N59 ) );
  XOR U5025 ( .A(n5019), .B(n5020), .Z(n2469) );
  ANDN U5026 ( .A(n4110), .B(n2415), .Z(\modmult_1/N589 ) );
  XOR U5027 ( .A(n5021), .B(n5022), .Z(n2415) );
  ANDN U5028 ( .A(n4110), .B(n2418), .Z(\modmult_1/N588 ) );
  XOR U5029 ( .A(n5023), .B(n5024), .Z(n2418) );
  ANDN U5030 ( .A(n4110), .B(n2421), .Z(\modmult_1/N587 ) );
  XOR U5031 ( .A(n5025), .B(n5026), .Z(n2421) );
  ANDN U5032 ( .A(n4110), .B(n2424), .Z(\modmult_1/N586 ) );
  XOR U5033 ( .A(n5027), .B(n5028), .Z(n2424) );
  ANDN U5034 ( .A(n4110), .B(n2427), .Z(\modmult_1/N585 ) );
  XOR U5035 ( .A(n5029), .B(n5030), .Z(n2427) );
  ANDN U5036 ( .A(n4110), .B(n2430), .Z(\modmult_1/N584 ) );
  XOR U5037 ( .A(n5031), .B(n5032), .Z(n2430) );
  ANDN U5038 ( .A(n4110), .B(n2433), .Z(\modmult_1/N583 ) );
  XOR U5039 ( .A(n5033), .B(n5034), .Z(n2433) );
  ANDN U5040 ( .A(n4110), .B(n2439), .Z(\modmult_1/N582 ) );
  XOR U5041 ( .A(n5035), .B(n5036), .Z(n2439) );
  ANDN U5042 ( .A(n4110), .B(n2442), .Z(\modmult_1/N581 ) );
  XOR U5043 ( .A(n5037), .B(n5038), .Z(n2442) );
  ANDN U5044 ( .A(n4110), .B(n2445), .Z(\modmult_1/N580 ) );
  XOR U5045 ( .A(n5039), .B(n5040), .Z(n2445) );
  ANDN U5046 ( .A(n4110), .B(n2502), .Z(\modmult_1/N58 ) );
  XOR U5047 ( .A(n5041), .B(n5042), .Z(n2502) );
  ANDN U5048 ( .A(n4110), .B(n2448), .Z(\modmult_1/N579 ) );
  XOR U5049 ( .A(n5043), .B(n5044), .Z(n2448) );
  ANDN U5050 ( .A(n4110), .B(n2451), .Z(\modmult_1/N578 ) );
  XOR U5051 ( .A(n5045), .B(n5046), .Z(n2451) );
  ANDN U5052 ( .A(n4110), .B(n2454), .Z(\modmult_1/N577 ) );
  XOR U5053 ( .A(n5047), .B(n5048), .Z(n2454) );
  ANDN U5054 ( .A(n4110), .B(n2457), .Z(\modmult_1/N576 ) );
  XOR U5055 ( .A(n5049), .B(n5050), .Z(n2457) );
  ANDN U5056 ( .A(n4110), .B(n2460), .Z(\modmult_1/N575 ) );
  XOR U5057 ( .A(n5051), .B(n5052), .Z(n2460) );
  ANDN U5058 ( .A(n4110), .B(n2463), .Z(\modmult_1/N574 ) );
  XOR U5059 ( .A(n5053), .B(n5054), .Z(n2463) );
  ANDN U5060 ( .A(n4110), .B(n2466), .Z(\modmult_1/N573 ) );
  XOR U5061 ( .A(n5055), .B(n5056), .Z(n2466) );
  ANDN U5062 ( .A(n4110), .B(n2472), .Z(\modmult_1/N572 ) );
  XOR U5063 ( .A(n5057), .B(n5058), .Z(n2472) );
  ANDN U5064 ( .A(n4110), .B(n2475), .Z(\modmult_1/N571 ) );
  XOR U5065 ( .A(n5059), .B(n5060), .Z(n2475) );
  ANDN U5066 ( .A(n4110), .B(n2478), .Z(\modmult_1/N570 ) );
  XOR U5067 ( .A(n5061), .B(n5062), .Z(n2478) );
  ANDN U5068 ( .A(n4110), .B(n2535), .Z(\modmult_1/N57 ) );
  XOR U5069 ( .A(n5063), .B(n5064), .Z(n2535) );
  ANDN U5070 ( .A(n4110), .B(n2481), .Z(\modmult_1/N569 ) );
  XOR U5071 ( .A(n5065), .B(n5066), .Z(n2481) );
  ANDN U5072 ( .A(n4110), .B(n2484), .Z(\modmult_1/N568 ) );
  XOR U5073 ( .A(n5067), .B(n5068), .Z(n2484) );
  ANDN U5074 ( .A(n4110), .B(n2487), .Z(\modmult_1/N567 ) );
  XOR U5075 ( .A(n5069), .B(n5070), .Z(n2487) );
  ANDN U5076 ( .A(n4110), .B(n2490), .Z(\modmult_1/N566 ) );
  XOR U5077 ( .A(n5071), .B(n5072), .Z(n2490) );
  ANDN U5078 ( .A(n4110), .B(n2493), .Z(\modmult_1/N565 ) );
  XOR U5079 ( .A(n5073), .B(n5074), .Z(n2493) );
  ANDN U5080 ( .A(n4110), .B(n2496), .Z(\modmult_1/N564 ) );
  XOR U5081 ( .A(n5075), .B(n5076), .Z(n2496) );
  ANDN U5082 ( .A(n4110), .B(n2499), .Z(\modmult_1/N563 ) );
  XOR U5083 ( .A(n5077), .B(n5078), .Z(n2499) );
  ANDN U5084 ( .A(n4110), .B(n2505), .Z(\modmult_1/N562 ) );
  XOR U5085 ( .A(n5079), .B(n5080), .Z(n2505) );
  ANDN U5086 ( .A(n4110), .B(n2508), .Z(\modmult_1/N561 ) );
  XOR U5087 ( .A(n5081), .B(n5082), .Z(n2508) );
  ANDN U5088 ( .A(n4110), .B(n2511), .Z(\modmult_1/N560 ) );
  XOR U5089 ( .A(n5083), .B(n5084), .Z(n2511) );
  ANDN U5090 ( .A(n4110), .B(n2568), .Z(\modmult_1/N56 ) );
  XOR U5091 ( .A(n5085), .B(n5086), .Z(n2568) );
  ANDN U5092 ( .A(n4110), .B(n2514), .Z(\modmult_1/N559 ) );
  XOR U5093 ( .A(n5087), .B(n5088), .Z(n2514) );
  ANDN U5094 ( .A(n4110), .B(n2517), .Z(\modmult_1/N558 ) );
  XOR U5095 ( .A(n5089), .B(n5090), .Z(n2517) );
  ANDN U5096 ( .A(n4110), .B(n2520), .Z(\modmult_1/N557 ) );
  XOR U5097 ( .A(n5091), .B(n5092), .Z(n2520) );
  ANDN U5098 ( .A(n4110), .B(n2523), .Z(\modmult_1/N556 ) );
  XOR U5099 ( .A(n5093), .B(n5094), .Z(n2523) );
  ANDN U5100 ( .A(n4110), .B(n2526), .Z(\modmult_1/N555 ) );
  XOR U5101 ( .A(n5095), .B(n5096), .Z(n2526) );
  ANDN U5102 ( .A(n4110), .B(n2529), .Z(\modmult_1/N554 ) );
  XOR U5103 ( .A(n5097), .B(n5098), .Z(n2529) );
  ANDN U5104 ( .A(n4110), .B(n2532), .Z(\modmult_1/N553 ) );
  XOR U5105 ( .A(n5099), .B(n5100), .Z(n2532) );
  ANDN U5106 ( .A(n4110), .B(n2538), .Z(\modmult_1/N552 ) );
  XOR U5107 ( .A(n5101), .B(n5102), .Z(n2538) );
  ANDN U5108 ( .A(n4110), .B(n2541), .Z(\modmult_1/N551 ) );
  XOR U5109 ( .A(n5103), .B(n5104), .Z(n2541) );
  ANDN U5110 ( .A(n4110), .B(n2544), .Z(\modmult_1/N550 ) );
  XOR U5111 ( .A(n5105), .B(n5106), .Z(n2544) );
  ANDN U5112 ( .A(n4110), .B(n2601), .Z(\modmult_1/N55 ) );
  XOR U5113 ( .A(n5107), .B(n5108), .Z(n2601) );
  ANDN U5114 ( .A(n4110), .B(n2547), .Z(\modmult_1/N549 ) );
  XOR U5115 ( .A(n5109), .B(n5110), .Z(n2547) );
  ANDN U5116 ( .A(n4110), .B(n2550), .Z(\modmult_1/N548 ) );
  XOR U5117 ( .A(n5111), .B(n5112), .Z(n2550) );
  ANDN U5118 ( .A(n4110), .B(n2553), .Z(\modmult_1/N547 ) );
  XOR U5119 ( .A(n5113), .B(n5114), .Z(n2553) );
  ANDN U5120 ( .A(n4110), .B(n2556), .Z(\modmult_1/N546 ) );
  XOR U5121 ( .A(n5115), .B(n5116), .Z(n2556) );
  ANDN U5122 ( .A(n4110), .B(n2559), .Z(\modmult_1/N545 ) );
  XOR U5123 ( .A(n5117), .B(n5118), .Z(n2559) );
  ANDN U5124 ( .A(n4110), .B(n2562), .Z(\modmult_1/N544 ) );
  XOR U5125 ( .A(n5119), .B(n5120), .Z(n2562) );
  ANDN U5126 ( .A(n4110), .B(n2565), .Z(\modmult_1/N543 ) );
  XOR U5127 ( .A(n5121), .B(n5122), .Z(n2565) );
  ANDN U5128 ( .A(n4110), .B(n2571), .Z(\modmult_1/N542 ) );
  XOR U5129 ( .A(n5123), .B(n5124), .Z(n2571) );
  ANDN U5130 ( .A(n4110), .B(n2574), .Z(\modmult_1/N541 ) );
  XOR U5131 ( .A(n5125), .B(n5126), .Z(n2574) );
  ANDN U5132 ( .A(n4110), .B(n2577), .Z(\modmult_1/N540 ) );
  XOR U5133 ( .A(n5127), .B(n5128), .Z(n2577) );
  ANDN U5134 ( .A(n4110), .B(n2634), .Z(\modmult_1/N54 ) );
  XOR U5135 ( .A(n5129), .B(n5130), .Z(n2634) );
  ANDN U5136 ( .A(n4110), .B(n2580), .Z(\modmult_1/N539 ) );
  XOR U5137 ( .A(n5131), .B(n5132), .Z(n2580) );
  ANDN U5138 ( .A(n4110), .B(n2583), .Z(\modmult_1/N538 ) );
  XOR U5139 ( .A(n5133), .B(n5134), .Z(n2583) );
  ANDN U5140 ( .A(n4110), .B(n2586), .Z(\modmult_1/N537 ) );
  XOR U5141 ( .A(n5135), .B(n5136), .Z(n2586) );
  ANDN U5142 ( .A(n4110), .B(n2589), .Z(\modmult_1/N536 ) );
  XOR U5143 ( .A(n5137), .B(n5138), .Z(n2589) );
  ANDN U5144 ( .A(n4110), .B(n2592), .Z(\modmult_1/N535 ) );
  XOR U5145 ( .A(n5139), .B(n5140), .Z(n2592) );
  ANDN U5146 ( .A(n4110), .B(n2595), .Z(\modmult_1/N534 ) );
  XOR U5147 ( .A(n5141), .B(n5142), .Z(n2595) );
  ANDN U5148 ( .A(n4110), .B(n2598), .Z(\modmult_1/N533 ) );
  XOR U5149 ( .A(n5143), .B(n5144), .Z(n2598) );
  ANDN U5150 ( .A(n4110), .B(n2604), .Z(\modmult_1/N532 ) );
  XOR U5151 ( .A(n5145), .B(n5146), .Z(n2604) );
  ANDN U5152 ( .A(n4110), .B(n2607), .Z(\modmult_1/N531 ) );
  XOR U5153 ( .A(n5147), .B(n5148), .Z(n2607) );
  ANDN U5154 ( .A(n4110), .B(n2610), .Z(\modmult_1/N530 ) );
  XOR U5155 ( .A(n5149), .B(n5150), .Z(n2610) );
  ANDN U5156 ( .A(n4110), .B(n2667), .Z(\modmult_1/N53 ) );
  XOR U5157 ( .A(n5151), .B(n5152), .Z(n2667) );
  ANDN U5158 ( .A(n4110), .B(n2613), .Z(\modmult_1/N529 ) );
  XOR U5159 ( .A(n5153), .B(n5154), .Z(n2613) );
  ANDN U5160 ( .A(n4110), .B(n2616), .Z(\modmult_1/N528 ) );
  XOR U5161 ( .A(n5155), .B(n5156), .Z(n2616) );
  ANDN U5162 ( .A(n4110), .B(n2619), .Z(\modmult_1/N527 ) );
  XOR U5163 ( .A(n5157), .B(n5158), .Z(n2619) );
  ANDN U5164 ( .A(n4110), .B(n2622), .Z(\modmult_1/N526 ) );
  XOR U5165 ( .A(n5159), .B(n5160), .Z(n2622) );
  ANDN U5166 ( .A(n4110), .B(n2625), .Z(\modmult_1/N525 ) );
  XOR U5167 ( .A(n5161), .B(n5162), .Z(n2625) );
  ANDN U5168 ( .A(n4110), .B(n2628), .Z(\modmult_1/N524 ) );
  XOR U5169 ( .A(n5163), .B(n5164), .Z(n2628) );
  ANDN U5170 ( .A(n4110), .B(n2631), .Z(\modmult_1/N523 ) );
  XOR U5171 ( .A(n5165), .B(n5166), .Z(n2631) );
  ANDN U5172 ( .A(n4110), .B(n2637), .Z(\modmult_1/N522 ) );
  XOR U5173 ( .A(n5167), .B(n5168), .Z(n2637) );
  ANDN U5174 ( .A(n4110), .B(n2640), .Z(\modmult_1/N521 ) );
  XOR U5175 ( .A(n5169), .B(n5170), .Z(n2640) );
  ANDN U5176 ( .A(n4110), .B(n2643), .Z(\modmult_1/N520 ) );
  XOR U5177 ( .A(n5171), .B(n5172), .Z(n2643) );
  ANDN U5178 ( .A(n4110), .B(n2703), .Z(\modmult_1/N52 ) );
  XOR U5179 ( .A(n5173), .B(n5174), .Z(n2703) );
  ANDN U5180 ( .A(n4110), .B(n2646), .Z(\modmult_1/N519 ) );
  XOR U5181 ( .A(n5175), .B(n5176), .Z(n2646) );
  ANDN U5182 ( .A(n4110), .B(n2649), .Z(\modmult_1/N518 ) );
  XOR U5183 ( .A(n5177), .B(n5178), .Z(n2649) );
  ANDN U5184 ( .A(n4110), .B(n2652), .Z(\modmult_1/N517 ) );
  XOR U5185 ( .A(n5179), .B(n5180), .Z(n2652) );
  ANDN U5186 ( .A(n4110), .B(n2655), .Z(\modmult_1/N516 ) );
  XOR U5187 ( .A(n5181), .B(n5182), .Z(n2655) );
  ANDN U5188 ( .A(n4110), .B(n2658), .Z(\modmult_1/N515 ) );
  XOR U5189 ( .A(n5183), .B(n5184), .Z(n2658) );
  ANDN U5190 ( .A(n4110), .B(n2661), .Z(\modmult_1/N514 ) );
  XOR U5191 ( .A(n5185), .B(n5186), .Z(n2661) );
  ANDN U5192 ( .A(n4110), .B(n2664), .Z(\modmult_1/N513 ) );
  XOR U5193 ( .A(n5187), .B(n5188), .Z(n2664) );
  ANDN U5194 ( .A(n4110), .B(n2670), .Z(\modmult_1/N512 ) );
  XOR U5195 ( .A(n5189), .B(n5190), .Z(n2670) );
  ANDN U5196 ( .A(n4110), .B(n2673), .Z(\modmult_1/N511 ) );
  XOR U5197 ( .A(n5191), .B(n5192), .Z(n2673) );
  ANDN U5198 ( .A(n4110), .B(n2676), .Z(\modmult_1/N510 ) );
  XOR U5199 ( .A(n5193), .B(n5194), .Z(n2676) );
  ANDN U5200 ( .A(n4110), .B(n2736), .Z(\modmult_1/N51 ) );
  XOR U5201 ( .A(n5195), .B(n5196), .Z(n2736) );
  ANDN U5202 ( .A(n4110), .B(n2679), .Z(\modmult_1/N509 ) );
  XOR U5203 ( .A(n5197), .B(n5198), .Z(n2679) );
  ANDN U5204 ( .A(n4110), .B(n2682), .Z(\modmult_1/N508 ) );
  XOR U5205 ( .A(n5199), .B(n5200), .Z(n2682) );
  ANDN U5206 ( .A(n4110), .B(n2685), .Z(\modmult_1/N507 ) );
  XOR U5207 ( .A(n5201), .B(n5202), .Z(n2685) );
  ANDN U5208 ( .A(n4110), .B(n2688), .Z(\modmult_1/N506 ) );
  XOR U5209 ( .A(n5203), .B(n5204), .Z(n2688) );
  ANDN U5210 ( .A(n4110), .B(n2691), .Z(\modmult_1/N505 ) );
  XOR U5211 ( .A(n5205), .B(n5206), .Z(n2691) );
  ANDN U5212 ( .A(n4110), .B(n2694), .Z(\modmult_1/N504 ) );
  XOR U5213 ( .A(n5207), .B(n5208), .Z(n2694) );
  ANDN U5214 ( .A(n4110), .B(n2697), .Z(\modmult_1/N503 ) );
  XOR U5215 ( .A(n5209), .B(n5210), .Z(n2697) );
  ANDN U5216 ( .A(n4110), .B(n2706), .Z(\modmult_1/N502 ) );
  XOR U5217 ( .A(n5211), .B(n5212), .Z(n2706) );
  ANDN U5218 ( .A(n4110), .B(n2709), .Z(\modmult_1/N501 ) );
  XOR U5219 ( .A(n5213), .B(n5214), .Z(n2709) );
  ANDN U5220 ( .A(n4110), .B(n2712), .Z(\modmult_1/N500 ) );
  XOR U5221 ( .A(n5215), .B(n5216), .Z(n2712) );
  ANDN U5222 ( .A(n4110), .B(n2769), .Z(\modmult_1/N50 ) );
  XOR U5223 ( .A(n5217), .B(n5218), .Z(n2769) );
  ANDN U5224 ( .A(n4110), .B(n3366), .Z(\modmult_1/N5 ) );
  XOR U5225 ( .A(n5219), .B(n5220), .Z(n3366) );
  ANDN U5226 ( .A(n4110), .B(n2715), .Z(\modmult_1/N499 ) );
  XOR U5227 ( .A(n5221), .B(n5222), .Z(n2715) );
  ANDN U5228 ( .A(n4110), .B(n2718), .Z(\modmult_1/N498 ) );
  XOR U5229 ( .A(n5223), .B(n5224), .Z(n2718) );
  ANDN U5230 ( .A(n4110), .B(n2721), .Z(\modmult_1/N497 ) );
  XOR U5231 ( .A(n5225), .B(n5226), .Z(n2721) );
  ANDN U5232 ( .A(n4110), .B(n2724), .Z(\modmult_1/N496 ) );
  XOR U5233 ( .A(n5227), .B(n5228), .Z(n2724) );
  ANDN U5234 ( .A(n4110), .B(n2727), .Z(\modmult_1/N495 ) );
  XOR U5235 ( .A(n5229), .B(n5230), .Z(n2727) );
  ANDN U5236 ( .A(n4110), .B(n2730), .Z(\modmult_1/N494 ) );
  XOR U5237 ( .A(n5231), .B(n5232), .Z(n2730) );
  ANDN U5238 ( .A(n4110), .B(n2733), .Z(\modmult_1/N493 ) );
  XOR U5239 ( .A(n5233), .B(n5234), .Z(n2733) );
  ANDN U5240 ( .A(n4110), .B(n2739), .Z(\modmult_1/N492 ) );
  XOR U5241 ( .A(n5235), .B(n5236), .Z(n2739) );
  ANDN U5242 ( .A(n4110), .B(n2742), .Z(\modmult_1/N491 ) );
  XOR U5243 ( .A(n5237), .B(n5238), .Z(n2742) );
  ANDN U5244 ( .A(n4110), .B(n2745), .Z(\modmult_1/N490 ) );
  XOR U5245 ( .A(n5239), .B(n5240), .Z(n2745) );
  ANDN U5246 ( .A(n4110), .B(n2802), .Z(\modmult_1/N49 ) );
  XOR U5247 ( .A(n5241), .B(n5242), .Z(n2802) );
  ANDN U5248 ( .A(n4110), .B(n2748), .Z(\modmult_1/N489 ) );
  XOR U5249 ( .A(n5243), .B(n5244), .Z(n2748) );
  ANDN U5250 ( .A(n4110), .B(n2751), .Z(\modmult_1/N488 ) );
  XOR U5251 ( .A(n5245), .B(n5246), .Z(n2751) );
  ANDN U5252 ( .A(n4110), .B(n2754), .Z(\modmult_1/N487 ) );
  XOR U5253 ( .A(n5247), .B(n5248), .Z(n2754) );
  ANDN U5254 ( .A(n4110), .B(n2757), .Z(\modmult_1/N486 ) );
  XOR U5255 ( .A(n5249), .B(n5250), .Z(n2757) );
  ANDN U5256 ( .A(n4110), .B(n2760), .Z(\modmult_1/N485 ) );
  XOR U5257 ( .A(n5251), .B(n5252), .Z(n2760) );
  ANDN U5258 ( .A(n4110), .B(n2763), .Z(\modmult_1/N484 ) );
  XOR U5259 ( .A(n5253), .B(n5254), .Z(n2763) );
  ANDN U5260 ( .A(n4110), .B(n2766), .Z(\modmult_1/N483 ) );
  XOR U5261 ( .A(n5255), .B(n5256), .Z(n2766) );
  ANDN U5262 ( .A(n4110), .B(n2772), .Z(\modmult_1/N482 ) );
  XOR U5263 ( .A(n5257), .B(n5258), .Z(n2772) );
  ANDN U5264 ( .A(n4110), .B(n2775), .Z(\modmult_1/N481 ) );
  XOR U5265 ( .A(n5259), .B(n5260), .Z(n2775) );
  ANDN U5266 ( .A(n4110), .B(n2778), .Z(\modmult_1/N480 ) );
  XOR U5267 ( .A(n5261), .B(n5262), .Z(n2778) );
  ANDN U5268 ( .A(n4110), .B(n2835), .Z(\modmult_1/N48 ) );
  XOR U5269 ( .A(n5263), .B(n5264), .Z(n2835) );
  ANDN U5270 ( .A(n4110), .B(n2781), .Z(\modmult_1/N479 ) );
  XOR U5271 ( .A(n5265), .B(n5266), .Z(n2781) );
  ANDN U5272 ( .A(n4110), .B(n2784), .Z(\modmult_1/N478 ) );
  XOR U5273 ( .A(n5267), .B(n5268), .Z(n2784) );
  ANDN U5274 ( .A(n4110), .B(n2787), .Z(\modmult_1/N477 ) );
  XOR U5275 ( .A(n5269), .B(n5270), .Z(n2787) );
  ANDN U5276 ( .A(n4110), .B(n2790), .Z(\modmult_1/N476 ) );
  XOR U5277 ( .A(n5271), .B(n5272), .Z(n2790) );
  ANDN U5278 ( .A(n4110), .B(n2793), .Z(\modmult_1/N475 ) );
  XOR U5279 ( .A(n5273), .B(n5274), .Z(n2793) );
  ANDN U5280 ( .A(n4110), .B(n2796), .Z(\modmult_1/N474 ) );
  XOR U5281 ( .A(n5275), .B(n5276), .Z(n2796) );
  ANDN U5282 ( .A(n4110), .B(n2799), .Z(\modmult_1/N473 ) );
  XOR U5283 ( .A(n5277), .B(n5278), .Z(n2799) );
  ANDN U5284 ( .A(n4110), .B(n2805), .Z(\modmult_1/N472 ) );
  XOR U5285 ( .A(n5279), .B(n5280), .Z(n2805) );
  ANDN U5286 ( .A(n4110), .B(n2808), .Z(\modmult_1/N471 ) );
  XOR U5287 ( .A(n5281), .B(n5282), .Z(n2808) );
  ANDN U5288 ( .A(n4110), .B(n2811), .Z(\modmult_1/N470 ) );
  XOR U5289 ( .A(n5283), .B(n5284), .Z(n2811) );
  ANDN U5290 ( .A(n4110), .B(n2868), .Z(\modmult_1/N47 ) );
  XOR U5291 ( .A(n5285), .B(n5286), .Z(n2868) );
  ANDN U5292 ( .A(n4110), .B(n2814), .Z(\modmult_1/N469 ) );
  XOR U5293 ( .A(n5287), .B(n5288), .Z(n2814) );
  ANDN U5294 ( .A(n4110), .B(n2817), .Z(\modmult_1/N468 ) );
  XOR U5295 ( .A(n5289), .B(n5290), .Z(n2817) );
  ANDN U5296 ( .A(n4110), .B(n2820), .Z(\modmult_1/N467 ) );
  XOR U5297 ( .A(n5291), .B(n5292), .Z(n2820) );
  ANDN U5298 ( .A(n4110), .B(n2823), .Z(\modmult_1/N466 ) );
  XOR U5299 ( .A(n5293), .B(n5294), .Z(n2823) );
  ANDN U5300 ( .A(n4110), .B(n2826), .Z(\modmult_1/N465 ) );
  XOR U5301 ( .A(n5295), .B(n5296), .Z(n2826) );
  ANDN U5302 ( .A(n4110), .B(n2829), .Z(\modmult_1/N464 ) );
  XOR U5303 ( .A(n5297), .B(n5298), .Z(n2829) );
  ANDN U5304 ( .A(n4110), .B(n2832), .Z(\modmult_1/N463 ) );
  XOR U5305 ( .A(n5299), .B(n5300), .Z(n2832) );
  ANDN U5306 ( .A(n4110), .B(n2838), .Z(\modmult_1/N462 ) );
  XOR U5307 ( .A(n5301), .B(n5302), .Z(n2838) );
  ANDN U5308 ( .A(n4110), .B(n2841), .Z(\modmult_1/N461 ) );
  XOR U5309 ( .A(n5303), .B(n5304), .Z(n2841) );
  ANDN U5310 ( .A(n4110), .B(n2844), .Z(\modmult_1/N460 ) );
  XOR U5311 ( .A(n5305), .B(n5306), .Z(n2844) );
  ANDN U5312 ( .A(n4110), .B(n2901), .Z(\modmult_1/N46 ) );
  XOR U5313 ( .A(n5307), .B(n5308), .Z(n2901) );
  ANDN U5314 ( .A(n4110), .B(n2847), .Z(\modmult_1/N459 ) );
  XOR U5315 ( .A(n5309), .B(n5310), .Z(n2847) );
  ANDN U5316 ( .A(n4110), .B(n2850), .Z(\modmult_1/N458 ) );
  XOR U5317 ( .A(n5311), .B(n5312), .Z(n2850) );
  ANDN U5318 ( .A(n4110), .B(n2853), .Z(\modmult_1/N457 ) );
  XOR U5319 ( .A(n5313), .B(n5314), .Z(n2853) );
  ANDN U5320 ( .A(n4110), .B(n2856), .Z(\modmult_1/N456 ) );
  XOR U5321 ( .A(n5315), .B(n5316), .Z(n2856) );
  ANDN U5322 ( .A(n4110), .B(n2859), .Z(\modmult_1/N455 ) );
  XOR U5323 ( .A(n5317), .B(n5318), .Z(n2859) );
  ANDN U5324 ( .A(n4110), .B(n2862), .Z(\modmult_1/N454 ) );
  XOR U5325 ( .A(n5319), .B(n5320), .Z(n2862) );
  ANDN U5326 ( .A(n4110), .B(n2865), .Z(\modmult_1/N453 ) );
  XOR U5327 ( .A(n5321), .B(n5322), .Z(n2865) );
  ANDN U5328 ( .A(n4110), .B(n2871), .Z(\modmult_1/N452 ) );
  XOR U5329 ( .A(n5323), .B(n5324), .Z(n2871) );
  ANDN U5330 ( .A(n4110), .B(n2874), .Z(\modmult_1/N451 ) );
  XOR U5331 ( .A(n5325), .B(n5326), .Z(n2874) );
  ANDN U5332 ( .A(n4110), .B(n2877), .Z(\modmult_1/N450 ) );
  XOR U5333 ( .A(n5327), .B(n5328), .Z(n2877) );
  ANDN U5334 ( .A(n4110), .B(n2934), .Z(\modmult_1/N45 ) );
  XOR U5335 ( .A(n5329), .B(n5330), .Z(n2934) );
  ANDN U5336 ( .A(n4110), .B(n2880), .Z(\modmult_1/N449 ) );
  XOR U5337 ( .A(n5331), .B(n5332), .Z(n2880) );
  ANDN U5338 ( .A(n4110), .B(n2883), .Z(\modmult_1/N448 ) );
  XOR U5339 ( .A(n5333), .B(n5334), .Z(n2883) );
  ANDN U5340 ( .A(n4110), .B(n2886), .Z(\modmult_1/N447 ) );
  XOR U5341 ( .A(n5335), .B(n5336), .Z(n2886) );
  ANDN U5342 ( .A(n4110), .B(n2889), .Z(\modmult_1/N446 ) );
  XOR U5343 ( .A(n5337), .B(n5338), .Z(n2889) );
  ANDN U5344 ( .A(n4110), .B(n2892), .Z(\modmult_1/N445 ) );
  XOR U5345 ( .A(n5339), .B(n5340), .Z(n2892) );
  ANDN U5346 ( .A(n4110), .B(n2895), .Z(\modmult_1/N444 ) );
  XOR U5347 ( .A(n5341), .B(n5342), .Z(n2895) );
  ANDN U5348 ( .A(n4110), .B(n2898), .Z(\modmult_1/N443 ) );
  XOR U5349 ( .A(n5343), .B(n5344), .Z(n2898) );
  ANDN U5350 ( .A(n4110), .B(n2904), .Z(\modmult_1/N442 ) );
  XOR U5351 ( .A(n5345), .B(n5346), .Z(n2904) );
  ANDN U5352 ( .A(n4110), .B(n2907), .Z(\modmult_1/N441 ) );
  XOR U5353 ( .A(n5347), .B(n5348), .Z(n2907) );
  ANDN U5354 ( .A(n4110), .B(n2910), .Z(\modmult_1/N440 ) );
  XOR U5355 ( .A(n5349), .B(n5350), .Z(n2910) );
  ANDN U5356 ( .A(n4110), .B(n2967), .Z(\modmult_1/N44 ) );
  XOR U5357 ( .A(n5351), .B(n5352), .Z(n2967) );
  ANDN U5358 ( .A(n4110), .B(n2913), .Z(\modmult_1/N439 ) );
  XOR U5359 ( .A(n5353), .B(n5354), .Z(n2913) );
  ANDN U5360 ( .A(n4110), .B(n2916), .Z(\modmult_1/N438 ) );
  XOR U5361 ( .A(n5355), .B(n5356), .Z(n2916) );
  ANDN U5362 ( .A(n4110), .B(n2919), .Z(\modmult_1/N437 ) );
  XOR U5363 ( .A(n5357), .B(n5358), .Z(n2919) );
  ANDN U5364 ( .A(n4110), .B(n2922), .Z(\modmult_1/N436 ) );
  XOR U5365 ( .A(n5359), .B(n5360), .Z(n2922) );
  ANDN U5366 ( .A(n4110), .B(n2925), .Z(\modmult_1/N435 ) );
  XOR U5367 ( .A(n5361), .B(n5362), .Z(n2925) );
  ANDN U5368 ( .A(n4110), .B(n2928), .Z(\modmult_1/N434 ) );
  XOR U5369 ( .A(n5363), .B(n5364), .Z(n2928) );
  ANDN U5370 ( .A(n4110), .B(n2931), .Z(\modmult_1/N433 ) );
  XOR U5371 ( .A(n5365), .B(n5366), .Z(n2931) );
  ANDN U5372 ( .A(n4110), .B(n2937), .Z(\modmult_1/N432 ) );
  XOR U5373 ( .A(n5367), .B(n5368), .Z(n2937) );
  ANDN U5374 ( .A(n4110), .B(n2940), .Z(\modmult_1/N431 ) );
  XOR U5375 ( .A(n5369), .B(n5370), .Z(n2940) );
  ANDN U5376 ( .A(n4110), .B(n2943), .Z(\modmult_1/N430 ) );
  XOR U5377 ( .A(n5371), .B(n5372), .Z(n2943) );
  ANDN U5378 ( .A(n4110), .B(n3000), .Z(\modmult_1/N43 ) );
  XOR U5379 ( .A(n5373), .B(n5374), .Z(n3000) );
  ANDN U5380 ( .A(n4110), .B(n2946), .Z(\modmult_1/N429 ) );
  XOR U5381 ( .A(n5375), .B(n5376), .Z(n2946) );
  ANDN U5382 ( .A(n4110), .B(n2949), .Z(\modmult_1/N428 ) );
  XOR U5383 ( .A(n5377), .B(n5378), .Z(n2949) );
  ANDN U5384 ( .A(n4110), .B(n2952), .Z(\modmult_1/N427 ) );
  XOR U5385 ( .A(n5379), .B(n5380), .Z(n2952) );
  ANDN U5386 ( .A(n4110), .B(n2955), .Z(\modmult_1/N426 ) );
  XOR U5387 ( .A(n5381), .B(n5382), .Z(n2955) );
  ANDN U5388 ( .A(n4110), .B(n2958), .Z(\modmult_1/N425 ) );
  XOR U5389 ( .A(n5383), .B(n5384), .Z(n2958) );
  ANDN U5390 ( .A(n4110), .B(n2961), .Z(\modmult_1/N424 ) );
  XOR U5391 ( .A(n5385), .B(n5386), .Z(n2961) );
  ANDN U5392 ( .A(n4110), .B(n2964), .Z(\modmult_1/N423 ) );
  XOR U5393 ( .A(n5387), .B(n5388), .Z(n2964) );
  ANDN U5394 ( .A(n4110), .B(n2970), .Z(\modmult_1/N422 ) );
  XOR U5395 ( .A(n5389), .B(n5390), .Z(n2970) );
  ANDN U5396 ( .A(n4110), .B(n2973), .Z(\modmult_1/N421 ) );
  XOR U5397 ( .A(n5391), .B(n5392), .Z(n2973) );
  ANDN U5398 ( .A(n4110), .B(n2976), .Z(\modmult_1/N420 ) );
  XOR U5399 ( .A(n5393), .B(n5394), .Z(n2976) );
  ANDN U5400 ( .A(n4110), .B(n3036), .Z(\modmult_1/N42 ) );
  XOR U5401 ( .A(n5395), .B(n5396), .Z(n3036) );
  ANDN U5402 ( .A(n4110), .B(n2979), .Z(\modmult_1/N419 ) );
  XOR U5403 ( .A(n5397), .B(n5398), .Z(n2979) );
  ANDN U5404 ( .A(n4110), .B(n2982), .Z(\modmult_1/N418 ) );
  XOR U5405 ( .A(n5399), .B(n5400), .Z(n2982) );
  ANDN U5406 ( .A(n4110), .B(n2985), .Z(\modmult_1/N417 ) );
  XOR U5407 ( .A(n5401), .B(n5402), .Z(n2985) );
  ANDN U5408 ( .A(n4110), .B(n2988), .Z(\modmult_1/N416 ) );
  XOR U5409 ( .A(n5403), .B(n5404), .Z(n2988) );
  ANDN U5410 ( .A(n4110), .B(n2991), .Z(\modmult_1/N415 ) );
  XOR U5411 ( .A(n5405), .B(n5406), .Z(n2991) );
  ANDN U5412 ( .A(n4110), .B(n2994), .Z(\modmult_1/N414 ) );
  XOR U5413 ( .A(n5407), .B(n5408), .Z(n2994) );
  ANDN U5414 ( .A(n4110), .B(n2997), .Z(\modmult_1/N413 ) );
  XOR U5415 ( .A(n5409), .B(n5410), .Z(n2997) );
  ANDN U5416 ( .A(n4110), .B(n3003), .Z(\modmult_1/N412 ) );
  XOR U5417 ( .A(n5411), .B(n5412), .Z(n3003) );
  ANDN U5418 ( .A(n4110), .B(n3006), .Z(\modmult_1/N411 ) );
  XOR U5419 ( .A(n5413), .B(n5414), .Z(n3006) );
  ANDN U5420 ( .A(n4110), .B(n3009), .Z(\modmult_1/N410 ) );
  XOR U5421 ( .A(n5415), .B(n5416), .Z(n3009) );
  ANDN U5422 ( .A(n4110), .B(n3069), .Z(\modmult_1/N41 ) );
  XOR U5423 ( .A(n5417), .B(n5418), .Z(n3069) );
  ANDN U5424 ( .A(n4110), .B(n3012), .Z(\modmult_1/N409 ) );
  XOR U5425 ( .A(n5419), .B(n5420), .Z(n3012) );
  ANDN U5426 ( .A(n4110), .B(n3015), .Z(\modmult_1/N408 ) );
  XOR U5427 ( .A(n5421), .B(n5422), .Z(n3015) );
  ANDN U5428 ( .A(n4110), .B(n3018), .Z(\modmult_1/N407 ) );
  XOR U5429 ( .A(n5423), .B(n5424), .Z(n3018) );
  ANDN U5430 ( .A(n4110), .B(n3021), .Z(\modmult_1/N406 ) );
  XOR U5431 ( .A(n5425), .B(n5426), .Z(n3021) );
  ANDN U5432 ( .A(n4110), .B(n3024), .Z(\modmult_1/N405 ) );
  XOR U5433 ( .A(n5427), .B(n5428), .Z(n3024) );
  ANDN U5434 ( .A(n4110), .B(n3027), .Z(\modmult_1/N404 ) );
  XOR U5435 ( .A(n5429), .B(n5430), .Z(n3027) );
  ANDN U5436 ( .A(n4110), .B(n3030), .Z(\modmult_1/N403 ) );
  XOR U5437 ( .A(n5431), .B(n5432), .Z(n3030) );
  ANDN U5438 ( .A(n4110), .B(n3039), .Z(\modmult_1/N402 ) );
  XOR U5439 ( .A(n5433), .B(n5434), .Z(n3039) );
  ANDN U5440 ( .A(n4110), .B(n3042), .Z(\modmult_1/N401 ) );
  XOR U5441 ( .A(n5435), .B(n5436), .Z(n3042) );
  ANDN U5442 ( .A(n4110), .B(n3045), .Z(\modmult_1/N400 ) );
  XOR U5443 ( .A(n5437), .B(n5438), .Z(n3045) );
  ANDN U5444 ( .A(n4110), .B(n3102), .Z(\modmult_1/N40 ) );
  XOR U5445 ( .A(n5439), .B(n5440), .Z(n3102) );
  ANDN U5446 ( .A(n4110), .B(n3699), .Z(\modmult_1/N4 ) );
  XOR U5447 ( .A(n5441), .B(n5442), .Z(n3699) );
  ANDN U5448 ( .A(n4110), .B(n3048), .Z(\modmult_1/N399 ) );
  XOR U5449 ( .A(n5443), .B(n5444), .Z(n3048) );
  ANDN U5450 ( .A(n4110), .B(n3051), .Z(\modmult_1/N398 ) );
  XOR U5451 ( .A(n5445), .B(n5446), .Z(n3051) );
  ANDN U5452 ( .A(n4110), .B(n3054), .Z(\modmult_1/N397 ) );
  XOR U5453 ( .A(n5447), .B(n5448), .Z(n3054) );
  ANDN U5454 ( .A(n4110), .B(n3057), .Z(\modmult_1/N396 ) );
  XOR U5455 ( .A(n5449), .B(n5450), .Z(n3057) );
  ANDN U5456 ( .A(n4110), .B(n3060), .Z(\modmult_1/N395 ) );
  XOR U5457 ( .A(n5451), .B(n5452), .Z(n3060) );
  ANDN U5458 ( .A(n4110), .B(n3063), .Z(\modmult_1/N394 ) );
  XOR U5459 ( .A(n5453), .B(n5454), .Z(n3063) );
  ANDN U5460 ( .A(n4110), .B(n3066), .Z(\modmult_1/N393 ) );
  XOR U5461 ( .A(n5455), .B(n5456), .Z(n3066) );
  ANDN U5462 ( .A(n4110), .B(n3072), .Z(\modmult_1/N392 ) );
  XOR U5463 ( .A(n5457), .B(n5458), .Z(n3072) );
  ANDN U5464 ( .A(n4110), .B(n3075), .Z(\modmult_1/N391 ) );
  XOR U5465 ( .A(n5459), .B(n5460), .Z(n3075) );
  ANDN U5466 ( .A(n4110), .B(n3078), .Z(\modmult_1/N390 ) );
  XOR U5467 ( .A(n5461), .B(n5462), .Z(n3078) );
  ANDN U5468 ( .A(n4110), .B(n3135), .Z(\modmult_1/N39 ) );
  XOR U5469 ( .A(n5463), .B(n5464), .Z(n3135) );
  ANDN U5470 ( .A(n4110), .B(n3081), .Z(\modmult_1/N389 ) );
  XOR U5471 ( .A(n5465), .B(n5466), .Z(n3081) );
  ANDN U5472 ( .A(n4110), .B(n3084), .Z(\modmult_1/N388 ) );
  XOR U5473 ( .A(n5467), .B(n5468), .Z(n3084) );
  ANDN U5474 ( .A(n4110), .B(n3087), .Z(\modmult_1/N387 ) );
  XOR U5475 ( .A(n5469), .B(n5470), .Z(n3087) );
  ANDN U5476 ( .A(n4110), .B(n3090), .Z(\modmult_1/N386 ) );
  XOR U5477 ( .A(n5471), .B(n5472), .Z(n3090) );
  ANDN U5478 ( .A(n4110), .B(n3093), .Z(\modmult_1/N385 ) );
  XOR U5479 ( .A(n5473), .B(n5474), .Z(n3093) );
  ANDN U5480 ( .A(n4110), .B(n3096), .Z(\modmult_1/N384 ) );
  XOR U5481 ( .A(n5475), .B(n5476), .Z(n3096) );
  ANDN U5482 ( .A(n4110), .B(n3099), .Z(\modmult_1/N383 ) );
  XOR U5483 ( .A(n5477), .B(n5478), .Z(n3099) );
  ANDN U5484 ( .A(n4110), .B(n3105), .Z(\modmult_1/N382 ) );
  XOR U5485 ( .A(n5479), .B(n5480), .Z(n3105) );
  ANDN U5486 ( .A(n4110), .B(n3108), .Z(\modmult_1/N381 ) );
  XOR U5487 ( .A(n5481), .B(n5482), .Z(n3108) );
  ANDN U5488 ( .A(n4110), .B(n3111), .Z(\modmult_1/N380 ) );
  XOR U5489 ( .A(n5483), .B(n5484), .Z(n3111) );
  ANDN U5490 ( .A(n4110), .B(n3168), .Z(\modmult_1/N38 ) );
  XOR U5491 ( .A(n5485), .B(n5486), .Z(n3168) );
  ANDN U5492 ( .A(n4110), .B(n3114), .Z(\modmult_1/N379 ) );
  XOR U5493 ( .A(n5487), .B(n5488), .Z(n3114) );
  ANDN U5494 ( .A(n4110), .B(n3117), .Z(\modmult_1/N378 ) );
  XOR U5495 ( .A(n5489), .B(n5490), .Z(n3117) );
  ANDN U5496 ( .A(n4110), .B(n3120), .Z(\modmult_1/N377 ) );
  XOR U5497 ( .A(n5491), .B(n5492), .Z(n3120) );
  ANDN U5498 ( .A(n4110), .B(n3123), .Z(\modmult_1/N376 ) );
  XOR U5499 ( .A(n5493), .B(n5494), .Z(n3123) );
  ANDN U5500 ( .A(n4110), .B(n3126), .Z(\modmult_1/N375 ) );
  XOR U5501 ( .A(n5495), .B(n5496), .Z(n3126) );
  ANDN U5502 ( .A(n4110), .B(n3129), .Z(\modmult_1/N374 ) );
  XOR U5503 ( .A(n5497), .B(n5498), .Z(n3129) );
  ANDN U5504 ( .A(n4110), .B(n3132), .Z(\modmult_1/N373 ) );
  XOR U5505 ( .A(n5499), .B(n5500), .Z(n3132) );
  ANDN U5506 ( .A(n4110), .B(n3138), .Z(\modmult_1/N372 ) );
  XOR U5507 ( .A(n5501), .B(n5502), .Z(n3138) );
  ANDN U5508 ( .A(n4110), .B(n3141), .Z(\modmult_1/N371 ) );
  XOR U5509 ( .A(n5503), .B(n5504), .Z(n3141) );
  ANDN U5510 ( .A(n4110), .B(n3144), .Z(\modmult_1/N370 ) );
  XOR U5511 ( .A(n5505), .B(n5506), .Z(n3144) );
  ANDN U5512 ( .A(n4110), .B(n3201), .Z(\modmult_1/N37 ) );
  XOR U5513 ( .A(n5507), .B(n5508), .Z(n3201) );
  ANDN U5514 ( .A(n4110), .B(n3147), .Z(\modmult_1/N369 ) );
  XOR U5515 ( .A(n5509), .B(n5510), .Z(n3147) );
  ANDN U5516 ( .A(n4110), .B(n3150), .Z(\modmult_1/N368 ) );
  XOR U5517 ( .A(n5511), .B(n5512), .Z(n3150) );
  ANDN U5518 ( .A(n4110), .B(n3153), .Z(\modmult_1/N367 ) );
  XOR U5519 ( .A(n5513), .B(n5514), .Z(n3153) );
  ANDN U5520 ( .A(n4110), .B(n3156), .Z(\modmult_1/N366 ) );
  XOR U5521 ( .A(n5515), .B(n5516), .Z(n3156) );
  ANDN U5522 ( .A(n4110), .B(n3159), .Z(\modmult_1/N365 ) );
  XOR U5523 ( .A(n5517), .B(n5518), .Z(n3159) );
  ANDN U5524 ( .A(n4110), .B(n3162), .Z(\modmult_1/N364 ) );
  XOR U5525 ( .A(n5519), .B(n5520), .Z(n3162) );
  ANDN U5526 ( .A(n4110), .B(n3165), .Z(\modmult_1/N363 ) );
  XOR U5527 ( .A(n5521), .B(n5522), .Z(n3165) );
  ANDN U5528 ( .A(n4110), .B(n3171), .Z(\modmult_1/N362 ) );
  XOR U5529 ( .A(n5523), .B(n5524), .Z(n3171) );
  ANDN U5530 ( .A(n4110), .B(n3174), .Z(\modmult_1/N361 ) );
  XOR U5531 ( .A(n5525), .B(n5526), .Z(n3174) );
  ANDN U5532 ( .A(n4110), .B(n3177), .Z(\modmult_1/N360 ) );
  XOR U5533 ( .A(n5527), .B(n5528), .Z(n3177) );
  ANDN U5534 ( .A(n4110), .B(n3234), .Z(\modmult_1/N36 ) );
  XOR U5535 ( .A(n5529), .B(n5530), .Z(n3234) );
  ANDN U5536 ( .A(n4110), .B(n3180), .Z(\modmult_1/N359 ) );
  XOR U5537 ( .A(n5531), .B(n5532), .Z(n3180) );
  ANDN U5538 ( .A(n4110), .B(n3183), .Z(\modmult_1/N358 ) );
  XOR U5539 ( .A(n5533), .B(n5534), .Z(n3183) );
  ANDN U5540 ( .A(n4110), .B(n3186), .Z(\modmult_1/N357 ) );
  XOR U5541 ( .A(n5535), .B(n5536), .Z(n3186) );
  ANDN U5542 ( .A(n4110), .B(n3189), .Z(\modmult_1/N356 ) );
  XOR U5543 ( .A(n5537), .B(n5538), .Z(n3189) );
  ANDN U5544 ( .A(n4110), .B(n3192), .Z(\modmult_1/N355 ) );
  XOR U5545 ( .A(n5539), .B(n5540), .Z(n3192) );
  ANDN U5546 ( .A(n4110), .B(n3195), .Z(\modmult_1/N354 ) );
  XOR U5547 ( .A(n5541), .B(n5542), .Z(n3195) );
  ANDN U5548 ( .A(n4110), .B(n3198), .Z(\modmult_1/N353 ) );
  XOR U5549 ( .A(n5543), .B(n5544), .Z(n3198) );
  ANDN U5550 ( .A(n4110), .B(n3204), .Z(\modmult_1/N352 ) );
  XOR U5551 ( .A(n5545), .B(n5546), .Z(n3204) );
  ANDN U5552 ( .A(n4110), .B(n3207), .Z(\modmult_1/N351 ) );
  XOR U5553 ( .A(n5547), .B(n5548), .Z(n3207) );
  ANDN U5554 ( .A(n4110), .B(n3210), .Z(\modmult_1/N350 ) );
  XOR U5555 ( .A(n5549), .B(n5550), .Z(n3210) );
  ANDN U5556 ( .A(n4110), .B(n3267), .Z(\modmult_1/N35 ) );
  XOR U5557 ( .A(n5551), .B(n5552), .Z(n3267) );
  ANDN U5558 ( .A(n4110), .B(n3213), .Z(\modmult_1/N349 ) );
  XOR U5559 ( .A(n5553), .B(n5554), .Z(n3213) );
  ANDN U5560 ( .A(n4110), .B(n3216), .Z(\modmult_1/N348 ) );
  XOR U5561 ( .A(n5555), .B(n5556), .Z(n3216) );
  ANDN U5562 ( .A(n4110), .B(n3219), .Z(\modmult_1/N347 ) );
  XOR U5563 ( .A(n5557), .B(n5558), .Z(n3219) );
  ANDN U5564 ( .A(n4110), .B(n3222), .Z(\modmult_1/N346 ) );
  XOR U5565 ( .A(n5559), .B(n5560), .Z(n3222) );
  ANDN U5566 ( .A(n4110), .B(n3225), .Z(\modmult_1/N345 ) );
  XOR U5567 ( .A(n5561), .B(n5562), .Z(n3225) );
  ANDN U5568 ( .A(n4110), .B(n3228), .Z(\modmult_1/N344 ) );
  XOR U5569 ( .A(n5563), .B(n5564), .Z(n3228) );
  ANDN U5570 ( .A(n4110), .B(n3231), .Z(\modmult_1/N343 ) );
  XOR U5571 ( .A(n5565), .B(n5566), .Z(n3231) );
  ANDN U5572 ( .A(n4110), .B(n3237), .Z(\modmult_1/N342 ) );
  XOR U5573 ( .A(n5567), .B(n5568), .Z(n3237) );
  ANDN U5574 ( .A(n4110), .B(n3240), .Z(\modmult_1/N341 ) );
  XOR U5575 ( .A(n5569), .B(n5570), .Z(n3240) );
  ANDN U5576 ( .A(n4110), .B(n3243), .Z(\modmult_1/N340 ) );
  XOR U5577 ( .A(n5571), .B(n5572), .Z(n3243) );
  ANDN U5578 ( .A(n4110), .B(n3300), .Z(\modmult_1/N34 ) );
  XOR U5579 ( .A(n5573), .B(n5574), .Z(n3300) );
  ANDN U5580 ( .A(n4110), .B(n3246), .Z(\modmult_1/N339 ) );
  XOR U5581 ( .A(n5575), .B(n5576), .Z(n3246) );
  ANDN U5582 ( .A(n4110), .B(n3249), .Z(\modmult_1/N338 ) );
  XOR U5583 ( .A(n5577), .B(n5578), .Z(n3249) );
  ANDN U5584 ( .A(n4110), .B(n3252), .Z(\modmult_1/N337 ) );
  XOR U5585 ( .A(n5579), .B(n5580), .Z(n3252) );
  ANDN U5586 ( .A(n4110), .B(n3255), .Z(\modmult_1/N336 ) );
  XOR U5587 ( .A(n5581), .B(n5582), .Z(n3255) );
  ANDN U5588 ( .A(n4110), .B(n3258), .Z(\modmult_1/N335 ) );
  XOR U5589 ( .A(n5583), .B(n5584), .Z(n3258) );
  ANDN U5590 ( .A(n4110), .B(n3261), .Z(\modmult_1/N334 ) );
  XOR U5591 ( .A(n5585), .B(n5586), .Z(n3261) );
  ANDN U5592 ( .A(n4110), .B(n3264), .Z(\modmult_1/N333 ) );
  XOR U5593 ( .A(n5587), .B(n5588), .Z(n3264) );
  ANDN U5594 ( .A(n4110), .B(n3270), .Z(\modmult_1/N332 ) );
  XOR U5595 ( .A(n5589), .B(n5590), .Z(n3270) );
  ANDN U5596 ( .A(n4110), .B(n3273), .Z(\modmult_1/N331 ) );
  XOR U5597 ( .A(n5591), .B(n5592), .Z(n3273) );
  ANDN U5598 ( .A(n4110), .B(n3276), .Z(\modmult_1/N330 ) );
  XOR U5599 ( .A(n5593), .B(n5594), .Z(n3276) );
  ANDN U5600 ( .A(n4110), .B(n3333), .Z(\modmult_1/N33 ) );
  XOR U5601 ( .A(n5595), .B(n5596), .Z(n3333) );
  ANDN U5602 ( .A(n4110), .B(n3279), .Z(\modmult_1/N329 ) );
  XOR U5603 ( .A(n5597), .B(n5598), .Z(n3279) );
  ANDN U5604 ( .A(n4110), .B(n3282), .Z(\modmult_1/N328 ) );
  XOR U5605 ( .A(n5599), .B(n5600), .Z(n3282) );
  ANDN U5606 ( .A(n4110), .B(n3285), .Z(\modmult_1/N327 ) );
  XOR U5607 ( .A(n5601), .B(n5602), .Z(n3285) );
  ANDN U5608 ( .A(n4110), .B(n3288), .Z(\modmult_1/N326 ) );
  XOR U5609 ( .A(n5603), .B(n5604), .Z(n3288) );
  ANDN U5610 ( .A(n4110), .B(n3291), .Z(\modmult_1/N325 ) );
  XOR U5611 ( .A(n5605), .B(n5606), .Z(n3291) );
  ANDN U5612 ( .A(n4110), .B(n3294), .Z(\modmult_1/N324 ) );
  XOR U5613 ( .A(n5607), .B(n5608), .Z(n3294) );
  ANDN U5614 ( .A(n4110), .B(n3297), .Z(\modmult_1/N323 ) );
  XOR U5615 ( .A(n5609), .B(n5610), .Z(n3297) );
  ANDN U5616 ( .A(n4110), .B(n3303), .Z(\modmult_1/N322 ) );
  XOR U5617 ( .A(n5611), .B(n5612), .Z(n3303) );
  ANDN U5618 ( .A(n4110), .B(n3306), .Z(\modmult_1/N321 ) );
  XOR U5619 ( .A(n5613), .B(n5614), .Z(n3306) );
  ANDN U5620 ( .A(n4110), .B(n3309), .Z(\modmult_1/N320 ) );
  XOR U5621 ( .A(n5615), .B(n5616), .Z(n3309) );
  ANDN U5622 ( .A(n4110), .B(n3369), .Z(\modmult_1/N32 ) );
  XOR U5623 ( .A(n5617), .B(n5618), .Z(n3369) );
  ANDN U5624 ( .A(n4110), .B(n3312), .Z(\modmult_1/N319 ) );
  XOR U5625 ( .A(n5619), .B(n5620), .Z(n3312) );
  ANDN U5626 ( .A(n4110), .B(n3315), .Z(\modmult_1/N318 ) );
  XOR U5627 ( .A(n5621), .B(n5622), .Z(n3315) );
  ANDN U5628 ( .A(n4110), .B(n3318), .Z(\modmult_1/N317 ) );
  XOR U5629 ( .A(n5623), .B(n5624), .Z(n3318) );
  ANDN U5630 ( .A(n4110), .B(n3321), .Z(\modmult_1/N316 ) );
  XOR U5631 ( .A(n5625), .B(n5626), .Z(n3321) );
  ANDN U5632 ( .A(n4110), .B(n3324), .Z(\modmult_1/N315 ) );
  XOR U5633 ( .A(n5627), .B(n5628), .Z(n3324) );
  ANDN U5634 ( .A(n4110), .B(n3327), .Z(\modmult_1/N314 ) );
  XOR U5635 ( .A(n5629), .B(n5630), .Z(n3327) );
  ANDN U5636 ( .A(n4110), .B(n3330), .Z(\modmult_1/N313 ) );
  XOR U5637 ( .A(n5631), .B(n5632), .Z(n3330) );
  ANDN U5638 ( .A(n4110), .B(n3336), .Z(\modmult_1/N312 ) );
  XOR U5639 ( .A(n5633), .B(n5634), .Z(n3336) );
  ANDN U5640 ( .A(n4110), .B(n3339), .Z(\modmult_1/N311 ) );
  XOR U5641 ( .A(n5635), .B(n5636), .Z(n3339) );
  ANDN U5642 ( .A(n4110), .B(n3342), .Z(\modmult_1/N310 ) );
  XOR U5643 ( .A(n5637), .B(n5638), .Z(n3342) );
  ANDN U5644 ( .A(n4110), .B(n3402), .Z(\modmult_1/N31 ) );
  XOR U5645 ( .A(n5639), .B(n5640), .Z(n3402) );
  ANDN U5646 ( .A(n4110), .B(n3345), .Z(\modmult_1/N309 ) );
  XOR U5647 ( .A(n5641), .B(n5642), .Z(n3345) );
  ANDN U5648 ( .A(n4110), .B(n3348), .Z(\modmult_1/N308 ) );
  XOR U5649 ( .A(n5643), .B(n5644), .Z(n3348) );
  ANDN U5650 ( .A(n4110), .B(n3351), .Z(\modmult_1/N307 ) );
  XOR U5651 ( .A(n5645), .B(n5646), .Z(n3351) );
  ANDN U5652 ( .A(n4110), .B(n3354), .Z(\modmult_1/N306 ) );
  XOR U5653 ( .A(n5647), .B(n5648), .Z(n3354) );
  ANDN U5654 ( .A(n4110), .B(n3357), .Z(\modmult_1/N305 ) );
  XOR U5655 ( .A(n5649), .B(n5650), .Z(n3357) );
  ANDN U5656 ( .A(n4110), .B(n3360), .Z(\modmult_1/N304 ) );
  XOR U5657 ( .A(n5651), .B(n5652), .Z(n3360) );
  ANDN U5658 ( .A(n4110), .B(n3363), .Z(\modmult_1/N303 ) );
  XOR U5659 ( .A(n5653), .B(n5654), .Z(n3363) );
  ANDN U5660 ( .A(n4110), .B(n3372), .Z(\modmult_1/N302 ) );
  XOR U5661 ( .A(n5655), .B(n5656), .Z(n3372) );
  ANDN U5662 ( .A(n4110), .B(n3375), .Z(\modmult_1/N301 ) );
  XOR U5663 ( .A(n5657), .B(n5658), .Z(n3375) );
  ANDN U5664 ( .A(n4110), .B(n3378), .Z(\modmult_1/N300 ) );
  XOR U5665 ( .A(n5659), .B(n5660), .Z(n3378) );
  ANDN U5666 ( .A(n4110), .B(n3435), .Z(\modmult_1/N30 ) );
  XOR U5667 ( .A(n5661), .B(n5662), .Z(n3435) );
  AND U5668 ( .A(n4104), .B(n4110), .Z(\modmult_1/N3 ) );
  XOR U5669 ( .A(n5663), .B(n5664), .Z(n4104) );
  ANDN U5670 ( .A(n4110), .B(n3381), .Z(\modmult_1/N299 ) );
  XOR U5671 ( .A(n5665), .B(n5666), .Z(n3381) );
  ANDN U5672 ( .A(n4110), .B(n3384), .Z(\modmult_1/N298 ) );
  XOR U5673 ( .A(n5667), .B(n5668), .Z(n3384) );
  ANDN U5674 ( .A(n4110), .B(n3387), .Z(\modmult_1/N297 ) );
  XOR U5675 ( .A(n5669), .B(n5670), .Z(n3387) );
  ANDN U5676 ( .A(n4110), .B(n3390), .Z(\modmult_1/N296 ) );
  XOR U5677 ( .A(n5671), .B(n5672), .Z(n3390) );
  ANDN U5678 ( .A(n4110), .B(n3393), .Z(\modmult_1/N295 ) );
  XOR U5679 ( .A(n5673), .B(n5674), .Z(n3393) );
  ANDN U5680 ( .A(n4110), .B(n3396), .Z(\modmult_1/N294 ) );
  XOR U5681 ( .A(n5675), .B(n5676), .Z(n3396) );
  ANDN U5682 ( .A(n4110), .B(n3399), .Z(\modmult_1/N293 ) );
  XOR U5683 ( .A(n5677), .B(n5678), .Z(n3399) );
  ANDN U5684 ( .A(n4110), .B(n3405), .Z(\modmult_1/N292 ) );
  XOR U5685 ( .A(n5679), .B(n5680), .Z(n3405) );
  ANDN U5686 ( .A(n4110), .B(n3408), .Z(\modmult_1/N291 ) );
  XOR U5687 ( .A(n5681), .B(n5682), .Z(n3408) );
  ANDN U5688 ( .A(n4110), .B(n3411), .Z(\modmult_1/N290 ) );
  XOR U5689 ( .A(n5683), .B(n5684), .Z(n3411) );
  ANDN U5690 ( .A(n4110), .B(n3468), .Z(\modmult_1/N29 ) );
  XOR U5691 ( .A(n5685), .B(n5686), .Z(n3468) );
  ANDN U5692 ( .A(n4110), .B(n3414), .Z(\modmult_1/N289 ) );
  XOR U5693 ( .A(n5687), .B(n5688), .Z(n3414) );
  ANDN U5694 ( .A(n4110), .B(n3417), .Z(\modmult_1/N288 ) );
  XOR U5695 ( .A(n5689), .B(n5690), .Z(n3417) );
  ANDN U5696 ( .A(n4110), .B(n3420), .Z(\modmult_1/N287 ) );
  XOR U5697 ( .A(n5691), .B(n5692), .Z(n3420) );
  ANDN U5698 ( .A(n4110), .B(n3423), .Z(\modmult_1/N286 ) );
  XOR U5699 ( .A(n5693), .B(n5694), .Z(n3423) );
  ANDN U5700 ( .A(n4110), .B(n3426), .Z(\modmult_1/N285 ) );
  XOR U5701 ( .A(n5695), .B(n5696), .Z(n3426) );
  ANDN U5702 ( .A(n4110), .B(n3429), .Z(\modmult_1/N284 ) );
  XOR U5703 ( .A(n5697), .B(n5698), .Z(n3429) );
  ANDN U5704 ( .A(n4110), .B(n3432), .Z(\modmult_1/N283 ) );
  XOR U5705 ( .A(n5699), .B(n5700), .Z(n3432) );
  ANDN U5706 ( .A(n4110), .B(n3438), .Z(\modmult_1/N282 ) );
  XOR U5707 ( .A(n5701), .B(n5702), .Z(n3438) );
  ANDN U5708 ( .A(n4110), .B(n3441), .Z(\modmult_1/N281 ) );
  XOR U5709 ( .A(n5703), .B(n5704), .Z(n3441) );
  ANDN U5710 ( .A(n4110), .B(n3444), .Z(\modmult_1/N280 ) );
  XOR U5711 ( .A(n5705), .B(n5706), .Z(n3444) );
  ANDN U5712 ( .A(n4110), .B(n3501), .Z(\modmult_1/N28 ) );
  XOR U5713 ( .A(n5707), .B(n5708), .Z(n3501) );
  ANDN U5714 ( .A(n4110), .B(n3447), .Z(\modmult_1/N279 ) );
  XOR U5715 ( .A(n5709), .B(n5710), .Z(n3447) );
  ANDN U5716 ( .A(n4110), .B(n3450), .Z(\modmult_1/N278 ) );
  XOR U5717 ( .A(n5711), .B(n5712), .Z(n3450) );
  ANDN U5718 ( .A(n4110), .B(n3453), .Z(\modmult_1/N277 ) );
  XOR U5719 ( .A(n5713), .B(n5714), .Z(n3453) );
  ANDN U5720 ( .A(n4110), .B(n3456), .Z(\modmult_1/N276 ) );
  XOR U5721 ( .A(n5715), .B(n5716), .Z(n3456) );
  ANDN U5722 ( .A(n4110), .B(n3459), .Z(\modmult_1/N275 ) );
  XOR U5723 ( .A(n5717), .B(n5718), .Z(n3459) );
  ANDN U5724 ( .A(n4110), .B(n3462), .Z(\modmult_1/N274 ) );
  XOR U5725 ( .A(n5719), .B(n5720), .Z(n3462) );
  ANDN U5726 ( .A(n4110), .B(n3465), .Z(\modmult_1/N273 ) );
  XOR U5727 ( .A(n5721), .B(n5722), .Z(n3465) );
  ANDN U5728 ( .A(n4110), .B(n3471), .Z(\modmult_1/N272 ) );
  XOR U5729 ( .A(n5723), .B(n5724), .Z(n3471) );
  ANDN U5730 ( .A(n4110), .B(n3474), .Z(\modmult_1/N271 ) );
  XOR U5731 ( .A(n5725), .B(n5726), .Z(n3474) );
  ANDN U5732 ( .A(n4110), .B(n3477), .Z(\modmult_1/N270 ) );
  XOR U5733 ( .A(n5727), .B(n5728), .Z(n3477) );
  ANDN U5734 ( .A(n4110), .B(n3534), .Z(\modmult_1/N27 ) );
  XOR U5735 ( .A(n5729), .B(n5730), .Z(n3534) );
  ANDN U5736 ( .A(n4110), .B(n3480), .Z(\modmult_1/N269 ) );
  XOR U5737 ( .A(n5731), .B(n5732), .Z(n3480) );
  ANDN U5738 ( .A(n4110), .B(n3483), .Z(\modmult_1/N268 ) );
  XOR U5739 ( .A(n5733), .B(n5734), .Z(n3483) );
  ANDN U5740 ( .A(n4110), .B(n3486), .Z(\modmult_1/N267 ) );
  XOR U5741 ( .A(n5735), .B(n5736), .Z(n3486) );
  ANDN U5742 ( .A(n4110), .B(n3489), .Z(\modmult_1/N266 ) );
  XOR U5743 ( .A(n5737), .B(n5738), .Z(n3489) );
  ANDN U5744 ( .A(n4110), .B(n3492), .Z(\modmult_1/N265 ) );
  XOR U5745 ( .A(n5739), .B(n5740), .Z(n3492) );
  ANDN U5746 ( .A(n4110), .B(n3495), .Z(\modmult_1/N264 ) );
  XOR U5747 ( .A(n5741), .B(n5742), .Z(n3495) );
  ANDN U5748 ( .A(n4110), .B(n3498), .Z(\modmult_1/N263 ) );
  XOR U5749 ( .A(n5743), .B(n5744), .Z(n3498) );
  ANDN U5750 ( .A(n4110), .B(n3504), .Z(\modmult_1/N262 ) );
  XOR U5751 ( .A(n5745), .B(n5746), .Z(n3504) );
  ANDN U5752 ( .A(n4110), .B(n3507), .Z(\modmult_1/N261 ) );
  XOR U5753 ( .A(n5747), .B(n5748), .Z(n3507) );
  ANDN U5754 ( .A(n4110), .B(n3510), .Z(\modmult_1/N260 ) );
  XOR U5755 ( .A(n5749), .B(n5750), .Z(n3510) );
  ANDN U5756 ( .A(n4110), .B(n3567), .Z(\modmult_1/N26 ) );
  XOR U5757 ( .A(n5751), .B(n5752), .Z(n3567) );
  ANDN U5758 ( .A(n4110), .B(n3513), .Z(\modmult_1/N259 ) );
  XOR U5759 ( .A(n5753), .B(n5754), .Z(n3513) );
  ANDN U5760 ( .A(n4110), .B(n3516), .Z(\modmult_1/N258 ) );
  XOR U5761 ( .A(n5755), .B(n5756), .Z(n3516) );
  ANDN U5762 ( .A(n4110), .B(n3519), .Z(\modmult_1/N257 ) );
  XOR U5763 ( .A(n5757), .B(n5758), .Z(n3519) );
  ANDN U5764 ( .A(n4110), .B(n3522), .Z(\modmult_1/N256 ) );
  XOR U5765 ( .A(n5759), .B(n5760), .Z(n3522) );
  ANDN U5766 ( .A(n4110), .B(n3525), .Z(\modmult_1/N255 ) );
  XOR U5767 ( .A(n5761), .B(n5762), .Z(n3525) );
  ANDN U5768 ( .A(n4110), .B(n3528), .Z(\modmult_1/N254 ) );
  XOR U5769 ( .A(n5763), .B(n5764), .Z(n3528) );
  ANDN U5770 ( .A(n4110), .B(n3531), .Z(\modmult_1/N253 ) );
  XOR U5771 ( .A(n5765), .B(n5766), .Z(n3531) );
  ANDN U5772 ( .A(n4110), .B(n3537), .Z(\modmult_1/N252 ) );
  XOR U5773 ( .A(n5767), .B(n5768), .Z(n3537) );
  ANDN U5774 ( .A(n4110), .B(n3540), .Z(\modmult_1/N251 ) );
  XOR U5775 ( .A(n5769), .B(n5770), .Z(n3540) );
  ANDN U5776 ( .A(n4110), .B(n3543), .Z(\modmult_1/N250 ) );
  XOR U5777 ( .A(n5771), .B(n5772), .Z(n3543) );
  ANDN U5778 ( .A(n4110), .B(n3600), .Z(\modmult_1/N25 ) );
  XOR U5779 ( .A(n5773), .B(n5774), .Z(n3600) );
  ANDN U5780 ( .A(n4110), .B(n3546), .Z(\modmult_1/N249 ) );
  XOR U5781 ( .A(n5775), .B(n5776), .Z(n3546) );
  ANDN U5782 ( .A(n4110), .B(n3549), .Z(\modmult_1/N248 ) );
  XOR U5783 ( .A(n5777), .B(n5778), .Z(n3549) );
  ANDN U5784 ( .A(n4110), .B(n3552), .Z(\modmult_1/N247 ) );
  XOR U5785 ( .A(n5779), .B(n5780), .Z(n3552) );
  ANDN U5786 ( .A(n4110), .B(n3555), .Z(\modmult_1/N246 ) );
  XOR U5787 ( .A(n5781), .B(n5782), .Z(n3555) );
  ANDN U5788 ( .A(n4110), .B(n3558), .Z(\modmult_1/N245 ) );
  XOR U5789 ( .A(n5783), .B(n5784), .Z(n3558) );
  ANDN U5790 ( .A(n4110), .B(n3561), .Z(\modmult_1/N244 ) );
  XOR U5791 ( .A(n5785), .B(n5786), .Z(n3561) );
  ANDN U5792 ( .A(n4110), .B(n3564), .Z(\modmult_1/N243 ) );
  XOR U5793 ( .A(n5787), .B(n5788), .Z(n3564) );
  ANDN U5794 ( .A(n4110), .B(n3570), .Z(\modmult_1/N242 ) );
  XOR U5795 ( .A(n5789), .B(n5790), .Z(n3570) );
  ANDN U5796 ( .A(n4110), .B(n3573), .Z(\modmult_1/N241 ) );
  XOR U5797 ( .A(n5791), .B(n5792), .Z(n3573) );
  ANDN U5798 ( .A(n4110), .B(n3576), .Z(\modmult_1/N240 ) );
  XOR U5799 ( .A(n5793), .B(n5794), .Z(n3576) );
  ANDN U5800 ( .A(n4110), .B(n3633), .Z(\modmult_1/N24 ) );
  XOR U5801 ( .A(n5795), .B(n5796), .Z(n3633) );
  ANDN U5802 ( .A(n4110), .B(n3579), .Z(\modmult_1/N239 ) );
  XOR U5803 ( .A(n5797), .B(n5798), .Z(n3579) );
  ANDN U5804 ( .A(n4110), .B(n3582), .Z(\modmult_1/N238 ) );
  XOR U5805 ( .A(n5799), .B(n5800), .Z(n3582) );
  ANDN U5806 ( .A(n4110), .B(n3585), .Z(\modmult_1/N237 ) );
  XOR U5807 ( .A(n5801), .B(n5802), .Z(n3585) );
  ANDN U5808 ( .A(n4110), .B(n3588), .Z(\modmult_1/N236 ) );
  XOR U5809 ( .A(n5803), .B(n5804), .Z(n3588) );
  ANDN U5810 ( .A(n4110), .B(n3591), .Z(\modmult_1/N235 ) );
  XOR U5811 ( .A(n5805), .B(n5806), .Z(n3591) );
  ANDN U5812 ( .A(n4110), .B(n3594), .Z(\modmult_1/N234 ) );
  XOR U5813 ( .A(n5807), .B(n5808), .Z(n3594) );
  ANDN U5814 ( .A(n4110), .B(n3597), .Z(\modmult_1/N233 ) );
  XOR U5815 ( .A(n5809), .B(n5810), .Z(n3597) );
  ANDN U5816 ( .A(n4110), .B(n3603), .Z(\modmult_1/N232 ) );
  XOR U5817 ( .A(n5811), .B(n5812), .Z(n3603) );
  ANDN U5818 ( .A(n4110), .B(n3606), .Z(\modmult_1/N231 ) );
  XOR U5819 ( .A(n5813), .B(n5814), .Z(n3606) );
  ANDN U5820 ( .A(n4110), .B(n3609), .Z(\modmult_1/N230 ) );
  XOR U5821 ( .A(n5815), .B(n5816), .Z(n3609) );
  ANDN U5822 ( .A(n4110), .B(n3666), .Z(\modmult_1/N23 ) );
  XOR U5823 ( .A(n5817), .B(n5818), .Z(n3666) );
  ANDN U5824 ( .A(n4110), .B(n3612), .Z(\modmult_1/N229 ) );
  XOR U5825 ( .A(n5819), .B(n5820), .Z(n3612) );
  ANDN U5826 ( .A(n4110), .B(n3615), .Z(\modmult_1/N228 ) );
  XOR U5827 ( .A(n5821), .B(n5822), .Z(n3615) );
  ANDN U5828 ( .A(n4110), .B(n3618), .Z(\modmult_1/N227 ) );
  XOR U5829 ( .A(n5823), .B(n5824), .Z(n3618) );
  ANDN U5830 ( .A(n4110), .B(n3621), .Z(\modmult_1/N226 ) );
  XOR U5831 ( .A(n5825), .B(n5826), .Z(n3621) );
  ANDN U5832 ( .A(n4110), .B(n3624), .Z(\modmult_1/N225 ) );
  XOR U5833 ( .A(n5827), .B(n5828), .Z(n3624) );
  ANDN U5834 ( .A(n4110), .B(n3627), .Z(\modmult_1/N224 ) );
  XOR U5835 ( .A(n5829), .B(n5830), .Z(n3627) );
  ANDN U5836 ( .A(n4110), .B(n3630), .Z(\modmult_1/N223 ) );
  XOR U5837 ( .A(n5831), .B(n5832), .Z(n3630) );
  ANDN U5838 ( .A(n4110), .B(n3636), .Z(\modmult_1/N222 ) );
  XOR U5839 ( .A(n5833), .B(n5834), .Z(n3636) );
  ANDN U5840 ( .A(n4110), .B(n3639), .Z(\modmult_1/N221 ) );
  XOR U5841 ( .A(n5835), .B(n5836), .Z(n3639) );
  ANDN U5842 ( .A(n4110), .B(n3642), .Z(\modmult_1/N220 ) );
  XOR U5843 ( .A(n5837), .B(n5838), .Z(n3642) );
  ANDN U5844 ( .A(n4110), .B(n3702), .Z(\modmult_1/N22 ) );
  XOR U5845 ( .A(n5839), .B(n5840), .Z(n3702) );
  ANDN U5846 ( .A(n4110), .B(n3645), .Z(\modmult_1/N219 ) );
  XOR U5847 ( .A(n5841), .B(n5842), .Z(n3645) );
  ANDN U5848 ( .A(n4110), .B(n3648), .Z(\modmult_1/N218 ) );
  XOR U5849 ( .A(n5843), .B(n5844), .Z(n3648) );
  ANDN U5850 ( .A(n4110), .B(n3651), .Z(\modmult_1/N217 ) );
  XOR U5851 ( .A(n5845), .B(n5846), .Z(n3651) );
  ANDN U5852 ( .A(n4110), .B(n3654), .Z(\modmult_1/N216 ) );
  XOR U5853 ( .A(n5847), .B(n5848), .Z(n3654) );
  ANDN U5854 ( .A(n4110), .B(n3657), .Z(\modmult_1/N215 ) );
  XOR U5855 ( .A(n5849), .B(n5850), .Z(n3657) );
  ANDN U5856 ( .A(n4110), .B(n3660), .Z(\modmult_1/N214 ) );
  XOR U5857 ( .A(n5851), .B(n5852), .Z(n3660) );
  ANDN U5858 ( .A(n4110), .B(n3663), .Z(\modmult_1/N213 ) );
  XOR U5859 ( .A(n5853), .B(n5854), .Z(n3663) );
  ANDN U5860 ( .A(n4110), .B(n3669), .Z(\modmult_1/N212 ) );
  XOR U5861 ( .A(n5855), .B(n5856), .Z(n3669) );
  ANDN U5862 ( .A(n4110), .B(n3672), .Z(\modmult_1/N211 ) );
  XOR U5863 ( .A(n5857), .B(n5858), .Z(n3672) );
  ANDN U5864 ( .A(n4110), .B(n3675), .Z(\modmult_1/N210 ) );
  XOR U5865 ( .A(n5859), .B(n5860), .Z(n3675) );
  ANDN U5866 ( .A(n4110), .B(n3735), .Z(\modmult_1/N21 ) );
  XOR U5867 ( .A(n5861), .B(n5862), .Z(n3735) );
  ANDN U5868 ( .A(n4110), .B(n3678), .Z(\modmult_1/N209 ) );
  XOR U5869 ( .A(n5863), .B(n5864), .Z(n3678) );
  ANDN U5870 ( .A(n4110), .B(n3681), .Z(\modmult_1/N208 ) );
  XOR U5871 ( .A(n5865), .B(n5866), .Z(n3681) );
  ANDN U5872 ( .A(n4110), .B(n3684), .Z(\modmult_1/N207 ) );
  XOR U5873 ( .A(n5867), .B(n5868), .Z(n3684) );
  ANDN U5874 ( .A(n4110), .B(n3687), .Z(\modmult_1/N206 ) );
  XOR U5875 ( .A(n5869), .B(n5870), .Z(n3687) );
  MUX U5876 ( .IN0(\modmult_1/xin[1022] ), .IN1(creg[1023]), .SEL(start_in[0]), 
        .F(\modmult_1/N2052 ) );
  MUX U5877 ( .IN0(\modmult_1/xin[1021] ), .IN1(creg[1022]), .SEL(start_in[0]), 
        .F(\modmult_1/N2051 ) );
  MUX U5878 ( .IN0(\modmult_1/xin[1020] ), .IN1(creg[1021]), .SEL(start_in[0]), 
        .F(\modmult_1/N2050 ) );
  ANDN U5879 ( .A(n4110), .B(n3690), .Z(\modmult_1/N205 ) );
  XOR U5880 ( .A(n5871), .B(n5872), .Z(n3690) );
  MUX U5881 ( .IN0(\modmult_1/xin[1019] ), .IN1(creg[1020]), .SEL(start_in[0]), 
        .F(\modmult_1/N2049 ) );
  MUX U5882 ( .IN0(\modmult_1/xin[1018] ), .IN1(creg[1019]), .SEL(start_in[0]), 
        .F(\modmult_1/N2048 ) );
  MUX U5883 ( .IN0(\modmult_1/xin[1017] ), .IN1(creg[1018]), .SEL(start_in[0]), 
        .F(\modmult_1/N2047 ) );
  MUX U5884 ( .IN0(\modmult_1/xin[1016] ), .IN1(creg[1017]), .SEL(start_in[0]), 
        .F(\modmult_1/N2046 ) );
  MUX U5885 ( .IN0(\modmult_1/xin[1015] ), .IN1(creg[1016]), .SEL(start_in[0]), 
        .F(\modmult_1/N2045 ) );
  MUX U5886 ( .IN0(\modmult_1/xin[1014] ), .IN1(creg[1015]), .SEL(start_in[0]), 
        .F(\modmult_1/N2044 ) );
  MUX U5887 ( .IN0(\modmult_1/xin[1013] ), .IN1(creg[1014]), .SEL(start_in[0]), 
        .F(\modmult_1/N2043 ) );
  MUX U5888 ( .IN0(\modmult_1/xin[1012] ), .IN1(creg[1013]), .SEL(start_in[0]), 
        .F(\modmult_1/N2042 ) );
  MUX U5889 ( .IN0(\modmult_1/xin[1011] ), .IN1(creg[1012]), .SEL(start_in[0]), 
        .F(\modmult_1/N2041 ) );
  MUX U5890 ( .IN0(\modmult_1/xin[1010] ), .IN1(creg[1011]), .SEL(start_in[0]), 
        .F(\modmult_1/N2040 ) );
  ANDN U5891 ( .A(n4110), .B(n3693), .Z(\modmult_1/N204 ) );
  XOR U5892 ( .A(n5873), .B(n5874), .Z(n3693) );
  MUX U5893 ( .IN0(\modmult_1/xin[1009] ), .IN1(creg[1010]), .SEL(start_in[0]), 
        .F(\modmult_1/N2039 ) );
  MUX U5894 ( .IN0(\modmult_1/xin[1008] ), .IN1(creg[1009]), .SEL(start_in[0]), 
        .F(\modmult_1/N2038 ) );
  MUX U5895 ( .IN0(\modmult_1/xin[1007] ), .IN1(creg[1008]), .SEL(start_in[0]), 
        .F(\modmult_1/N2037 ) );
  MUX U5896 ( .IN0(\modmult_1/xin[1006] ), .IN1(creg[1007]), .SEL(start_in[0]), 
        .F(\modmult_1/N2036 ) );
  MUX U5897 ( .IN0(\modmult_1/xin[1005] ), .IN1(creg[1006]), .SEL(start_in[0]), 
        .F(\modmult_1/N2035 ) );
  MUX U5898 ( .IN0(\modmult_1/xin[1004] ), .IN1(creg[1005]), .SEL(start_in[0]), 
        .F(\modmult_1/N2034 ) );
  MUX U5899 ( .IN0(\modmult_1/xin[1003] ), .IN1(creg[1004]), .SEL(start_in[0]), 
        .F(\modmult_1/N2033 ) );
  MUX U5900 ( .IN0(\modmult_1/xin[1002] ), .IN1(creg[1003]), .SEL(start_in[0]), 
        .F(\modmult_1/N2032 ) );
  MUX U5901 ( .IN0(\modmult_1/xin[1001] ), .IN1(creg[1002]), .SEL(start_in[0]), 
        .F(\modmult_1/N2031 ) );
  MUX U5902 ( .IN0(\modmult_1/xin[1000] ), .IN1(creg[1001]), .SEL(start_in[0]), 
        .F(\modmult_1/N2030 ) );
  ANDN U5903 ( .A(n4110), .B(n3696), .Z(\modmult_1/N203 ) );
  XOR U5904 ( .A(n5875), .B(n5876), .Z(n3696) );
  MUX U5905 ( .IN0(\modmult_1/xin[999] ), .IN1(creg[1000]), .SEL(start_in[0]), 
        .F(\modmult_1/N2029 ) );
  MUX U5906 ( .IN0(\modmult_1/xin[998] ), .IN1(creg[999]), .SEL(start_in[0]), 
        .F(\modmult_1/N2028 ) );
  MUX U5907 ( .IN0(\modmult_1/xin[997] ), .IN1(creg[998]), .SEL(start_in[0]), 
        .F(\modmult_1/N2027 ) );
  MUX U5908 ( .IN0(\modmult_1/xin[996] ), .IN1(creg[997]), .SEL(start_in[0]), 
        .F(\modmult_1/N2026 ) );
  MUX U5909 ( .IN0(\modmult_1/xin[995] ), .IN1(creg[996]), .SEL(start_in[0]), 
        .F(\modmult_1/N2025 ) );
  MUX U5910 ( .IN0(\modmult_1/xin[994] ), .IN1(creg[995]), .SEL(start_in[0]), 
        .F(\modmult_1/N2024 ) );
  MUX U5911 ( .IN0(\modmult_1/xin[993] ), .IN1(creg[994]), .SEL(start_in[0]), 
        .F(\modmult_1/N2023 ) );
  MUX U5912 ( .IN0(\modmult_1/xin[992] ), .IN1(creg[993]), .SEL(start_in[0]), 
        .F(\modmult_1/N2022 ) );
  MUX U5913 ( .IN0(\modmult_1/xin[991] ), .IN1(creg[992]), .SEL(start_in[0]), 
        .F(\modmult_1/N2021 ) );
  MUX U5914 ( .IN0(\modmult_1/xin[990] ), .IN1(creg[991]), .SEL(start_in[0]), 
        .F(\modmult_1/N2020 ) );
  ANDN U5915 ( .A(n4110), .B(n3705), .Z(\modmult_1/N202 ) );
  XOR U5916 ( .A(n5877), .B(n5878), .Z(n3705) );
  MUX U5917 ( .IN0(\modmult_1/xin[989] ), .IN1(creg[990]), .SEL(start_in[0]), 
        .F(\modmult_1/N2019 ) );
  MUX U5918 ( .IN0(\modmult_1/xin[988] ), .IN1(creg[989]), .SEL(start_in[0]), 
        .F(\modmult_1/N2018 ) );
  MUX U5919 ( .IN0(\modmult_1/xin[987] ), .IN1(creg[988]), .SEL(start_in[0]), 
        .F(\modmult_1/N2017 ) );
  MUX U5920 ( .IN0(\modmult_1/xin[986] ), .IN1(creg[987]), .SEL(start_in[0]), 
        .F(\modmult_1/N2016 ) );
  MUX U5921 ( .IN0(\modmult_1/xin[985] ), .IN1(creg[986]), .SEL(start_in[0]), 
        .F(\modmult_1/N2015 ) );
  MUX U5922 ( .IN0(\modmult_1/xin[984] ), .IN1(creg[985]), .SEL(start_in[0]), 
        .F(\modmult_1/N2014 ) );
  MUX U5923 ( .IN0(\modmult_1/xin[983] ), .IN1(creg[984]), .SEL(start_in[0]), 
        .F(\modmult_1/N2013 ) );
  MUX U5924 ( .IN0(\modmult_1/xin[982] ), .IN1(creg[983]), .SEL(start_in[0]), 
        .F(\modmult_1/N2012 ) );
  MUX U5925 ( .IN0(\modmult_1/xin[981] ), .IN1(creg[982]), .SEL(start_in[0]), 
        .F(\modmult_1/N2011 ) );
  MUX U5926 ( .IN0(\modmult_1/xin[980] ), .IN1(creg[981]), .SEL(start_in[0]), 
        .F(\modmult_1/N2010 ) );
  ANDN U5927 ( .A(n4110), .B(n3708), .Z(\modmult_1/N201 ) );
  XOR U5928 ( .A(n5879), .B(n5880), .Z(n3708) );
  MUX U5929 ( .IN0(\modmult_1/xin[979] ), .IN1(creg[980]), .SEL(start_in[0]), 
        .F(\modmult_1/N2009 ) );
  MUX U5930 ( .IN0(\modmult_1/xin[978] ), .IN1(creg[979]), .SEL(start_in[0]), 
        .F(\modmult_1/N2008 ) );
  MUX U5931 ( .IN0(\modmult_1/xin[977] ), .IN1(creg[978]), .SEL(start_in[0]), 
        .F(\modmult_1/N2007 ) );
  MUX U5932 ( .IN0(\modmult_1/xin[976] ), .IN1(creg[977]), .SEL(start_in[0]), 
        .F(\modmult_1/N2006 ) );
  MUX U5933 ( .IN0(\modmult_1/xin[975] ), .IN1(creg[976]), .SEL(start_in[0]), 
        .F(\modmult_1/N2005 ) );
  MUX U5934 ( .IN0(\modmult_1/xin[974] ), .IN1(creg[975]), .SEL(start_in[0]), 
        .F(\modmult_1/N2004 ) );
  MUX U5935 ( .IN0(\modmult_1/xin[973] ), .IN1(creg[974]), .SEL(start_in[0]), 
        .F(\modmult_1/N2003 ) );
  MUX U5936 ( .IN0(\modmult_1/xin[972] ), .IN1(creg[973]), .SEL(start_in[0]), 
        .F(\modmult_1/N2002 ) );
  MUX U5937 ( .IN0(\modmult_1/xin[971] ), .IN1(creg[972]), .SEL(start_in[0]), 
        .F(\modmult_1/N2001 ) );
  MUX U5938 ( .IN0(\modmult_1/xin[970] ), .IN1(creg[971]), .SEL(start_in[0]), 
        .F(\modmult_1/N2000 ) );
  ANDN U5939 ( .A(n4110), .B(n3711), .Z(\modmult_1/N200 ) );
  XOR U5940 ( .A(n5881), .B(n5882), .Z(n3711) );
  ANDN U5941 ( .A(n4110), .B(n3768), .Z(\modmult_1/N20 ) );
  XOR U5942 ( .A(n5883), .B(n5884), .Z(n3768) );
  MUX U5943 ( .IN0(\modmult_1/xin[969] ), .IN1(creg[970]), .SEL(start_in[0]), 
        .F(\modmult_1/N1999 ) );
  MUX U5944 ( .IN0(\modmult_1/xin[968] ), .IN1(creg[969]), .SEL(start_in[0]), 
        .F(\modmult_1/N1998 ) );
  MUX U5945 ( .IN0(\modmult_1/xin[967] ), .IN1(creg[968]), .SEL(start_in[0]), 
        .F(\modmult_1/N1997 ) );
  MUX U5946 ( .IN0(\modmult_1/xin[966] ), .IN1(creg[967]), .SEL(start_in[0]), 
        .F(\modmult_1/N1996 ) );
  MUX U5947 ( .IN0(\modmult_1/xin[965] ), .IN1(creg[966]), .SEL(start_in[0]), 
        .F(\modmult_1/N1995 ) );
  MUX U5948 ( .IN0(\modmult_1/xin[964] ), .IN1(creg[965]), .SEL(start_in[0]), 
        .F(\modmult_1/N1994 ) );
  MUX U5949 ( .IN0(\modmult_1/xin[963] ), .IN1(creg[964]), .SEL(start_in[0]), 
        .F(\modmult_1/N1993 ) );
  MUX U5950 ( .IN0(\modmult_1/xin[962] ), .IN1(creg[963]), .SEL(start_in[0]), 
        .F(\modmult_1/N1992 ) );
  MUX U5951 ( .IN0(\modmult_1/xin[961] ), .IN1(creg[962]), .SEL(start_in[0]), 
        .F(\modmult_1/N1991 ) );
  MUX U5952 ( .IN0(\modmult_1/xin[960] ), .IN1(creg[961]), .SEL(start_in[0]), 
        .F(\modmult_1/N1990 ) );
  ANDN U5953 ( .A(n4110), .B(n3714), .Z(\modmult_1/N199 ) );
  XOR U5954 ( .A(n5885), .B(n5886), .Z(n3714) );
  MUX U5955 ( .IN0(\modmult_1/xin[959] ), .IN1(creg[960]), .SEL(start_in[0]), 
        .F(\modmult_1/N1989 ) );
  MUX U5956 ( .IN0(\modmult_1/xin[958] ), .IN1(creg[959]), .SEL(start_in[0]), 
        .F(\modmult_1/N1988 ) );
  MUX U5957 ( .IN0(\modmult_1/xin[957] ), .IN1(creg[958]), .SEL(start_in[0]), 
        .F(\modmult_1/N1987 ) );
  MUX U5958 ( .IN0(\modmult_1/xin[956] ), .IN1(creg[957]), .SEL(start_in[0]), 
        .F(\modmult_1/N1986 ) );
  MUX U5959 ( .IN0(\modmult_1/xin[955] ), .IN1(creg[956]), .SEL(start_in[0]), 
        .F(\modmult_1/N1985 ) );
  MUX U5960 ( .IN0(\modmult_1/xin[954] ), .IN1(creg[955]), .SEL(start_in[0]), 
        .F(\modmult_1/N1984 ) );
  MUX U5961 ( .IN0(\modmult_1/xin[953] ), .IN1(creg[954]), .SEL(start_in[0]), 
        .F(\modmult_1/N1983 ) );
  MUX U5962 ( .IN0(\modmult_1/xin[952] ), .IN1(creg[953]), .SEL(start_in[0]), 
        .F(\modmult_1/N1982 ) );
  MUX U5963 ( .IN0(\modmult_1/xin[951] ), .IN1(creg[952]), .SEL(start_in[0]), 
        .F(\modmult_1/N1981 ) );
  MUX U5964 ( .IN0(\modmult_1/xin[950] ), .IN1(creg[951]), .SEL(start_in[0]), 
        .F(\modmult_1/N1980 ) );
  ANDN U5965 ( .A(n4110), .B(n3717), .Z(\modmult_1/N198 ) );
  XOR U5966 ( .A(n5887), .B(n5888), .Z(n3717) );
  MUX U5967 ( .IN0(\modmult_1/xin[949] ), .IN1(creg[950]), .SEL(start_in[0]), 
        .F(\modmult_1/N1979 ) );
  MUX U5968 ( .IN0(\modmult_1/xin[948] ), .IN1(creg[949]), .SEL(start_in[0]), 
        .F(\modmult_1/N1978 ) );
  MUX U5969 ( .IN0(\modmult_1/xin[947] ), .IN1(creg[948]), .SEL(start_in[0]), 
        .F(\modmult_1/N1977 ) );
  MUX U5970 ( .IN0(\modmult_1/xin[946] ), .IN1(creg[947]), .SEL(start_in[0]), 
        .F(\modmult_1/N1976 ) );
  MUX U5971 ( .IN0(\modmult_1/xin[945] ), .IN1(creg[946]), .SEL(start_in[0]), 
        .F(\modmult_1/N1975 ) );
  MUX U5972 ( .IN0(\modmult_1/xin[944] ), .IN1(creg[945]), .SEL(start_in[0]), 
        .F(\modmult_1/N1974 ) );
  MUX U5973 ( .IN0(\modmult_1/xin[943] ), .IN1(creg[944]), .SEL(start_in[0]), 
        .F(\modmult_1/N1973 ) );
  MUX U5974 ( .IN0(\modmult_1/xin[942] ), .IN1(creg[943]), .SEL(start_in[0]), 
        .F(\modmult_1/N1972 ) );
  MUX U5975 ( .IN0(\modmult_1/xin[941] ), .IN1(creg[942]), .SEL(start_in[0]), 
        .F(\modmult_1/N1971 ) );
  MUX U5976 ( .IN0(\modmult_1/xin[940] ), .IN1(creg[941]), .SEL(start_in[0]), 
        .F(\modmult_1/N1970 ) );
  ANDN U5977 ( .A(n4110), .B(n3720), .Z(\modmult_1/N197 ) );
  XOR U5978 ( .A(n5889), .B(n5890), .Z(n3720) );
  MUX U5979 ( .IN0(\modmult_1/xin[939] ), .IN1(creg[940]), .SEL(start_in[0]), 
        .F(\modmult_1/N1969 ) );
  MUX U5980 ( .IN0(\modmult_1/xin[938] ), .IN1(creg[939]), .SEL(start_in[0]), 
        .F(\modmult_1/N1968 ) );
  MUX U5981 ( .IN0(\modmult_1/xin[937] ), .IN1(creg[938]), .SEL(start_in[0]), 
        .F(\modmult_1/N1967 ) );
  MUX U5982 ( .IN0(\modmult_1/xin[936] ), .IN1(creg[937]), .SEL(start_in[0]), 
        .F(\modmult_1/N1966 ) );
  MUX U5983 ( .IN0(\modmult_1/xin[935] ), .IN1(creg[936]), .SEL(start_in[0]), 
        .F(\modmult_1/N1965 ) );
  MUX U5984 ( .IN0(\modmult_1/xin[934] ), .IN1(creg[935]), .SEL(start_in[0]), 
        .F(\modmult_1/N1964 ) );
  MUX U5985 ( .IN0(\modmult_1/xin[933] ), .IN1(creg[934]), .SEL(start_in[0]), 
        .F(\modmult_1/N1963 ) );
  MUX U5986 ( .IN0(\modmult_1/xin[932] ), .IN1(creg[933]), .SEL(start_in[0]), 
        .F(\modmult_1/N1962 ) );
  MUX U5987 ( .IN0(\modmult_1/xin[931] ), .IN1(creg[932]), .SEL(start_in[0]), 
        .F(\modmult_1/N1961 ) );
  MUX U5988 ( .IN0(\modmult_1/xin[930] ), .IN1(creg[931]), .SEL(start_in[0]), 
        .F(\modmult_1/N1960 ) );
  ANDN U5989 ( .A(n4110), .B(n3723), .Z(\modmult_1/N196 ) );
  XOR U5990 ( .A(n5891), .B(n5892), .Z(n3723) );
  MUX U5991 ( .IN0(\modmult_1/xin[929] ), .IN1(creg[930]), .SEL(start_in[0]), 
        .F(\modmult_1/N1959 ) );
  MUX U5992 ( .IN0(\modmult_1/xin[928] ), .IN1(creg[929]), .SEL(start_in[0]), 
        .F(\modmult_1/N1958 ) );
  MUX U5993 ( .IN0(\modmult_1/xin[927] ), .IN1(creg[928]), .SEL(start_in[0]), 
        .F(\modmult_1/N1957 ) );
  MUX U5994 ( .IN0(\modmult_1/xin[926] ), .IN1(creg[927]), .SEL(start_in[0]), 
        .F(\modmult_1/N1956 ) );
  MUX U5995 ( .IN0(\modmult_1/xin[925] ), .IN1(creg[926]), .SEL(start_in[0]), 
        .F(\modmult_1/N1955 ) );
  MUX U5996 ( .IN0(\modmult_1/xin[924] ), .IN1(creg[925]), .SEL(start_in[0]), 
        .F(\modmult_1/N1954 ) );
  MUX U5997 ( .IN0(\modmult_1/xin[923] ), .IN1(creg[924]), .SEL(start_in[0]), 
        .F(\modmult_1/N1953 ) );
  MUX U5998 ( .IN0(\modmult_1/xin[922] ), .IN1(creg[923]), .SEL(start_in[0]), 
        .F(\modmult_1/N1952 ) );
  MUX U5999 ( .IN0(\modmult_1/xin[921] ), .IN1(creg[922]), .SEL(start_in[0]), 
        .F(\modmult_1/N1951 ) );
  MUX U6000 ( .IN0(\modmult_1/xin[920] ), .IN1(creg[921]), .SEL(start_in[0]), 
        .F(\modmult_1/N1950 ) );
  ANDN U6001 ( .A(n4110), .B(n3726), .Z(\modmult_1/N195 ) );
  XOR U6002 ( .A(n5893), .B(n5894), .Z(n3726) );
  MUX U6003 ( .IN0(\modmult_1/xin[919] ), .IN1(creg[920]), .SEL(start_in[0]), 
        .F(\modmult_1/N1949 ) );
  MUX U6004 ( .IN0(\modmult_1/xin[918] ), .IN1(creg[919]), .SEL(start_in[0]), 
        .F(\modmult_1/N1948 ) );
  MUX U6005 ( .IN0(\modmult_1/xin[917] ), .IN1(creg[918]), .SEL(start_in[0]), 
        .F(\modmult_1/N1947 ) );
  MUX U6006 ( .IN0(\modmult_1/xin[916] ), .IN1(creg[917]), .SEL(start_in[0]), 
        .F(\modmult_1/N1946 ) );
  MUX U6007 ( .IN0(\modmult_1/xin[915] ), .IN1(creg[916]), .SEL(start_in[0]), 
        .F(\modmult_1/N1945 ) );
  MUX U6008 ( .IN0(\modmult_1/xin[914] ), .IN1(creg[915]), .SEL(start_in[0]), 
        .F(\modmult_1/N1944 ) );
  MUX U6009 ( .IN0(\modmult_1/xin[913] ), .IN1(creg[914]), .SEL(start_in[0]), 
        .F(\modmult_1/N1943 ) );
  MUX U6010 ( .IN0(\modmult_1/xin[912] ), .IN1(creg[913]), .SEL(start_in[0]), 
        .F(\modmult_1/N1942 ) );
  MUX U6011 ( .IN0(\modmult_1/xin[911] ), .IN1(creg[912]), .SEL(start_in[0]), 
        .F(\modmult_1/N1941 ) );
  MUX U6012 ( .IN0(\modmult_1/xin[910] ), .IN1(creg[911]), .SEL(start_in[0]), 
        .F(\modmult_1/N1940 ) );
  ANDN U6013 ( .A(n4110), .B(n3729), .Z(\modmult_1/N194 ) );
  XOR U6014 ( .A(n5895), .B(n5896), .Z(n3729) );
  MUX U6015 ( .IN0(\modmult_1/xin[909] ), .IN1(creg[910]), .SEL(start_in[0]), 
        .F(\modmult_1/N1939 ) );
  MUX U6016 ( .IN0(\modmult_1/xin[908] ), .IN1(creg[909]), .SEL(start_in[0]), 
        .F(\modmult_1/N1938 ) );
  MUX U6017 ( .IN0(\modmult_1/xin[907] ), .IN1(creg[908]), .SEL(start_in[0]), 
        .F(\modmult_1/N1937 ) );
  MUX U6018 ( .IN0(\modmult_1/xin[906] ), .IN1(creg[907]), .SEL(start_in[0]), 
        .F(\modmult_1/N1936 ) );
  MUX U6019 ( .IN0(\modmult_1/xin[905] ), .IN1(creg[906]), .SEL(start_in[0]), 
        .F(\modmult_1/N1935 ) );
  MUX U6020 ( .IN0(\modmult_1/xin[904] ), .IN1(creg[905]), .SEL(start_in[0]), 
        .F(\modmult_1/N1934 ) );
  MUX U6021 ( .IN0(\modmult_1/xin[903] ), .IN1(creg[904]), .SEL(start_in[0]), 
        .F(\modmult_1/N1933 ) );
  MUX U6022 ( .IN0(\modmult_1/xin[902] ), .IN1(creg[903]), .SEL(start_in[0]), 
        .F(\modmult_1/N1932 ) );
  MUX U6023 ( .IN0(\modmult_1/xin[901] ), .IN1(creg[902]), .SEL(start_in[0]), 
        .F(\modmult_1/N1931 ) );
  MUX U6024 ( .IN0(\modmult_1/xin[900] ), .IN1(creg[901]), .SEL(start_in[0]), 
        .F(\modmult_1/N1930 ) );
  ANDN U6025 ( .A(n4110), .B(n3732), .Z(\modmult_1/N193 ) );
  XOR U6026 ( .A(n5897), .B(n5898), .Z(n3732) );
  MUX U6027 ( .IN0(\modmult_1/xin[899] ), .IN1(creg[900]), .SEL(start_in[0]), 
        .F(\modmult_1/N1929 ) );
  MUX U6028 ( .IN0(\modmult_1/xin[898] ), .IN1(creg[899]), .SEL(start_in[0]), 
        .F(\modmult_1/N1928 ) );
  MUX U6029 ( .IN0(\modmult_1/xin[897] ), .IN1(creg[898]), .SEL(start_in[0]), 
        .F(\modmult_1/N1927 ) );
  MUX U6030 ( .IN0(\modmult_1/xin[896] ), .IN1(creg[897]), .SEL(start_in[0]), 
        .F(\modmult_1/N1926 ) );
  MUX U6031 ( .IN0(\modmult_1/xin[895] ), .IN1(creg[896]), .SEL(start_in[0]), 
        .F(\modmult_1/N1925 ) );
  MUX U6032 ( .IN0(\modmult_1/xin[894] ), .IN1(creg[895]), .SEL(start_in[0]), 
        .F(\modmult_1/N1924 ) );
  MUX U6033 ( .IN0(\modmult_1/xin[893] ), .IN1(creg[894]), .SEL(start_in[0]), 
        .F(\modmult_1/N1923 ) );
  MUX U6034 ( .IN0(\modmult_1/xin[892] ), .IN1(creg[893]), .SEL(start_in[0]), 
        .F(\modmult_1/N1922 ) );
  MUX U6035 ( .IN0(\modmult_1/xin[891] ), .IN1(creg[892]), .SEL(start_in[0]), 
        .F(\modmult_1/N1921 ) );
  MUX U6036 ( .IN0(\modmult_1/xin[890] ), .IN1(creg[891]), .SEL(start_in[0]), 
        .F(\modmult_1/N1920 ) );
  ANDN U6037 ( .A(n4110), .B(n3738), .Z(\modmult_1/N192 ) );
  XOR U6038 ( .A(n5899), .B(n5900), .Z(n3738) );
  MUX U6039 ( .IN0(\modmult_1/xin[889] ), .IN1(creg[890]), .SEL(start_in[0]), 
        .F(\modmult_1/N1919 ) );
  MUX U6040 ( .IN0(\modmult_1/xin[888] ), .IN1(creg[889]), .SEL(start_in[0]), 
        .F(\modmult_1/N1918 ) );
  MUX U6041 ( .IN0(\modmult_1/xin[887] ), .IN1(creg[888]), .SEL(start_in[0]), 
        .F(\modmult_1/N1917 ) );
  MUX U6042 ( .IN0(\modmult_1/xin[886] ), .IN1(creg[887]), .SEL(start_in[0]), 
        .F(\modmult_1/N1916 ) );
  MUX U6043 ( .IN0(\modmult_1/xin[885] ), .IN1(creg[886]), .SEL(start_in[0]), 
        .F(\modmult_1/N1915 ) );
  MUX U6044 ( .IN0(\modmult_1/xin[884] ), .IN1(creg[885]), .SEL(start_in[0]), 
        .F(\modmult_1/N1914 ) );
  MUX U6045 ( .IN0(\modmult_1/xin[883] ), .IN1(creg[884]), .SEL(start_in[0]), 
        .F(\modmult_1/N1913 ) );
  MUX U6046 ( .IN0(\modmult_1/xin[882] ), .IN1(creg[883]), .SEL(start_in[0]), 
        .F(\modmult_1/N1912 ) );
  MUX U6047 ( .IN0(\modmult_1/xin[881] ), .IN1(creg[882]), .SEL(start_in[0]), 
        .F(\modmult_1/N1911 ) );
  MUX U6048 ( .IN0(\modmult_1/xin[880] ), .IN1(creg[881]), .SEL(start_in[0]), 
        .F(\modmult_1/N1910 ) );
  ANDN U6049 ( .A(n4110), .B(n3741), .Z(\modmult_1/N191 ) );
  XOR U6050 ( .A(n5901), .B(n5902), .Z(n3741) );
  MUX U6051 ( .IN0(\modmult_1/xin[879] ), .IN1(creg[880]), .SEL(start_in[0]), 
        .F(\modmult_1/N1909 ) );
  MUX U6052 ( .IN0(\modmult_1/xin[878] ), .IN1(creg[879]), .SEL(start_in[0]), 
        .F(\modmult_1/N1908 ) );
  MUX U6053 ( .IN0(\modmult_1/xin[877] ), .IN1(creg[878]), .SEL(start_in[0]), 
        .F(\modmult_1/N1907 ) );
  MUX U6054 ( .IN0(\modmult_1/xin[876] ), .IN1(creg[877]), .SEL(start_in[0]), 
        .F(\modmult_1/N1906 ) );
  MUX U6055 ( .IN0(\modmult_1/xin[875] ), .IN1(creg[876]), .SEL(start_in[0]), 
        .F(\modmult_1/N1905 ) );
  MUX U6056 ( .IN0(\modmult_1/xin[874] ), .IN1(creg[875]), .SEL(start_in[0]), 
        .F(\modmult_1/N1904 ) );
  MUX U6057 ( .IN0(\modmult_1/xin[873] ), .IN1(creg[874]), .SEL(start_in[0]), 
        .F(\modmult_1/N1903 ) );
  MUX U6058 ( .IN0(\modmult_1/xin[872] ), .IN1(creg[873]), .SEL(start_in[0]), 
        .F(\modmult_1/N1902 ) );
  MUX U6059 ( .IN0(\modmult_1/xin[871] ), .IN1(creg[872]), .SEL(start_in[0]), 
        .F(\modmult_1/N1901 ) );
  MUX U6060 ( .IN0(\modmult_1/xin[870] ), .IN1(creg[871]), .SEL(start_in[0]), 
        .F(\modmult_1/N1900 ) );
  ANDN U6061 ( .A(n4110), .B(n3744), .Z(\modmult_1/N190 ) );
  XOR U6062 ( .A(n5903), .B(n5904), .Z(n3744) );
  ANDN U6063 ( .A(n4110), .B(n3801), .Z(\modmult_1/N19 ) );
  XOR U6064 ( .A(n5905), .B(n5906), .Z(n3801) );
  MUX U6065 ( .IN0(\modmult_1/xin[869] ), .IN1(creg[870]), .SEL(start_in[0]), 
        .F(\modmult_1/N1899 ) );
  MUX U6066 ( .IN0(\modmult_1/xin[868] ), .IN1(creg[869]), .SEL(start_in[0]), 
        .F(\modmult_1/N1898 ) );
  MUX U6067 ( .IN0(\modmult_1/xin[867] ), .IN1(creg[868]), .SEL(start_in[0]), 
        .F(\modmult_1/N1897 ) );
  MUX U6068 ( .IN0(\modmult_1/xin[866] ), .IN1(creg[867]), .SEL(start_in[0]), 
        .F(\modmult_1/N1896 ) );
  MUX U6069 ( .IN0(\modmult_1/xin[865] ), .IN1(creg[866]), .SEL(start_in[0]), 
        .F(\modmult_1/N1895 ) );
  MUX U6070 ( .IN0(\modmult_1/xin[864] ), .IN1(creg[865]), .SEL(start_in[0]), 
        .F(\modmult_1/N1894 ) );
  MUX U6071 ( .IN0(\modmult_1/xin[863] ), .IN1(creg[864]), .SEL(start_in[0]), 
        .F(\modmult_1/N1893 ) );
  MUX U6072 ( .IN0(\modmult_1/xin[862] ), .IN1(creg[863]), .SEL(start_in[0]), 
        .F(\modmult_1/N1892 ) );
  MUX U6073 ( .IN0(\modmult_1/xin[861] ), .IN1(creg[862]), .SEL(start_in[0]), 
        .F(\modmult_1/N1891 ) );
  MUX U6074 ( .IN0(\modmult_1/xin[860] ), .IN1(creg[861]), .SEL(start_in[0]), 
        .F(\modmult_1/N1890 ) );
  ANDN U6075 ( .A(n4110), .B(n3747), .Z(\modmult_1/N189 ) );
  XOR U6076 ( .A(n5907), .B(n5908), .Z(n3747) );
  MUX U6077 ( .IN0(\modmult_1/xin[859] ), .IN1(creg[860]), .SEL(start_in[0]), 
        .F(\modmult_1/N1889 ) );
  MUX U6078 ( .IN0(\modmult_1/xin[858] ), .IN1(creg[859]), .SEL(start_in[0]), 
        .F(\modmult_1/N1888 ) );
  MUX U6079 ( .IN0(\modmult_1/xin[857] ), .IN1(creg[858]), .SEL(start_in[0]), 
        .F(\modmult_1/N1887 ) );
  MUX U6080 ( .IN0(\modmult_1/xin[856] ), .IN1(creg[857]), .SEL(start_in[0]), 
        .F(\modmult_1/N1886 ) );
  MUX U6081 ( .IN0(\modmult_1/xin[855] ), .IN1(creg[856]), .SEL(start_in[0]), 
        .F(\modmult_1/N1885 ) );
  MUX U6082 ( .IN0(\modmult_1/xin[854] ), .IN1(creg[855]), .SEL(start_in[0]), 
        .F(\modmult_1/N1884 ) );
  MUX U6083 ( .IN0(\modmult_1/xin[853] ), .IN1(creg[854]), .SEL(start_in[0]), 
        .F(\modmult_1/N1883 ) );
  MUX U6084 ( .IN0(\modmult_1/xin[852] ), .IN1(creg[853]), .SEL(start_in[0]), 
        .F(\modmult_1/N1882 ) );
  MUX U6085 ( .IN0(\modmult_1/xin[851] ), .IN1(creg[852]), .SEL(start_in[0]), 
        .F(\modmult_1/N1881 ) );
  MUX U6086 ( .IN0(\modmult_1/xin[850] ), .IN1(creg[851]), .SEL(start_in[0]), 
        .F(\modmult_1/N1880 ) );
  ANDN U6087 ( .A(n4110), .B(n3750), .Z(\modmult_1/N188 ) );
  XOR U6088 ( .A(n5909), .B(n5910), .Z(n3750) );
  MUX U6089 ( .IN0(\modmult_1/xin[849] ), .IN1(creg[850]), .SEL(start_in[0]), 
        .F(\modmult_1/N1879 ) );
  MUX U6090 ( .IN0(\modmult_1/xin[848] ), .IN1(creg[849]), .SEL(start_in[0]), 
        .F(\modmult_1/N1878 ) );
  MUX U6091 ( .IN0(\modmult_1/xin[847] ), .IN1(creg[848]), .SEL(start_in[0]), 
        .F(\modmult_1/N1877 ) );
  MUX U6092 ( .IN0(\modmult_1/xin[846] ), .IN1(creg[847]), .SEL(start_in[0]), 
        .F(\modmult_1/N1876 ) );
  MUX U6093 ( .IN0(\modmult_1/xin[845] ), .IN1(creg[846]), .SEL(start_in[0]), 
        .F(\modmult_1/N1875 ) );
  MUX U6094 ( .IN0(\modmult_1/xin[844] ), .IN1(creg[845]), .SEL(start_in[0]), 
        .F(\modmult_1/N1874 ) );
  MUX U6095 ( .IN0(\modmult_1/xin[843] ), .IN1(creg[844]), .SEL(start_in[0]), 
        .F(\modmult_1/N1873 ) );
  MUX U6096 ( .IN0(\modmult_1/xin[842] ), .IN1(creg[843]), .SEL(start_in[0]), 
        .F(\modmult_1/N1872 ) );
  MUX U6097 ( .IN0(\modmult_1/xin[841] ), .IN1(creg[842]), .SEL(start_in[0]), 
        .F(\modmult_1/N1871 ) );
  MUX U6098 ( .IN0(\modmult_1/xin[840] ), .IN1(creg[841]), .SEL(start_in[0]), 
        .F(\modmult_1/N1870 ) );
  ANDN U6099 ( .A(n4110), .B(n3753), .Z(\modmult_1/N187 ) );
  XOR U6100 ( .A(n5911), .B(n5912), .Z(n3753) );
  MUX U6101 ( .IN0(\modmult_1/xin[839] ), .IN1(creg[840]), .SEL(start_in[0]), 
        .F(\modmult_1/N1869 ) );
  MUX U6102 ( .IN0(\modmult_1/xin[838] ), .IN1(creg[839]), .SEL(start_in[0]), 
        .F(\modmult_1/N1868 ) );
  MUX U6103 ( .IN0(\modmult_1/xin[837] ), .IN1(creg[838]), .SEL(start_in[0]), 
        .F(\modmult_1/N1867 ) );
  MUX U6104 ( .IN0(\modmult_1/xin[836] ), .IN1(creg[837]), .SEL(start_in[0]), 
        .F(\modmult_1/N1866 ) );
  MUX U6105 ( .IN0(\modmult_1/xin[835] ), .IN1(creg[836]), .SEL(start_in[0]), 
        .F(\modmult_1/N1865 ) );
  MUX U6106 ( .IN0(\modmult_1/xin[834] ), .IN1(creg[835]), .SEL(start_in[0]), 
        .F(\modmult_1/N1864 ) );
  MUX U6107 ( .IN0(\modmult_1/xin[833] ), .IN1(creg[834]), .SEL(start_in[0]), 
        .F(\modmult_1/N1863 ) );
  MUX U6108 ( .IN0(\modmult_1/xin[832] ), .IN1(creg[833]), .SEL(start_in[0]), 
        .F(\modmult_1/N1862 ) );
  MUX U6109 ( .IN0(\modmult_1/xin[831] ), .IN1(creg[832]), .SEL(start_in[0]), 
        .F(\modmult_1/N1861 ) );
  MUX U6110 ( .IN0(\modmult_1/xin[830] ), .IN1(creg[831]), .SEL(start_in[0]), 
        .F(\modmult_1/N1860 ) );
  ANDN U6111 ( .A(n4110), .B(n3756), .Z(\modmult_1/N186 ) );
  XOR U6112 ( .A(n5913), .B(n5914), .Z(n3756) );
  MUX U6113 ( .IN0(\modmult_1/xin[829] ), .IN1(creg[830]), .SEL(start_in[0]), 
        .F(\modmult_1/N1859 ) );
  MUX U6114 ( .IN0(\modmult_1/xin[828] ), .IN1(creg[829]), .SEL(start_in[0]), 
        .F(\modmult_1/N1858 ) );
  MUX U6115 ( .IN0(\modmult_1/xin[827] ), .IN1(creg[828]), .SEL(start_in[0]), 
        .F(\modmult_1/N1857 ) );
  MUX U6116 ( .IN0(\modmult_1/xin[826] ), .IN1(creg[827]), .SEL(start_in[0]), 
        .F(\modmult_1/N1856 ) );
  MUX U6117 ( .IN0(\modmult_1/xin[825] ), .IN1(creg[826]), .SEL(start_in[0]), 
        .F(\modmult_1/N1855 ) );
  MUX U6118 ( .IN0(\modmult_1/xin[824] ), .IN1(creg[825]), .SEL(start_in[0]), 
        .F(\modmult_1/N1854 ) );
  MUX U6119 ( .IN0(\modmult_1/xin[823] ), .IN1(creg[824]), .SEL(start_in[0]), 
        .F(\modmult_1/N1853 ) );
  MUX U6120 ( .IN0(\modmult_1/xin[822] ), .IN1(creg[823]), .SEL(start_in[0]), 
        .F(\modmult_1/N1852 ) );
  MUX U6121 ( .IN0(\modmult_1/xin[821] ), .IN1(creg[822]), .SEL(start_in[0]), 
        .F(\modmult_1/N1851 ) );
  MUX U6122 ( .IN0(\modmult_1/xin[820] ), .IN1(creg[821]), .SEL(start_in[0]), 
        .F(\modmult_1/N1850 ) );
  ANDN U6123 ( .A(n4110), .B(n3759), .Z(\modmult_1/N185 ) );
  XOR U6124 ( .A(n5915), .B(n5916), .Z(n3759) );
  MUX U6125 ( .IN0(\modmult_1/xin[819] ), .IN1(creg[820]), .SEL(start_in[0]), 
        .F(\modmult_1/N1849 ) );
  MUX U6126 ( .IN0(\modmult_1/xin[818] ), .IN1(creg[819]), .SEL(start_in[0]), 
        .F(\modmult_1/N1848 ) );
  MUX U6127 ( .IN0(\modmult_1/xin[817] ), .IN1(creg[818]), .SEL(start_in[0]), 
        .F(\modmult_1/N1847 ) );
  MUX U6128 ( .IN0(\modmult_1/xin[816] ), .IN1(creg[817]), .SEL(start_in[0]), 
        .F(\modmult_1/N1846 ) );
  MUX U6129 ( .IN0(\modmult_1/xin[815] ), .IN1(creg[816]), .SEL(start_in[0]), 
        .F(\modmult_1/N1845 ) );
  MUX U6130 ( .IN0(\modmult_1/xin[814] ), .IN1(creg[815]), .SEL(start_in[0]), 
        .F(\modmult_1/N1844 ) );
  MUX U6131 ( .IN0(\modmult_1/xin[813] ), .IN1(creg[814]), .SEL(start_in[0]), 
        .F(\modmult_1/N1843 ) );
  MUX U6132 ( .IN0(\modmult_1/xin[812] ), .IN1(creg[813]), .SEL(start_in[0]), 
        .F(\modmult_1/N1842 ) );
  MUX U6133 ( .IN0(\modmult_1/xin[811] ), .IN1(creg[812]), .SEL(start_in[0]), 
        .F(\modmult_1/N1841 ) );
  MUX U6134 ( .IN0(\modmult_1/xin[810] ), .IN1(creg[811]), .SEL(start_in[0]), 
        .F(\modmult_1/N1840 ) );
  ANDN U6135 ( .A(n4110), .B(n3762), .Z(\modmult_1/N184 ) );
  XOR U6136 ( .A(n5917), .B(n5918), .Z(n3762) );
  MUX U6137 ( .IN0(\modmult_1/xin[809] ), .IN1(creg[810]), .SEL(start_in[0]), 
        .F(\modmult_1/N1839 ) );
  MUX U6138 ( .IN0(\modmult_1/xin[808] ), .IN1(creg[809]), .SEL(start_in[0]), 
        .F(\modmult_1/N1838 ) );
  MUX U6139 ( .IN0(\modmult_1/xin[807] ), .IN1(creg[808]), .SEL(start_in[0]), 
        .F(\modmult_1/N1837 ) );
  MUX U6140 ( .IN0(\modmult_1/xin[806] ), .IN1(creg[807]), .SEL(start_in[0]), 
        .F(\modmult_1/N1836 ) );
  MUX U6141 ( .IN0(\modmult_1/xin[805] ), .IN1(creg[806]), .SEL(start_in[0]), 
        .F(\modmult_1/N1835 ) );
  MUX U6142 ( .IN0(\modmult_1/xin[804] ), .IN1(creg[805]), .SEL(start_in[0]), 
        .F(\modmult_1/N1834 ) );
  MUX U6143 ( .IN0(\modmult_1/xin[803] ), .IN1(creg[804]), .SEL(start_in[0]), 
        .F(\modmult_1/N1833 ) );
  MUX U6144 ( .IN0(\modmult_1/xin[802] ), .IN1(creg[803]), .SEL(start_in[0]), 
        .F(\modmult_1/N1832 ) );
  MUX U6145 ( .IN0(\modmult_1/xin[801] ), .IN1(creg[802]), .SEL(start_in[0]), 
        .F(\modmult_1/N1831 ) );
  MUX U6146 ( .IN0(\modmult_1/xin[800] ), .IN1(creg[801]), .SEL(start_in[0]), 
        .F(\modmult_1/N1830 ) );
  ANDN U6147 ( .A(n4110), .B(n3765), .Z(\modmult_1/N183 ) );
  XOR U6148 ( .A(n5919), .B(n5920), .Z(n3765) );
  MUX U6149 ( .IN0(\modmult_1/xin[799] ), .IN1(creg[800]), .SEL(start_in[0]), 
        .F(\modmult_1/N1829 ) );
  MUX U6150 ( .IN0(\modmult_1/xin[798] ), .IN1(creg[799]), .SEL(start_in[0]), 
        .F(\modmult_1/N1828 ) );
  MUX U6151 ( .IN0(\modmult_1/xin[797] ), .IN1(creg[798]), .SEL(start_in[0]), 
        .F(\modmult_1/N1827 ) );
  MUX U6152 ( .IN0(\modmult_1/xin[796] ), .IN1(creg[797]), .SEL(start_in[0]), 
        .F(\modmult_1/N1826 ) );
  MUX U6153 ( .IN0(\modmult_1/xin[795] ), .IN1(creg[796]), .SEL(start_in[0]), 
        .F(\modmult_1/N1825 ) );
  MUX U6154 ( .IN0(\modmult_1/xin[794] ), .IN1(creg[795]), .SEL(start_in[0]), 
        .F(\modmult_1/N1824 ) );
  MUX U6155 ( .IN0(\modmult_1/xin[793] ), .IN1(creg[794]), .SEL(start_in[0]), 
        .F(\modmult_1/N1823 ) );
  MUX U6156 ( .IN0(\modmult_1/xin[792] ), .IN1(creg[793]), .SEL(start_in[0]), 
        .F(\modmult_1/N1822 ) );
  MUX U6157 ( .IN0(\modmult_1/xin[791] ), .IN1(creg[792]), .SEL(start_in[0]), 
        .F(\modmult_1/N1821 ) );
  MUX U6158 ( .IN0(\modmult_1/xin[790] ), .IN1(creg[791]), .SEL(start_in[0]), 
        .F(\modmult_1/N1820 ) );
  ANDN U6159 ( .A(n4110), .B(n3771), .Z(\modmult_1/N182 ) );
  XOR U6160 ( .A(n5921), .B(n5922), .Z(n3771) );
  MUX U6161 ( .IN0(\modmult_1/xin[789] ), .IN1(creg[790]), .SEL(start_in[0]), 
        .F(\modmult_1/N1819 ) );
  MUX U6162 ( .IN0(\modmult_1/xin[788] ), .IN1(creg[789]), .SEL(start_in[0]), 
        .F(\modmult_1/N1818 ) );
  MUX U6163 ( .IN0(\modmult_1/xin[787] ), .IN1(creg[788]), .SEL(start_in[0]), 
        .F(\modmult_1/N1817 ) );
  MUX U6164 ( .IN0(\modmult_1/xin[786] ), .IN1(creg[787]), .SEL(start_in[0]), 
        .F(\modmult_1/N1816 ) );
  MUX U6165 ( .IN0(\modmult_1/xin[785] ), .IN1(creg[786]), .SEL(start_in[0]), 
        .F(\modmult_1/N1815 ) );
  MUX U6166 ( .IN0(\modmult_1/xin[784] ), .IN1(creg[785]), .SEL(start_in[0]), 
        .F(\modmult_1/N1814 ) );
  MUX U6167 ( .IN0(\modmult_1/xin[783] ), .IN1(creg[784]), .SEL(start_in[0]), 
        .F(\modmult_1/N1813 ) );
  MUX U6168 ( .IN0(\modmult_1/xin[782] ), .IN1(creg[783]), .SEL(start_in[0]), 
        .F(\modmult_1/N1812 ) );
  MUX U6169 ( .IN0(\modmult_1/xin[781] ), .IN1(creg[782]), .SEL(start_in[0]), 
        .F(\modmult_1/N1811 ) );
  MUX U6170 ( .IN0(\modmult_1/xin[780] ), .IN1(creg[781]), .SEL(start_in[0]), 
        .F(\modmult_1/N1810 ) );
  ANDN U6171 ( .A(n4110), .B(n3774), .Z(\modmult_1/N181 ) );
  XOR U6172 ( .A(n5923), .B(n5924), .Z(n3774) );
  MUX U6173 ( .IN0(\modmult_1/xin[779] ), .IN1(creg[780]), .SEL(start_in[0]), 
        .F(\modmult_1/N1809 ) );
  MUX U6174 ( .IN0(\modmult_1/xin[778] ), .IN1(creg[779]), .SEL(start_in[0]), 
        .F(\modmult_1/N1808 ) );
  MUX U6175 ( .IN0(\modmult_1/xin[777] ), .IN1(creg[778]), .SEL(start_in[0]), 
        .F(\modmult_1/N1807 ) );
  MUX U6176 ( .IN0(\modmult_1/xin[776] ), .IN1(creg[777]), .SEL(start_in[0]), 
        .F(\modmult_1/N1806 ) );
  MUX U6177 ( .IN0(\modmult_1/xin[775] ), .IN1(creg[776]), .SEL(start_in[0]), 
        .F(\modmult_1/N1805 ) );
  MUX U6178 ( .IN0(\modmult_1/xin[774] ), .IN1(creg[775]), .SEL(start_in[0]), 
        .F(\modmult_1/N1804 ) );
  MUX U6179 ( .IN0(\modmult_1/xin[773] ), .IN1(creg[774]), .SEL(start_in[0]), 
        .F(\modmult_1/N1803 ) );
  MUX U6180 ( .IN0(\modmult_1/xin[772] ), .IN1(creg[773]), .SEL(start_in[0]), 
        .F(\modmult_1/N1802 ) );
  MUX U6181 ( .IN0(\modmult_1/xin[771] ), .IN1(creg[772]), .SEL(start_in[0]), 
        .F(\modmult_1/N1801 ) );
  MUX U6182 ( .IN0(\modmult_1/xin[770] ), .IN1(creg[771]), .SEL(start_in[0]), 
        .F(\modmult_1/N1800 ) );
  ANDN U6183 ( .A(n4110), .B(n3777), .Z(\modmult_1/N180 ) );
  XOR U6184 ( .A(n5925), .B(n5926), .Z(n3777) );
  ANDN U6185 ( .A(n4110), .B(n3834), .Z(\modmult_1/N18 ) );
  XOR U6186 ( .A(n5927), .B(n5928), .Z(n3834) );
  MUX U6187 ( .IN0(\modmult_1/xin[769] ), .IN1(creg[770]), .SEL(start_in[0]), 
        .F(\modmult_1/N1799 ) );
  MUX U6188 ( .IN0(\modmult_1/xin[768] ), .IN1(creg[769]), .SEL(start_in[0]), 
        .F(\modmult_1/N1798 ) );
  MUX U6189 ( .IN0(\modmult_1/xin[767] ), .IN1(creg[768]), .SEL(start_in[0]), 
        .F(\modmult_1/N1797 ) );
  MUX U6190 ( .IN0(\modmult_1/xin[766] ), .IN1(creg[767]), .SEL(start_in[0]), 
        .F(\modmult_1/N1796 ) );
  MUX U6191 ( .IN0(\modmult_1/xin[765] ), .IN1(creg[766]), .SEL(start_in[0]), 
        .F(\modmult_1/N1795 ) );
  MUX U6192 ( .IN0(\modmult_1/xin[764] ), .IN1(creg[765]), .SEL(start_in[0]), 
        .F(\modmult_1/N1794 ) );
  MUX U6193 ( .IN0(\modmult_1/xin[763] ), .IN1(creg[764]), .SEL(start_in[0]), 
        .F(\modmult_1/N1793 ) );
  MUX U6194 ( .IN0(\modmult_1/xin[762] ), .IN1(creg[763]), .SEL(start_in[0]), 
        .F(\modmult_1/N1792 ) );
  MUX U6195 ( .IN0(\modmult_1/xin[761] ), .IN1(creg[762]), .SEL(start_in[0]), 
        .F(\modmult_1/N1791 ) );
  MUX U6196 ( .IN0(\modmult_1/xin[760] ), .IN1(creg[761]), .SEL(start_in[0]), 
        .F(\modmult_1/N1790 ) );
  ANDN U6197 ( .A(n4110), .B(n3780), .Z(\modmult_1/N179 ) );
  XOR U6198 ( .A(n5929), .B(n5930), .Z(n3780) );
  MUX U6199 ( .IN0(\modmult_1/xin[759] ), .IN1(creg[760]), .SEL(start_in[0]), 
        .F(\modmult_1/N1789 ) );
  MUX U6200 ( .IN0(\modmult_1/xin[758] ), .IN1(creg[759]), .SEL(start_in[0]), 
        .F(\modmult_1/N1788 ) );
  MUX U6201 ( .IN0(\modmult_1/xin[757] ), .IN1(creg[758]), .SEL(start_in[0]), 
        .F(\modmult_1/N1787 ) );
  MUX U6202 ( .IN0(\modmult_1/xin[756] ), .IN1(creg[757]), .SEL(start_in[0]), 
        .F(\modmult_1/N1786 ) );
  MUX U6203 ( .IN0(\modmult_1/xin[755] ), .IN1(creg[756]), .SEL(start_in[0]), 
        .F(\modmult_1/N1785 ) );
  MUX U6204 ( .IN0(\modmult_1/xin[754] ), .IN1(creg[755]), .SEL(start_in[0]), 
        .F(\modmult_1/N1784 ) );
  MUX U6205 ( .IN0(\modmult_1/xin[753] ), .IN1(creg[754]), .SEL(start_in[0]), 
        .F(\modmult_1/N1783 ) );
  MUX U6206 ( .IN0(\modmult_1/xin[752] ), .IN1(creg[753]), .SEL(start_in[0]), 
        .F(\modmult_1/N1782 ) );
  MUX U6207 ( .IN0(\modmult_1/xin[751] ), .IN1(creg[752]), .SEL(start_in[0]), 
        .F(\modmult_1/N1781 ) );
  MUX U6208 ( .IN0(\modmult_1/xin[750] ), .IN1(creg[751]), .SEL(start_in[0]), 
        .F(\modmult_1/N1780 ) );
  ANDN U6209 ( .A(n4110), .B(n3783), .Z(\modmult_1/N178 ) );
  XOR U6210 ( .A(n5931), .B(n5932), .Z(n3783) );
  MUX U6211 ( .IN0(\modmult_1/xin[749] ), .IN1(creg[750]), .SEL(start_in[0]), 
        .F(\modmult_1/N1779 ) );
  MUX U6212 ( .IN0(\modmult_1/xin[748] ), .IN1(creg[749]), .SEL(start_in[0]), 
        .F(\modmult_1/N1778 ) );
  MUX U6213 ( .IN0(\modmult_1/xin[747] ), .IN1(creg[748]), .SEL(start_in[0]), 
        .F(\modmult_1/N1777 ) );
  MUX U6214 ( .IN0(\modmult_1/xin[746] ), .IN1(creg[747]), .SEL(start_in[0]), 
        .F(\modmult_1/N1776 ) );
  MUX U6215 ( .IN0(\modmult_1/xin[745] ), .IN1(creg[746]), .SEL(start_in[0]), 
        .F(\modmult_1/N1775 ) );
  MUX U6216 ( .IN0(\modmult_1/xin[744] ), .IN1(creg[745]), .SEL(start_in[0]), 
        .F(\modmult_1/N1774 ) );
  MUX U6217 ( .IN0(\modmult_1/xin[743] ), .IN1(creg[744]), .SEL(start_in[0]), 
        .F(\modmult_1/N1773 ) );
  MUX U6218 ( .IN0(\modmult_1/xin[742] ), .IN1(creg[743]), .SEL(start_in[0]), 
        .F(\modmult_1/N1772 ) );
  MUX U6219 ( .IN0(\modmult_1/xin[741] ), .IN1(creg[742]), .SEL(start_in[0]), 
        .F(\modmult_1/N1771 ) );
  MUX U6220 ( .IN0(\modmult_1/xin[740] ), .IN1(creg[741]), .SEL(start_in[0]), 
        .F(\modmult_1/N1770 ) );
  ANDN U6221 ( .A(n4110), .B(n3786), .Z(\modmult_1/N177 ) );
  XOR U6222 ( .A(n5933), .B(n5934), .Z(n3786) );
  MUX U6223 ( .IN0(\modmult_1/xin[739] ), .IN1(creg[740]), .SEL(start_in[0]), 
        .F(\modmult_1/N1769 ) );
  MUX U6224 ( .IN0(\modmult_1/xin[738] ), .IN1(creg[739]), .SEL(start_in[0]), 
        .F(\modmult_1/N1768 ) );
  MUX U6225 ( .IN0(\modmult_1/xin[737] ), .IN1(creg[738]), .SEL(start_in[0]), 
        .F(\modmult_1/N1767 ) );
  MUX U6226 ( .IN0(\modmult_1/xin[736] ), .IN1(creg[737]), .SEL(start_in[0]), 
        .F(\modmult_1/N1766 ) );
  MUX U6227 ( .IN0(\modmult_1/xin[735] ), .IN1(creg[736]), .SEL(start_in[0]), 
        .F(\modmult_1/N1765 ) );
  MUX U6228 ( .IN0(\modmult_1/xin[734] ), .IN1(creg[735]), .SEL(start_in[0]), 
        .F(\modmult_1/N1764 ) );
  MUX U6229 ( .IN0(\modmult_1/xin[733] ), .IN1(creg[734]), .SEL(start_in[0]), 
        .F(\modmult_1/N1763 ) );
  MUX U6230 ( .IN0(\modmult_1/xin[732] ), .IN1(creg[733]), .SEL(start_in[0]), 
        .F(\modmult_1/N1762 ) );
  MUX U6231 ( .IN0(\modmult_1/xin[731] ), .IN1(creg[732]), .SEL(start_in[0]), 
        .F(\modmult_1/N1761 ) );
  MUX U6232 ( .IN0(\modmult_1/xin[730] ), .IN1(creg[731]), .SEL(start_in[0]), 
        .F(\modmult_1/N1760 ) );
  ANDN U6233 ( .A(n4110), .B(n3789), .Z(\modmult_1/N176 ) );
  XOR U6234 ( .A(n5935), .B(n5936), .Z(n3789) );
  MUX U6235 ( .IN0(\modmult_1/xin[729] ), .IN1(creg[730]), .SEL(start_in[0]), 
        .F(\modmult_1/N1759 ) );
  MUX U6236 ( .IN0(\modmult_1/xin[728] ), .IN1(creg[729]), .SEL(start_in[0]), 
        .F(\modmult_1/N1758 ) );
  MUX U6237 ( .IN0(\modmult_1/xin[727] ), .IN1(creg[728]), .SEL(start_in[0]), 
        .F(\modmult_1/N1757 ) );
  MUX U6238 ( .IN0(\modmult_1/xin[726] ), .IN1(creg[727]), .SEL(start_in[0]), 
        .F(\modmult_1/N1756 ) );
  MUX U6239 ( .IN0(\modmult_1/xin[725] ), .IN1(creg[726]), .SEL(start_in[0]), 
        .F(\modmult_1/N1755 ) );
  MUX U6240 ( .IN0(\modmult_1/xin[724] ), .IN1(creg[725]), .SEL(start_in[0]), 
        .F(\modmult_1/N1754 ) );
  MUX U6241 ( .IN0(\modmult_1/xin[723] ), .IN1(creg[724]), .SEL(start_in[0]), 
        .F(\modmult_1/N1753 ) );
  MUX U6242 ( .IN0(\modmult_1/xin[722] ), .IN1(creg[723]), .SEL(start_in[0]), 
        .F(\modmult_1/N1752 ) );
  MUX U6243 ( .IN0(\modmult_1/xin[721] ), .IN1(creg[722]), .SEL(start_in[0]), 
        .F(\modmult_1/N1751 ) );
  MUX U6244 ( .IN0(\modmult_1/xin[720] ), .IN1(creg[721]), .SEL(start_in[0]), 
        .F(\modmult_1/N1750 ) );
  ANDN U6245 ( .A(n4110), .B(n3792), .Z(\modmult_1/N175 ) );
  XOR U6246 ( .A(n5937), .B(n5938), .Z(n3792) );
  MUX U6247 ( .IN0(\modmult_1/xin[719] ), .IN1(creg[720]), .SEL(start_in[0]), 
        .F(\modmult_1/N1749 ) );
  MUX U6248 ( .IN0(\modmult_1/xin[718] ), .IN1(creg[719]), .SEL(start_in[0]), 
        .F(\modmult_1/N1748 ) );
  MUX U6249 ( .IN0(\modmult_1/xin[717] ), .IN1(creg[718]), .SEL(start_in[0]), 
        .F(\modmult_1/N1747 ) );
  MUX U6250 ( .IN0(\modmult_1/xin[716] ), .IN1(creg[717]), .SEL(start_in[0]), 
        .F(\modmult_1/N1746 ) );
  MUX U6251 ( .IN0(\modmult_1/xin[715] ), .IN1(creg[716]), .SEL(start_in[0]), 
        .F(\modmult_1/N1745 ) );
  MUX U6252 ( .IN0(\modmult_1/xin[714] ), .IN1(creg[715]), .SEL(start_in[0]), 
        .F(\modmult_1/N1744 ) );
  MUX U6253 ( .IN0(\modmult_1/xin[713] ), .IN1(creg[714]), .SEL(start_in[0]), 
        .F(\modmult_1/N1743 ) );
  MUX U6254 ( .IN0(\modmult_1/xin[712] ), .IN1(creg[713]), .SEL(start_in[0]), 
        .F(\modmult_1/N1742 ) );
  MUX U6255 ( .IN0(\modmult_1/xin[711] ), .IN1(creg[712]), .SEL(start_in[0]), 
        .F(\modmult_1/N1741 ) );
  MUX U6256 ( .IN0(\modmult_1/xin[710] ), .IN1(creg[711]), .SEL(start_in[0]), 
        .F(\modmult_1/N1740 ) );
  ANDN U6257 ( .A(n4110), .B(n3795), .Z(\modmult_1/N174 ) );
  XOR U6258 ( .A(n5939), .B(n5940), .Z(n3795) );
  MUX U6259 ( .IN0(\modmult_1/xin[709] ), .IN1(creg[710]), .SEL(start_in[0]), 
        .F(\modmult_1/N1739 ) );
  MUX U6260 ( .IN0(\modmult_1/xin[708] ), .IN1(creg[709]), .SEL(start_in[0]), 
        .F(\modmult_1/N1738 ) );
  MUX U6261 ( .IN0(\modmult_1/xin[707] ), .IN1(creg[708]), .SEL(start_in[0]), 
        .F(\modmult_1/N1737 ) );
  MUX U6262 ( .IN0(\modmult_1/xin[706] ), .IN1(creg[707]), .SEL(start_in[0]), 
        .F(\modmult_1/N1736 ) );
  MUX U6263 ( .IN0(\modmult_1/xin[705] ), .IN1(creg[706]), .SEL(start_in[0]), 
        .F(\modmult_1/N1735 ) );
  MUX U6264 ( .IN0(\modmult_1/xin[704] ), .IN1(creg[705]), .SEL(start_in[0]), 
        .F(\modmult_1/N1734 ) );
  MUX U6265 ( .IN0(\modmult_1/xin[703] ), .IN1(creg[704]), .SEL(start_in[0]), 
        .F(\modmult_1/N1733 ) );
  MUX U6266 ( .IN0(\modmult_1/xin[702] ), .IN1(creg[703]), .SEL(start_in[0]), 
        .F(\modmult_1/N1732 ) );
  MUX U6267 ( .IN0(\modmult_1/xin[701] ), .IN1(creg[702]), .SEL(start_in[0]), 
        .F(\modmult_1/N1731 ) );
  MUX U6268 ( .IN0(\modmult_1/xin[700] ), .IN1(creg[701]), .SEL(start_in[0]), 
        .F(\modmult_1/N1730 ) );
  ANDN U6269 ( .A(n4110), .B(n3798), .Z(\modmult_1/N173 ) );
  XOR U6270 ( .A(n5941), .B(n5942), .Z(n3798) );
  MUX U6271 ( .IN0(\modmult_1/xin[699] ), .IN1(creg[700]), .SEL(start_in[0]), 
        .F(\modmult_1/N1729 ) );
  MUX U6272 ( .IN0(\modmult_1/xin[698] ), .IN1(creg[699]), .SEL(start_in[0]), 
        .F(\modmult_1/N1728 ) );
  MUX U6273 ( .IN0(\modmult_1/xin[697] ), .IN1(creg[698]), .SEL(start_in[0]), 
        .F(\modmult_1/N1727 ) );
  MUX U6274 ( .IN0(\modmult_1/xin[696] ), .IN1(creg[697]), .SEL(start_in[0]), 
        .F(\modmult_1/N1726 ) );
  MUX U6275 ( .IN0(\modmult_1/xin[695] ), .IN1(creg[696]), .SEL(start_in[0]), 
        .F(\modmult_1/N1725 ) );
  MUX U6276 ( .IN0(\modmult_1/xin[694] ), .IN1(creg[695]), .SEL(start_in[0]), 
        .F(\modmult_1/N1724 ) );
  MUX U6277 ( .IN0(\modmult_1/xin[693] ), .IN1(creg[694]), .SEL(start_in[0]), 
        .F(\modmult_1/N1723 ) );
  MUX U6278 ( .IN0(\modmult_1/xin[692] ), .IN1(creg[693]), .SEL(start_in[0]), 
        .F(\modmult_1/N1722 ) );
  MUX U6279 ( .IN0(\modmult_1/xin[691] ), .IN1(creg[692]), .SEL(start_in[0]), 
        .F(\modmult_1/N1721 ) );
  MUX U6280 ( .IN0(\modmult_1/xin[690] ), .IN1(creg[691]), .SEL(start_in[0]), 
        .F(\modmult_1/N1720 ) );
  ANDN U6281 ( .A(n4110), .B(n3804), .Z(\modmult_1/N172 ) );
  XOR U6282 ( .A(n5943), .B(n5944), .Z(n3804) );
  MUX U6283 ( .IN0(\modmult_1/xin[689] ), .IN1(creg[690]), .SEL(start_in[0]), 
        .F(\modmult_1/N1719 ) );
  MUX U6284 ( .IN0(\modmult_1/xin[688] ), .IN1(creg[689]), .SEL(start_in[0]), 
        .F(\modmult_1/N1718 ) );
  MUX U6285 ( .IN0(\modmult_1/xin[687] ), .IN1(creg[688]), .SEL(start_in[0]), 
        .F(\modmult_1/N1717 ) );
  MUX U6286 ( .IN0(\modmult_1/xin[686] ), .IN1(creg[687]), .SEL(start_in[0]), 
        .F(\modmult_1/N1716 ) );
  MUX U6287 ( .IN0(\modmult_1/xin[685] ), .IN1(creg[686]), .SEL(start_in[0]), 
        .F(\modmult_1/N1715 ) );
  MUX U6288 ( .IN0(\modmult_1/xin[684] ), .IN1(creg[685]), .SEL(start_in[0]), 
        .F(\modmult_1/N1714 ) );
  MUX U6289 ( .IN0(\modmult_1/xin[683] ), .IN1(creg[684]), .SEL(start_in[0]), 
        .F(\modmult_1/N1713 ) );
  MUX U6290 ( .IN0(\modmult_1/xin[682] ), .IN1(creg[683]), .SEL(start_in[0]), 
        .F(\modmult_1/N1712 ) );
  MUX U6291 ( .IN0(\modmult_1/xin[681] ), .IN1(creg[682]), .SEL(start_in[0]), 
        .F(\modmult_1/N1711 ) );
  MUX U6292 ( .IN0(\modmult_1/xin[680] ), .IN1(creg[681]), .SEL(start_in[0]), 
        .F(\modmult_1/N1710 ) );
  ANDN U6293 ( .A(n4110), .B(n3807), .Z(\modmult_1/N171 ) );
  XOR U6294 ( .A(n5945), .B(n5946), .Z(n3807) );
  MUX U6295 ( .IN0(\modmult_1/xin[679] ), .IN1(creg[680]), .SEL(start_in[0]), 
        .F(\modmult_1/N1709 ) );
  MUX U6296 ( .IN0(\modmult_1/xin[678] ), .IN1(creg[679]), .SEL(start_in[0]), 
        .F(\modmult_1/N1708 ) );
  MUX U6297 ( .IN0(\modmult_1/xin[677] ), .IN1(creg[678]), .SEL(start_in[0]), 
        .F(\modmult_1/N1707 ) );
  MUX U6298 ( .IN0(\modmult_1/xin[676] ), .IN1(creg[677]), .SEL(start_in[0]), 
        .F(\modmult_1/N1706 ) );
  MUX U6299 ( .IN0(\modmult_1/xin[675] ), .IN1(creg[676]), .SEL(start_in[0]), 
        .F(\modmult_1/N1705 ) );
  MUX U6300 ( .IN0(\modmult_1/xin[674] ), .IN1(creg[675]), .SEL(start_in[0]), 
        .F(\modmult_1/N1704 ) );
  MUX U6301 ( .IN0(\modmult_1/xin[673] ), .IN1(creg[674]), .SEL(start_in[0]), 
        .F(\modmult_1/N1703 ) );
  MUX U6302 ( .IN0(\modmult_1/xin[672] ), .IN1(creg[673]), .SEL(start_in[0]), 
        .F(\modmult_1/N1702 ) );
  MUX U6303 ( .IN0(\modmult_1/xin[671] ), .IN1(creg[672]), .SEL(start_in[0]), 
        .F(\modmult_1/N1701 ) );
  MUX U6304 ( .IN0(\modmult_1/xin[670] ), .IN1(creg[671]), .SEL(start_in[0]), 
        .F(\modmult_1/N1700 ) );
  ANDN U6305 ( .A(n4110), .B(n3810), .Z(\modmult_1/N170 ) );
  XOR U6306 ( .A(n5947), .B(n5948), .Z(n3810) );
  ANDN U6307 ( .A(n4110), .B(n3867), .Z(\modmult_1/N17 ) );
  XOR U6308 ( .A(n5949), .B(n5950), .Z(n3867) );
  MUX U6309 ( .IN0(\modmult_1/xin[669] ), .IN1(creg[670]), .SEL(start_in[0]), 
        .F(\modmult_1/N1699 ) );
  MUX U6310 ( .IN0(\modmult_1/xin[668] ), .IN1(creg[669]), .SEL(start_in[0]), 
        .F(\modmult_1/N1698 ) );
  MUX U6311 ( .IN0(\modmult_1/xin[667] ), .IN1(creg[668]), .SEL(start_in[0]), 
        .F(\modmult_1/N1697 ) );
  MUX U6312 ( .IN0(\modmult_1/xin[666] ), .IN1(creg[667]), .SEL(start_in[0]), 
        .F(\modmult_1/N1696 ) );
  MUX U6313 ( .IN0(\modmult_1/xin[665] ), .IN1(creg[666]), .SEL(start_in[0]), 
        .F(\modmult_1/N1695 ) );
  MUX U6314 ( .IN0(\modmult_1/xin[664] ), .IN1(creg[665]), .SEL(start_in[0]), 
        .F(\modmult_1/N1694 ) );
  MUX U6315 ( .IN0(\modmult_1/xin[663] ), .IN1(creg[664]), .SEL(start_in[0]), 
        .F(\modmult_1/N1693 ) );
  MUX U6316 ( .IN0(\modmult_1/xin[662] ), .IN1(creg[663]), .SEL(start_in[0]), 
        .F(\modmult_1/N1692 ) );
  MUX U6317 ( .IN0(\modmult_1/xin[661] ), .IN1(creg[662]), .SEL(start_in[0]), 
        .F(\modmult_1/N1691 ) );
  MUX U6318 ( .IN0(\modmult_1/xin[660] ), .IN1(creg[661]), .SEL(start_in[0]), 
        .F(\modmult_1/N1690 ) );
  ANDN U6319 ( .A(n4110), .B(n3813), .Z(\modmult_1/N169 ) );
  XOR U6320 ( .A(n5951), .B(n5952), .Z(n3813) );
  MUX U6321 ( .IN0(\modmult_1/xin[659] ), .IN1(creg[660]), .SEL(start_in[0]), 
        .F(\modmult_1/N1689 ) );
  MUX U6322 ( .IN0(\modmult_1/xin[658] ), .IN1(creg[659]), .SEL(start_in[0]), 
        .F(\modmult_1/N1688 ) );
  MUX U6323 ( .IN0(\modmult_1/xin[657] ), .IN1(creg[658]), .SEL(start_in[0]), 
        .F(\modmult_1/N1687 ) );
  MUX U6324 ( .IN0(\modmult_1/xin[656] ), .IN1(creg[657]), .SEL(start_in[0]), 
        .F(\modmult_1/N1686 ) );
  MUX U6325 ( .IN0(\modmult_1/xin[655] ), .IN1(creg[656]), .SEL(start_in[0]), 
        .F(\modmult_1/N1685 ) );
  MUX U6326 ( .IN0(\modmult_1/xin[654] ), .IN1(creg[655]), .SEL(start_in[0]), 
        .F(\modmult_1/N1684 ) );
  MUX U6327 ( .IN0(\modmult_1/xin[653] ), .IN1(creg[654]), .SEL(start_in[0]), 
        .F(\modmult_1/N1683 ) );
  MUX U6328 ( .IN0(\modmult_1/xin[652] ), .IN1(creg[653]), .SEL(start_in[0]), 
        .F(\modmult_1/N1682 ) );
  MUX U6329 ( .IN0(\modmult_1/xin[651] ), .IN1(creg[652]), .SEL(start_in[0]), 
        .F(\modmult_1/N1681 ) );
  MUX U6330 ( .IN0(\modmult_1/xin[650] ), .IN1(creg[651]), .SEL(start_in[0]), 
        .F(\modmult_1/N1680 ) );
  ANDN U6331 ( .A(n4110), .B(n3816), .Z(\modmult_1/N168 ) );
  XOR U6332 ( .A(n5953), .B(n5954), .Z(n3816) );
  MUX U6333 ( .IN0(\modmult_1/xin[649] ), .IN1(creg[650]), .SEL(start_in[0]), 
        .F(\modmult_1/N1679 ) );
  MUX U6334 ( .IN0(\modmult_1/xin[648] ), .IN1(creg[649]), .SEL(start_in[0]), 
        .F(\modmult_1/N1678 ) );
  MUX U6335 ( .IN0(\modmult_1/xin[647] ), .IN1(creg[648]), .SEL(start_in[0]), 
        .F(\modmult_1/N1677 ) );
  MUX U6336 ( .IN0(\modmult_1/xin[646] ), .IN1(creg[647]), .SEL(start_in[0]), 
        .F(\modmult_1/N1676 ) );
  MUX U6337 ( .IN0(\modmult_1/xin[645] ), .IN1(creg[646]), .SEL(start_in[0]), 
        .F(\modmult_1/N1675 ) );
  MUX U6338 ( .IN0(\modmult_1/xin[644] ), .IN1(creg[645]), .SEL(start_in[0]), 
        .F(\modmult_1/N1674 ) );
  MUX U6339 ( .IN0(\modmult_1/xin[643] ), .IN1(creg[644]), .SEL(start_in[0]), 
        .F(\modmult_1/N1673 ) );
  MUX U6340 ( .IN0(\modmult_1/xin[642] ), .IN1(creg[643]), .SEL(start_in[0]), 
        .F(\modmult_1/N1672 ) );
  MUX U6341 ( .IN0(\modmult_1/xin[641] ), .IN1(creg[642]), .SEL(start_in[0]), 
        .F(\modmult_1/N1671 ) );
  MUX U6342 ( .IN0(\modmult_1/xin[640] ), .IN1(creg[641]), .SEL(start_in[0]), 
        .F(\modmult_1/N1670 ) );
  ANDN U6343 ( .A(n4110), .B(n3819), .Z(\modmult_1/N167 ) );
  XOR U6344 ( .A(n5955), .B(n5956), .Z(n3819) );
  MUX U6345 ( .IN0(\modmult_1/xin[639] ), .IN1(creg[640]), .SEL(start_in[0]), 
        .F(\modmult_1/N1669 ) );
  MUX U6346 ( .IN0(\modmult_1/xin[638] ), .IN1(creg[639]), .SEL(start_in[0]), 
        .F(\modmult_1/N1668 ) );
  MUX U6347 ( .IN0(\modmult_1/xin[637] ), .IN1(creg[638]), .SEL(start_in[0]), 
        .F(\modmult_1/N1667 ) );
  MUX U6348 ( .IN0(\modmult_1/xin[636] ), .IN1(creg[637]), .SEL(start_in[0]), 
        .F(\modmult_1/N1666 ) );
  MUX U6349 ( .IN0(\modmult_1/xin[635] ), .IN1(creg[636]), .SEL(start_in[0]), 
        .F(\modmult_1/N1665 ) );
  MUX U6350 ( .IN0(\modmult_1/xin[634] ), .IN1(creg[635]), .SEL(start_in[0]), 
        .F(\modmult_1/N1664 ) );
  MUX U6351 ( .IN0(\modmult_1/xin[633] ), .IN1(creg[634]), .SEL(start_in[0]), 
        .F(\modmult_1/N1663 ) );
  MUX U6352 ( .IN0(\modmult_1/xin[632] ), .IN1(creg[633]), .SEL(start_in[0]), 
        .F(\modmult_1/N1662 ) );
  MUX U6353 ( .IN0(\modmult_1/xin[631] ), .IN1(creg[632]), .SEL(start_in[0]), 
        .F(\modmult_1/N1661 ) );
  MUX U6354 ( .IN0(\modmult_1/xin[630] ), .IN1(creg[631]), .SEL(start_in[0]), 
        .F(\modmult_1/N1660 ) );
  ANDN U6355 ( .A(n4110), .B(n3822), .Z(\modmult_1/N166 ) );
  XOR U6356 ( .A(n5957), .B(n5958), .Z(n3822) );
  MUX U6357 ( .IN0(\modmult_1/xin[629] ), .IN1(creg[630]), .SEL(start_in[0]), 
        .F(\modmult_1/N1659 ) );
  MUX U6358 ( .IN0(\modmult_1/xin[628] ), .IN1(creg[629]), .SEL(start_in[0]), 
        .F(\modmult_1/N1658 ) );
  MUX U6359 ( .IN0(\modmult_1/xin[627] ), .IN1(creg[628]), .SEL(start_in[0]), 
        .F(\modmult_1/N1657 ) );
  MUX U6360 ( .IN0(\modmult_1/xin[626] ), .IN1(creg[627]), .SEL(start_in[0]), 
        .F(\modmult_1/N1656 ) );
  MUX U6361 ( .IN0(\modmult_1/xin[625] ), .IN1(creg[626]), .SEL(start_in[0]), 
        .F(\modmult_1/N1655 ) );
  MUX U6362 ( .IN0(\modmult_1/xin[624] ), .IN1(creg[625]), .SEL(start_in[0]), 
        .F(\modmult_1/N1654 ) );
  MUX U6363 ( .IN0(\modmult_1/xin[623] ), .IN1(creg[624]), .SEL(start_in[0]), 
        .F(\modmult_1/N1653 ) );
  MUX U6364 ( .IN0(\modmult_1/xin[622] ), .IN1(creg[623]), .SEL(start_in[0]), 
        .F(\modmult_1/N1652 ) );
  MUX U6365 ( .IN0(\modmult_1/xin[621] ), .IN1(creg[622]), .SEL(start_in[0]), 
        .F(\modmult_1/N1651 ) );
  MUX U6366 ( .IN0(\modmult_1/xin[620] ), .IN1(creg[621]), .SEL(start_in[0]), 
        .F(\modmult_1/N1650 ) );
  ANDN U6367 ( .A(n4110), .B(n3825), .Z(\modmult_1/N165 ) );
  XOR U6368 ( .A(n5959), .B(n5960), .Z(n3825) );
  MUX U6369 ( .IN0(\modmult_1/xin[619] ), .IN1(creg[620]), .SEL(start_in[0]), 
        .F(\modmult_1/N1649 ) );
  MUX U6370 ( .IN0(\modmult_1/xin[618] ), .IN1(creg[619]), .SEL(start_in[0]), 
        .F(\modmult_1/N1648 ) );
  MUX U6371 ( .IN0(\modmult_1/xin[617] ), .IN1(creg[618]), .SEL(start_in[0]), 
        .F(\modmult_1/N1647 ) );
  MUX U6372 ( .IN0(\modmult_1/xin[616] ), .IN1(creg[617]), .SEL(start_in[0]), 
        .F(\modmult_1/N1646 ) );
  MUX U6373 ( .IN0(\modmult_1/xin[615] ), .IN1(creg[616]), .SEL(start_in[0]), 
        .F(\modmult_1/N1645 ) );
  MUX U6374 ( .IN0(\modmult_1/xin[614] ), .IN1(creg[615]), .SEL(start_in[0]), 
        .F(\modmult_1/N1644 ) );
  MUX U6375 ( .IN0(\modmult_1/xin[613] ), .IN1(creg[614]), .SEL(start_in[0]), 
        .F(\modmult_1/N1643 ) );
  MUX U6376 ( .IN0(\modmult_1/xin[612] ), .IN1(creg[613]), .SEL(start_in[0]), 
        .F(\modmult_1/N1642 ) );
  MUX U6377 ( .IN0(\modmult_1/xin[611] ), .IN1(creg[612]), .SEL(start_in[0]), 
        .F(\modmult_1/N1641 ) );
  MUX U6378 ( .IN0(\modmult_1/xin[610] ), .IN1(creg[611]), .SEL(start_in[0]), 
        .F(\modmult_1/N1640 ) );
  ANDN U6379 ( .A(n4110), .B(n3828), .Z(\modmult_1/N164 ) );
  XOR U6380 ( .A(n5961), .B(n5962), .Z(n3828) );
  MUX U6381 ( .IN0(\modmult_1/xin[609] ), .IN1(creg[610]), .SEL(start_in[0]), 
        .F(\modmult_1/N1639 ) );
  MUX U6382 ( .IN0(\modmult_1/xin[608] ), .IN1(creg[609]), .SEL(start_in[0]), 
        .F(\modmult_1/N1638 ) );
  MUX U6383 ( .IN0(\modmult_1/xin[607] ), .IN1(creg[608]), .SEL(start_in[0]), 
        .F(\modmult_1/N1637 ) );
  MUX U6384 ( .IN0(\modmult_1/xin[606] ), .IN1(creg[607]), .SEL(start_in[0]), 
        .F(\modmult_1/N1636 ) );
  MUX U6385 ( .IN0(\modmult_1/xin[605] ), .IN1(creg[606]), .SEL(start_in[0]), 
        .F(\modmult_1/N1635 ) );
  MUX U6386 ( .IN0(\modmult_1/xin[604] ), .IN1(creg[605]), .SEL(start_in[0]), 
        .F(\modmult_1/N1634 ) );
  MUX U6387 ( .IN0(\modmult_1/xin[603] ), .IN1(creg[604]), .SEL(start_in[0]), 
        .F(\modmult_1/N1633 ) );
  MUX U6388 ( .IN0(\modmult_1/xin[602] ), .IN1(creg[603]), .SEL(start_in[0]), 
        .F(\modmult_1/N1632 ) );
  MUX U6389 ( .IN0(\modmult_1/xin[601] ), .IN1(creg[602]), .SEL(start_in[0]), 
        .F(\modmult_1/N1631 ) );
  MUX U6390 ( .IN0(\modmult_1/xin[600] ), .IN1(creg[601]), .SEL(start_in[0]), 
        .F(\modmult_1/N1630 ) );
  ANDN U6391 ( .A(n4110), .B(n3831), .Z(\modmult_1/N163 ) );
  XOR U6392 ( .A(n5963), .B(n5964), .Z(n3831) );
  MUX U6393 ( .IN0(\modmult_1/xin[599] ), .IN1(creg[600]), .SEL(start_in[0]), 
        .F(\modmult_1/N1629 ) );
  MUX U6394 ( .IN0(\modmult_1/xin[598] ), .IN1(creg[599]), .SEL(start_in[0]), 
        .F(\modmult_1/N1628 ) );
  MUX U6395 ( .IN0(\modmult_1/xin[597] ), .IN1(creg[598]), .SEL(start_in[0]), 
        .F(\modmult_1/N1627 ) );
  MUX U6396 ( .IN0(\modmult_1/xin[596] ), .IN1(creg[597]), .SEL(start_in[0]), 
        .F(\modmult_1/N1626 ) );
  MUX U6397 ( .IN0(\modmult_1/xin[595] ), .IN1(creg[596]), .SEL(start_in[0]), 
        .F(\modmult_1/N1625 ) );
  MUX U6398 ( .IN0(\modmult_1/xin[594] ), .IN1(creg[595]), .SEL(start_in[0]), 
        .F(\modmult_1/N1624 ) );
  MUX U6399 ( .IN0(\modmult_1/xin[593] ), .IN1(creg[594]), .SEL(start_in[0]), 
        .F(\modmult_1/N1623 ) );
  MUX U6400 ( .IN0(\modmult_1/xin[592] ), .IN1(creg[593]), .SEL(start_in[0]), 
        .F(\modmult_1/N1622 ) );
  MUX U6401 ( .IN0(\modmult_1/xin[591] ), .IN1(creg[592]), .SEL(start_in[0]), 
        .F(\modmult_1/N1621 ) );
  MUX U6402 ( .IN0(\modmult_1/xin[590] ), .IN1(creg[591]), .SEL(start_in[0]), 
        .F(\modmult_1/N1620 ) );
  ANDN U6403 ( .A(n4110), .B(n3837), .Z(\modmult_1/N162 ) );
  XOR U6404 ( .A(n5965), .B(n5966), .Z(n3837) );
  MUX U6405 ( .IN0(\modmult_1/xin[589] ), .IN1(creg[590]), .SEL(start_in[0]), 
        .F(\modmult_1/N1619 ) );
  MUX U6406 ( .IN0(\modmult_1/xin[588] ), .IN1(creg[589]), .SEL(start_in[0]), 
        .F(\modmult_1/N1618 ) );
  MUX U6407 ( .IN0(\modmult_1/xin[587] ), .IN1(creg[588]), .SEL(start_in[0]), 
        .F(\modmult_1/N1617 ) );
  MUX U6408 ( .IN0(\modmult_1/xin[586] ), .IN1(creg[587]), .SEL(start_in[0]), 
        .F(\modmult_1/N1616 ) );
  MUX U6409 ( .IN0(\modmult_1/xin[585] ), .IN1(creg[586]), .SEL(start_in[0]), 
        .F(\modmult_1/N1615 ) );
  MUX U6410 ( .IN0(\modmult_1/xin[584] ), .IN1(creg[585]), .SEL(start_in[0]), 
        .F(\modmult_1/N1614 ) );
  MUX U6411 ( .IN0(\modmult_1/xin[583] ), .IN1(creg[584]), .SEL(start_in[0]), 
        .F(\modmult_1/N1613 ) );
  MUX U6412 ( .IN0(\modmult_1/xin[582] ), .IN1(creg[583]), .SEL(start_in[0]), 
        .F(\modmult_1/N1612 ) );
  MUX U6413 ( .IN0(\modmult_1/xin[581] ), .IN1(creg[582]), .SEL(start_in[0]), 
        .F(\modmult_1/N1611 ) );
  MUX U6414 ( .IN0(\modmult_1/xin[580] ), .IN1(creg[581]), .SEL(start_in[0]), 
        .F(\modmult_1/N1610 ) );
  ANDN U6415 ( .A(n4110), .B(n3840), .Z(\modmult_1/N161 ) );
  XOR U6416 ( .A(n5967), .B(n5968), .Z(n3840) );
  MUX U6417 ( .IN0(\modmult_1/xin[579] ), .IN1(creg[580]), .SEL(start_in[0]), 
        .F(\modmult_1/N1609 ) );
  MUX U6418 ( .IN0(\modmult_1/xin[578] ), .IN1(creg[579]), .SEL(start_in[0]), 
        .F(\modmult_1/N1608 ) );
  MUX U6419 ( .IN0(\modmult_1/xin[577] ), .IN1(creg[578]), .SEL(start_in[0]), 
        .F(\modmult_1/N1607 ) );
  MUX U6420 ( .IN0(\modmult_1/xin[576] ), .IN1(creg[577]), .SEL(start_in[0]), 
        .F(\modmult_1/N1606 ) );
  MUX U6421 ( .IN0(\modmult_1/xin[575] ), .IN1(creg[576]), .SEL(start_in[0]), 
        .F(\modmult_1/N1605 ) );
  MUX U6422 ( .IN0(\modmult_1/xin[574] ), .IN1(creg[575]), .SEL(start_in[0]), 
        .F(\modmult_1/N1604 ) );
  MUX U6423 ( .IN0(\modmult_1/xin[573] ), .IN1(creg[574]), .SEL(start_in[0]), 
        .F(\modmult_1/N1603 ) );
  MUX U6424 ( .IN0(\modmult_1/xin[572] ), .IN1(creg[573]), .SEL(start_in[0]), 
        .F(\modmult_1/N1602 ) );
  MUX U6425 ( .IN0(\modmult_1/xin[571] ), .IN1(creg[572]), .SEL(start_in[0]), 
        .F(\modmult_1/N1601 ) );
  MUX U6426 ( .IN0(\modmult_1/xin[570] ), .IN1(creg[571]), .SEL(start_in[0]), 
        .F(\modmult_1/N1600 ) );
  ANDN U6427 ( .A(n4110), .B(n3843), .Z(\modmult_1/N160 ) );
  XOR U6428 ( .A(n5969), .B(n5970), .Z(n3843) );
  ANDN U6429 ( .A(n4110), .B(n3900), .Z(\modmult_1/N16 ) );
  XOR U6430 ( .A(n5971), .B(n5972), .Z(n3900) );
  MUX U6431 ( .IN0(\modmult_1/xin[569] ), .IN1(creg[570]), .SEL(start_in[0]), 
        .F(\modmult_1/N1599 ) );
  MUX U6432 ( .IN0(\modmult_1/xin[568] ), .IN1(creg[569]), .SEL(start_in[0]), 
        .F(\modmult_1/N1598 ) );
  MUX U6433 ( .IN0(\modmult_1/xin[567] ), .IN1(creg[568]), .SEL(start_in[0]), 
        .F(\modmult_1/N1597 ) );
  MUX U6434 ( .IN0(\modmult_1/xin[566] ), .IN1(creg[567]), .SEL(start_in[0]), 
        .F(\modmult_1/N1596 ) );
  MUX U6435 ( .IN0(\modmult_1/xin[565] ), .IN1(creg[566]), .SEL(start_in[0]), 
        .F(\modmult_1/N1595 ) );
  MUX U6436 ( .IN0(\modmult_1/xin[564] ), .IN1(creg[565]), .SEL(start_in[0]), 
        .F(\modmult_1/N1594 ) );
  MUX U6437 ( .IN0(\modmult_1/xin[563] ), .IN1(creg[564]), .SEL(start_in[0]), 
        .F(\modmult_1/N1593 ) );
  MUX U6438 ( .IN0(\modmult_1/xin[562] ), .IN1(creg[563]), .SEL(start_in[0]), 
        .F(\modmult_1/N1592 ) );
  MUX U6439 ( .IN0(\modmult_1/xin[561] ), .IN1(creg[562]), .SEL(start_in[0]), 
        .F(\modmult_1/N1591 ) );
  MUX U6440 ( .IN0(\modmult_1/xin[560] ), .IN1(creg[561]), .SEL(start_in[0]), 
        .F(\modmult_1/N1590 ) );
  ANDN U6441 ( .A(n4110), .B(n3846), .Z(\modmult_1/N159 ) );
  XOR U6442 ( .A(n5973), .B(n5974), .Z(n3846) );
  MUX U6443 ( .IN0(\modmult_1/xin[559] ), .IN1(creg[560]), .SEL(start_in[0]), 
        .F(\modmult_1/N1589 ) );
  MUX U6444 ( .IN0(\modmult_1/xin[558] ), .IN1(creg[559]), .SEL(start_in[0]), 
        .F(\modmult_1/N1588 ) );
  MUX U6445 ( .IN0(\modmult_1/xin[557] ), .IN1(creg[558]), .SEL(start_in[0]), 
        .F(\modmult_1/N1587 ) );
  MUX U6446 ( .IN0(\modmult_1/xin[556] ), .IN1(creg[557]), .SEL(start_in[0]), 
        .F(\modmult_1/N1586 ) );
  MUX U6447 ( .IN0(\modmult_1/xin[555] ), .IN1(creg[556]), .SEL(start_in[0]), 
        .F(\modmult_1/N1585 ) );
  MUX U6448 ( .IN0(\modmult_1/xin[554] ), .IN1(creg[555]), .SEL(start_in[0]), 
        .F(\modmult_1/N1584 ) );
  MUX U6449 ( .IN0(\modmult_1/xin[553] ), .IN1(creg[554]), .SEL(start_in[0]), 
        .F(\modmult_1/N1583 ) );
  MUX U6450 ( .IN0(\modmult_1/xin[552] ), .IN1(creg[553]), .SEL(start_in[0]), 
        .F(\modmult_1/N1582 ) );
  MUX U6451 ( .IN0(\modmult_1/xin[551] ), .IN1(creg[552]), .SEL(start_in[0]), 
        .F(\modmult_1/N1581 ) );
  MUX U6452 ( .IN0(\modmult_1/xin[550] ), .IN1(creg[551]), .SEL(start_in[0]), 
        .F(\modmult_1/N1580 ) );
  ANDN U6453 ( .A(n4110), .B(n3849), .Z(\modmult_1/N158 ) );
  XOR U6454 ( .A(n5975), .B(n5976), .Z(n3849) );
  MUX U6455 ( .IN0(\modmult_1/xin[549] ), .IN1(creg[550]), .SEL(start_in[0]), 
        .F(\modmult_1/N1579 ) );
  MUX U6456 ( .IN0(\modmult_1/xin[548] ), .IN1(creg[549]), .SEL(start_in[0]), 
        .F(\modmult_1/N1578 ) );
  MUX U6457 ( .IN0(\modmult_1/xin[547] ), .IN1(creg[548]), .SEL(start_in[0]), 
        .F(\modmult_1/N1577 ) );
  MUX U6458 ( .IN0(\modmult_1/xin[546] ), .IN1(creg[547]), .SEL(start_in[0]), 
        .F(\modmult_1/N1576 ) );
  MUX U6459 ( .IN0(\modmult_1/xin[545] ), .IN1(creg[546]), .SEL(start_in[0]), 
        .F(\modmult_1/N1575 ) );
  MUX U6460 ( .IN0(\modmult_1/xin[544] ), .IN1(creg[545]), .SEL(start_in[0]), 
        .F(\modmult_1/N1574 ) );
  MUX U6461 ( .IN0(\modmult_1/xin[543] ), .IN1(creg[544]), .SEL(start_in[0]), 
        .F(\modmult_1/N1573 ) );
  MUX U6462 ( .IN0(\modmult_1/xin[542] ), .IN1(creg[543]), .SEL(start_in[0]), 
        .F(\modmult_1/N1572 ) );
  MUX U6463 ( .IN0(\modmult_1/xin[541] ), .IN1(creg[542]), .SEL(start_in[0]), 
        .F(\modmult_1/N1571 ) );
  MUX U6464 ( .IN0(\modmult_1/xin[540] ), .IN1(creg[541]), .SEL(start_in[0]), 
        .F(\modmult_1/N1570 ) );
  ANDN U6465 ( .A(n4110), .B(n3852), .Z(\modmult_1/N157 ) );
  XOR U6466 ( .A(n5977), .B(n5978), .Z(n3852) );
  MUX U6467 ( .IN0(\modmult_1/xin[539] ), .IN1(creg[540]), .SEL(start_in[0]), 
        .F(\modmult_1/N1569 ) );
  MUX U6468 ( .IN0(\modmult_1/xin[538] ), .IN1(creg[539]), .SEL(start_in[0]), 
        .F(\modmult_1/N1568 ) );
  MUX U6469 ( .IN0(\modmult_1/xin[537] ), .IN1(creg[538]), .SEL(start_in[0]), 
        .F(\modmult_1/N1567 ) );
  MUX U6470 ( .IN0(\modmult_1/xin[536] ), .IN1(creg[537]), .SEL(start_in[0]), 
        .F(\modmult_1/N1566 ) );
  MUX U6471 ( .IN0(\modmult_1/xin[535] ), .IN1(creg[536]), .SEL(start_in[0]), 
        .F(\modmult_1/N1565 ) );
  MUX U6472 ( .IN0(\modmult_1/xin[534] ), .IN1(creg[535]), .SEL(start_in[0]), 
        .F(\modmult_1/N1564 ) );
  MUX U6473 ( .IN0(\modmult_1/xin[533] ), .IN1(creg[534]), .SEL(start_in[0]), 
        .F(\modmult_1/N1563 ) );
  MUX U6474 ( .IN0(\modmult_1/xin[532] ), .IN1(creg[533]), .SEL(start_in[0]), 
        .F(\modmult_1/N1562 ) );
  MUX U6475 ( .IN0(\modmult_1/xin[531] ), .IN1(creg[532]), .SEL(start_in[0]), 
        .F(\modmult_1/N1561 ) );
  MUX U6476 ( .IN0(\modmult_1/xin[530] ), .IN1(creg[531]), .SEL(start_in[0]), 
        .F(\modmult_1/N1560 ) );
  ANDN U6477 ( .A(n4110), .B(n3855), .Z(\modmult_1/N156 ) );
  XOR U6478 ( .A(n5979), .B(n5980), .Z(n3855) );
  MUX U6479 ( .IN0(\modmult_1/xin[529] ), .IN1(creg[530]), .SEL(start_in[0]), 
        .F(\modmult_1/N1559 ) );
  MUX U6480 ( .IN0(\modmult_1/xin[528] ), .IN1(creg[529]), .SEL(start_in[0]), 
        .F(\modmult_1/N1558 ) );
  MUX U6481 ( .IN0(\modmult_1/xin[527] ), .IN1(creg[528]), .SEL(start_in[0]), 
        .F(\modmult_1/N1557 ) );
  MUX U6482 ( .IN0(\modmult_1/xin[526] ), .IN1(creg[527]), .SEL(start_in[0]), 
        .F(\modmult_1/N1556 ) );
  MUX U6483 ( .IN0(\modmult_1/xin[525] ), .IN1(creg[526]), .SEL(start_in[0]), 
        .F(\modmult_1/N1555 ) );
  MUX U6484 ( .IN0(\modmult_1/xin[524] ), .IN1(creg[525]), .SEL(start_in[0]), 
        .F(\modmult_1/N1554 ) );
  MUX U6485 ( .IN0(\modmult_1/xin[523] ), .IN1(creg[524]), .SEL(start_in[0]), 
        .F(\modmult_1/N1553 ) );
  MUX U6486 ( .IN0(\modmult_1/xin[522] ), .IN1(creg[523]), .SEL(start_in[0]), 
        .F(\modmult_1/N1552 ) );
  MUX U6487 ( .IN0(\modmult_1/xin[521] ), .IN1(creg[522]), .SEL(start_in[0]), 
        .F(\modmult_1/N1551 ) );
  MUX U6488 ( .IN0(\modmult_1/xin[520] ), .IN1(creg[521]), .SEL(start_in[0]), 
        .F(\modmult_1/N1550 ) );
  ANDN U6489 ( .A(n4110), .B(n3858), .Z(\modmult_1/N155 ) );
  XOR U6490 ( .A(n5981), .B(n5982), .Z(n3858) );
  MUX U6491 ( .IN0(\modmult_1/xin[519] ), .IN1(creg[520]), .SEL(start_in[0]), 
        .F(\modmult_1/N1549 ) );
  MUX U6492 ( .IN0(\modmult_1/xin[518] ), .IN1(creg[519]), .SEL(start_in[0]), 
        .F(\modmult_1/N1548 ) );
  MUX U6493 ( .IN0(\modmult_1/xin[517] ), .IN1(creg[518]), .SEL(start_in[0]), 
        .F(\modmult_1/N1547 ) );
  MUX U6494 ( .IN0(\modmult_1/xin[516] ), .IN1(creg[517]), .SEL(start_in[0]), 
        .F(\modmult_1/N1546 ) );
  MUX U6495 ( .IN0(\modmult_1/xin[515] ), .IN1(creg[516]), .SEL(start_in[0]), 
        .F(\modmult_1/N1545 ) );
  MUX U6496 ( .IN0(\modmult_1/xin[514] ), .IN1(creg[515]), .SEL(start_in[0]), 
        .F(\modmult_1/N1544 ) );
  MUX U6497 ( .IN0(\modmult_1/xin[513] ), .IN1(creg[514]), .SEL(start_in[0]), 
        .F(\modmult_1/N1543 ) );
  MUX U6498 ( .IN0(\modmult_1/xin[512] ), .IN1(creg[513]), .SEL(start_in[0]), 
        .F(\modmult_1/N1542 ) );
  MUX U6499 ( .IN0(\modmult_1/xin[511] ), .IN1(creg[512]), .SEL(start_in[0]), 
        .F(\modmult_1/N1541 ) );
  MUX U6500 ( .IN0(\modmult_1/xin[510] ), .IN1(creg[511]), .SEL(start_in[0]), 
        .F(\modmult_1/N1540 ) );
  ANDN U6501 ( .A(n4110), .B(n3861), .Z(\modmult_1/N154 ) );
  XOR U6502 ( .A(n5983), .B(n5984), .Z(n3861) );
  MUX U6503 ( .IN0(\modmult_1/xin[509] ), .IN1(creg[510]), .SEL(start_in[0]), 
        .F(\modmult_1/N1539 ) );
  MUX U6504 ( .IN0(\modmult_1/xin[508] ), .IN1(creg[509]), .SEL(start_in[0]), 
        .F(\modmult_1/N1538 ) );
  MUX U6505 ( .IN0(\modmult_1/xin[507] ), .IN1(creg[508]), .SEL(start_in[0]), 
        .F(\modmult_1/N1537 ) );
  MUX U6506 ( .IN0(\modmult_1/xin[506] ), .IN1(creg[507]), .SEL(start_in[0]), 
        .F(\modmult_1/N1536 ) );
  MUX U6507 ( .IN0(\modmult_1/xin[505] ), .IN1(creg[506]), .SEL(start_in[0]), 
        .F(\modmult_1/N1535 ) );
  MUX U6508 ( .IN0(\modmult_1/xin[504] ), .IN1(creg[505]), .SEL(start_in[0]), 
        .F(\modmult_1/N1534 ) );
  MUX U6509 ( .IN0(\modmult_1/xin[503] ), .IN1(creg[504]), .SEL(start_in[0]), 
        .F(\modmult_1/N1533 ) );
  MUX U6510 ( .IN0(\modmult_1/xin[502] ), .IN1(creg[503]), .SEL(start_in[0]), 
        .F(\modmult_1/N1532 ) );
  MUX U6511 ( .IN0(\modmult_1/xin[501] ), .IN1(creg[502]), .SEL(start_in[0]), 
        .F(\modmult_1/N1531 ) );
  MUX U6512 ( .IN0(\modmult_1/xin[500] ), .IN1(creg[501]), .SEL(start_in[0]), 
        .F(\modmult_1/N1530 ) );
  ANDN U6513 ( .A(n4110), .B(n3864), .Z(\modmult_1/N153 ) );
  XOR U6514 ( .A(n5985), .B(n5986), .Z(n3864) );
  MUX U6515 ( .IN0(\modmult_1/xin[499] ), .IN1(creg[500]), .SEL(start_in[0]), 
        .F(\modmult_1/N1529 ) );
  MUX U6516 ( .IN0(\modmult_1/xin[498] ), .IN1(creg[499]), .SEL(start_in[0]), 
        .F(\modmult_1/N1528 ) );
  MUX U6517 ( .IN0(\modmult_1/xin[497] ), .IN1(creg[498]), .SEL(start_in[0]), 
        .F(\modmult_1/N1527 ) );
  MUX U6518 ( .IN0(\modmult_1/xin[496] ), .IN1(creg[497]), .SEL(start_in[0]), 
        .F(\modmult_1/N1526 ) );
  MUX U6519 ( .IN0(\modmult_1/xin[495] ), .IN1(creg[496]), .SEL(start_in[0]), 
        .F(\modmult_1/N1525 ) );
  MUX U6520 ( .IN0(\modmult_1/xin[494] ), .IN1(creg[495]), .SEL(start_in[0]), 
        .F(\modmult_1/N1524 ) );
  MUX U6521 ( .IN0(\modmult_1/xin[493] ), .IN1(creg[494]), .SEL(start_in[0]), 
        .F(\modmult_1/N1523 ) );
  MUX U6522 ( .IN0(\modmult_1/xin[492] ), .IN1(creg[493]), .SEL(start_in[0]), 
        .F(\modmult_1/N1522 ) );
  MUX U6523 ( .IN0(\modmult_1/xin[491] ), .IN1(creg[492]), .SEL(start_in[0]), 
        .F(\modmult_1/N1521 ) );
  MUX U6524 ( .IN0(\modmult_1/xin[490] ), .IN1(creg[491]), .SEL(start_in[0]), 
        .F(\modmult_1/N1520 ) );
  ANDN U6525 ( .A(n4110), .B(n3870), .Z(\modmult_1/N152 ) );
  XOR U6526 ( .A(n5987), .B(n5988), .Z(n3870) );
  MUX U6527 ( .IN0(\modmult_1/xin[489] ), .IN1(creg[490]), .SEL(start_in[0]), 
        .F(\modmult_1/N1519 ) );
  MUX U6528 ( .IN0(\modmult_1/xin[488] ), .IN1(creg[489]), .SEL(start_in[0]), 
        .F(\modmult_1/N1518 ) );
  MUX U6529 ( .IN0(\modmult_1/xin[487] ), .IN1(creg[488]), .SEL(start_in[0]), 
        .F(\modmult_1/N1517 ) );
  MUX U6530 ( .IN0(\modmult_1/xin[486] ), .IN1(creg[487]), .SEL(start_in[0]), 
        .F(\modmult_1/N1516 ) );
  MUX U6531 ( .IN0(\modmult_1/xin[485] ), .IN1(creg[486]), .SEL(start_in[0]), 
        .F(\modmult_1/N1515 ) );
  MUX U6532 ( .IN0(\modmult_1/xin[484] ), .IN1(creg[485]), .SEL(start_in[0]), 
        .F(\modmult_1/N1514 ) );
  MUX U6533 ( .IN0(\modmult_1/xin[483] ), .IN1(creg[484]), .SEL(start_in[0]), 
        .F(\modmult_1/N1513 ) );
  MUX U6534 ( .IN0(\modmult_1/xin[482] ), .IN1(creg[483]), .SEL(start_in[0]), 
        .F(\modmult_1/N1512 ) );
  MUX U6535 ( .IN0(\modmult_1/xin[481] ), .IN1(creg[482]), .SEL(start_in[0]), 
        .F(\modmult_1/N1511 ) );
  MUX U6536 ( .IN0(\modmult_1/xin[480] ), .IN1(creg[481]), .SEL(start_in[0]), 
        .F(\modmult_1/N1510 ) );
  ANDN U6537 ( .A(n4110), .B(n3873), .Z(\modmult_1/N151 ) );
  XOR U6538 ( .A(n5989), .B(n5990), .Z(n3873) );
  MUX U6539 ( .IN0(\modmult_1/xin[479] ), .IN1(creg[480]), .SEL(start_in[0]), 
        .F(\modmult_1/N1509 ) );
  MUX U6540 ( .IN0(\modmult_1/xin[478] ), .IN1(creg[479]), .SEL(start_in[0]), 
        .F(\modmult_1/N1508 ) );
  MUX U6541 ( .IN0(\modmult_1/xin[477] ), .IN1(creg[478]), .SEL(start_in[0]), 
        .F(\modmult_1/N1507 ) );
  MUX U6542 ( .IN0(\modmult_1/xin[476] ), .IN1(creg[477]), .SEL(start_in[0]), 
        .F(\modmult_1/N1506 ) );
  MUX U6543 ( .IN0(\modmult_1/xin[475] ), .IN1(creg[476]), .SEL(start_in[0]), 
        .F(\modmult_1/N1505 ) );
  MUX U6544 ( .IN0(\modmult_1/xin[474] ), .IN1(creg[475]), .SEL(start_in[0]), 
        .F(\modmult_1/N1504 ) );
  MUX U6545 ( .IN0(\modmult_1/xin[473] ), .IN1(creg[474]), .SEL(start_in[0]), 
        .F(\modmult_1/N1503 ) );
  MUX U6546 ( .IN0(\modmult_1/xin[472] ), .IN1(creg[473]), .SEL(start_in[0]), 
        .F(\modmult_1/N1502 ) );
  MUX U6547 ( .IN0(\modmult_1/xin[471] ), .IN1(creg[472]), .SEL(start_in[0]), 
        .F(\modmult_1/N1501 ) );
  MUX U6548 ( .IN0(\modmult_1/xin[470] ), .IN1(creg[471]), .SEL(start_in[0]), 
        .F(\modmult_1/N1500 ) );
  ANDN U6549 ( .A(n4110), .B(n3876), .Z(\modmult_1/N150 ) );
  XOR U6550 ( .A(n5991), .B(n5992), .Z(n3876) );
  ANDN U6551 ( .A(n4110), .B(n3933), .Z(\modmult_1/N15 ) );
  XOR U6552 ( .A(n5993), .B(n5994), .Z(n3933) );
  MUX U6553 ( .IN0(\modmult_1/xin[469] ), .IN1(creg[470]), .SEL(start_in[0]), 
        .F(\modmult_1/N1499 ) );
  MUX U6554 ( .IN0(\modmult_1/xin[468] ), .IN1(creg[469]), .SEL(start_in[0]), 
        .F(\modmult_1/N1498 ) );
  MUX U6555 ( .IN0(\modmult_1/xin[467] ), .IN1(creg[468]), .SEL(start_in[0]), 
        .F(\modmult_1/N1497 ) );
  MUX U6556 ( .IN0(\modmult_1/xin[466] ), .IN1(creg[467]), .SEL(start_in[0]), 
        .F(\modmult_1/N1496 ) );
  MUX U6557 ( .IN0(\modmult_1/xin[465] ), .IN1(creg[466]), .SEL(start_in[0]), 
        .F(\modmult_1/N1495 ) );
  MUX U6558 ( .IN0(\modmult_1/xin[464] ), .IN1(creg[465]), .SEL(start_in[0]), 
        .F(\modmult_1/N1494 ) );
  MUX U6559 ( .IN0(\modmult_1/xin[463] ), .IN1(creg[464]), .SEL(start_in[0]), 
        .F(\modmult_1/N1493 ) );
  MUX U6560 ( .IN0(\modmult_1/xin[462] ), .IN1(creg[463]), .SEL(start_in[0]), 
        .F(\modmult_1/N1492 ) );
  MUX U6561 ( .IN0(\modmult_1/xin[461] ), .IN1(creg[462]), .SEL(start_in[0]), 
        .F(\modmult_1/N1491 ) );
  MUX U6562 ( .IN0(\modmult_1/xin[460] ), .IN1(creg[461]), .SEL(start_in[0]), 
        .F(\modmult_1/N1490 ) );
  ANDN U6563 ( .A(n4110), .B(n3879), .Z(\modmult_1/N149 ) );
  XOR U6564 ( .A(n5995), .B(n5996), .Z(n3879) );
  MUX U6565 ( .IN0(\modmult_1/xin[459] ), .IN1(creg[460]), .SEL(start_in[0]), 
        .F(\modmult_1/N1489 ) );
  MUX U6566 ( .IN0(\modmult_1/xin[458] ), .IN1(creg[459]), .SEL(start_in[0]), 
        .F(\modmult_1/N1488 ) );
  MUX U6567 ( .IN0(\modmult_1/xin[457] ), .IN1(creg[458]), .SEL(start_in[0]), 
        .F(\modmult_1/N1487 ) );
  MUX U6568 ( .IN0(\modmult_1/xin[456] ), .IN1(creg[457]), .SEL(start_in[0]), 
        .F(\modmult_1/N1486 ) );
  MUX U6569 ( .IN0(\modmult_1/xin[455] ), .IN1(creg[456]), .SEL(start_in[0]), 
        .F(\modmult_1/N1485 ) );
  MUX U6570 ( .IN0(\modmult_1/xin[454] ), .IN1(creg[455]), .SEL(start_in[0]), 
        .F(\modmult_1/N1484 ) );
  MUX U6571 ( .IN0(\modmult_1/xin[453] ), .IN1(creg[454]), .SEL(start_in[0]), 
        .F(\modmult_1/N1483 ) );
  MUX U6572 ( .IN0(\modmult_1/xin[452] ), .IN1(creg[453]), .SEL(start_in[0]), 
        .F(\modmult_1/N1482 ) );
  MUX U6573 ( .IN0(\modmult_1/xin[451] ), .IN1(creg[452]), .SEL(start_in[0]), 
        .F(\modmult_1/N1481 ) );
  MUX U6574 ( .IN0(\modmult_1/xin[450] ), .IN1(creg[451]), .SEL(start_in[0]), 
        .F(\modmult_1/N1480 ) );
  ANDN U6575 ( .A(n4110), .B(n3882), .Z(\modmult_1/N148 ) );
  XOR U6576 ( .A(n5997), .B(n5998), .Z(n3882) );
  MUX U6577 ( .IN0(\modmult_1/xin[449] ), .IN1(creg[450]), .SEL(start_in[0]), 
        .F(\modmult_1/N1479 ) );
  MUX U6578 ( .IN0(\modmult_1/xin[448] ), .IN1(creg[449]), .SEL(start_in[0]), 
        .F(\modmult_1/N1478 ) );
  MUX U6579 ( .IN0(\modmult_1/xin[447] ), .IN1(creg[448]), .SEL(start_in[0]), 
        .F(\modmult_1/N1477 ) );
  MUX U6580 ( .IN0(\modmult_1/xin[446] ), .IN1(creg[447]), .SEL(start_in[0]), 
        .F(\modmult_1/N1476 ) );
  MUX U6581 ( .IN0(\modmult_1/xin[445] ), .IN1(creg[446]), .SEL(start_in[0]), 
        .F(\modmult_1/N1475 ) );
  MUX U6582 ( .IN0(\modmult_1/xin[444] ), .IN1(creg[445]), .SEL(start_in[0]), 
        .F(\modmult_1/N1474 ) );
  MUX U6583 ( .IN0(\modmult_1/xin[443] ), .IN1(creg[444]), .SEL(start_in[0]), 
        .F(\modmult_1/N1473 ) );
  MUX U6584 ( .IN0(\modmult_1/xin[442] ), .IN1(creg[443]), .SEL(start_in[0]), 
        .F(\modmult_1/N1472 ) );
  MUX U6585 ( .IN0(\modmult_1/xin[441] ), .IN1(creg[442]), .SEL(start_in[0]), 
        .F(\modmult_1/N1471 ) );
  MUX U6586 ( .IN0(\modmult_1/xin[440] ), .IN1(creg[441]), .SEL(start_in[0]), 
        .F(\modmult_1/N1470 ) );
  ANDN U6587 ( .A(n4110), .B(n3885), .Z(\modmult_1/N147 ) );
  XOR U6588 ( .A(n5999), .B(n6000), .Z(n3885) );
  MUX U6589 ( .IN0(\modmult_1/xin[439] ), .IN1(creg[440]), .SEL(start_in[0]), 
        .F(\modmult_1/N1469 ) );
  MUX U6590 ( .IN0(\modmult_1/xin[438] ), .IN1(creg[439]), .SEL(start_in[0]), 
        .F(\modmult_1/N1468 ) );
  MUX U6591 ( .IN0(\modmult_1/xin[437] ), .IN1(creg[438]), .SEL(start_in[0]), 
        .F(\modmult_1/N1467 ) );
  MUX U6592 ( .IN0(\modmult_1/xin[436] ), .IN1(creg[437]), .SEL(start_in[0]), 
        .F(\modmult_1/N1466 ) );
  MUX U6593 ( .IN0(\modmult_1/xin[435] ), .IN1(creg[436]), .SEL(start_in[0]), 
        .F(\modmult_1/N1465 ) );
  MUX U6594 ( .IN0(\modmult_1/xin[434] ), .IN1(creg[435]), .SEL(start_in[0]), 
        .F(\modmult_1/N1464 ) );
  MUX U6595 ( .IN0(\modmult_1/xin[433] ), .IN1(creg[434]), .SEL(start_in[0]), 
        .F(\modmult_1/N1463 ) );
  MUX U6596 ( .IN0(\modmult_1/xin[432] ), .IN1(creg[433]), .SEL(start_in[0]), 
        .F(\modmult_1/N1462 ) );
  MUX U6597 ( .IN0(\modmult_1/xin[431] ), .IN1(creg[432]), .SEL(start_in[0]), 
        .F(\modmult_1/N1461 ) );
  MUX U6598 ( .IN0(\modmult_1/xin[430] ), .IN1(creg[431]), .SEL(start_in[0]), 
        .F(\modmult_1/N1460 ) );
  ANDN U6599 ( .A(n4110), .B(n3888), .Z(\modmult_1/N146 ) );
  XOR U6600 ( .A(n6001), .B(n6002), .Z(n3888) );
  MUX U6601 ( .IN0(\modmult_1/xin[429] ), .IN1(creg[430]), .SEL(start_in[0]), 
        .F(\modmult_1/N1459 ) );
  MUX U6602 ( .IN0(\modmult_1/xin[428] ), .IN1(creg[429]), .SEL(start_in[0]), 
        .F(\modmult_1/N1458 ) );
  MUX U6603 ( .IN0(\modmult_1/xin[427] ), .IN1(creg[428]), .SEL(start_in[0]), 
        .F(\modmult_1/N1457 ) );
  MUX U6604 ( .IN0(\modmult_1/xin[426] ), .IN1(creg[427]), .SEL(start_in[0]), 
        .F(\modmult_1/N1456 ) );
  MUX U6605 ( .IN0(\modmult_1/xin[425] ), .IN1(creg[426]), .SEL(start_in[0]), 
        .F(\modmult_1/N1455 ) );
  MUX U6606 ( .IN0(\modmult_1/xin[424] ), .IN1(creg[425]), .SEL(start_in[0]), 
        .F(\modmult_1/N1454 ) );
  MUX U6607 ( .IN0(\modmult_1/xin[423] ), .IN1(creg[424]), .SEL(start_in[0]), 
        .F(\modmult_1/N1453 ) );
  MUX U6608 ( .IN0(\modmult_1/xin[422] ), .IN1(creg[423]), .SEL(start_in[0]), 
        .F(\modmult_1/N1452 ) );
  MUX U6609 ( .IN0(\modmult_1/xin[421] ), .IN1(creg[422]), .SEL(start_in[0]), 
        .F(\modmult_1/N1451 ) );
  MUX U6610 ( .IN0(\modmult_1/xin[420] ), .IN1(creg[421]), .SEL(start_in[0]), 
        .F(\modmult_1/N1450 ) );
  ANDN U6611 ( .A(n4110), .B(n3891), .Z(\modmult_1/N145 ) );
  XOR U6612 ( .A(n6003), .B(n6004), .Z(n3891) );
  MUX U6613 ( .IN0(\modmult_1/xin[419] ), .IN1(creg[420]), .SEL(start_in[0]), 
        .F(\modmult_1/N1449 ) );
  MUX U6614 ( .IN0(\modmult_1/xin[418] ), .IN1(creg[419]), .SEL(start_in[0]), 
        .F(\modmult_1/N1448 ) );
  MUX U6615 ( .IN0(\modmult_1/xin[417] ), .IN1(creg[418]), .SEL(start_in[0]), 
        .F(\modmult_1/N1447 ) );
  MUX U6616 ( .IN0(\modmult_1/xin[416] ), .IN1(creg[417]), .SEL(start_in[0]), 
        .F(\modmult_1/N1446 ) );
  MUX U6617 ( .IN0(\modmult_1/xin[415] ), .IN1(creg[416]), .SEL(start_in[0]), 
        .F(\modmult_1/N1445 ) );
  MUX U6618 ( .IN0(\modmult_1/xin[414] ), .IN1(creg[415]), .SEL(start_in[0]), 
        .F(\modmult_1/N1444 ) );
  MUX U6619 ( .IN0(\modmult_1/xin[413] ), .IN1(creg[414]), .SEL(start_in[0]), 
        .F(\modmult_1/N1443 ) );
  MUX U6620 ( .IN0(\modmult_1/xin[412] ), .IN1(creg[413]), .SEL(start_in[0]), 
        .F(\modmult_1/N1442 ) );
  MUX U6621 ( .IN0(\modmult_1/xin[411] ), .IN1(creg[412]), .SEL(start_in[0]), 
        .F(\modmult_1/N1441 ) );
  MUX U6622 ( .IN0(\modmult_1/xin[410] ), .IN1(creg[411]), .SEL(start_in[0]), 
        .F(\modmult_1/N1440 ) );
  ANDN U6623 ( .A(n4110), .B(n3894), .Z(\modmult_1/N144 ) );
  XOR U6624 ( .A(n6005), .B(n6006), .Z(n3894) );
  MUX U6625 ( .IN0(\modmult_1/xin[409] ), .IN1(creg[410]), .SEL(start_in[0]), 
        .F(\modmult_1/N1439 ) );
  MUX U6626 ( .IN0(\modmult_1/xin[408] ), .IN1(creg[409]), .SEL(start_in[0]), 
        .F(\modmult_1/N1438 ) );
  MUX U6627 ( .IN0(\modmult_1/xin[407] ), .IN1(creg[408]), .SEL(start_in[0]), 
        .F(\modmult_1/N1437 ) );
  MUX U6628 ( .IN0(\modmult_1/xin[406] ), .IN1(creg[407]), .SEL(start_in[0]), 
        .F(\modmult_1/N1436 ) );
  MUX U6629 ( .IN0(\modmult_1/xin[405] ), .IN1(creg[406]), .SEL(start_in[0]), 
        .F(\modmult_1/N1435 ) );
  MUX U6630 ( .IN0(\modmult_1/xin[404] ), .IN1(creg[405]), .SEL(start_in[0]), 
        .F(\modmult_1/N1434 ) );
  MUX U6631 ( .IN0(\modmult_1/xin[403] ), .IN1(creg[404]), .SEL(start_in[0]), 
        .F(\modmult_1/N1433 ) );
  MUX U6632 ( .IN0(\modmult_1/xin[402] ), .IN1(creg[403]), .SEL(start_in[0]), 
        .F(\modmult_1/N1432 ) );
  MUX U6633 ( .IN0(\modmult_1/xin[401] ), .IN1(creg[402]), .SEL(start_in[0]), 
        .F(\modmult_1/N1431 ) );
  MUX U6634 ( .IN0(\modmult_1/xin[400] ), .IN1(creg[401]), .SEL(start_in[0]), 
        .F(\modmult_1/N1430 ) );
  ANDN U6635 ( .A(n4110), .B(n3897), .Z(\modmult_1/N143 ) );
  XOR U6636 ( .A(n6007), .B(n6008), .Z(n3897) );
  MUX U6637 ( .IN0(\modmult_1/xin[399] ), .IN1(creg[400]), .SEL(start_in[0]), 
        .F(\modmult_1/N1429 ) );
  MUX U6638 ( .IN0(\modmult_1/xin[398] ), .IN1(creg[399]), .SEL(start_in[0]), 
        .F(\modmult_1/N1428 ) );
  MUX U6639 ( .IN0(\modmult_1/xin[397] ), .IN1(creg[398]), .SEL(start_in[0]), 
        .F(\modmult_1/N1427 ) );
  MUX U6640 ( .IN0(\modmult_1/xin[396] ), .IN1(creg[397]), .SEL(start_in[0]), 
        .F(\modmult_1/N1426 ) );
  MUX U6641 ( .IN0(\modmult_1/xin[395] ), .IN1(creg[396]), .SEL(start_in[0]), 
        .F(\modmult_1/N1425 ) );
  MUX U6642 ( .IN0(\modmult_1/xin[394] ), .IN1(creg[395]), .SEL(start_in[0]), 
        .F(\modmult_1/N1424 ) );
  MUX U6643 ( .IN0(\modmult_1/xin[393] ), .IN1(creg[394]), .SEL(start_in[0]), 
        .F(\modmult_1/N1423 ) );
  MUX U6644 ( .IN0(\modmult_1/xin[392] ), .IN1(creg[393]), .SEL(start_in[0]), 
        .F(\modmult_1/N1422 ) );
  MUX U6645 ( .IN0(\modmult_1/xin[391] ), .IN1(creg[392]), .SEL(start_in[0]), 
        .F(\modmult_1/N1421 ) );
  MUX U6646 ( .IN0(\modmult_1/xin[390] ), .IN1(creg[391]), .SEL(start_in[0]), 
        .F(\modmult_1/N1420 ) );
  ANDN U6647 ( .A(n4110), .B(n3903), .Z(\modmult_1/N142 ) );
  XOR U6648 ( .A(n6009), .B(n6010), .Z(n3903) );
  MUX U6649 ( .IN0(\modmult_1/xin[389] ), .IN1(creg[390]), .SEL(start_in[0]), 
        .F(\modmult_1/N1419 ) );
  MUX U6650 ( .IN0(\modmult_1/xin[388] ), .IN1(creg[389]), .SEL(start_in[0]), 
        .F(\modmult_1/N1418 ) );
  MUX U6651 ( .IN0(\modmult_1/xin[387] ), .IN1(creg[388]), .SEL(start_in[0]), 
        .F(\modmult_1/N1417 ) );
  MUX U6652 ( .IN0(\modmult_1/xin[386] ), .IN1(creg[387]), .SEL(start_in[0]), 
        .F(\modmult_1/N1416 ) );
  MUX U6653 ( .IN0(\modmult_1/xin[385] ), .IN1(creg[386]), .SEL(start_in[0]), 
        .F(\modmult_1/N1415 ) );
  MUX U6654 ( .IN0(\modmult_1/xin[384] ), .IN1(creg[385]), .SEL(start_in[0]), 
        .F(\modmult_1/N1414 ) );
  MUX U6655 ( .IN0(\modmult_1/xin[383] ), .IN1(creg[384]), .SEL(start_in[0]), 
        .F(\modmult_1/N1413 ) );
  MUX U6656 ( .IN0(\modmult_1/xin[382] ), .IN1(creg[383]), .SEL(start_in[0]), 
        .F(\modmult_1/N1412 ) );
  MUX U6657 ( .IN0(\modmult_1/xin[381] ), .IN1(creg[382]), .SEL(start_in[0]), 
        .F(\modmult_1/N1411 ) );
  MUX U6658 ( .IN0(\modmult_1/xin[380] ), .IN1(creg[381]), .SEL(start_in[0]), 
        .F(\modmult_1/N1410 ) );
  ANDN U6659 ( .A(n4110), .B(n3906), .Z(\modmult_1/N141 ) );
  XOR U6660 ( .A(n6011), .B(n6012), .Z(n3906) );
  MUX U6661 ( .IN0(\modmult_1/xin[379] ), .IN1(creg[380]), .SEL(start_in[0]), 
        .F(\modmult_1/N1409 ) );
  MUX U6662 ( .IN0(\modmult_1/xin[378] ), .IN1(creg[379]), .SEL(start_in[0]), 
        .F(\modmult_1/N1408 ) );
  MUX U6663 ( .IN0(\modmult_1/xin[377] ), .IN1(creg[378]), .SEL(start_in[0]), 
        .F(\modmult_1/N1407 ) );
  MUX U6664 ( .IN0(\modmult_1/xin[376] ), .IN1(creg[377]), .SEL(start_in[0]), 
        .F(\modmult_1/N1406 ) );
  MUX U6665 ( .IN0(\modmult_1/xin[375] ), .IN1(creg[376]), .SEL(start_in[0]), 
        .F(\modmult_1/N1405 ) );
  MUX U6666 ( .IN0(\modmult_1/xin[374] ), .IN1(creg[375]), .SEL(start_in[0]), 
        .F(\modmult_1/N1404 ) );
  MUX U6667 ( .IN0(\modmult_1/xin[373] ), .IN1(creg[374]), .SEL(start_in[0]), 
        .F(\modmult_1/N1403 ) );
  MUX U6668 ( .IN0(\modmult_1/xin[372] ), .IN1(creg[373]), .SEL(start_in[0]), 
        .F(\modmult_1/N1402 ) );
  MUX U6669 ( .IN0(\modmult_1/xin[371] ), .IN1(creg[372]), .SEL(start_in[0]), 
        .F(\modmult_1/N1401 ) );
  MUX U6670 ( .IN0(\modmult_1/xin[370] ), .IN1(creg[371]), .SEL(start_in[0]), 
        .F(\modmult_1/N1400 ) );
  ANDN U6671 ( .A(n4110), .B(n3909), .Z(\modmult_1/N140 ) );
  XOR U6672 ( .A(n6013), .B(n6014), .Z(n3909) );
  ANDN U6673 ( .A(n4110), .B(n3966), .Z(\modmult_1/N14 ) );
  XOR U6674 ( .A(n6015), .B(n6016), .Z(n3966) );
  MUX U6675 ( .IN0(\modmult_1/xin[369] ), .IN1(creg[370]), .SEL(start_in[0]), 
        .F(\modmult_1/N1399 ) );
  MUX U6676 ( .IN0(\modmult_1/xin[368] ), .IN1(creg[369]), .SEL(start_in[0]), 
        .F(\modmult_1/N1398 ) );
  MUX U6677 ( .IN0(\modmult_1/xin[367] ), .IN1(creg[368]), .SEL(start_in[0]), 
        .F(\modmult_1/N1397 ) );
  MUX U6678 ( .IN0(\modmult_1/xin[366] ), .IN1(creg[367]), .SEL(start_in[0]), 
        .F(\modmult_1/N1396 ) );
  MUX U6679 ( .IN0(\modmult_1/xin[365] ), .IN1(creg[366]), .SEL(start_in[0]), 
        .F(\modmult_1/N1395 ) );
  MUX U6680 ( .IN0(\modmult_1/xin[364] ), .IN1(creg[365]), .SEL(start_in[0]), 
        .F(\modmult_1/N1394 ) );
  MUX U6681 ( .IN0(\modmult_1/xin[363] ), .IN1(creg[364]), .SEL(start_in[0]), 
        .F(\modmult_1/N1393 ) );
  MUX U6682 ( .IN0(\modmult_1/xin[362] ), .IN1(creg[363]), .SEL(start_in[0]), 
        .F(\modmult_1/N1392 ) );
  MUX U6683 ( .IN0(\modmult_1/xin[361] ), .IN1(creg[362]), .SEL(start_in[0]), 
        .F(\modmult_1/N1391 ) );
  MUX U6684 ( .IN0(\modmult_1/xin[360] ), .IN1(creg[361]), .SEL(start_in[0]), 
        .F(\modmult_1/N1390 ) );
  ANDN U6685 ( .A(n4110), .B(n3912), .Z(\modmult_1/N139 ) );
  XOR U6686 ( .A(n6017), .B(n6018), .Z(n3912) );
  MUX U6687 ( .IN0(\modmult_1/xin[359] ), .IN1(creg[360]), .SEL(start_in[0]), 
        .F(\modmult_1/N1389 ) );
  MUX U6688 ( .IN0(\modmult_1/xin[358] ), .IN1(creg[359]), .SEL(start_in[0]), 
        .F(\modmult_1/N1388 ) );
  MUX U6689 ( .IN0(\modmult_1/xin[357] ), .IN1(creg[358]), .SEL(start_in[0]), 
        .F(\modmult_1/N1387 ) );
  MUX U6690 ( .IN0(\modmult_1/xin[356] ), .IN1(creg[357]), .SEL(start_in[0]), 
        .F(\modmult_1/N1386 ) );
  MUX U6691 ( .IN0(\modmult_1/xin[355] ), .IN1(creg[356]), .SEL(start_in[0]), 
        .F(\modmult_1/N1385 ) );
  MUX U6692 ( .IN0(\modmult_1/xin[354] ), .IN1(creg[355]), .SEL(start_in[0]), 
        .F(\modmult_1/N1384 ) );
  MUX U6693 ( .IN0(\modmult_1/xin[353] ), .IN1(creg[354]), .SEL(start_in[0]), 
        .F(\modmult_1/N1383 ) );
  MUX U6694 ( .IN0(\modmult_1/xin[352] ), .IN1(creg[353]), .SEL(start_in[0]), 
        .F(\modmult_1/N1382 ) );
  MUX U6695 ( .IN0(\modmult_1/xin[351] ), .IN1(creg[352]), .SEL(start_in[0]), 
        .F(\modmult_1/N1381 ) );
  MUX U6696 ( .IN0(\modmult_1/xin[350] ), .IN1(creg[351]), .SEL(start_in[0]), 
        .F(\modmult_1/N1380 ) );
  ANDN U6697 ( .A(n4110), .B(n3915), .Z(\modmult_1/N138 ) );
  XOR U6698 ( .A(n6019), .B(n6020), .Z(n3915) );
  MUX U6699 ( .IN0(\modmult_1/xin[349] ), .IN1(creg[350]), .SEL(start_in[0]), 
        .F(\modmult_1/N1379 ) );
  MUX U6700 ( .IN0(\modmult_1/xin[348] ), .IN1(creg[349]), .SEL(start_in[0]), 
        .F(\modmult_1/N1378 ) );
  MUX U6701 ( .IN0(\modmult_1/xin[347] ), .IN1(creg[348]), .SEL(start_in[0]), 
        .F(\modmult_1/N1377 ) );
  MUX U6702 ( .IN0(\modmult_1/xin[346] ), .IN1(creg[347]), .SEL(start_in[0]), 
        .F(\modmult_1/N1376 ) );
  MUX U6703 ( .IN0(\modmult_1/xin[345] ), .IN1(creg[346]), .SEL(start_in[0]), 
        .F(\modmult_1/N1375 ) );
  MUX U6704 ( .IN0(\modmult_1/xin[344] ), .IN1(creg[345]), .SEL(start_in[0]), 
        .F(\modmult_1/N1374 ) );
  MUX U6705 ( .IN0(\modmult_1/xin[343] ), .IN1(creg[344]), .SEL(start_in[0]), 
        .F(\modmult_1/N1373 ) );
  MUX U6706 ( .IN0(\modmult_1/xin[342] ), .IN1(creg[343]), .SEL(start_in[0]), 
        .F(\modmult_1/N1372 ) );
  MUX U6707 ( .IN0(\modmult_1/xin[341] ), .IN1(creg[342]), .SEL(start_in[0]), 
        .F(\modmult_1/N1371 ) );
  MUX U6708 ( .IN0(\modmult_1/xin[340] ), .IN1(creg[341]), .SEL(start_in[0]), 
        .F(\modmult_1/N1370 ) );
  ANDN U6709 ( .A(n4110), .B(n3918), .Z(\modmult_1/N137 ) );
  XOR U6710 ( .A(n6021), .B(n6022), .Z(n3918) );
  MUX U6711 ( .IN0(\modmult_1/xin[339] ), .IN1(creg[340]), .SEL(start_in[0]), 
        .F(\modmult_1/N1369 ) );
  MUX U6712 ( .IN0(\modmult_1/xin[338] ), .IN1(creg[339]), .SEL(start_in[0]), 
        .F(\modmult_1/N1368 ) );
  MUX U6713 ( .IN0(\modmult_1/xin[337] ), .IN1(creg[338]), .SEL(start_in[0]), 
        .F(\modmult_1/N1367 ) );
  MUX U6714 ( .IN0(\modmult_1/xin[336] ), .IN1(creg[337]), .SEL(start_in[0]), 
        .F(\modmult_1/N1366 ) );
  MUX U6715 ( .IN0(\modmult_1/xin[335] ), .IN1(creg[336]), .SEL(start_in[0]), 
        .F(\modmult_1/N1365 ) );
  MUX U6716 ( .IN0(\modmult_1/xin[334] ), .IN1(creg[335]), .SEL(start_in[0]), 
        .F(\modmult_1/N1364 ) );
  MUX U6717 ( .IN0(\modmult_1/xin[333] ), .IN1(creg[334]), .SEL(start_in[0]), 
        .F(\modmult_1/N1363 ) );
  MUX U6718 ( .IN0(\modmult_1/xin[332] ), .IN1(creg[333]), .SEL(start_in[0]), 
        .F(\modmult_1/N1362 ) );
  MUX U6719 ( .IN0(\modmult_1/xin[331] ), .IN1(creg[332]), .SEL(start_in[0]), 
        .F(\modmult_1/N1361 ) );
  MUX U6720 ( .IN0(\modmult_1/xin[330] ), .IN1(creg[331]), .SEL(start_in[0]), 
        .F(\modmult_1/N1360 ) );
  ANDN U6721 ( .A(n4110), .B(n3921), .Z(\modmult_1/N136 ) );
  XOR U6722 ( .A(n6023), .B(n6024), .Z(n3921) );
  MUX U6723 ( .IN0(\modmult_1/xin[329] ), .IN1(creg[330]), .SEL(start_in[0]), 
        .F(\modmult_1/N1359 ) );
  MUX U6724 ( .IN0(\modmult_1/xin[328] ), .IN1(creg[329]), .SEL(start_in[0]), 
        .F(\modmult_1/N1358 ) );
  MUX U6725 ( .IN0(\modmult_1/xin[327] ), .IN1(creg[328]), .SEL(start_in[0]), 
        .F(\modmult_1/N1357 ) );
  MUX U6726 ( .IN0(\modmult_1/xin[326] ), .IN1(creg[327]), .SEL(start_in[0]), 
        .F(\modmult_1/N1356 ) );
  MUX U6727 ( .IN0(\modmult_1/xin[325] ), .IN1(creg[326]), .SEL(start_in[0]), 
        .F(\modmult_1/N1355 ) );
  MUX U6728 ( .IN0(\modmult_1/xin[324] ), .IN1(creg[325]), .SEL(start_in[0]), 
        .F(\modmult_1/N1354 ) );
  MUX U6729 ( .IN0(\modmult_1/xin[323] ), .IN1(creg[324]), .SEL(start_in[0]), 
        .F(\modmult_1/N1353 ) );
  MUX U6730 ( .IN0(\modmult_1/xin[322] ), .IN1(creg[323]), .SEL(start_in[0]), 
        .F(\modmult_1/N1352 ) );
  MUX U6731 ( .IN0(\modmult_1/xin[321] ), .IN1(creg[322]), .SEL(start_in[0]), 
        .F(\modmult_1/N1351 ) );
  MUX U6732 ( .IN0(\modmult_1/xin[320] ), .IN1(creg[321]), .SEL(start_in[0]), 
        .F(\modmult_1/N1350 ) );
  ANDN U6733 ( .A(n4110), .B(n3924), .Z(\modmult_1/N135 ) );
  XOR U6734 ( .A(n6025), .B(n6026), .Z(n3924) );
  MUX U6735 ( .IN0(\modmult_1/xin[319] ), .IN1(creg[320]), .SEL(start_in[0]), 
        .F(\modmult_1/N1349 ) );
  MUX U6736 ( .IN0(\modmult_1/xin[318] ), .IN1(creg[319]), .SEL(start_in[0]), 
        .F(\modmult_1/N1348 ) );
  MUX U6737 ( .IN0(\modmult_1/xin[317] ), .IN1(creg[318]), .SEL(start_in[0]), 
        .F(\modmult_1/N1347 ) );
  MUX U6738 ( .IN0(\modmult_1/xin[316] ), .IN1(creg[317]), .SEL(start_in[0]), 
        .F(\modmult_1/N1346 ) );
  MUX U6739 ( .IN0(\modmult_1/xin[315] ), .IN1(creg[316]), .SEL(start_in[0]), 
        .F(\modmult_1/N1345 ) );
  MUX U6740 ( .IN0(\modmult_1/xin[314] ), .IN1(creg[315]), .SEL(start_in[0]), 
        .F(\modmult_1/N1344 ) );
  MUX U6741 ( .IN0(\modmult_1/xin[313] ), .IN1(creg[314]), .SEL(start_in[0]), 
        .F(\modmult_1/N1343 ) );
  MUX U6742 ( .IN0(\modmult_1/xin[312] ), .IN1(creg[313]), .SEL(start_in[0]), 
        .F(\modmult_1/N1342 ) );
  MUX U6743 ( .IN0(\modmult_1/xin[311] ), .IN1(creg[312]), .SEL(start_in[0]), 
        .F(\modmult_1/N1341 ) );
  MUX U6744 ( .IN0(\modmult_1/xin[310] ), .IN1(creg[311]), .SEL(start_in[0]), 
        .F(\modmult_1/N1340 ) );
  ANDN U6745 ( .A(n4110), .B(n3927), .Z(\modmult_1/N134 ) );
  XOR U6746 ( .A(n6027), .B(n6028), .Z(n3927) );
  MUX U6747 ( .IN0(\modmult_1/xin[309] ), .IN1(creg[310]), .SEL(start_in[0]), 
        .F(\modmult_1/N1339 ) );
  MUX U6748 ( .IN0(\modmult_1/xin[308] ), .IN1(creg[309]), .SEL(start_in[0]), 
        .F(\modmult_1/N1338 ) );
  MUX U6749 ( .IN0(\modmult_1/xin[307] ), .IN1(creg[308]), .SEL(start_in[0]), 
        .F(\modmult_1/N1337 ) );
  MUX U6750 ( .IN0(\modmult_1/xin[306] ), .IN1(creg[307]), .SEL(start_in[0]), 
        .F(\modmult_1/N1336 ) );
  MUX U6751 ( .IN0(\modmult_1/xin[305] ), .IN1(creg[306]), .SEL(start_in[0]), 
        .F(\modmult_1/N1335 ) );
  MUX U6752 ( .IN0(\modmult_1/xin[304] ), .IN1(creg[305]), .SEL(start_in[0]), 
        .F(\modmult_1/N1334 ) );
  MUX U6753 ( .IN0(\modmult_1/xin[303] ), .IN1(creg[304]), .SEL(start_in[0]), 
        .F(\modmult_1/N1333 ) );
  MUX U6754 ( .IN0(\modmult_1/xin[302] ), .IN1(creg[303]), .SEL(start_in[0]), 
        .F(\modmult_1/N1332 ) );
  MUX U6755 ( .IN0(\modmult_1/xin[301] ), .IN1(creg[302]), .SEL(start_in[0]), 
        .F(\modmult_1/N1331 ) );
  MUX U6756 ( .IN0(\modmult_1/xin[300] ), .IN1(creg[301]), .SEL(start_in[0]), 
        .F(\modmult_1/N1330 ) );
  ANDN U6757 ( .A(n4110), .B(n3930), .Z(\modmult_1/N133 ) );
  XOR U6758 ( .A(n6029), .B(n6030), .Z(n3930) );
  MUX U6759 ( .IN0(\modmult_1/xin[299] ), .IN1(creg[300]), .SEL(start_in[0]), 
        .F(\modmult_1/N1329 ) );
  MUX U6760 ( .IN0(\modmult_1/xin[298] ), .IN1(creg[299]), .SEL(start_in[0]), 
        .F(\modmult_1/N1328 ) );
  MUX U6761 ( .IN0(\modmult_1/xin[297] ), .IN1(creg[298]), .SEL(start_in[0]), 
        .F(\modmult_1/N1327 ) );
  MUX U6762 ( .IN0(\modmult_1/xin[296] ), .IN1(creg[297]), .SEL(start_in[0]), 
        .F(\modmult_1/N1326 ) );
  MUX U6763 ( .IN0(\modmult_1/xin[295] ), .IN1(creg[296]), .SEL(start_in[0]), 
        .F(\modmult_1/N1325 ) );
  MUX U6764 ( .IN0(\modmult_1/xin[294] ), .IN1(creg[295]), .SEL(start_in[0]), 
        .F(\modmult_1/N1324 ) );
  MUX U6765 ( .IN0(\modmult_1/xin[293] ), .IN1(creg[294]), .SEL(start_in[0]), 
        .F(\modmult_1/N1323 ) );
  MUX U6766 ( .IN0(\modmult_1/xin[292] ), .IN1(creg[293]), .SEL(start_in[0]), 
        .F(\modmult_1/N1322 ) );
  MUX U6767 ( .IN0(\modmult_1/xin[291] ), .IN1(creg[292]), .SEL(start_in[0]), 
        .F(\modmult_1/N1321 ) );
  MUX U6768 ( .IN0(\modmult_1/xin[290] ), .IN1(creg[291]), .SEL(start_in[0]), 
        .F(\modmult_1/N1320 ) );
  ANDN U6769 ( .A(n4110), .B(n3936), .Z(\modmult_1/N132 ) );
  XOR U6770 ( .A(n6031), .B(n6032), .Z(n3936) );
  MUX U6771 ( .IN0(\modmult_1/xin[289] ), .IN1(creg[290]), .SEL(start_in[0]), 
        .F(\modmult_1/N1319 ) );
  MUX U6772 ( .IN0(\modmult_1/xin[288] ), .IN1(creg[289]), .SEL(start_in[0]), 
        .F(\modmult_1/N1318 ) );
  MUX U6773 ( .IN0(\modmult_1/xin[287] ), .IN1(creg[288]), .SEL(start_in[0]), 
        .F(\modmult_1/N1317 ) );
  MUX U6774 ( .IN0(\modmult_1/xin[286] ), .IN1(creg[287]), .SEL(start_in[0]), 
        .F(\modmult_1/N1316 ) );
  MUX U6775 ( .IN0(\modmult_1/xin[285] ), .IN1(creg[286]), .SEL(start_in[0]), 
        .F(\modmult_1/N1315 ) );
  MUX U6776 ( .IN0(\modmult_1/xin[284] ), .IN1(creg[285]), .SEL(start_in[0]), 
        .F(\modmult_1/N1314 ) );
  MUX U6777 ( .IN0(\modmult_1/xin[283] ), .IN1(creg[284]), .SEL(start_in[0]), 
        .F(\modmult_1/N1313 ) );
  MUX U6778 ( .IN0(\modmult_1/xin[282] ), .IN1(creg[283]), .SEL(start_in[0]), 
        .F(\modmult_1/N1312 ) );
  MUX U6779 ( .IN0(\modmult_1/xin[281] ), .IN1(creg[282]), .SEL(start_in[0]), 
        .F(\modmult_1/N1311 ) );
  MUX U6780 ( .IN0(\modmult_1/xin[280] ), .IN1(creg[281]), .SEL(start_in[0]), 
        .F(\modmult_1/N1310 ) );
  ANDN U6781 ( .A(n4110), .B(n3939), .Z(\modmult_1/N131 ) );
  XOR U6782 ( .A(n6033), .B(n6034), .Z(n3939) );
  MUX U6783 ( .IN0(\modmult_1/xin[279] ), .IN1(creg[280]), .SEL(start_in[0]), 
        .F(\modmult_1/N1309 ) );
  MUX U6784 ( .IN0(\modmult_1/xin[278] ), .IN1(creg[279]), .SEL(start_in[0]), 
        .F(\modmult_1/N1308 ) );
  MUX U6785 ( .IN0(\modmult_1/xin[277] ), .IN1(creg[278]), .SEL(start_in[0]), 
        .F(\modmult_1/N1307 ) );
  MUX U6786 ( .IN0(\modmult_1/xin[276] ), .IN1(creg[277]), .SEL(start_in[0]), 
        .F(\modmult_1/N1306 ) );
  MUX U6787 ( .IN0(\modmult_1/xin[275] ), .IN1(creg[276]), .SEL(start_in[0]), 
        .F(\modmult_1/N1305 ) );
  MUX U6788 ( .IN0(\modmult_1/xin[274] ), .IN1(creg[275]), .SEL(start_in[0]), 
        .F(\modmult_1/N1304 ) );
  MUX U6789 ( .IN0(\modmult_1/xin[273] ), .IN1(creg[274]), .SEL(start_in[0]), 
        .F(\modmult_1/N1303 ) );
  MUX U6790 ( .IN0(\modmult_1/xin[272] ), .IN1(creg[273]), .SEL(start_in[0]), 
        .F(\modmult_1/N1302 ) );
  MUX U6791 ( .IN0(\modmult_1/xin[271] ), .IN1(creg[272]), .SEL(start_in[0]), 
        .F(\modmult_1/N1301 ) );
  MUX U6792 ( .IN0(\modmult_1/xin[270] ), .IN1(creg[271]), .SEL(start_in[0]), 
        .F(\modmult_1/N1300 ) );
  ANDN U6793 ( .A(n4110), .B(n3942), .Z(\modmult_1/N130 ) );
  XOR U6794 ( .A(n6035), .B(n6036), .Z(n3942) );
  ANDN U6795 ( .A(n4110), .B(n3999), .Z(\modmult_1/N13 ) );
  XOR U6796 ( .A(n6037), .B(n6038), .Z(n3999) );
  MUX U6797 ( .IN0(\modmult_1/xin[269] ), .IN1(creg[270]), .SEL(start_in[0]), 
        .F(\modmult_1/N1299 ) );
  MUX U6798 ( .IN0(\modmult_1/xin[268] ), .IN1(creg[269]), .SEL(start_in[0]), 
        .F(\modmult_1/N1298 ) );
  MUX U6799 ( .IN0(\modmult_1/xin[267] ), .IN1(creg[268]), .SEL(start_in[0]), 
        .F(\modmult_1/N1297 ) );
  MUX U6800 ( .IN0(\modmult_1/xin[266] ), .IN1(creg[267]), .SEL(start_in[0]), 
        .F(\modmult_1/N1296 ) );
  MUX U6801 ( .IN0(\modmult_1/xin[265] ), .IN1(creg[266]), .SEL(start_in[0]), 
        .F(\modmult_1/N1295 ) );
  MUX U6802 ( .IN0(\modmult_1/xin[264] ), .IN1(creg[265]), .SEL(start_in[0]), 
        .F(\modmult_1/N1294 ) );
  MUX U6803 ( .IN0(\modmult_1/xin[263] ), .IN1(creg[264]), .SEL(start_in[0]), 
        .F(\modmult_1/N1293 ) );
  MUX U6804 ( .IN0(\modmult_1/xin[262] ), .IN1(creg[263]), .SEL(start_in[0]), 
        .F(\modmult_1/N1292 ) );
  MUX U6805 ( .IN0(\modmult_1/xin[261] ), .IN1(creg[262]), .SEL(start_in[0]), 
        .F(\modmult_1/N1291 ) );
  MUX U6806 ( .IN0(\modmult_1/xin[260] ), .IN1(creg[261]), .SEL(start_in[0]), 
        .F(\modmult_1/N1290 ) );
  ANDN U6807 ( .A(n4110), .B(n3945), .Z(\modmult_1/N129 ) );
  XOR U6808 ( .A(n6039), .B(n6040), .Z(n3945) );
  MUX U6809 ( .IN0(\modmult_1/xin[259] ), .IN1(creg[260]), .SEL(start_in[0]), 
        .F(\modmult_1/N1289 ) );
  MUX U6810 ( .IN0(\modmult_1/xin[258] ), .IN1(creg[259]), .SEL(start_in[0]), 
        .F(\modmult_1/N1288 ) );
  MUX U6811 ( .IN0(\modmult_1/xin[257] ), .IN1(creg[258]), .SEL(start_in[0]), 
        .F(\modmult_1/N1287 ) );
  MUX U6812 ( .IN0(\modmult_1/xin[256] ), .IN1(creg[257]), .SEL(start_in[0]), 
        .F(\modmult_1/N1286 ) );
  MUX U6813 ( .IN0(\modmult_1/xin[255] ), .IN1(creg[256]), .SEL(start_in[0]), 
        .F(\modmult_1/N1285 ) );
  MUX U6814 ( .IN0(\modmult_1/xin[254] ), .IN1(creg[255]), .SEL(start_in[0]), 
        .F(\modmult_1/N1284 ) );
  MUX U6815 ( .IN0(\modmult_1/xin[253] ), .IN1(creg[254]), .SEL(start_in[0]), 
        .F(\modmult_1/N1283 ) );
  MUX U6816 ( .IN0(\modmult_1/xin[252] ), .IN1(creg[253]), .SEL(start_in[0]), 
        .F(\modmult_1/N1282 ) );
  MUX U6817 ( .IN0(\modmult_1/xin[251] ), .IN1(creg[252]), .SEL(start_in[0]), 
        .F(\modmult_1/N1281 ) );
  MUX U6818 ( .IN0(\modmult_1/xin[250] ), .IN1(creg[251]), .SEL(start_in[0]), 
        .F(\modmult_1/N1280 ) );
  ANDN U6819 ( .A(n4110), .B(n3948), .Z(\modmult_1/N128 ) );
  XOR U6820 ( .A(n6041), .B(n6042), .Z(n3948) );
  MUX U6821 ( .IN0(\modmult_1/xin[249] ), .IN1(creg[250]), .SEL(start_in[0]), 
        .F(\modmult_1/N1279 ) );
  MUX U6822 ( .IN0(\modmult_1/xin[248] ), .IN1(creg[249]), .SEL(start_in[0]), 
        .F(\modmult_1/N1278 ) );
  MUX U6823 ( .IN0(\modmult_1/xin[247] ), .IN1(creg[248]), .SEL(start_in[0]), 
        .F(\modmult_1/N1277 ) );
  MUX U6824 ( .IN0(\modmult_1/xin[246] ), .IN1(creg[247]), .SEL(start_in[0]), 
        .F(\modmult_1/N1276 ) );
  MUX U6825 ( .IN0(\modmult_1/xin[245] ), .IN1(creg[246]), .SEL(start_in[0]), 
        .F(\modmult_1/N1275 ) );
  MUX U6826 ( .IN0(\modmult_1/xin[244] ), .IN1(creg[245]), .SEL(start_in[0]), 
        .F(\modmult_1/N1274 ) );
  MUX U6827 ( .IN0(\modmult_1/xin[243] ), .IN1(creg[244]), .SEL(start_in[0]), 
        .F(\modmult_1/N1273 ) );
  MUX U6828 ( .IN0(\modmult_1/xin[242] ), .IN1(creg[243]), .SEL(start_in[0]), 
        .F(\modmult_1/N1272 ) );
  MUX U6829 ( .IN0(\modmult_1/xin[241] ), .IN1(creg[242]), .SEL(start_in[0]), 
        .F(\modmult_1/N1271 ) );
  MUX U6830 ( .IN0(\modmult_1/xin[240] ), .IN1(creg[241]), .SEL(start_in[0]), 
        .F(\modmult_1/N1270 ) );
  ANDN U6831 ( .A(n4110), .B(n3951), .Z(\modmult_1/N127 ) );
  XOR U6832 ( .A(n6043), .B(n6044), .Z(n3951) );
  MUX U6833 ( .IN0(\modmult_1/xin[239] ), .IN1(creg[240]), .SEL(start_in[0]), 
        .F(\modmult_1/N1269 ) );
  MUX U6834 ( .IN0(\modmult_1/xin[238] ), .IN1(creg[239]), .SEL(start_in[0]), 
        .F(\modmult_1/N1268 ) );
  MUX U6835 ( .IN0(\modmult_1/xin[237] ), .IN1(creg[238]), .SEL(start_in[0]), 
        .F(\modmult_1/N1267 ) );
  MUX U6836 ( .IN0(\modmult_1/xin[236] ), .IN1(creg[237]), .SEL(start_in[0]), 
        .F(\modmult_1/N1266 ) );
  MUX U6837 ( .IN0(\modmult_1/xin[235] ), .IN1(creg[236]), .SEL(start_in[0]), 
        .F(\modmult_1/N1265 ) );
  MUX U6838 ( .IN0(\modmult_1/xin[234] ), .IN1(creg[235]), .SEL(start_in[0]), 
        .F(\modmult_1/N1264 ) );
  MUX U6839 ( .IN0(\modmult_1/xin[233] ), .IN1(creg[234]), .SEL(start_in[0]), 
        .F(\modmult_1/N1263 ) );
  MUX U6840 ( .IN0(\modmult_1/xin[232] ), .IN1(creg[233]), .SEL(start_in[0]), 
        .F(\modmult_1/N1262 ) );
  MUX U6841 ( .IN0(\modmult_1/xin[231] ), .IN1(creg[232]), .SEL(start_in[0]), 
        .F(\modmult_1/N1261 ) );
  MUX U6842 ( .IN0(\modmult_1/xin[230] ), .IN1(creg[231]), .SEL(start_in[0]), 
        .F(\modmult_1/N1260 ) );
  ANDN U6843 ( .A(n4110), .B(n3954), .Z(\modmult_1/N126 ) );
  XOR U6844 ( .A(n6045), .B(n6046), .Z(n3954) );
  MUX U6845 ( .IN0(\modmult_1/xin[229] ), .IN1(creg[230]), .SEL(start_in[0]), 
        .F(\modmult_1/N1259 ) );
  MUX U6846 ( .IN0(\modmult_1/xin[228] ), .IN1(creg[229]), .SEL(start_in[0]), 
        .F(\modmult_1/N1258 ) );
  MUX U6847 ( .IN0(\modmult_1/xin[227] ), .IN1(creg[228]), .SEL(start_in[0]), 
        .F(\modmult_1/N1257 ) );
  MUX U6848 ( .IN0(\modmult_1/xin[226] ), .IN1(creg[227]), .SEL(start_in[0]), 
        .F(\modmult_1/N1256 ) );
  MUX U6849 ( .IN0(\modmult_1/xin[225] ), .IN1(creg[226]), .SEL(start_in[0]), 
        .F(\modmult_1/N1255 ) );
  MUX U6850 ( .IN0(\modmult_1/xin[224] ), .IN1(creg[225]), .SEL(start_in[0]), 
        .F(\modmult_1/N1254 ) );
  MUX U6851 ( .IN0(\modmult_1/xin[223] ), .IN1(creg[224]), .SEL(start_in[0]), 
        .F(\modmult_1/N1253 ) );
  MUX U6852 ( .IN0(\modmult_1/xin[222] ), .IN1(creg[223]), .SEL(start_in[0]), 
        .F(\modmult_1/N1252 ) );
  MUX U6853 ( .IN0(\modmult_1/xin[221] ), .IN1(creg[222]), .SEL(start_in[0]), 
        .F(\modmult_1/N1251 ) );
  MUX U6854 ( .IN0(\modmult_1/xin[220] ), .IN1(creg[221]), .SEL(start_in[0]), 
        .F(\modmult_1/N1250 ) );
  ANDN U6855 ( .A(n4110), .B(n3957), .Z(\modmult_1/N125 ) );
  XOR U6856 ( .A(n6047), .B(n6048), .Z(n3957) );
  MUX U6857 ( .IN0(\modmult_1/xin[219] ), .IN1(creg[220]), .SEL(start_in[0]), 
        .F(\modmult_1/N1249 ) );
  MUX U6858 ( .IN0(\modmult_1/xin[218] ), .IN1(creg[219]), .SEL(start_in[0]), 
        .F(\modmult_1/N1248 ) );
  MUX U6859 ( .IN0(\modmult_1/xin[217] ), .IN1(creg[218]), .SEL(start_in[0]), 
        .F(\modmult_1/N1247 ) );
  MUX U6860 ( .IN0(\modmult_1/xin[216] ), .IN1(creg[217]), .SEL(start_in[0]), 
        .F(\modmult_1/N1246 ) );
  MUX U6861 ( .IN0(\modmult_1/xin[215] ), .IN1(creg[216]), .SEL(start_in[0]), 
        .F(\modmult_1/N1245 ) );
  MUX U6862 ( .IN0(\modmult_1/xin[214] ), .IN1(creg[215]), .SEL(start_in[0]), 
        .F(\modmult_1/N1244 ) );
  MUX U6863 ( .IN0(\modmult_1/xin[213] ), .IN1(creg[214]), .SEL(start_in[0]), 
        .F(\modmult_1/N1243 ) );
  MUX U6864 ( .IN0(\modmult_1/xin[212] ), .IN1(creg[213]), .SEL(start_in[0]), 
        .F(\modmult_1/N1242 ) );
  MUX U6865 ( .IN0(\modmult_1/xin[211] ), .IN1(creg[212]), .SEL(start_in[0]), 
        .F(\modmult_1/N1241 ) );
  MUX U6866 ( .IN0(\modmult_1/xin[210] ), .IN1(creg[211]), .SEL(start_in[0]), 
        .F(\modmult_1/N1240 ) );
  ANDN U6867 ( .A(n4110), .B(n3960), .Z(\modmult_1/N124 ) );
  XOR U6868 ( .A(n6049), .B(n6050), .Z(n3960) );
  MUX U6869 ( .IN0(\modmult_1/xin[209] ), .IN1(creg[210]), .SEL(start_in[0]), 
        .F(\modmult_1/N1239 ) );
  MUX U6870 ( .IN0(\modmult_1/xin[208] ), .IN1(creg[209]), .SEL(start_in[0]), 
        .F(\modmult_1/N1238 ) );
  MUX U6871 ( .IN0(\modmult_1/xin[207] ), .IN1(creg[208]), .SEL(start_in[0]), 
        .F(\modmult_1/N1237 ) );
  MUX U6872 ( .IN0(\modmult_1/xin[206] ), .IN1(creg[207]), .SEL(start_in[0]), 
        .F(\modmult_1/N1236 ) );
  MUX U6873 ( .IN0(\modmult_1/xin[205] ), .IN1(creg[206]), .SEL(start_in[0]), 
        .F(\modmult_1/N1235 ) );
  MUX U6874 ( .IN0(\modmult_1/xin[204] ), .IN1(creg[205]), .SEL(start_in[0]), 
        .F(\modmult_1/N1234 ) );
  MUX U6875 ( .IN0(\modmult_1/xin[203] ), .IN1(creg[204]), .SEL(start_in[0]), 
        .F(\modmult_1/N1233 ) );
  MUX U6876 ( .IN0(\modmult_1/xin[202] ), .IN1(creg[203]), .SEL(start_in[0]), 
        .F(\modmult_1/N1232 ) );
  MUX U6877 ( .IN0(\modmult_1/xin[201] ), .IN1(creg[202]), .SEL(start_in[0]), 
        .F(\modmult_1/N1231 ) );
  MUX U6878 ( .IN0(\modmult_1/xin[200] ), .IN1(creg[201]), .SEL(start_in[0]), 
        .F(\modmult_1/N1230 ) );
  ANDN U6879 ( .A(n4110), .B(n3963), .Z(\modmult_1/N123 ) );
  XOR U6880 ( .A(n6051), .B(n6052), .Z(n3963) );
  MUX U6881 ( .IN0(\modmult_1/xin[199] ), .IN1(creg[200]), .SEL(start_in[0]), 
        .F(\modmult_1/N1229 ) );
  MUX U6882 ( .IN0(\modmult_1/xin[198] ), .IN1(creg[199]), .SEL(start_in[0]), 
        .F(\modmult_1/N1228 ) );
  MUX U6883 ( .IN0(\modmult_1/xin[197] ), .IN1(creg[198]), .SEL(start_in[0]), 
        .F(\modmult_1/N1227 ) );
  MUX U6884 ( .IN0(\modmult_1/xin[196] ), .IN1(creg[197]), .SEL(start_in[0]), 
        .F(\modmult_1/N1226 ) );
  MUX U6885 ( .IN0(\modmult_1/xin[195] ), .IN1(creg[196]), .SEL(start_in[0]), 
        .F(\modmult_1/N1225 ) );
  MUX U6886 ( .IN0(\modmult_1/xin[194] ), .IN1(creg[195]), .SEL(start_in[0]), 
        .F(\modmult_1/N1224 ) );
  MUX U6887 ( .IN0(\modmult_1/xin[193] ), .IN1(creg[194]), .SEL(start_in[0]), 
        .F(\modmult_1/N1223 ) );
  MUX U6888 ( .IN0(\modmult_1/xin[192] ), .IN1(creg[193]), .SEL(start_in[0]), 
        .F(\modmult_1/N1222 ) );
  MUX U6889 ( .IN0(\modmult_1/xin[191] ), .IN1(creg[192]), .SEL(start_in[0]), 
        .F(\modmult_1/N1221 ) );
  MUX U6890 ( .IN0(\modmult_1/xin[190] ), .IN1(creg[191]), .SEL(start_in[0]), 
        .F(\modmult_1/N1220 ) );
  ANDN U6891 ( .A(n4110), .B(n3969), .Z(\modmult_1/N122 ) );
  XOR U6892 ( .A(n6053), .B(n6054), .Z(n3969) );
  MUX U6893 ( .IN0(\modmult_1/xin[189] ), .IN1(creg[190]), .SEL(start_in[0]), 
        .F(\modmult_1/N1219 ) );
  MUX U6894 ( .IN0(\modmult_1/xin[188] ), .IN1(creg[189]), .SEL(start_in[0]), 
        .F(\modmult_1/N1218 ) );
  MUX U6895 ( .IN0(\modmult_1/xin[187] ), .IN1(creg[188]), .SEL(start_in[0]), 
        .F(\modmult_1/N1217 ) );
  MUX U6896 ( .IN0(\modmult_1/xin[186] ), .IN1(creg[187]), .SEL(start_in[0]), 
        .F(\modmult_1/N1216 ) );
  MUX U6897 ( .IN0(\modmult_1/xin[185] ), .IN1(creg[186]), .SEL(start_in[0]), 
        .F(\modmult_1/N1215 ) );
  MUX U6898 ( .IN0(\modmult_1/xin[184] ), .IN1(creg[185]), .SEL(start_in[0]), 
        .F(\modmult_1/N1214 ) );
  MUX U6899 ( .IN0(\modmult_1/xin[183] ), .IN1(creg[184]), .SEL(start_in[0]), 
        .F(\modmult_1/N1213 ) );
  MUX U6900 ( .IN0(\modmult_1/xin[182] ), .IN1(creg[183]), .SEL(start_in[0]), 
        .F(\modmult_1/N1212 ) );
  MUX U6901 ( .IN0(\modmult_1/xin[181] ), .IN1(creg[182]), .SEL(start_in[0]), 
        .F(\modmult_1/N1211 ) );
  MUX U6902 ( .IN0(\modmult_1/xin[180] ), .IN1(creg[181]), .SEL(start_in[0]), 
        .F(\modmult_1/N1210 ) );
  ANDN U6903 ( .A(n4110), .B(n3972), .Z(\modmult_1/N121 ) );
  XOR U6904 ( .A(n6055), .B(n6056), .Z(n3972) );
  MUX U6905 ( .IN0(\modmult_1/xin[179] ), .IN1(creg[180]), .SEL(start_in[0]), 
        .F(\modmult_1/N1209 ) );
  MUX U6906 ( .IN0(\modmult_1/xin[178] ), .IN1(creg[179]), .SEL(start_in[0]), 
        .F(\modmult_1/N1208 ) );
  MUX U6907 ( .IN0(\modmult_1/xin[177] ), .IN1(creg[178]), .SEL(start_in[0]), 
        .F(\modmult_1/N1207 ) );
  MUX U6908 ( .IN0(\modmult_1/xin[176] ), .IN1(creg[177]), .SEL(start_in[0]), 
        .F(\modmult_1/N1206 ) );
  MUX U6909 ( .IN0(\modmult_1/xin[175] ), .IN1(creg[176]), .SEL(start_in[0]), 
        .F(\modmult_1/N1205 ) );
  MUX U6910 ( .IN0(\modmult_1/xin[174] ), .IN1(creg[175]), .SEL(start_in[0]), 
        .F(\modmult_1/N1204 ) );
  MUX U6911 ( .IN0(\modmult_1/xin[173] ), .IN1(creg[174]), .SEL(start_in[0]), 
        .F(\modmult_1/N1203 ) );
  MUX U6912 ( .IN0(\modmult_1/xin[172] ), .IN1(creg[173]), .SEL(start_in[0]), 
        .F(\modmult_1/N1202 ) );
  MUX U6913 ( .IN0(\modmult_1/xin[171] ), .IN1(creg[172]), .SEL(start_in[0]), 
        .F(\modmult_1/N1201 ) );
  MUX U6914 ( .IN0(\modmult_1/xin[170] ), .IN1(creg[171]), .SEL(start_in[0]), 
        .F(\modmult_1/N1200 ) );
  ANDN U6915 ( .A(n4110), .B(n3975), .Z(\modmult_1/N120 ) );
  XOR U6916 ( .A(n6057), .B(n6058), .Z(n3975) );
  ANDN U6917 ( .A(n4110), .B(n1034), .Z(\modmult_1/N12 ) );
  XOR U6918 ( .A(n6059), .B(n6060), .Z(n1034) );
  MUX U6919 ( .IN0(\modmult_1/xin[169] ), .IN1(creg[170]), .SEL(start_in[0]), 
        .F(\modmult_1/N1199 ) );
  MUX U6920 ( .IN0(\modmult_1/xin[168] ), .IN1(creg[169]), .SEL(start_in[0]), 
        .F(\modmult_1/N1198 ) );
  MUX U6921 ( .IN0(\modmult_1/xin[167] ), .IN1(creg[168]), .SEL(start_in[0]), 
        .F(\modmult_1/N1197 ) );
  MUX U6922 ( .IN0(\modmult_1/xin[166] ), .IN1(creg[167]), .SEL(start_in[0]), 
        .F(\modmult_1/N1196 ) );
  MUX U6923 ( .IN0(\modmult_1/xin[165] ), .IN1(creg[166]), .SEL(start_in[0]), 
        .F(\modmult_1/N1195 ) );
  MUX U6924 ( .IN0(\modmult_1/xin[164] ), .IN1(creg[165]), .SEL(start_in[0]), 
        .F(\modmult_1/N1194 ) );
  MUX U6925 ( .IN0(\modmult_1/xin[163] ), .IN1(creg[164]), .SEL(start_in[0]), 
        .F(\modmult_1/N1193 ) );
  MUX U6926 ( .IN0(\modmult_1/xin[162] ), .IN1(creg[163]), .SEL(start_in[0]), 
        .F(\modmult_1/N1192 ) );
  MUX U6927 ( .IN0(\modmult_1/xin[161] ), .IN1(creg[162]), .SEL(start_in[0]), 
        .F(\modmult_1/N1191 ) );
  MUX U6928 ( .IN0(\modmult_1/xin[160] ), .IN1(creg[161]), .SEL(start_in[0]), 
        .F(\modmult_1/N1190 ) );
  ANDN U6929 ( .A(n4110), .B(n3978), .Z(\modmult_1/N119 ) );
  XOR U6930 ( .A(n6061), .B(n6062), .Z(n3978) );
  MUX U6931 ( .IN0(\modmult_1/xin[159] ), .IN1(creg[160]), .SEL(start_in[0]), 
        .F(\modmult_1/N1189 ) );
  MUX U6932 ( .IN0(\modmult_1/xin[158] ), .IN1(creg[159]), .SEL(start_in[0]), 
        .F(\modmult_1/N1188 ) );
  MUX U6933 ( .IN0(\modmult_1/xin[157] ), .IN1(creg[158]), .SEL(start_in[0]), 
        .F(\modmult_1/N1187 ) );
  MUX U6934 ( .IN0(\modmult_1/xin[156] ), .IN1(creg[157]), .SEL(start_in[0]), 
        .F(\modmult_1/N1186 ) );
  MUX U6935 ( .IN0(\modmult_1/xin[155] ), .IN1(creg[156]), .SEL(start_in[0]), 
        .F(\modmult_1/N1185 ) );
  MUX U6936 ( .IN0(\modmult_1/xin[154] ), .IN1(creg[155]), .SEL(start_in[0]), 
        .F(\modmult_1/N1184 ) );
  MUX U6937 ( .IN0(\modmult_1/xin[153] ), .IN1(creg[154]), .SEL(start_in[0]), 
        .F(\modmult_1/N1183 ) );
  MUX U6938 ( .IN0(\modmult_1/xin[152] ), .IN1(creg[153]), .SEL(start_in[0]), 
        .F(\modmult_1/N1182 ) );
  MUX U6939 ( .IN0(\modmult_1/xin[151] ), .IN1(creg[152]), .SEL(start_in[0]), 
        .F(\modmult_1/N1181 ) );
  MUX U6940 ( .IN0(\modmult_1/xin[150] ), .IN1(creg[151]), .SEL(start_in[0]), 
        .F(\modmult_1/N1180 ) );
  ANDN U6941 ( .A(n4110), .B(n3981), .Z(\modmult_1/N118 ) );
  XOR U6942 ( .A(n6063), .B(n6064), .Z(n3981) );
  MUX U6943 ( .IN0(\modmult_1/xin[149] ), .IN1(creg[150]), .SEL(start_in[0]), 
        .F(\modmult_1/N1179 ) );
  MUX U6944 ( .IN0(\modmult_1/xin[148] ), .IN1(creg[149]), .SEL(start_in[0]), 
        .F(\modmult_1/N1178 ) );
  MUX U6945 ( .IN0(\modmult_1/xin[147] ), .IN1(creg[148]), .SEL(start_in[0]), 
        .F(\modmult_1/N1177 ) );
  MUX U6946 ( .IN0(\modmult_1/xin[146] ), .IN1(creg[147]), .SEL(start_in[0]), 
        .F(\modmult_1/N1176 ) );
  MUX U6947 ( .IN0(\modmult_1/xin[145] ), .IN1(creg[146]), .SEL(start_in[0]), 
        .F(\modmult_1/N1175 ) );
  MUX U6948 ( .IN0(\modmult_1/xin[144] ), .IN1(creg[145]), .SEL(start_in[0]), 
        .F(\modmult_1/N1174 ) );
  MUX U6949 ( .IN0(\modmult_1/xin[143] ), .IN1(creg[144]), .SEL(start_in[0]), 
        .F(\modmult_1/N1173 ) );
  MUX U6950 ( .IN0(\modmult_1/xin[142] ), .IN1(creg[143]), .SEL(start_in[0]), 
        .F(\modmult_1/N1172 ) );
  MUX U6951 ( .IN0(\modmult_1/xin[141] ), .IN1(creg[142]), .SEL(start_in[0]), 
        .F(\modmult_1/N1171 ) );
  MUX U6952 ( .IN0(\modmult_1/xin[140] ), .IN1(creg[141]), .SEL(start_in[0]), 
        .F(\modmult_1/N1170 ) );
  ANDN U6953 ( .A(n4110), .B(n3984), .Z(\modmult_1/N117 ) );
  XOR U6954 ( .A(n6065), .B(n6066), .Z(n3984) );
  MUX U6955 ( .IN0(\modmult_1/xin[139] ), .IN1(creg[140]), .SEL(start_in[0]), 
        .F(\modmult_1/N1169 ) );
  MUX U6956 ( .IN0(\modmult_1/xin[138] ), .IN1(creg[139]), .SEL(start_in[0]), 
        .F(\modmult_1/N1168 ) );
  MUX U6957 ( .IN0(\modmult_1/xin[137] ), .IN1(creg[138]), .SEL(start_in[0]), 
        .F(\modmult_1/N1167 ) );
  MUX U6958 ( .IN0(\modmult_1/xin[136] ), .IN1(creg[137]), .SEL(start_in[0]), 
        .F(\modmult_1/N1166 ) );
  MUX U6959 ( .IN0(\modmult_1/xin[135] ), .IN1(creg[136]), .SEL(start_in[0]), 
        .F(\modmult_1/N1165 ) );
  MUX U6960 ( .IN0(\modmult_1/xin[134] ), .IN1(creg[135]), .SEL(start_in[0]), 
        .F(\modmult_1/N1164 ) );
  MUX U6961 ( .IN0(\modmult_1/xin[133] ), .IN1(creg[134]), .SEL(start_in[0]), 
        .F(\modmult_1/N1163 ) );
  MUX U6962 ( .IN0(\modmult_1/xin[132] ), .IN1(creg[133]), .SEL(start_in[0]), 
        .F(\modmult_1/N1162 ) );
  MUX U6963 ( .IN0(\modmult_1/xin[131] ), .IN1(creg[132]), .SEL(start_in[0]), 
        .F(\modmult_1/N1161 ) );
  MUX U6964 ( .IN0(\modmult_1/xin[130] ), .IN1(creg[131]), .SEL(start_in[0]), 
        .F(\modmult_1/N1160 ) );
  ANDN U6965 ( .A(n4110), .B(n3987), .Z(\modmult_1/N116 ) );
  XOR U6966 ( .A(n6067), .B(n6068), .Z(n3987) );
  MUX U6967 ( .IN0(\modmult_1/xin[129] ), .IN1(creg[130]), .SEL(start_in[0]), 
        .F(\modmult_1/N1159 ) );
  MUX U6968 ( .IN0(\modmult_1/xin[128] ), .IN1(creg[129]), .SEL(start_in[0]), 
        .F(\modmult_1/N1158 ) );
  MUX U6969 ( .IN0(\modmult_1/xin[127] ), .IN1(creg[128]), .SEL(start_in[0]), 
        .F(\modmult_1/N1157 ) );
  MUX U6970 ( .IN0(\modmult_1/xin[126] ), .IN1(creg[127]), .SEL(start_in[0]), 
        .F(\modmult_1/N1156 ) );
  MUX U6971 ( .IN0(\modmult_1/xin[125] ), .IN1(creg[126]), .SEL(start_in[0]), 
        .F(\modmult_1/N1155 ) );
  MUX U6972 ( .IN0(\modmult_1/xin[124] ), .IN1(creg[125]), .SEL(start_in[0]), 
        .F(\modmult_1/N1154 ) );
  MUX U6973 ( .IN0(\modmult_1/xin[123] ), .IN1(creg[124]), .SEL(start_in[0]), 
        .F(\modmult_1/N1153 ) );
  MUX U6974 ( .IN0(\modmult_1/xin[122] ), .IN1(creg[123]), .SEL(start_in[0]), 
        .F(\modmult_1/N1152 ) );
  MUX U6975 ( .IN0(\modmult_1/xin[121] ), .IN1(creg[122]), .SEL(start_in[0]), 
        .F(\modmult_1/N1151 ) );
  MUX U6976 ( .IN0(\modmult_1/xin[120] ), .IN1(creg[121]), .SEL(start_in[0]), 
        .F(\modmult_1/N1150 ) );
  ANDN U6977 ( .A(n4110), .B(n3990), .Z(\modmult_1/N115 ) );
  XOR U6978 ( .A(n6069), .B(n6070), .Z(n3990) );
  MUX U6979 ( .IN0(\modmult_1/xin[119] ), .IN1(creg[120]), .SEL(start_in[0]), 
        .F(\modmult_1/N1149 ) );
  MUX U6980 ( .IN0(\modmult_1/xin[118] ), .IN1(creg[119]), .SEL(start_in[0]), 
        .F(\modmult_1/N1148 ) );
  MUX U6981 ( .IN0(\modmult_1/xin[117] ), .IN1(creg[118]), .SEL(start_in[0]), 
        .F(\modmult_1/N1147 ) );
  MUX U6982 ( .IN0(\modmult_1/xin[116] ), .IN1(creg[117]), .SEL(start_in[0]), 
        .F(\modmult_1/N1146 ) );
  MUX U6983 ( .IN0(\modmult_1/xin[115] ), .IN1(creg[116]), .SEL(start_in[0]), 
        .F(\modmult_1/N1145 ) );
  MUX U6984 ( .IN0(\modmult_1/xin[114] ), .IN1(creg[115]), .SEL(start_in[0]), 
        .F(\modmult_1/N1144 ) );
  MUX U6985 ( .IN0(\modmult_1/xin[113] ), .IN1(creg[114]), .SEL(start_in[0]), 
        .F(\modmult_1/N1143 ) );
  MUX U6986 ( .IN0(\modmult_1/xin[112] ), .IN1(creg[113]), .SEL(start_in[0]), 
        .F(\modmult_1/N1142 ) );
  MUX U6987 ( .IN0(\modmult_1/xin[111] ), .IN1(creg[112]), .SEL(start_in[0]), 
        .F(\modmult_1/N1141 ) );
  MUX U6988 ( .IN0(\modmult_1/xin[110] ), .IN1(creg[111]), .SEL(start_in[0]), 
        .F(\modmult_1/N1140 ) );
  ANDN U6989 ( .A(n4110), .B(n3993), .Z(\modmult_1/N114 ) );
  XOR U6990 ( .A(n6071), .B(n6072), .Z(n3993) );
  MUX U6991 ( .IN0(\modmult_1/xin[109] ), .IN1(creg[110]), .SEL(start_in[0]), 
        .F(\modmult_1/N1139 ) );
  MUX U6992 ( .IN0(\modmult_1/xin[108] ), .IN1(creg[109]), .SEL(start_in[0]), 
        .F(\modmult_1/N1138 ) );
  MUX U6993 ( .IN0(\modmult_1/xin[107] ), .IN1(creg[108]), .SEL(start_in[0]), 
        .F(\modmult_1/N1137 ) );
  MUX U6994 ( .IN0(\modmult_1/xin[106] ), .IN1(creg[107]), .SEL(start_in[0]), 
        .F(\modmult_1/N1136 ) );
  MUX U6995 ( .IN0(\modmult_1/xin[105] ), .IN1(creg[106]), .SEL(start_in[0]), 
        .F(\modmult_1/N1135 ) );
  MUX U6996 ( .IN0(\modmult_1/xin[104] ), .IN1(creg[105]), .SEL(start_in[0]), 
        .F(\modmult_1/N1134 ) );
  MUX U6997 ( .IN0(\modmult_1/xin[103] ), .IN1(creg[104]), .SEL(start_in[0]), 
        .F(\modmult_1/N1133 ) );
  MUX U6998 ( .IN0(\modmult_1/xin[102] ), .IN1(creg[103]), .SEL(start_in[0]), 
        .F(\modmult_1/N1132 ) );
  MUX U6999 ( .IN0(\modmult_1/xin[101] ), .IN1(creg[102]), .SEL(start_in[0]), 
        .F(\modmult_1/N1131 ) );
  MUX U7000 ( .IN0(\modmult_1/xin[100] ), .IN1(creg[101]), .SEL(start_in[0]), 
        .F(\modmult_1/N1130 ) );
  ANDN U7001 ( .A(n4110), .B(n3996), .Z(\modmult_1/N113 ) );
  XOR U7002 ( .A(n6073), .B(n6074), .Z(n3996) );
  MUX U7003 ( .IN0(\modmult_1/xin[99] ), .IN1(creg[100]), .SEL(start_in[0]), 
        .F(\modmult_1/N1129 ) );
  MUX U7004 ( .IN0(\modmult_1/xin[98] ), .IN1(creg[99]), .SEL(start_in[0]), 
        .F(\modmult_1/N1128 ) );
  MUX U7005 ( .IN0(\modmult_1/xin[97] ), .IN1(creg[98]), .SEL(start_in[0]), 
        .F(\modmult_1/N1127 ) );
  MUX U7006 ( .IN0(\modmult_1/xin[96] ), .IN1(creg[97]), .SEL(start_in[0]), 
        .F(\modmult_1/N1126 ) );
  MUX U7007 ( .IN0(\modmult_1/xin[95] ), .IN1(creg[96]), .SEL(start_in[0]), 
        .F(\modmult_1/N1125 ) );
  MUX U7008 ( .IN0(\modmult_1/xin[94] ), .IN1(creg[95]), .SEL(start_in[0]), 
        .F(\modmult_1/N1124 ) );
  MUX U7009 ( .IN0(\modmult_1/xin[93] ), .IN1(creg[94]), .SEL(start_in[0]), 
        .F(\modmult_1/N1123 ) );
  MUX U7010 ( .IN0(\modmult_1/xin[92] ), .IN1(creg[93]), .SEL(start_in[0]), 
        .F(\modmult_1/N1122 ) );
  MUX U7011 ( .IN0(\modmult_1/xin[91] ), .IN1(creg[92]), .SEL(start_in[0]), 
        .F(\modmult_1/N1121 ) );
  MUX U7012 ( .IN0(\modmult_1/xin[90] ), .IN1(creg[91]), .SEL(start_in[0]), 
        .F(\modmult_1/N1120 ) );
  ANDN U7013 ( .A(n4110), .B(n4002), .Z(\modmult_1/N112 ) );
  XOR U7014 ( .A(n6075), .B(n6076), .Z(n4002) );
  MUX U7015 ( .IN0(\modmult_1/xin[89] ), .IN1(creg[90]), .SEL(start_in[0]), 
        .F(\modmult_1/N1119 ) );
  MUX U7016 ( .IN0(\modmult_1/xin[88] ), .IN1(creg[89]), .SEL(start_in[0]), 
        .F(\modmult_1/N1118 ) );
  MUX U7017 ( .IN0(\modmult_1/xin[87] ), .IN1(creg[88]), .SEL(start_in[0]), 
        .F(\modmult_1/N1117 ) );
  MUX U7018 ( .IN0(\modmult_1/xin[86] ), .IN1(creg[87]), .SEL(start_in[0]), 
        .F(\modmult_1/N1116 ) );
  MUX U7019 ( .IN0(\modmult_1/xin[85] ), .IN1(creg[86]), .SEL(start_in[0]), 
        .F(\modmult_1/N1115 ) );
  MUX U7020 ( .IN0(\modmult_1/xin[84] ), .IN1(creg[85]), .SEL(start_in[0]), 
        .F(\modmult_1/N1114 ) );
  MUX U7021 ( .IN0(\modmult_1/xin[83] ), .IN1(creg[84]), .SEL(start_in[0]), 
        .F(\modmult_1/N1113 ) );
  MUX U7022 ( .IN0(\modmult_1/xin[82] ), .IN1(creg[83]), .SEL(start_in[0]), 
        .F(\modmult_1/N1112 ) );
  MUX U7023 ( .IN0(\modmult_1/xin[81] ), .IN1(creg[82]), .SEL(start_in[0]), 
        .F(\modmult_1/N1111 ) );
  MUX U7024 ( .IN0(\modmult_1/xin[80] ), .IN1(creg[81]), .SEL(start_in[0]), 
        .F(\modmult_1/N1110 ) );
  ANDN U7025 ( .A(n4110), .B(n4005), .Z(\modmult_1/N111 ) );
  XOR U7026 ( .A(n6077), .B(n6078), .Z(n4005) );
  MUX U7027 ( .IN0(\modmult_1/xin[79] ), .IN1(creg[80]), .SEL(start_in[0]), 
        .F(\modmult_1/N1109 ) );
  MUX U7028 ( .IN0(\modmult_1/xin[78] ), .IN1(creg[79]), .SEL(start_in[0]), 
        .F(\modmult_1/N1108 ) );
  MUX U7029 ( .IN0(\modmult_1/xin[77] ), .IN1(creg[78]), .SEL(start_in[0]), 
        .F(\modmult_1/N1107 ) );
  MUX U7030 ( .IN0(\modmult_1/xin[76] ), .IN1(creg[77]), .SEL(start_in[0]), 
        .F(\modmult_1/N1106 ) );
  MUX U7031 ( .IN0(\modmult_1/xin[75] ), .IN1(creg[76]), .SEL(start_in[0]), 
        .F(\modmult_1/N1105 ) );
  MUX U7032 ( .IN0(\modmult_1/xin[74] ), .IN1(creg[75]), .SEL(start_in[0]), 
        .F(\modmult_1/N1104 ) );
  MUX U7033 ( .IN0(\modmult_1/xin[73] ), .IN1(creg[74]), .SEL(start_in[0]), 
        .F(\modmult_1/N1103 ) );
  MUX U7034 ( .IN0(\modmult_1/xin[72] ), .IN1(creg[73]), .SEL(start_in[0]), 
        .F(\modmult_1/N1102 ) );
  MUX U7035 ( .IN0(\modmult_1/xin[71] ), .IN1(creg[72]), .SEL(start_in[0]), 
        .F(\modmult_1/N1101 ) );
  MUX U7036 ( .IN0(\modmult_1/xin[70] ), .IN1(creg[71]), .SEL(start_in[0]), 
        .F(\modmult_1/N1100 ) );
  ANDN U7037 ( .A(n4110), .B(n4008), .Z(\modmult_1/N110 ) );
  XOR U7038 ( .A(n6079), .B(n6080), .Z(n4008) );
  ANDN U7039 ( .A(n4110), .B(n1368), .Z(\modmult_1/N11 ) );
  XOR U7040 ( .A(n6081), .B(n6082), .Z(n1368) );
  MUX U7041 ( .IN0(\modmult_1/xin[69] ), .IN1(creg[70]), .SEL(start_in[0]), 
        .F(\modmult_1/N1099 ) );
  MUX U7042 ( .IN0(\modmult_1/xin[68] ), .IN1(creg[69]), .SEL(start_in[0]), 
        .F(\modmult_1/N1098 ) );
  MUX U7043 ( .IN0(\modmult_1/xin[67] ), .IN1(creg[68]), .SEL(start_in[0]), 
        .F(\modmult_1/N1097 ) );
  MUX U7044 ( .IN0(\modmult_1/xin[66] ), .IN1(creg[67]), .SEL(start_in[0]), 
        .F(\modmult_1/N1096 ) );
  MUX U7045 ( .IN0(\modmult_1/xin[65] ), .IN1(creg[66]), .SEL(start_in[0]), 
        .F(\modmult_1/N1095 ) );
  MUX U7046 ( .IN0(\modmult_1/xin[64] ), .IN1(creg[65]), .SEL(start_in[0]), 
        .F(\modmult_1/N1094 ) );
  MUX U7047 ( .IN0(\modmult_1/xin[63] ), .IN1(creg[64]), .SEL(start_in[0]), 
        .F(\modmult_1/N1093 ) );
  MUX U7048 ( .IN0(\modmult_1/xin[62] ), .IN1(creg[63]), .SEL(start_in[0]), 
        .F(\modmult_1/N1092 ) );
  MUX U7049 ( .IN0(\modmult_1/xin[61] ), .IN1(creg[62]), .SEL(start_in[0]), 
        .F(\modmult_1/N1091 ) );
  MUX U7050 ( .IN0(\modmult_1/xin[60] ), .IN1(creg[61]), .SEL(start_in[0]), 
        .F(\modmult_1/N1090 ) );
  ANDN U7051 ( .A(n4110), .B(n4011), .Z(\modmult_1/N109 ) );
  XOR U7052 ( .A(n6083), .B(n6084), .Z(n4011) );
  MUX U7053 ( .IN0(\modmult_1/xin[59] ), .IN1(creg[60]), .SEL(start_in[0]), 
        .F(\modmult_1/N1089 ) );
  MUX U7054 ( .IN0(\modmult_1/xin[58] ), .IN1(creg[59]), .SEL(start_in[0]), 
        .F(\modmult_1/N1088 ) );
  MUX U7055 ( .IN0(\modmult_1/xin[57] ), .IN1(creg[58]), .SEL(start_in[0]), 
        .F(\modmult_1/N1087 ) );
  MUX U7056 ( .IN0(\modmult_1/xin[56] ), .IN1(creg[57]), .SEL(start_in[0]), 
        .F(\modmult_1/N1086 ) );
  MUX U7057 ( .IN0(\modmult_1/xin[55] ), .IN1(creg[56]), .SEL(start_in[0]), 
        .F(\modmult_1/N1085 ) );
  MUX U7058 ( .IN0(\modmult_1/xin[54] ), .IN1(creg[55]), .SEL(start_in[0]), 
        .F(\modmult_1/N1084 ) );
  MUX U7059 ( .IN0(\modmult_1/xin[53] ), .IN1(creg[54]), .SEL(start_in[0]), 
        .F(\modmult_1/N1083 ) );
  MUX U7060 ( .IN0(\modmult_1/xin[52] ), .IN1(creg[53]), .SEL(start_in[0]), 
        .F(\modmult_1/N1082 ) );
  MUX U7061 ( .IN0(\modmult_1/xin[51] ), .IN1(creg[52]), .SEL(start_in[0]), 
        .F(\modmult_1/N1081 ) );
  MUX U7062 ( .IN0(\modmult_1/xin[50] ), .IN1(creg[51]), .SEL(start_in[0]), 
        .F(\modmult_1/N1080 ) );
  ANDN U7063 ( .A(n4110), .B(n4014), .Z(\modmult_1/N108 ) );
  XOR U7064 ( .A(n6085), .B(n6086), .Z(n4014) );
  MUX U7065 ( .IN0(\modmult_1/xin[49] ), .IN1(creg[50]), .SEL(start_in[0]), 
        .F(\modmult_1/N1079 ) );
  MUX U7066 ( .IN0(\modmult_1/xin[48] ), .IN1(creg[49]), .SEL(start_in[0]), 
        .F(\modmult_1/N1078 ) );
  MUX U7067 ( .IN0(\modmult_1/xin[47] ), .IN1(creg[48]), .SEL(start_in[0]), 
        .F(\modmult_1/N1077 ) );
  MUX U7068 ( .IN0(\modmult_1/xin[46] ), .IN1(creg[47]), .SEL(start_in[0]), 
        .F(\modmult_1/N1076 ) );
  MUX U7069 ( .IN0(\modmult_1/xin[45] ), .IN1(creg[46]), .SEL(start_in[0]), 
        .F(\modmult_1/N1075 ) );
  MUX U7070 ( .IN0(\modmult_1/xin[44] ), .IN1(creg[45]), .SEL(start_in[0]), 
        .F(\modmult_1/N1074 ) );
  MUX U7071 ( .IN0(\modmult_1/xin[43] ), .IN1(creg[44]), .SEL(start_in[0]), 
        .F(\modmult_1/N1073 ) );
  MUX U7072 ( .IN0(\modmult_1/xin[42] ), .IN1(creg[43]), .SEL(start_in[0]), 
        .F(\modmult_1/N1072 ) );
  MUX U7073 ( .IN0(\modmult_1/xin[41] ), .IN1(creg[42]), .SEL(start_in[0]), 
        .F(\modmult_1/N1071 ) );
  MUX U7074 ( .IN0(\modmult_1/xin[40] ), .IN1(creg[41]), .SEL(start_in[0]), 
        .F(\modmult_1/N1070 ) );
  ANDN U7075 ( .A(n4110), .B(n4017), .Z(\modmult_1/N107 ) );
  XOR U7076 ( .A(n6087), .B(n6088), .Z(n4017) );
  MUX U7077 ( .IN0(\modmult_1/xin[39] ), .IN1(creg[40]), .SEL(start_in[0]), 
        .F(\modmult_1/N1069 ) );
  MUX U7078 ( .IN0(\modmult_1/xin[38] ), .IN1(creg[39]), .SEL(start_in[0]), 
        .F(\modmult_1/N1068 ) );
  MUX U7079 ( .IN0(\modmult_1/xin[37] ), .IN1(creg[38]), .SEL(start_in[0]), 
        .F(\modmult_1/N1067 ) );
  MUX U7080 ( .IN0(\modmult_1/xin[36] ), .IN1(creg[37]), .SEL(start_in[0]), 
        .F(\modmult_1/N1066 ) );
  MUX U7081 ( .IN0(\modmult_1/xin[35] ), .IN1(creg[36]), .SEL(start_in[0]), 
        .F(\modmult_1/N1065 ) );
  MUX U7082 ( .IN0(\modmult_1/xin[34] ), .IN1(creg[35]), .SEL(start_in[0]), 
        .F(\modmult_1/N1064 ) );
  MUX U7083 ( .IN0(\modmult_1/xin[33] ), .IN1(creg[34]), .SEL(start_in[0]), 
        .F(\modmult_1/N1063 ) );
  MUX U7084 ( .IN0(\modmult_1/xin[32] ), .IN1(creg[33]), .SEL(start_in[0]), 
        .F(\modmult_1/N1062 ) );
  MUX U7085 ( .IN0(\modmult_1/xin[31] ), .IN1(creg[32]), .SEL(start_in[0]), 
        .F(\modmult_1/N1061 ) );
  MUX U7086 ( .IN0(\modmult_1/xin[30] ), .IN1(creg[31]), .SEL(start_in[0]), 
        .F(\modmult_1/N1060 ) );
  ANDN U7087 ( .A(n4110), .B(n4020), .Z(\modmult_1/N106 ) );
  XOR U7088 ( .A(n6089), .B(n6090), .Z(n4020) );
  MUX U7089 ( .IN0(\modmult_1/xin[29] ), .IN1(creg[30]), .SEL(start_in[0]), 
        .F(\modmult_1/N1059 ) );
  MUX U7090 ( .IN0(\modmult_1/xin[28] ), .IN1(creg[29]), .SEL(start_in[0]), 
        .F(\modmult_1/N1058 ) );
  MUX U7091 ( .IN0(\modmult_1/xin[27] ), .IN1(creg[28]), .SEL(start_in[0]), 
        .F(\modmult_1/N1057 ) );
  MUX U7092 ( .IN0(\modmult_1/xin[26] ), .IN1(creg[27]), .SEL(start_in[0]), 
        .F(\modmult_1/N1056 ) );
  MUX U7093 ( .IN0(\modmult_1/xin[25] ), .IN1(creg[26]), .SEL(start_in[0]), 
        .F(\modmult_1/N1055 ) );
  MUX U7094 ( .IN0(\modmult_1/xin[24] ), .IN1(creg[25]), .SEL(start_in[0]), 
        .F(\modmult_1/N1054 ) );
  MUX U7095 ( .IN0(\modmult_1/xin[23] ), .IN1(creg[24]), .SEL(start_in[0]), 
        .F(\modmult_1/N1053 ) );
  MUX U7096 ( .IN0(\modmult_1/xin[22] ), .IN1(creg[23]), .SEL(start_in[0]), 
        .F(\modmult_1/N1052 ) );
  MUX U7097 ( .IN0(\modmult_1/xin[21] ), .IN1(creg[22]), .SEL(start_in[0]), 
        .F(\modmult_1/N1051 ) );
  MUX U7098 ( .IN0(\modmult_1/xin[20] ), .IN1(creg[21]), .SEL(start_in[0]), 
        .F(\modmult_1/N1050 ) );
  ANDN U7099 ( .A(n4110), .B(n4023), .Z(\modmult_1/N105 ) );
  XOR U7100 ( .A(n6091), .B(n6092), .Z(n4023) );
  MUX U7101 ( .IN0(\modmult_1/xin[19] ), .IN1(creg[20]), .SEL(start_in[0]), 
        .F(\modmult_1/N1049 ) );
  MUX U7102 ( .IN0(\modmult_1/xin[18] ), .IN1(creg[19]), .SEL(start_in[0]), 
        .F(\modmult_1/N1048 ) );
  MUX U7103 ( .IN0(\modmult_1/xin[17] ), .IN1(creg[18]), .SEL(start_in[0]), 
        .F(\modmult_1/N1047 ) );
  MUX U7104 ( .IN0(\modmult_1/xin[16] ), .IN1(creg[17]), .SEL(start_in[0]), 
        .F(\modmult_1/N1046 ) );
  MUX U7105 ( .IN0(\modmult_1/xin[15] ), .IN1(creg[16]), .SEL(start_in[0]), 
        .F(\modmult_1/N1045 ) );
  MUX U7106 ( .IN0(\modmult_1/xin[14] ), .IN1(creg[15]), .SEL(start_in[0]), 
        .F(\modmult_1/N1044 ) );
  MUX U7107 ( .IN0(\modmult_1/xin[13] ), .IN1(creg[14]), .SEL(start_in[0]), 
        .F(\modmult_1/N1043 ) );
  MUX U7108 ( .IN0(\modmult_1/xin[12] ), .IN1(creg[13]), .SEL(start_in[0]), 
        .F(\modmult_1/N1042 ) );
  MUX U7109 ( .IN0(\modmult_1/xin[11] ), .IN1(creg[12]), .SEL(start_in[0]), 
        .F(\modmult_1/N1041 ) );
  MUX U7110 ( .IN0(\modmult_1/xin[10] ), .IN1(creg[11]), .SEL(start_in[0]), 
        .F(\modmult_1/N1040 ) );
  ANDN U7111 ( .A(n4110), .B(n4038), .Z(\modmult_1/N104 ) );
  XOR U7112 ( .A(n6093), .B(n6094), .Z(n4038) );
  MUX U7113 ( .IN0(\modmult_1/xin[9] ), .IN1(creg[10]), .SEL(start_in[0]), .F(
        \modmult_1/N1039 ) );
  MUX U7114 ( .IN0(\modmult_1/xin[8] ), .IN1(creg[9]), .SEL(start_in[0]), .F(
        \modmult_1/N1038 ) );
  MUX U7115 ( .IN0(\modmult_1/xin[7] ), .IN1(creg[8]), .SEL(start_in[0]), .F(
        \modmult_1/N1037 ) );
  MUX U7116 ( .IN0(\modmult_1/xin[6] ), .IN1(creg[7]), .SEL(start_in[0]), .F(
        \modmult_1/N1036 ) );
  MUX U7117 ( .IN0(\modmult_1/xin[5] ), .IN1(creg[6]), .SEL(start_in[0]), .F(
        \modmult_1/N1035 ) );
  MUX U7118 ( .IN0(\modmult_1/xin[4] ), .IN1(creg[5]), .SEL(start_in[0]), .F(
        \modmult_1/N1034 ) );
  MUX U7119 ( .IN0(\modmult_1/xin[3] ), .IN1(creg[4]), .SEL(start_in[0]), .F(
        \modmult_1/N1033 ) );
  MUX U7120 ( .IN0(\modmult_1/xin[2] ), .IN1(creg[3]), .SEL(start_in[0]), .F(
        \modmult_1/N1032 ) );
  MUX U7121 ( .IN0(\modmult_1/xin[1] ), .IN1(creg[2]), .SEL(start_in[0]), .F(
        \modmult_1/N1031 ) );
  MUX U7122 ( .IN0(\modmult_1/xin[0] ), .IN1(creg[1]), .SEL(start_in[0]), .F(
        \modmult_1/N1030 ) );
  ANDN U7123 ( .A(n4110), .B(n4071), .Z(\modmult_1/N103 ) );
  XOR U7124 ( .A(n6095), .B(n6096), .Z(n4071) );
  AND U7125 ( .A(creg[0]), .B(start_in[0]), .Z(\modmult_1/N1029 ) );
  AND U7126 ( .A(n6097), .B(n4110), .Z(\modmult_1/N1027 ) );
  XNOR U7127 ( .A(n6098), .B(n6099), .Z(n6097) );
  XOR U7128 ( .A(n6100), .B(n6101), .Z(n6099) );
  ANDN U7129 ( .A(n6102), .B(n6103), .Z(n6100) );
  XNOR U7130 ( .A(n6104), .B(n6105), .Z(n6102) );
  ANDN U7131 ( .A(n4110), .B(n4026), .Z(\modmult_1/N1026 ) );
  XOR U7132 ( .A(n6103), .B(n6104), .Z(n4026) );
  NAND U7133 ( .A(n6106), .B(nreg[1023]), .Z(n6104) );
  NAND U7134 ( .A(n6107), .B(nreg[1023]), .Z(n6106) );
  XOR U7135 ( .A(n6098), .B(n6108), .Z(n6103) );
  IV U7136 ( .A(n6105), .Z(n6098) );
  XOR U7137 ( .A(n6109), .B(n6110), .Z(n6105) );
  ANDN U7138 ( .A(n6111), .B(n6112), .Z(n6110) );
  XNOR U7139 ( .A(n6113), .B(n6109), .Z(n6111) );
  ANDN U7140 ( .A(n4110), .B(n4029), .Z(\modmult_1/N1025 ) );
  XOR U7141 ( .A(n6112), .B(n6113), .Z(n4029) );
  NAND U7142 ( .A(n6114), .B(nreg[1022]), .Z(n6113) );
  NAND U7143 ( .A(n6107), .B(nreg[1022]), .Z(n6114) );
  XOR U7144 ( .A(n6115), .B(n6116), .Z(n6112) );
  IV U7145 ( .A(n6109), .Z(n6115) );
  XOR U7146 ( .A(n6117), .B(n6118), .Z(n6109) );
  ANDN U7147 ( .A(n6119), .B(n6120), .Z(n6118) );
  XNOR U7148 ( .A(n6121), .B(n6117), .Z(n6119) );
  ANDN U7149 ( .A(n4110), .B(n4032), .Z(\modmult_1/N1024 ) );
  XOR U7150 ( .A(n6120), .B(n6121), .Z(n4032) );
  NAND U7151 ( .A(n6122), .B(nreg[1021]), .Z(n6121) );
  NAND U7152 ( .A(n6107), .B(nreg[1021]), .Z(n6122) );
  XOR U7153 ( .A(n6123), .B(n6124), .Z(n6120) );
  IV U7154 ( .A(n6117), .Z(n6123) );
  XOR U7155 ( .A(n6125), .B(n6126), .Z(n6117) );
  ANDN U7156 ( .A(n6127), .B(n6128), .Z(n6126) );
  XNOR U7157 ( .A(n6129), .B(n6125), .Z(n6127) );
  ANDN U7158 ( .A(n4110), .B(n4035), .Z(\modmult_1/N1023 ) );
  XOR U7159 ( .A(n6128), .B(n6129), .Z(n4035) );
  NAND U7160 ( .A(n6130), .B(nreg[1020]), .Z(n6129) );
  NAND U7161 ( .A(n6107), .B(nreg[1020]), .Z(n6130) );
  XOR U7162 ( .A(n6131), .B(n6132), .Z(n6128) );
  IV U7163 ( .A(n6125), .Z(n6131) );
  XOR U7164 ( .A(n6133), .B(n6134), .Z(n6125) );
  ANDN U7165 ( .A(n6135), .B(n6136), .Z(n6134) );
  XNOR U7166 ( .A(n6137), .B(n6133), .Z(n6135) );
  ANDN U7167 ( .A(n4110), .B(n4041), .Z(\modmult_1/N1022 ) );
  XOR U7168 ( .A(n6136), .B(n6137), .Z(n4041) );
  NAND U7169 ( .A(n6138), .B(nreg[1019]), .Z(n6137) );
  NAND U7170 ( .A(n6107), .B(nreg[1019]), .Z(n6138) );
  XOR U7171 ( .A(n6139), .B(n6140), .Z(n6136) );
  IV U7172 ( .A(n6133), .Z(n6139) );
  XOR U7173 ( .A(n6141), .B(n6142), .Z(n6133) );
  ANDN U7174 ( .A(n6143), .B(n6144), .Z(n6142) );
  XNOR U7175 ( .A(n6145), .B(n6141), .Z(n6143) );
  ANDN U7176 ( .A(n4110), .B(n4044), .Z(\modmult_1/N1021 ) );
  XOR U7177 ( .A(n6144), .B(n6145), .Z(n4044) );
  NAND U7178 ( .A(n6146), .B(nreg[1018]), .Z(n6145) );
  NAND U7179 ( .A(n6107), .B(nreg[1018]), .Z(n6146) );
  XOR U7180 ( .A(n6147), .B(n6148), .Z(n6144) );
  IV U7181 ( .A(n6141), .Z(n6147) );
  XOR U7182 ( .A(n6149), .B(n6150), .Z(n6141) );
  ANDN U7183 ( .A(n6151), .B(n6152), .Z(n6150) );
  XNOR U7184 ( .A(n6153), .B(n6149), .Z(n6151) );
  ANDN U7185 ( .A(n4110), .B(n4047), .Z(\modmult_1/N1020 ) );
  XOR U7186 ( .A(n6152), .B(n6153), .Z(n4047) );
  NAND U7187 ( .A(n6154), .B(nreg[1017]), .Z(n6153) );
  NAND U7188 ( .A(n6107), .B(nreg[1017]), .Z(n6154) );
  XOR U7189 ( .A(n6155), .B(n6156), .Z(n6152) );
  IV U7190 ( .A(n6149), .Z(n6155) );
  XOR U7191 ( .A(n6157), .B(n6158), .Z(n6149) );
  ANDN U7192 ( .A(n6159), .B(n6160), .Z(n6158) );
  XNOR U7193 ( .A(n6161), .B(n6157), .Z(n6159) );
  ANDN U7194 ( .A(n4110), .B(n1038), .Z(\modmult_1/N102 ) );
  XOR U7195 ( .A(n6162), .B(n6163), .Z(n1038) );
  ANDN U7196 ( .A(n4110), .B(n4050), .Z(\modmult_1/N1019 ) );
  XOR U7197 ( .A(n6160), .B(n6161), .Z(n4050) );
  NAND U7198 ( .A(n6164), .B(nreg[1016]), .Z(n6161) );
  NAND U7199 ( .A(n6107), .B(nreg[1016]), .Z(n6164) );
  XOR U7200 ( .A(n6165), .B(n6166), .Z(n6160) );
  IV U7201 ( .A(n6157), .Z(n6165) );
  XOR U7202 ( .A(n6167), .B(n6168), .Z(n6157) );
  ANDN U7203 ( .A(n6169), .B(n6170), .Z(n6168) );
  XNOR U7204 ( .A(n6171), .B(n6167), .Z(n6169) );
  ANDN U7205 ( .A(n4110), .B(n4053), .Z(\modmult_1/N1018 ) );
  XOR U7206 ( .A(n6170), .B(n6171), .Z(n4053) );
  NAND U7207 ( .A(n6172), .B(nreg[1015]), .Z(n6171) );
  NAND U7208 ( .A(n6107), .B(nreg[1015]), .Z(n6172) );
  XOR U7209 ( .A(n6173), .B(n6174), .Z(n6170) );
  IV U7210 ( .A(n6167), .Z(n6173) );
  XOR U7211 ( .A(n6175), .B(n6176), .Z(n6167) );
  ANDN U7212 ( .A(n6177), .B(n6178), .Z(n6176) );
  XNOR U7213 ( .A(n6179), .B(n6175), .Z(n6177) );
  ANDN U7214 ( .A(n4110), .B(n4056), .Z(\modmult_1/N1017 ) );
  XOR U7215 ( .A(n6178), .B(n6179), .Z(n4056) );
  NAND U7216 ( .A(n6180), .B(nreg[1014]), .Z(n6179) );
  NAND U7217 ( .A(n6107), .B(nreg[1014]), .Z(n6180) );
  XOR U7218 ( .A(n6181), .B(n6182), .Z(n6178) );
  IV U7219 ( .A(n6175), .Z(n6181) );
  XOR U7220 ( .A(n6183), .B(n6184), .Z(n6175) );
  ANDN U7221 ( .A(n6185), .B(n6186), .Z(n6184) );
  XNOR U7222 ( .A(n6187), .B(n6183), .Z(n6185) );
  ANDN U7223 ( .A(n4110), .B(n4059), .Z(\modmult_1/N1016 ) );
  XOR U7224 ( .A(n6186), .B(n6187), .Z(n4059) );
  NAND U7225 ( .A(n6188), .B(nreg[1013]), .Z(n6187) );
  NAND U7226 ( .A(n6107), .B(nreg[1013]), .Z(n6188) );
  XOR U7227 ( .A(n6189), .B(n6190), .Z(n6186) );
  IV U7228 ( .A(n6183), .Z(n6189) );
  XOR U7229 ( .A(n6191), .B(n6192), .Z(n6183) );
  ANDN U7230 ( .A(n6193), .B(n6194), .Z(n6192) );
  XNOR U7231 ( .A(n6195), .B(n6191), .Z(n6193) );
  ANDN U7232 ( .A(n4110), .B(n4062), .Z(\modmult_1/N1015 ) );
  XOR U7233 ( .A(n6194), .B(n6195), .Z(n4062) );
  NAND U7234 ( .A(n6196), .B(nreg[1012]), .Z(n6195) );
  NAND U7235 ( .A(n6107), .B(nreg[1012]), .Z(n6196) );
  XOR U7236 ( .A(n6197), .B(n6198), .Z(n6194) );
  IV U7237 ( .A(n6191), .Z(n6197) );
  XOR U7238 ( .A(n6199), .B(n6200), .Z(n6191) );
  ANDN U7239 ( .A(n6201), .B(n6202), .Z(n6200) );
  XNOR U7240 ( .A(n6203), .B(n6199), .Z(n6201) );
  ANDN U7241 ( .A(n4110), .B(n4065), .Z(\modmult_1/N1014 ) );
  XOR U7242 ( .A(n6202), .B(n6203), .Z(n4065) );
  NAND U7243 ( .A(n6204), .B(nreg[1011]), .Z(n6203) );
  NAND U7244 ( .A(n6107), .B(nreg[1011]), .Z(n6204) );
  XOR U7245 ( .A(n6205), .B(n6206), .Z(n6202) );
  IV U7246 ( .A(n6199), .Z(n6205) );
  XOR U7247 ( .A(n6207), .B(n6208), .Z(n6199) );
  ANDN U7248 ( .A(n6209), .B(n6210), .Z(n6208) );
  XNOR U7249 ( .A(n6211), .B(n6207), .Z(n6209) );
  ANDN U7250 ( .A(n4110), .B(n4068), .Z(\modmult_1/N1013 ) );
  XOR U7251 ( .A(n6210), .B(n6211), .Z(n4068) );
  NAND U7252 ( .A(n6212), .B(nreg[1010]), .Z(n6211) );
  NAND U7253 ( .A(n6107), .B(nreg[1010]), .Z(n6212) );
  XOR U7254 ( .A(n6213), .B(n6214), .Z(n6210) );
  IV U7255 ( .A(n6207), .Z(n6213) );
  XOR U7256 ( .A(n6215), .B(n6216), .Z(n6207) );
  ANDN U7257 ( .A(n6217), .B(n6218), .Z(n6216) );
  XNOR U7258 ( .A(n6219), .B(n6215), .Z(n6217) );
  ANDN U7259 ( .A(n4110), .B(n4074), .Z(\modmult_1/N1012 ) );
  XOR U7260 ( .A(n6218), .B(n6219), .Z(n4074) );
  NAND U7261 ( .A(n6220), .B(nreg[1009]), .Z(n6219) );
  NAND U7262 ( .A(n6107), .B(nreg[1009]), .Z(n6220) );
  XOR U7263 ( .A(n6221), .B(n6222), .Z(n6218) );
  IV U7264 ( .A(n6215), .Z(n6221) );
  XOR U7265 ( .A(n6223), .B(n6224), .Z(n6215) );
  ANDN U7266 ( .A(n6225), .B(n6226), .Z(n6224) );
  XNOR U7267 ( .A(n6227), .B(n6223), .Z(n6225) );
  ANDN U7268 ( .A(n4110), .B(n4077), .Z(\modmult_1/N1011 ) );
  XOR U7269 ( .A(n6226), .B(n6227), .Z(n4077) );
  NAND U7270 ( .A(n6228), .B(nreg[1008]), .Z(n6227) );
  NAND U7271 ( .A(n6107), .B(nreg[1008]), .Z(n6228) );
  XOR U7272 ( .A(n6229), .B(n6230), .Z(n6226) );
  IV U7273 ( .A(n6223), .Z(n6229) );
  XOR U7274 ( .A(n6231), .B(n6232), .Z(n6223) );
  ANDN U7275 ( .A(n6233), .B(n6234), .Z(n6232) );
  XNOR U7276 ( .A(n6235), .B(n6231), .Z(n6233) );
  ANDN U7277 ( .A(n4110), .B(n4080), .Z(\modmult_1/N1010 ) );
  XOR U7278 ( .A(n6234), .B(n6235), .Z(n4080) );
  NAND U7279 ( .A(n6236), .B(nreg[1007]), .Z(n6235) );
  NAND U7280 ( .A(n6107), .B(nreg[1007]), .Z(n6236) );
  XOR U7281 ( .A(n6237), .B(n6238), .Z(n6234) );
  IV U7282 ( .A(n6231), .Z(n6237) );
  XOR U7283 ( .A(n6239), .B(n6240), .Z(n6231) );
  ANDN U7284 ( .A(n6241), .B(n6242), .Z(n6240) );
  XNOR U7285 ( .A(n6243), .B(n6239), .Z(n6241) );
  ANDN U7286 ( .A(n4110), .B(n1071), .Z(\modmult_1/N101 ) );
  XOR U7287 ( .A(n6244), .B(n6245), .Z(n1071) );
  ANDN U7288 ( .A(n4110), .B(n4083), .Z(\modmult_1/N1009 ) );
  XOR U7289 ( .A(n6242), .B(n6243), .Z(n4083) );
  NAND U7290 ( .A(n6246), .B(nreg[1006]), .Z(n6243) );
  NAND U7291 ( .A(n6107), .B(nreg[1006]), .Z(n6246) );
  XOR U7292 ( .A(n6247), .B(n6248), .Z(n6242) );
  IV U7293 ( .A(n6239), .Z(n6247) );
  XOR U7294 ( .A(n6249), .B(n6250), .Z(n6239) );
  ANDN U7295 ( .A(n6251), .B(n6252), .Z(n6250) );
  XNOR U7296 ( .A(n6253), .B(n6249), .Z(n6251) );
  ANDN U7297 ( .A(n4110), .B(n4086), .Z(\modmult_1/N1008 ) );
  XOR U7298 ( .A(n6252), .B(n6253), .Z(n4086) );
  NAND U7299 ( .A(n6254), .B(nreg[1005]), .Z(n6253) );
  NAND U7300 ( .A(n6107), .B(nreg[1005]), .Z(n6254) );
  XOR U7301 ( .A(n6255), .B(n6256), .Z(n6252) );
  IV U7302 ( .A(n6249), .Z(n6255) );
  XOR U7303 ( .A(n6257), .B(n6258), .Z(n6249) );
  ANDN U7304 ( .A(n6259), .B(n6260), .Z(n6258) );
  XNOR U7305 ( .A(n6261), .B(n6257), .Z(n6259) );
  ANDN U7306 ( .A(n4110), .B(n4089), .Z(\modmult_1/N1007 ) );
  XOR U7307 ( .A(n6260), .B(n6261), .Z(n4089) );
  NAND U7308 ( .A(n6262), .B(nreg[1004]), .Z(n6261) );
  NAND U7309 ( .A(n6107), .B(nreg[1004]), .Z(n6262) );
  XOR U7310 ( .A(n6263), .B(n6264), .Z(n6260) );
  IV U7311 ( .A(n6257), .Z(n6263) );
  XOR U7312 ( .A(n6265), .B(n6266), .Z(n6257) );
  ANDN U7313 ( .A(n6267), .B(n6268), .Z(n6266) );
  XNOR U7314 ( .A(n6269), .B(n6265), .Z(n6267) );
  ANDN U7315 ( .A(n4110), .B(n4092), .Z(\modmult_1/N1006 ) );
  XOR U7316 ( .A(n6268), .B(n6269), .Z(n4092) );
  NAND U7317 ( .A(n6270), .B(nreg[1003]), .Z(n6269) );
  NAND U7318 ( .A(n6107), .B(nreg[1003]), .Z(n6270) );
  XOR U7319 ( .A(n6271), .B(n6272), .Z(n6268) );
  IV U7320 ( .A(n6265), .Z(n6271) );
  XOR U7321 ( .A(n6273), .B(n6274), .Z(n6265) );
  ANDN U7322 ( .A(n6275), .B(n6276), .Z(n6274) );
  XNOR U7323 ( .A(n6277), .B(n6273), .Z(n6275) );
  ANDN U7324 ( .A(n4110), .B(n4095), .Z(\modmult_1/N1005 ) );
  XOR U7325 ( .A(n6276), .B(n6277), .Z(n4095) );
  NAND U7326 ( .A(n6278), .B(nreg[1002]), .Z(n6277) );
  NAND U7327 ( .A(n6107), .B(nreg[1002]), .Z(n6278) );
  XOR U7328 ( .A(n6279), .B(n6280), .Z(n6276) );
  IV U7329 ( .A(n6273), .Z(n6279) );
  XOR U7330 ( .A(n6281), .B(n6282), .Z(n6273) );
  ANDN U7331 ( .A(n6283), .B(n6284), .Z(n6282) );
  XNOR U7332 ( .A(n6285), .B(n6281), .Z(n6283) );
  ANDN U7333 ( .A(n4110), .B(n4098), .Z(\modmult_1/N1004 ) );
  XOR U7334 ( .A(n6284), .B(n6285), .Z(n4098) );
  NAND U7335 ( .A(n6286), .B(nreg[1001]), .Z(n6285) );
  NAND U7336 ( .A(n6107), .B(nreg[1001]), .Z(n6286) );
  XOR U7337 ( .A(n6287), .B(n6288), .Z(n6284) );
  IV U7338 ( .A(n6281), .Z(n6287) );
  XOR U7339 ( .A(n6289), .B(n6290), .Z(n6281) );
  ANDN U7340 ( .A(n6291), .B(n6292), .Z(n6290) );
  XNOR U7341 ( .A(n6293), .B(n6289), .Z(n6291) );
  ANDN U7342 ( .A(n4110), .B(n4101), .Z(\modmult_1/N1003 ) );
  XOR U7343 ( .A(n6292), .B(n6293), .Z(n4101) );
  NAND U7344 ( .A(n6294), .B(nreg[1000]), .Z(n6293) );
  NAND U7345 ( .A(n6107), .B(nreg[1000]), .Z(n6294) );
  XOR U7346 ( .A(n6295), .B(n6296), .Z(n6292) );
  IV U7347 ( .A(n6289), .Z(n6295) );
  XOR U7348 ( .A(n6297), .B(n6298), .Z(n6289) );
  ANDN U7349 ( .A(n6299), .B(n6300), .Z(n6298) );
  XNOR U7350 ( .A(n6301), .B(n6297), .Z(n6299) );
  ANDN U7351 ( .A(n4110), .B(n1041), .Z(\modmult_1/N1002 ) );
  XOR U7352 ( .A(n6300), .B(n6301), .Z(n1041) );
  NAND U7353 ( .A(n6302), .B(nreg[999]), .Z(n6301) );
  NAND U7354 ( .A(n6107), .B(nreg[999]), .Z(n6302) );
  XOR U7355 ( .A(n6303), .B(n6304), .Z(n6300) );
  IV U7356 ( .A(n6297), .Z(n6303) );
  XOR U7357 ( .A(n6305), .B(n6306), .Z(n6297) );
  ANDN U7358 ( .A(n6307), .B(n6308), .Z(n6306) );
  XNOR U7359 ( .A(n6309), .B(n6305), .Z(n6307) );
  ANDN U7360 ( .A(n4110), .B(n1044), .Z(\modmult_1/N1001 ) );
  XOR U7361 ( .A(n6308), .B(n6309), .Z(n1044) );
  NAND U7362 ( .A(n6310), .B(nreg[998]), .Z(n6309) );
  NAND U7363 ( .A(n6107), .B(nreg[998]), .Z(n6310) );
  XOR U7364 ( .A(n6311), .B(n6312), .Z(n6308) );
  IV U7365 ( .A(n6305), .Z(n6311) );
  XOR U7366 ( .A(n6313), .B(n6314), .Z(n6305) );
  ANDN U7367 ( .A(n6315), .B(n6316), .Z(n6314) );
  XNOR U7368 ( .A(n6317), .B(n6313), .Z(n6315) );
  ANDN U7369 ( .A(n4110), .B(n1047), .Z(\modmult_1/N1000 ) );
  XOR U7370 ( .A(n6316), .B(n6317), .Z(n1047) );
  NAND U7371 ( .A(n6318), .B(nreg[997]), .Z(n6317) );
  NAND U7372 ( .A(n6107), .B(nreg[997]), .Z(n6318) );
  XOR U7373 ( .A(n6319), .B(n6320), .Z(n6316) );
  IV U7374 ( .A(n6313), .Z(n6319) );
  XOR U7375 ( .A(n6321), .B(n6322), .Z(n6313) );
  ANDN U7376 ( .A(n6323), .B(n4111), .Z(n6322) );
  XOR U7377 ( .A(n6324), .B(n6325), .Z(n4111) );
  IV U7378 ( .A(n6321), .Z(n6324) );
  XNOR U7379 ( .A(n4112), .B(n6321), .Z(n6323) );
  NAND U7380 ( .A(n6326), .B(nreg[996]), .Z(n4112) );
  NAND U7381 ( .A(n6107), .B(nreg[996]), .Z(n6326) );
  XOR U7382 ( .A(n6327), .B(n6328), .Z(n6321) );
  ANDN U7383 ( .A(n6329), .B(n4113), .Z(n6328) );
  XOR U7384 ( .A(n6330), .B(n6331), .Z(n4113) );
  IV U7385 ( .A(n6327), .Z(n6330) );
  XNOR U7386 ( .A(n4114), .B(n6327), .Z(n6329) );
  NAND U7387 ( .A(n6332), .B(nreg[995]), .Z(n4114) );
  NAND U7388 ( .A(n6107), .B(nreg[995]), .Z(n6332) );
  XOR U7389 ( .A(n6333), .B(n6334), .Z(n6327) );
  ANDN U7390 ( .A(n6335), .B(n4115), .Z(n6334) );
  XOR U7391 ( .A(n6336), .B(n6337), .Z(n4115) );
  IV U7392 ( .A(n6333), .Z(n6336) );
  XNOR U7393 ( .A(n4116), .B(n6333), .Z(n6335) );
  NAND U7394 ( .A(n6338), .B(nreg[994]), .Z(n4116) );
  NAND U7395 ( .A(n6107), .B(nreg[994]), .Z(n6338) );
  XOR U7396 ( .A(n6339), .B(n6340), .Z(n6333) );
  ANDN U7397 ( .A(n6341), .B(n4117), .Z(n6340) );
  XOR U7398 ( .A(n6342), .B(n6343), .Z(n4117) );
  IV U7399 ( .A(n6339), .Z(n6342) );
  XNOR U7400 ( .A(n4118), .B(n6339), .Z(n6341) );
  NAND U7401 ( .A(n6344), .B(nreg[993]), .Z(n4118) );
  NAND U7402 ( .A(n6107), .B(nreg[993]), .Z(n6344) );
  XOR U7403 ( .A(n6345), .B(n6346), .Z(n6339) );
  ANDN U7404 ( .A(n6347), .B(n4119), .Z(n6346) );
  XOR U7405 ( .A(n6348), .B(n6349), .Z(n4119) );
  IV U7406 ( .A(n6345), .Z(n6348) );
  XNOR U7407 ( .A(n4120), .B(n6345), .Z(n6347) );
  NAND U7408 ( .A(n6350), .B(nreg[992]), .Z(n4120) );
  NAND U7409 ( .A(n6107), .B(nreg[992]), .Z(n6350) );
  XOR U7410 ( .A(n6351), .B(n6352), .Z(n6345) );
  ANDN U7411 ( .A(n6353), .B(n4121), .Z(n6352) );
  XOR U7412 ( .A(n6354), .B(n6355), .Z(n4121) );
  IV U7413 ( .A(n6351), .Z(n6354) );
  XNOR U7414 ( .A(n4122), .B(n6351), .Z(n6353) );
  NAND U7415 ( .A(n6356), .B(nreg[991]), .Z(n4122) );
  NAND U7416 ( .A(n6107), .B(nreg[991]), .Z(n6356) );
  XOR U7417 ( .A(n6357), .B(n6358), .Z(n6351) );
  ANDN U7418 ( .A(n6359), .B(n4123), .Z(n6358) );
  XOR U7419 ( .A(n6360), .B(n6361), .Z(n4123) );
  IV U7420 ( .A(n6357), .Z(n6360) );
  XNOR U7421 ( .A(n4124), .B(n6357), .Z(n6359) );
  NAND U7422 ( .A(n6362), .B(nreg[990]), .Z(n4124) );
  NAND U7423 ( .A(n6107), .B(nreg[990]), .Z(n6362) );
  XOR U7424 ( .A(n6363), .B(n6364), .Z(n6357) );
  ANDN U7425 ( .A(n6365), .B(n4125), .Z(n6364) );
  XOR U7426 ( .A(n6366), .B(n6367), .Z(n4125) );
  IV U7427 ( .A(n6363), .Z(n6366) );
  XNOR U7428 ( .A(n4126), .B(n6363), .Z(n6365) );
  NAND U7429 ( .A(n6368), .B(nreg[989]), .Z(n4126) );
  NAND U7430 ( .A(n6107), .B(nreg[989]), .Z(n6368) );
  XOR U7431 ( .A(n6369), .B(n6370), .Z(n6363) );
  ANDN U7432 ( .A(n6371), .B(n4127), .Z(n6370) );
  XOR U7433 ( .A(n6372), .B(n6373), .Z(n4127) );
  IV U7434 ( .A(n6369), .Z(n6372) );
  XNOR U7435 ( .A(n4128), .B(n6369), .Z(n6371) );
  NAND U7436 ( .A(n6374), .B(nreg[988]), .Z(n4128) );
  NAND U7437 ( .A(n6107), .B(nreg[988]), .Z(n6374) );
  XOR U7438 ( .A(n6375), .B(n6376), .Z(n6369) );
  ANDN U7439 ( .A(n6377), .B(n4129), .Z(n6376) );
  XOR U7440 ( .A(n6378), .B(n6379), .Z(n4129) );
  IV U7441 ( .A(n6375), .Z(n6378) );
  XNOR U7442 ( .A(n4130), .B(n6375), .Z(n6377) );
  NAND U7443 ( .A(n6380), .B(nreg[987]), .Z(n4130) );
  NAND U7444 ( .A(n6107), .B(nreg[987]), .Z(n6380) );
  XOR U7445 ( .A(n6381), .B(n6382), .Z(n6375) );
  ANDN U7446 ( .A(n6383), .B(n4133), .Z(n6382) );
  XOR U7447 ( .A(n6384), .B(n6385), .Z(n4133) );
  IV U7448 ( .A(n6381), .Z(n6384) );
  XNOR U7449 ( .A(n4134), .B(n6381), .Z(n6383) );
  NAND U7450 ( .A(n6386), .B(nreg[986]), .Z(n4134) );
  NAND U7451 ( .A(n6107), .B(nreg[986]), .Z(n6386) );
  XOR U7452 ( .A(n6387), .B(n6388), .Z(n6381) );
  ANDN U7453 ( .A(n6389), .B(n4135), .Z(n6388) );
  XOR U7454 ( .A(n6390), .B(n6391), .Z(n4135) );
  IV U7455 ( .A(n6387), .Z(n6390) );
  XNOR U7456 ( .A(n4136), .B(n6387), .Z(n6389) );
  NAND U7457 ( .A(n6392), .B(nreg[985]), .Z(n4136) );
  NAND U7458 ( .A(n6107), .B(nreg[985]), .Z(n6392) );
  XOR U7459 ( .A(n6393), .B(n6394), .Z(n6387) );
  ANDN U7460 ( .A(n6395), .B(n4137), .Z(n6394) );
  XOR U7461 ( .A(n6396), .B(n6397), .Z(n4137) );
  IV U7462 ( .A(n6393), .Z(n6396) );
  XNOR U7463 ( .A(n4138), .B(n6393), .Z(n6395) );
  NAND U7464 ( .A(n6398), .B(nreg[984]), .Z(n4138) );
  NAND U7465 ( .A(n6107), .B(nreg[984]), .Z(n6398) );
  XOR U7466 ( .A(n6399), .B(n6400), .Z(n6393) );
  ANDN U7467 ( .A(n6401), .B(n4139), .Z(n6400) );
  XOR U7468 ( .A(n6402), .B(n6403), .Z(n4139) );
  IV U7469 ( .A(n6399), .Z(n6402) );
  XNOR U7470 ( .A(n4140), .B(n6399), .Z(n6401) );
  NAND U7471 ( .A(n6404), .B(nreg[983]), .Z(n4140) );
  NAND U7472 ( .A(n6107), .B(nreg[983]), .Z(n6404) );
  XOR U7473 ( .A(n6405), .B(n6406), .Z(n6399) );
  ANDN U7474 ( .A(n6407), .B(n4141), .Z(n6406) );
  XOR U7475 ( .A(n6408), .B(n6409), .Z(n4141) );
  IV U7476 ( .A(n6405), .Z(n6408) );
  XNOR U7477 ( .A(n4142), .B(n6405), .Z(n6407) );
  NAND U7478 ( .A(n6410), .B(nreg[982]), .Z(n4142) );
  NAND U7479 ( .A(n6107), .B(nreg[982]), .Z(n6410) );
  XOR U7480 ( .A(n6411), .B(n6412), .Z(n6405) );
  ANDN U7481 ( .A(n6413), .B(n4143), .Z(n6412) );
  XOR U7482 ( .A(n6414), .B(n6415), .Z(n4143) );
  IV U7483 ( .A(n6411), .Z(n6414) );
  XNOR U7484 ( .A(n4144), .B(n6411), .Z(n6413) );
  NAND U7485 ( .A(n6416), .B(nreg[981]), .Z(n4144) );
  NAND U7486 ( .A(n6107), .B(nreg[981]), .Z(n6416) );
  XOR U7487 ( .A(n6417), .B(n6418), .Z(n6411) );
  ANDN U7488 ( .A(n6419), .B(n4145), .Z(n6418) );
  XOR U7489 ( .A(n6420), .B(n6421), .Z(n4145) );
  IV U7490 ( .A(n6417), .Z(n6420) );
  XNOR U7491 ( .A(n4146), .B(n6417), .Z(n6419) );
  NAND U7492 ( .A(n6422), .B(nreg[980]), .Z(n4146) );
  NAND U7493 ( .A(n6107), .B(nreg[980]), .Z(n6422) );
  XOR U7494 ( .A(n6423), .B(n6424), .Z(n6417) );
  ANDN U7495 ( .A(n6425), .B(n4147), .Z(n6424) );
  XOR U7496 ( .A(n6426), .B(n6427), .Z(n4147) );
  IV U7497 ( .A(n6423), .Z(n6426) );
  XNOR U7498 ( .A(n4148), .B(n6423), .Z(n6425) );
  NAND U7499 ( .A(n6428), .B(nreg[979]), .Z(n4148) );
  NAND U7500 ( .A(n6107), .B(nreg[979]), .Z(n6428) );
  XOR U7501 ( .A(n6429), .B(n6430), .Z(n6423) );
  ANDN U7502 ( .A(n6431), .B(n4149), .Z(n6430) );
  XOR U7503 ( .A(n6432), .B(n6433), .Z(n4149) );
  IV U7504 ( .A(n6429), .Z(n6432) );
  XNOR U7505 ( .A(n4150), .B(n6429), .Z(n6431) );
  NAND U7506 ( .A(n6434), .B(nreg[978]), .Z(n4150) );
  NAND U7507 ( .A(n6107), .B(nreg[978]), .Z(n6434) );
  XOR U7508 ( .A(n6435), .B(n6436), .Z(n6429) );
  ANDN U7509 ( .A(n6437), .B(n4151), .Z(n6436) );
  XOR U7510 ( .A(n6438), .B(n6439), .Z(n4151) );
  IV U7511 ( .A(n6435), .Z(n6438) );
  XNOR U7512 ( .A(n4152), .B(n6435), .Z(n6437) );
  NAND U7513 ( .A(n6440), .B(nreg[977]), .Z(n4152) );
  NAND U7514 ( .A(n6107), .B(nreg[977]), .Z(n6440) );
  XOR U7515 ( .A(n6441), .B(n6442), .Z(n6435) );
  ANDN U7516 ( .A(n6443), .B(n4155), .Z(n6442) );
  XOR U7517 ( .A(n6444), .B(n6445), .Z(n4155) );
  IV U7518 ( .A(n6441), .Z(n6444) );
  XNOR U7519 ( .A(n4156), .B(n6441), .Z(n6443) );
  NAND U7520 ( .A(n6446), .B(nreg[976]), .Z(n4156) );
  NAND U7521 ( .A(n6107), .B(nreg[976]), .Z(n6446) );
  XOR U7522 ( .A(n6447), .B(n6448), .Z(n6441) );
  ANDN U7523 ( .A(n6449), .B(n4157), .Z(n6448) );
  XOR U7524 ( .A(n6450), .B(n6451), .Z(n4157) );
  IV U7525 ( .A(n6447), .Z(n6450) );
  XNOR U7526 ( .A(n4158), .B(n6447), .Z(n6449) );
  NAND U7527 ( .A(n6452), .B(nreg[975]), .Z(n4158) );
  NAND U7528 ( .A(n6107), .B(nreg[975]), .Z(n6452) );
  XOR U7529 ( .A(n6453), .B(n6454), .Z(n6447) );
  ANDN U7530 ( .A(n6455), .B(n4159), .Z(n6454) );
  XOR U7531 ( .A(n6456), .B(n6457), .Z(n4159) );
  IV U7532 ( .A(n6453), .Z(n6456) );
  XNOR U7533 ( .A(n4160), .B(n6453), .Z(n6455) );
  NAND U7534 ( .A(n6458), .B(nreg[974]), .Z(n4160) );
  NAND U7535 ( .A(n6107), .B(nreg[974]), .Z(n6458) );
  XOR U7536 ( .A(n6459), .B(n6460), .Z(n6453) );
  ANDN U7537 ( .A(n6461), .B(n4161), .Z(n6460) );
  XOR U7538 ( .A(n6462), .B(n6463), .Z(n4161) );
  IV U7539 ( .A(n6459), .Z(n6462) );
  XNOR U7540 ( .A(n4162), .B(n6459), .Z(n6461) );
  NAND U7541 ( .A(n6464), .B(nreg[973]), .Z(n4162) );
  NAND U7542 ( .A(n6107), .B(nreg[973]), .Z(n6464) );
  XOR U7543 ( .A(n6465), .B(n6466), .Z(n6459) );
  ANDN U7544 ( .A(n6467), .B(n4163), .Z(n6466) );
  XOR U7545 ( .A(n6468), .B(n6469), .Z(n4163) );
  IV U7546 ( .A(n6465), .Z(n6468) );
  XNOR U7547 ( .A(n4164), .B(n6465), .Z(n6467) );
  NAND U7548 ( .A(n6470), .B(nreg[972]), .Z(n4164) );
  NAND U7549 ( .A(n6107), .B(nreg[972]), .Z(n6470) );
  XOR U7550 ( .A(n6471), .B(n6472), .Z(n6465) );
  ANDN U7551 ( .A(n6473), .B(n4165), .Z(n6472) );
  XOR U7552 ( .A(n6474), .B(n6475), .Z(n4165) );
  IV U7553 ( .A(n6471), .Z(n6474) );
  XNOR U7554 ( .A(n4166), .B(n6471), .Z(n6473) );
  NAND U7555 ( .A(n6476), .B(nreg[971]), .Z(n4166) );
  NAND U7556 ( .A(n6107), .B(nreg[971]), .Z(n6476) );
  XOR U7557 ( .A(n6477), .B(n6478), .Z(n6471) );
  ANDN U7558 ( .A(n6479), .B(n4167), .Z(n6478) );
  XOR U7559 ( .A(n6480), .B(n6481), .Z(n4167) );
  IV U7560 ( .A(n6477), .Z(n6480) );
  XNOR U7561 ( .A(n4168), .B(n6477), .Z(n6479) );
  NAND U7562 ( .A(n6482), .B(nreg[970]), .Z(n4168) );
  NAND U7563 ( .A(n6107), .B(nreg[970]), .Z(n6482) );
  XOR U7564 ( .A(n6483), .B(n6484), .Z(n6477) );
  ANDN U7565 ( .A(n6485), .B(n4169), .Z(n6484) );
  XOR U7566 ( .A(n6486), .B(n6487), .Z(n4169) );
  IV U7567 ( .A(n6483), .Z(n6486) );
  XNOR U7568 ( .A(n4170), .B(n6483), .Z(n6485) );
  NAND U7569 ( .A(n6488), .B(nreg[969]), .Z(n4170) );
  NAND U7570 ( .A(n6107), .B(nreg[969]), .Z(n6488) );
  XOR U7571 ( .A(n6489), .B(n6490), .Z(n6483) );
  ANDN U7572 ( .A(n6491), .B(n4171), .Z(n6490) );
  XOR U7573 ( .A(n6492), .B(n6493), .Z(n4171) );
  IV U7574 ( .A(n6489), .Z(n6492) );
  XNOR U7575 ( .A(n4172), .B(n6489), .Z(n6491) );
  NAND U7576 ( .A(n6494), .B(nreg[968]), .Z(n4172) );
  NAND U7577 ( .A(n6107), .B(nreg[968]), .Z(n6494) );
  XOR U7578 ( .A(n6495), .B(n6496), .Z(n6489) );
  ANDN U7579 ( .A(n6497), .B(n4173), .Z(n6496) );
  XOR U7580 ( .A(n6498), .B(n6499), .Z(n4173) );
  IV U7581 ( .A(n6495), .Z(n6498) );
  XNOR U7582 ( .A(n4174), .B(n6495), .Z(n6497) );
  NAND U7583 ( .A(n6500), .B(nreg[967]), .Z(n4174) );
  NAND U7584 ( .A(n6107), .B(nreg[967]), .Z(n6500) );
  XOR U7585 ( .A(n6501), .B(n6502), .Z(n6495) );
  ANDN U7586 ( .A(n6503), .B(n4177), .Z(n6502) );
  XOR U7587 ( .A(n6504), .B(n6505), .Z(n4177) );
  IV U7588 ( .A(n6501), .Z(n6504) );
  XNOR U7589 ( .A(n4178), .B(n6501), .Z(n6503) );
  NAND U7590 ( .A(n6506), .B(nreg[966]), .Z(n4178) );
  NAND U7591 ( .A(n6107), .B(nreg[966]), .Z(n6506) );
  XOR U7592 ( .A(n6507), .B(n6508), .Z(n6501) );
  ANDN U7593 ( .A(n6509), .B(n4179), .Z(n6508) );
  XOR U7594 ( .A(n6510), .B(n6511), .Z(n4179) );
  IV U7595 ( .A(n6507), .Z(n6510) );
  XNOR U7596 ( .A(n4180), .B(n6507), .Z(n6509) );
  NAND U7597 ( .A(n6512), .B(nreg[965]), .Z(n4180) );
  NAND U7598 ( .A(n6107), .B(nreg[965]), .Z(n6512) );
  XOR U7599 ( .A(n6513), .B(n6514), .Z(n6507) );
  ANDN U7600 ( .A(n6515), .B(n4181), .Z(n6514) );
  XOR U7601 ( .A(n6516), .B(n6517), .Z(n4181) );
  IV U7602 ( .A(n6513), .Z(n6516) );
  XNOR U7603 ( .A(n4182), .B(n6513), .Z(n6515) );
  NAND U7604 ( .A(n6518), .B(nreg[964]), .Z(n4182) );
  NAND U7605 ( .A(n6107), .B(nreg[964]), .Z(n6518) );
  XOR U7606 ( .A(n6519), .B(n6520), .Z(n6513) );
  ANDN U7607 ( .A(n6521), .B(n4183), .Z(n6520) );
  XOR U7608 ( .A(n6522), .B(n6523), .Z(n4183) );
  IV U7609 ( .A(n6519), .Z(n6522) );
  XNOR U7610 ( .A(n4184), .B(n6519), .Z(n6521) );
  NAND U7611 ( .A(n6524), .B(nreg[963]), .Z(n4184) );
  NAND U7612 ( .A(n6107), .B(nreg[963]), .Z(n6524) );
  XOR U7613 ( .A(n6525), .B(n6526), .Z(n6519) );
  ANDN U7614 ( .A(n6527), .B(n4185), .Z(n6526) );
  XOR U7615 ( .A(n6528), .B(n6529), .Z(n4185) );
  IV U7616 ( .A(n6525), .Z(n6528) );
  XNOR U7617 ( .A(n4186), .B(n6525), .Z(n6527) );
  NAND U7618 ( .A(n6530), .B(nreg[962]), .Z(n4186) );
  NAND U7619 ( .A(n6107), .B(nreg[962]), .Z(n6530) );
  XOR U7620 ( .A(n6531), .B(n6532), .Z(n6525) );
  ANDN U7621 ( .A(n6533), .B(n4187), .Z(n6532) );
  XOR U7622 ( .A(n6534), .B(n6535), .Z(n4187) );
  IV U7623 ( .A(n6531), .Z(n6534) );
  XNOR U7624 ( .A(n4188), .B(n6531), .Z(n6533) );
  NAND U7625 ( .A(n6536), .B(nreg[961]), .Z(n4188) );
  NAND U7626 ( .A(n6107), .B(nreg[961]), .Z(n6536) );
  XOR U7627 ( .A(n6537), .B(n6538), .Z(n6531) );
  ANDN U7628 ( .A(n6539), .B(n4189), .Z(n6538) );
  XOR U7629 ( .A(n6540), .B(n6541), .Z(n4189) );
  IV U7630 ( .A(n6537), .Z(n6540) );
  XNOR U7631 ( .A(n4190), .B(n6537), .Z(n6539) );
  NAND U7632 ( .A(n6542), .B(nreg[960]), .Z(n4190) );
  NAND U7633 ( .A(n6107), .B(nreg[960]), .Z(n6542) );
  XOR U7634 ( .A(n6543), .B(n6544), .Z(n6537) );
  ANDN U7635 ( .A(n6545), .B(n4191), .Z(n6544) );
  XOR U7636 ( .A(n6546), .B(n6547), .Z(n4191) );
  IV U7637 ( .A(n6543), .Z(n6546) );
  XNOR U7638 ( .A(n4192), .B(n6543), .Z(n6545) );
  NAND U7639 ( .A(n6548), .B(nreg[959]), .Z(n4192) );
  NAND U7640 ( .A(n6107), .B(nreg[959]), .Z(n6548) );
  XOR U7641 ( .A(n6549), .B(n6550), .Z(n6543) );
  ANDN U7642 ( .A(n6551), .B(n4193), .Z(n6550) );
  XOR U7643 ( .A(n6552), .B(n6553), .Z(n4193) );
  IV U7644 ( .A(n6549), .Z(n6552) );
  XNOR U7645 ( .A(n4194), .B(n6549), .Z(n6551) );
  NAND U7646 ( .A(n6554), .B(nreg[958]), .Z(n4194) );
  NAND U7647 ( .A(n6107), .B(nreg[958]), .Z(n6554) );
  XOR U7648 ( .A(n6555), .B(n6556), .Z(n6549) );
  ANDN U7649 ( .A(n6557), .B(n4195), .Z(n6556) );
  XOR U7650 ( .A(n6558), .B(n6559), .Z(n4195) );
  IV U7651 ( .A(n6555), .Z(n6558) );
  XNOR U7652 ( .A(n4196), .B(n6555), .Z(n6557) );
  NAND U7653 ( .A(n6560), .B(nreg[957]), .Z(n4196) );
  NAND U7654 ( .A(n6107), .B(nreg[957]), .Z(n6560) );
  XOR U7655 ( .A(n6561), .B(n6562), .Z(n6555) );
  ANDN U7656 ( .A(n6563), .B(n4199), .Z(n6562) );
  XOR U7657 ( .A(n6564), .B(n6565), .Z(n4199) );
  IV U7658 ( .A(n6561), .Z(n6564) );
  XNOR U7659 ( .A(n4200), .B(n6561), .Z(n6563) );
  NAND U7660 ( .A(n6566), .B(nreg[956]), .Z(n4200) );
  NAND U7661 ( .A(n6107), .B(nreg[956]), .Z(n6566) );
  XOR U7662 ( .A(n6567), .B(n6568), .Z(n6561) );
  ANDN U7663 ( .A(n6569), .B(n4201), .Z(n6568) );
  XOR U7664 ( .A(n6570), .B(n6571), .Z(n4201) );
  IV U7665 ( .A(n6567), .Z(n6570) );
  XNOR U7666 ( .A(n4202), .B(n6567), .Z(n6569) );
  NAND U7667 ( .A(n6572), .B(nreg[955]), .Z(n4202) );
  NAND U7668 ( .A(n6107), .B(nreg[955]), .Z(n6572) );
  XOR U7669 ( .A(n6573), .B(n6574), .Z(n6567) );
  ANDN U7670 ( .A(n6575), .B(n4203), .Z(n6574) );
  XOR U7671 ( .A(n6576), .B(n6577), .Z(n4203) );
  IV U7672 ( .A(n6573), .Z(n6576) );
  XNOR U7673 ( .A(n4204), .B(n6573), .Z(n6575) );
  NAND U7674 ( .A(n6578), .B(nreg[954]), .Z(n4204) );
  NAND U7675 ( .A(n6107), .B(nreg[954]), .Z(n6578) );
  XOR U7676 ( .A(n6579), .B(n6580), .Z(n6573) );
  ANDN U7677 ( .A(n6581), .B(n4205), .Z(n6580) );
  XOR U7678 ( .A(n6582), .B(n6583), .Z(n4205) );
  IV U7679 ( .A(n6579), .Z(n6582) );
  XNOR U7680 ( .A(n4206), .B(n6579), .Z(n6581) );
  NAND U7681 ( .A(n6584), .B(nreg[953]), .Z(n4206) );
  NAND U7682 ( .A(n6107), .B(nreg[953]), .Z(n6584) );
  XOR U7683 ( .A(n6585), .B(n6586), .Z(n6579) );
  ANDN U7684 ( .A(n6587), .B(n4207), .Z(n6586) );
  XOR U7685 ( .A(n6588), .B(n6589), .Z(n4207) );
  IV U7686 ( .A(n6585), .Z(n6588) );
  XNOR U7687 ( .A(n4208), .B(n6585), .Z(n6587) );
  NAND U7688 ( .A(n6590), .B(nreg[952]), .Z(n4208) );
  NAND U7689 ( .A(n6107), .B(nreg[952]), .Z(n6590) );
  XOR U7690 ( .A(n6591), .B(n6592), .Z(n6585) );
  ANDN U7691 ( .A(n6593), .B(n4209), .Z(n6592) );
  XOR U7692 ( .A(n6594), .B(n6595), .Z(n4209) );
  IV U7693 ( .A(n6591), .Z(n6594) );
  XNOR U7694 ( .A(n4210), .B(n6591), .Z(n6593) );
  NAND U7695 ( .A(n6596), .B(nreg[951]), .Z(n4210) );
  NAND U7696 ( .A(n6107), .B(nreg[951]), .Z(n6596) );
  XOR U7697 ( .A(n6597), .B(n6598), .Z(n6591) );
  ANDN U7698 ( .A(n6599), .B(n4211), .Z(n6598) );
  XOR U7699 ( .A(n6600), .B(n6601), .Z(n4211) );
  IV U7700 ( .A(n6597), .Z(n6600) );
  XNOR U7701 ( .A(n4212), .B(n6597), .Z(n6599) );
  NAND U7702 ( .A(n6602), .B(nreg[950]), .Z(n4212) );
  NAND U7703 ( .A(n6107), .B(nreg[950]), .Z(n6602) );
  XOR U7704 ( .A(n6603), .B(n6604), .Z(n6597) );
  ANDN U7705 ( .A(n6605), .B(n4213), .Z(n6604) );
  XOR U7706 ( .A(n6606), .B(n6607), .Z(n4213) );
  IV U7707 ( .A(n6603), .Z(n6606) );
  XNOR U7708 ( .A(n4214), .B(n6603), .Z(n6605) );
  NAND U7709 ( .A(n6608), .B(nreg[949]), .Z(n4214) );
  NAND U7710 ( .A(n6107), .B(nreg[949]), .Z(n6608) );
  XOR U7711 ( .A(n6609), .B(n6610), .Z(n6603) );
  ANDN U7712 ( .A(n6611), .B(n4215), .Z(n6610) );
  XOR U7713 ( .A(n6612), .B(n6613), .Z(n4215) );
  IV U7714 ( .A(n6609), .Z(n6612) );
  XNOR U7715 ( .A(n4216), .B(n6609), .Z(n6611) );
  NAND U7716 ( .A(n6614), .B(nreg[948]), .Z(n4216) );
  NAND U7717 ( .A(n6107), .B(nreg[948]), .Z(n6614) );
  XOR U7718 ( .A(n6615), .B(n6616), .Z(n6609) );
  ANDN U7719 ( .A(n6617), .B(n4217), .Z(n6616) );
  XOR U7720 ( .A(n6618), .B(n6619), .Z(n4217) );
  IV U7721 ( .A(n6615), .Z(n6618) );
  XNOR U7722 ( .A(n4218), .B(n6615), .Z(n6617) );
  NAND U7723 ( .A(n6620), .B(nreg[947]), .Z(n4218) );
  NAND U7724 ( .A(n6107), .B(nreg[947]), .Z(n6620) );
  XOR U7725 ( .A(n6621), .B(n6622), .Z(n6615) );
  ANDN U7726 ( .A(n6623), .B(n4221), .Z(n6622) );
  XOR U7727 ( .A(n6624), .B(n6625), .Z(n4221) );
  IV U7728 ( .A(n6621), .Z(n6624) );
  XNOR U7729 ( .A(n4222), .B(n6621), .Z(n6623) );
  NAND U7730 ( .A(n6626), .B(nreg[946]), .Z(n4222) );
  NAND U7731 ( .A(n6107), .B(nreg[946]), .Z(n6626) );
  XOR U7732 ( .A(n6627), .B(n6628), .Z(n6621) );
  ANDN U7733 ( .A(n6629), .B(n4223), .Z(n6628) );
  XOR U7734 ( .A(n6630), .B(n6631), .Z(n4223) );
  IV U7735 ( .A(n6627), .Z(n6630) );
  XNOR U7736 ( .A(n4224), .B(n6627), .Z(n6629) );
  NAND U7737 ( .A(n6632), .B(nreg[945]), .Z(n4224) );
  NAND U7738 ( .A(n6107), .B(nreg[945]), .Z(n6632) );
  XOR U7739 ( .A(n6633), .B(n6634), .Z(n6627) );
  ANDN U7740 ( .A(n6635), .B(n4225), .Z(n6634) );
  XOR U7741 ( .A(n6636), .B(n6637), .Z(n4225) );
  IV U7742 ( .A(n6633), .Z(n6636) );
  XNOR U7743 ( .A(n4226), .B(n6633), .Z(n6635) );
  NAND U7744 ( .A(n6638), .B(nreg[944]), .Z(n4226) );
  NAND U7745 ( .A(n6107), .B(nreg[944]), .Z(n6638) );
  XOR U7746 ( .A(n6639), .B(n6640), .Z(n6633) );
  ANDN U7747 ( .A(n6641), .B(n4227), .Z(n6640) );
  XOR U7748 ( .A(n6642), .B(n6643), .Z(n4227) );
  IV U7749 ( .A(n6639), .Z(n6642) );
  XNOR U7750 ( .A(n4228), .B(n6639), .Z(n6641) );
  NAND U7751 ( .A(n6644), .B(nreg[943]), .Z(n4228) );
  NAND U7752 ( .A(n6107), .B(nreg[943]), .Z(n6644) );
  XOR U7753 ( .A(n6645), .B(n6646), .Z(n6639) );
  ANDN U7754 ( .A(n6647), .B(n4229), .Z(n6646) );
  XOR U7755 ( .A(n6648), .B(n6649), .Z(n4229) );
  IV U7756 ( .A(n6645), .Z(n6648) );
  XNOR U7757 ( .A(n4230), .B(n6645), .Z(n6647) );
  NAND U7758 ( .A(n6650), .B(nreg[942]), .Z(n4230) );
  NAND U7759 ( .A(n6107), .B(nreg[942]), .Z(n6650) );
  XOR U7760 ( .A(n6651), .B(n6652), .Z(n6645) );
  ANDN U7761 ( .A(n6653), .B(n4231), .Z(n6652) );
  XOR U7762 ( .A(n6654), .B(n6655), .Z(n4231) );
  IV U7763 ( .A(n6651), .Z(n6654) );
  XNOR U7764 ( .A(n4232), .B(n6651), .Z(n6653) );
  NAND U7765 ( .A(n6656), .B(nreg[941]), .Z(n4232) );
  NAND U7766 ( .A(n6107), .B(nreg[941]), .Z(n6656) );
  XOR U7767 ( .A(n6657), .B(n6658), .Z(n6651) );
  ANDN U7768 ( .A(n6659), .B(n4233), .Z(n6658) );
  XOR U7769 ( .A(n6660), .B(n6661), .Z(n4233) );
  IV U7770 ( .A(n6657), .Z(n6660) );
  XNOR U7771 ( .A(n4234), .B(n6657), .Z(n6659) );
  NAND U7772 ( .A(n6662), .B(nreg[940]), .Z(n4234) );
  NAND U7773 ( .A(n6107), .B(nreg[940]), .Z(n6662) );
  XOR U7774 ( .A(n6663), .B(n6664), .Z(n6657) );
  ANDN U7775 ( .A(n6665), .B(n4235), .Z(n6664) );
  XOR U7776 ( .A(n6666), .B(n6667), .Z(n4235) );
  IV U7777 ( .A(n6663), .Z(n6666) );
  XNOR U7778 ( .A(n4236), .B(n6663), .Z(n6665) );
  NAND U7779 ( .A(n6668), .B(nreg[939]), .Z(n4236) );
  NAND U7780 ( .A(n6107), .B(nreg[939]), .Z(n6668) );
  XOR U7781 ( .A(n6669), .B(n6670), .Z(n6663) );
  ANDN U7782 ( .A(n6671), .B(n4237), .Z(n6670) );
  XOR U7783 ( .A(n6672), .B(n6673), .Z(n4237) );
  IV U7784 ( .A(n6669), .Z(n6672) );
  XNOR U7785 ( .A(n4238), .B(n6669), .Z(n6671) );
  NAND U7786 ( .A(n6674), .B(nreg[938]), .Z(n4238) );
  NAND U7787 ( .A(n6107), .B(nreg[938]), .Z(n6674) );
  XOR U7788 ( .A(n6675), .B(n6676), .Z(n6669) );
  ANDN U7789 ( .A(n6677), .B(n4239), .Z(n6676) );
  XOR U7790 ( .A(n6678), .B(n6679), .Z(n4239) );
  IV U7791 ( .A(n6675), .Z(n6678) );
  XNOR U7792 ( .A(n4240), .B(n6675), .Z(n6677) );
  NAND U7793 ( .A(n6680), .B(nreg[937]), .Z(n4240) );
  NAND U7794 ( .A(n6107), .B(nreg[937]), .Z(n6680) );
  XOR U7795 ( .A(n6681), .B(n6682), .Z(n6675) );
  ANDN U7796 ( .A(n6683), .B(n4243), .Z(n6682) );
  XOR U7797 ( .A(n6684), .B(n6685), .Z(n4243) );
  IV U7798 ( .A(n6681), .Z(n6684) );
  XNOR U7799 ( .A(n4244), .B(n6681), .Z(n6683) );
  NAND U7800 ( .A(n6686), .B(nreg[936]), .Z(n4244) );
  NAND U7801 ( .A(n6107), .B(nreg[936]), .Z(n6686) );
  XOR U7802 ( .A(n6687), .B(n6688), .Z(n6681) );
  ANDN U7803 ( .A(n6689), .B(n4245), .Z(n6688) );
  XOR U7804 ( .A(n6690), .B(n6691), .Z(n4245) );
  IV U7805 ( .A(n6687), .Z(n6690) );
  XNOR U7806 ( .A(n4246), .B(n6687), .Z(n6689) );
  NAND U7807 ( .A(n6692), .B(nreg[935]), .Z(n4246) );
  NAND U7808 ( .A(n6107), .B(nreg[935]), .Z(n6692) );
  XOR U7809 ( .A(n6693), .B(n6694), .Z(n6687) );
  ANDN U7810 ( .A(n6695), .B(n4247), .Z(n6694) );
  XOR U7811 ( .A(n6696), .B(n6697), .Z(n4247) );
  IV U7812 ( .A(n6693), .Z(n6696) );
  XNOR U7813 ( .A(n4248), .B(n6693), .Z(n6695) );
  NAND U7814 ( .A(n6698), .B(nreg[934]), .Z(n4248) );
  NAND U7815 ( .A(n6107), .B(nreg[934]), .Z(n6698) );
  XOR U7816 ( .A(n6699), .B(n6700), .Z(n6693) );
  ANDN U7817 ( .A(n6701), .B(n4249), .Z(n6700) );
  XOR U7818 ( .A(n6702), .B(n6703), .Z(n4249) );
  IV U7819 ( .A(n6699), .Z(n6702) );
  XNOR U7820 ( .A(n4250), .B(n6699), .Z(n6701) );
  NAND U7821 ( .A(n6704), .B(nreg[933]), .Z(n4250) );
  NAND U7822 ( .A(n6107), .B(nreg[933]), .Z(n6704) );
  XOR U7823 ( .A(n6705), .B(n6706), .Z(n6699) );
  ANDN U7824 ( .A(n6707), .B(n4251), .Z(n6706) );
  XOR U7825 ( .A(n6708), .B(n6709), .Z(n4251) );
  IV U7826 ( .A(n6705), .Z(n6708) );
  XNOR U7827 ( .A(n4252), .B(n6705), .Z(n6707) );
  NAND U7828 ( .A(n6710), .B(nreg[932]), .Z(n4252) );
  NAND U7829 ( .A(n6107), .B(nreg[932]), .Z(n6710) );
  XOR U7830 ( .A(n6711), .B(n6712), .Z(n6705) );
  ANDN U7831 ( .A(n6713), .B(n4253), .Z(n6712) );
  XOR U7832 ( .A(n6714), .B(n6715), .Z(n4253) );
  IV U7833 ( .A(n6711), .Z(n6714) );
  XNOR U7834 ( .A(n4254), .B(n6711), .Z(n6713) );
  NAND U7835 ( .A(n6716), .B(nreg[931]), .Z(n4254) );
  NAND U7836 ( .A(n6107), .B(nreg[931]), .Z(n6716) );
  XOR U7837 ( .A(n6717), .B(n6718), .Z(n6711) );
  ANDN U7838 ( .A(n6719), .B(n4255), .Z(n6718) );
  XOR U7839 ( .A(n6720), .B(n6721), .Z(n4255) );
  IV U7840 ( .A(n6717), .Z(n6720) );
  XNOR U7841 ( .A(n4256), .B(n6717), .Z(n6719) );
  NAND U7842 ( .A(n6722), .B(nreg[930]), .Z(n4256) );
  NAND U7843 ( .A(n6107), .B(nreg[930]), .Z(n6722) );
  XOR U7844 ( .A(n6723), .B(n6724), .Z(n6717) );
  ANDN U7845 ( .A(n6725), .B(n4257), .Z(n6724) );
  XOR U7846 ( .A(n6726), .B(n6727), .Z(n4257) );
  IV U7847 ( .A(n6723), .Z(n6726) );
  XNOR U7848 ( .A(n4258), .B(n6723), .Z(n6725) );
  NAND U7849 ( .A(n6728), .B(nreg[929]), .Z(n4258) );
  NAND U7850 ( .A(n6107), .B(nreg[929]), .Z(n6728) );
  XOR U7851 ( .A(n6729), .B(n6730), .Z(n6723) );
  ANDN U7852 ( .A(n6731), .B(n4259), .Z(n6730) );
  XOR U7853 ( .A(n6732), .B(n6733), .Z(n4259) );
  IV U7854 ( .A(n6729), .Z(n6732) );
  XNOR U7855 ( .A(n4260), .B(n6729), .Z(n6731) );
  NAND U7856 ( .A(n6734), .B(nreg[928]), .Z(n4260) );
  NAND U7857 ( .A(n6107), .B(nreg[928]), .Z(n6734) );
  XOR U7858 ( .A(n6735), .B(n6736), .Z(n6729) );
  ANDN U7859 ( .A(n6737), .B(n4261), .Z(n6736) );
  XOR U7860 ( .A(n6738), .B(n6739), .Z(n4261) );
  IV U7861 ( .A(n6735), .Z(n6738) );
  XNOR U7862 ( .A(n4262), .B(n6735), .Z(n6737) );
  NAND U7863 ( .A(n6740), .B(nreg[927]), .Z(n4262) );
  NAND U7864 ( .A(n6107), .B(nreg[927]), .Z(n6740) );
  XOR U7865 ( .A(n6741), .B(n6742), .Z(n6735) );
  ANDN U7866 ( .A(n6743), .B(n4265), .Z(n6742) );
  XOR U7867 ( .A(n6744), .B(n6745), .Z(n4265) );
  IV U7868 ( .A(n6741), .Z(n6744) );
  XNOR U7869 ( .A(n4266), .B(n6741), .Z(n6743) );
  NAND U7870 ( .A(n6746), .B(nreg[926]), .Z(n4266) );
  NAND U7871 ( .A(n6107), .B(nreg[926]), .Z(n6746) );
  XOR U7872 ( .A(n6747), .B(n6748), .Z(n6741) );
  ANDN U7873 ( .A(n6749), .B(n4267), .Z(n6748) );
  XOR U7874 ( .A(n6750), .B(n6751), .Z(n4267) );
  IV U7875 ( .A(n6747), .Z(n6750) );
  XNOR U7876 ( .A(n4268), .B(n6747), .Z(n6749) );
  NAND U7877 ( .A(n6752), .B(nreg[925]), .Z(n4268) );
  NAND U7878 ( .A(n6107), .B(nreg[925]), .Z(n6752) );
  XOR U7879 ( .A(n6753), .B(n6754), .Z(n6747) );
  ANDN U7880 ( .A(n6755), .B(n4269), .Z(n6754) );
  XOR U7881 ( .A(n6756), .B(n6757), .Z(n4269) );
  IV U7882 ( .A(n6753), .Z(n6756) );
  XNOR U7883 ( .A(n4270), .B(n6753), .Z(n6755) );
  NAND U7884 ( .A(n6758), .B(nreg[924]), .Z(n4270) );
  NAND U7885 ( .A(n6107), .B(nreg[924]), .Z(n6758) );
  XOR U7886 ( .A(n6759), .B(n6760), .Z(n6753) );
  ANDN U7887 ( .A(n6761), .B(n4271), .Z(n6760) );
  XOR U7888 ( .A(n6762), .B(n6763), .Z(n4271) );
  IV U7889 ( .A(n6759), .Z(n6762) );
  XNOR U7890 ( .A(n4272), .B(n6759), .Z(n6761) );
  NAND U7891 ( .A(n6764), .B(nreg[923]), .Z(n4272) );
  NAND U7892 ( .A(n6107), .B(nreg[923]), .Z(n6764) );
  XOR U7893 ( .A(n6765), .B(n6766), .Z(n6759) );
  ANDN U7894 ( .A(n6767), .B(n4273), .Z(n6766) );
  XOR U7895 ( .A(n6768), .B(n6769), .Z(n4273) );
  IV U7896 ( .A(n6765), .Z(n6768) );
  XNOR U7897 ( .A(n4274), .B(n6765), .Z(n6767) );
  NAND U7898 ( .A(n6770), .B(nreg[922]), .Z(n4274) );
  NAND U7899 ( .A(n6107), .B(nreg[922]), .Z(n6770) );
  XOR U7900 ( .A(n6771), .B(n6772), .Z(n6765) );
  ANDN U7901 ( .A(n6773), .B(n4275), .Z(n6772) );
  XOR U7902 ( .A(n6774), .B(n6775), .Z(n4275) );
  IV U7903 ( .A(n6771), .Z(n6774) );
  XNOR U7904 ( .A(n4276), .B(n6771), .Z(n6773) );
  NAND U7905 ( .A(n6776), .B(nreg[921]), .Z(n4276) );
  NAND U7906 ( .A(n6107), .B(nreg[921]), .Z(n6776) );
  XOR U7907 ( .A(n6777), .B(n6778), .Z(n6771) );
  ANDN U7908 ( .A(n6779), .B(n4277), .Z(n6778) );
  XOR U7909 ( .A(n6780), .B(n6781), .Z(n4277) );
  IV U7910 ( .A(n6777), .Z(n6780) );
  XNOR U7911 ( .A(n4278), .B(n6777), .Z(n6779) );
  NAND U7912 ( .A(n6782), .B(nreg[920]), .Z(n4278) );
  NAND U7913 ( .A(n6107), .B(nreg[920]), .Z(n6782) );
  XOR U7914 ( .A(n6783), .B(n6784), .Z(n6777) );
  ANDN U7915 ( .A(n6785), .B(n4279), .Z(n6784) );
  XOR U7916 ( .A(n6786), .B(n6787), .Z(n4279) );
  IV U7917 ( .A(n6783), .Z(n6786) );
  XNOR U7918 ( .A(n4280), .B(n6783), .Z(n6785) );
  NAND U7919 ( .A(n6788), .B(nreg[919]), .Z(n4280) );
  NAND U7920 ( .A(n6107), .B(nreg[919]), .Z(n6788) );
  XOR U7921 ( .A(n6789), .B(n6790), .Z(n6783) );
  ANDN U7922 ( .A(n6791), .B(n4281), .Z(n6790) );
  XOR U7923 ( .A(n6792), .B(n6793), .Z(n4281) );
  IV U7924 ( .A(n6789), .Z(n6792) );
  XNOR U7925 ( .A(n4282), .B(n6789), .Z(n6791) );
  NAND U7926 ( .A(n6794), .B(nreg[918]), .Z(n4282) );
  NAND U7927 ( .A(n6107), .B(nreg[918]), .Z(n6794) );
  XOR U7928 ( .A(n6795), .B(n6796), .Z(n6789) );
  ANDN U7929 ( .A(n6797), .B(n4283), .Z(n6796) );
  XOR U7930 ( .A(n6798), .B(n6799), .Z(n4283) );
  IV U7931 ( .A(n6795), .Z(n6798) );
  XNOR U7932 ( .A(n4284), .B(n6795), .Z(n6797) );
  NAND U7933 ( .A(n6800), .B(nreg[917]), .Z(n4284) );
  NAND U7934 ( .A(n6107), .B(nreg[917]), .Z(n6800) );
  XOR U7935 ( .A(n6801), .B(n6802), .Z(n6795) );
  ANDN U7936 ( .A(n6803), .B(n4287), .Z(n6802) );
  XOR U7937 ( .A(n6804), .B(n6805), .Z(n4287) );
  IV U7938 ( .A(n6801), .Z(n6804) );
  XNOR U7939 ( .A(n4288), .B(n6801), .Z(n6803) );
  NAND U7940 ( .A(n6806), .B(nreg[916]), .Z(n4288) );
  NAND U7941 ( .A(n6107), .B(nreg[916]), .Z(n6806) );
  XOR U7942 ( .A(n6807), .B(n6808), .Z(n6801) );
  ANDN U7943 ( .A(n6809), .B(n4289), .Z(n6808) );
  XOR U7944 ( .A(n6810), .B(n6811), .Z(n4289) );
  IV U7945 ( .A(n6807), .Z(n6810) );
  XNOR U7946 ( .A(n4290), .B(n6807), .Z(n6809) );
  NAND U7947 ( .A(n6812), .B(nreg[915]), .Z(n4290) );
  NAND U7948 ( .A(n6107), .B(nreg[915]), .Z(n6812) );
  XOR U7949 ( .A(n6813), .B(n6814), .Z(n6807) );
  ANDN U7950 ( .A(n6815), .B(n4291), .Z(n6814) );
  XOR U7951 ( .A(n6816), .B(n6817), .Z(n4291) );
  IV U7952 ( .A(n6813), .Z(n6816) );
  XNOR U7953 ( .A(n4292), .B(n6813), .Z(n6815) );
  NAND U7954 ( .A(n6818), .B(nreg[914]), .Z(n4292) );
  NAND U7955 ( .A(n6107), .B(nreg[914]), .Z(n6818) );
  XOR U7956 ( .A(n6819), .B(n6820), .Z(n6813) );
  ANDN U7957 ( .A(n6821), .B(n4293), .Z(n6820) );
  XOR U7958 ( .A(n6822), .B(n6823), .Z(n4293) );
  IV U7959 ( .A(n6819), .Z(n6822) );
  XNOR U7960 ( .A(n4294), .B(n6819), .Z(n6821) );
  NAND U7961 ( .A(n6824), .B(nreg[913]), .Z(n4294) );
  NAND U7962 ( .A(n6107), .B(nreg[913]), .Z(n6824) );
  XOR U7963 ( .A(n6825), .B(n6826), .Z(n6819) );
  ANDN U7964 ( .A(n6827), .B(n4295), .Z(n6826) );
  XOR U7965 ( .A(n6828), .B(n6829), .Z(n4295) );
  IV U7966 ( .A(n6825), .Z(n6828) );
  XNOR U7967 ( .A(n4296), .B(n6825), .Z(n6827) );
  NAND U7968 ( .A(n6830), .B(nreg[912]), .Z(n4296) );
  NAND U7969 ( .A(n6107), .B(nreg[912]), .Z(n6830) );
  XOR U7970 ( .A(n6831), .B(n6832), .Z(n6825) );
  ANDN U7971 ( .A(n6833), .B(n4297), .Z(n6832) );
  XOR U7972 ( .A(n6834), .B(n6835), .Z(n4297) );
  IV U7973 ( .A(n6831), .Z(n6834) );
  XNOR U7974 ( .A(n4298), .B(n6831), .Z(n6833) );
  NAND U7975 ( .A(n6836), .B(nreg[911]), .Z(n4298) );
  NAND U7976 ( .A(n6107), .B(nreg[911]), .Z(n6836) );
  XOR U7977 ( .A(n6837), .B(n6838), .Z(n6831) );
  ANDN U7978 ( .A(n6839), .B(n4299), .Z(n6838) );
  XOR U7979 ( .A(n6840), .B(n6841), .Z(n4299) );
  IV U7980 ( .A(n6837), .Z(n6840) );
  XNOR U7981 ( .A(n4300), .B(n6837), .Z(n6839) );
  NAND U7982 ( .A(n6842), .B(nreg[910]), .Z(n4300) );
  NAND U7983 ( .A(n6107), .B(nreg[910]), .Z(n6842) );
  XOR U7984 ( .A(n6843), .B(n6844), .Z(n6837) );
  ANDN U7985 ( .A(n6845), .B(n4301), .Z(n6844) );
  XOR U7986 ( .A(n6846), .B(n6847), .Z(n4301) );
  IV U7987 ( .A(n6843), .Z(n6846) );
  XNOR U7988 ( .A(n4302), .B(n6843), .Z(n6845) );
  NAND U7989 ( .A(n6848), .B(nreg[909]), .Z(n4302) );
  NAND U7990 ( .A(n6107), .B(nreg[909]), .Z(n6848) );
  XOR U7991 ( .A(n6849), .B(n6850), .Z(n6843) );
  ANDN U7992 ( .A(n6851), .B(n4303), .Z(n6850) );
  XOR U7993 ( .A(n6852), .B(n6853), .Z(n4303) );
  IV U7994 ( .A(n6849), .Z(n6852) );
  XNOR U7995 ( .A(n4304), .B(n6849), .Z(n6851) );
  NAND U7996 ( .A(n6854), .B(nreg[908]), .Z(n4304) );
  NAND U7997 ( .A(n6107), .B(nreg[908]), .Z(n6854) );
  XOR U7998 ( .A(n6855), .B(n6856), .Z(n6849) );
  ANDN U7999 ( .A(n6857), .B(n4305), .Z(n6856) );
  XOR U8000 ( .A(n6858), .B(n6859), .Z(n4305) );
  IV U8001 ( .A(n6855), .Z(n6858) );
  XNOR U8002 ( .A(n4306), .B(n6855), .Z(n6857) );
  NAND U8003 ( .A(n6860), .B(nreg[907]), .Z(n4306) );
  NAND U8004 ( .A(n6107), .B(nreg[907]), .Z(n6860) );
  XOR U8005 ( .A(n6861), .B(n6862), .Z(n6855) );
  ANDN U8006 ( .A(n6863), .B(n4309), .Z(n6862) );
  XOR U8007 ( .A(n6864), .B(n6865), .Z(n4309) );
  IV U8008 ( .A(n6861), .Z(n6864) );
  XNOR U8009 ( .A(n4310), .B(n6861), .Z(n6863) );
  NAND U8010 ( .A(n6866), .B(nreg[906]), .Z(n4310) );
  NAND U8011 ( .A(n6107), .B(nreg[906]), .Z(n6866) );
  XOR U8012 ( .A(n6867), .B(n6868), .Z(n6861) );
  ANDN U8013 ( .A(n6869), .B(n4311), .Z(n6868) );
  XOR U8014 ( .A(n6870), .B(n6871), .Z(n4311) );
  IV U8015 ( .A(n6867), .Z(n6870) );
  XNOR U8016 ( .A(n4312), .B(n6867), .Z(n6869) );
  NAND U8017 ( .A(n6872), .B(nreg[905]), .Z(n4312) );
  NAND U8018 ( .A(n6107), .B(nreg[905]), .Z(n6872) );
  XOR U8019 ( .A(n6873), .B(n6874), .Z(n6867) );
  ANDN U8020 ( .A(n6875), .B(n4313), .Z(n6874) );
  XOR U8021 ( .A(n6876), .B(n6877), .Z(n4313) );
  IV U8022 ( .A(n6873), .Z(n6876) );
  XNOR U8023 ( .A(n4314), .B(n6873), .Z(n6875) );
  NAND U8024 ( .A(n6878), .B(nreg[904]), .Z(n4314) );
  NAND U8025 ( .A(n6107), .B(nreg[904]), .Z(n6878) );
  XOR U8026 ( .A(n6879), .B(n6880), .Z(n6873) );
  ANDN U8027 ( .A(n6881), .B(n4315), .Z(n6880) );
  XOR U8028 ( .A(n6882), .B(n6883), .Z(n4315) );
  IV U8029 ( .A(n6879), .Z(n6882) );
  XNOR U8030 ( .A(n4316), .B(n6879), .Z(n6881) );
  NAND U8031 ( .A(n6884), .B(nreg[903]), .Z(n4316) );
  NAND U8032 ( .A(n6107), .B(nreg[903]), .Z(n6884) );
  XOR U8033 ( .A(n6885), .B(n6886), .Z(n6879) );
  ANDN U8034 ( .A(n6887), .B(n4317), .Z(n6886) );
  XOR U8035 ( .A(n6888), .B(n6889), .Z(n4317) );
  IV U8036 ( .A(n6885), .Z(n6888) );
  XNOR U8037 ( .A(n4318), .B(n6885), .Z(n6887) );
  NAND U8038 ( .A(n6890), .B(nreg[902]), .Z(n4318) );
  NAND U8039 ( .A(n6107), .B(nreg[902]), .Z(n6890) );
  XOR U8040 ( .A(n6891), .B(n6892), .Z(n6885) );
  ANDN U8041 ( .A(n6893), .B(n4319), .Z(n6892) );
  XOR U8042 ( .A(n6894), .B(n6895), .Z(n4319) );
  IV U8043 ( .A(n6891), .Z(n6894) );
  XNOR U8044 ( .A(n4320), .B(n6891), .Z(n6893) );
  NAND U8045 ( .A(n6896), .B(nreg[901]), .Z(n4320) );
  NAND U8046 ( .A(n6107), .B(nreg[901]), .Z(n6896) );
  XOR U8047 ( .A(n6897), .B(n6898), .Z(n6891) );
  ANDN U8048 ( .A(n6899), .B(n4321), .Z(n6898) );
  XOR U8049 ( .A(n6900), .B(n6901), .Z(n4321) );
  IV U8050 ( .A(n6897), .Z(n6900) );
  XNOR U8051 ( .A(n4322), .B(n6897), .Z(n6899) );
  NAND U8052 ( .A(n6902), .B(nreg[900]), .Z(n4322) );
  NAND U8053 ( .A(n6107), .B(nreg[900]), .Z(n6902) );
  XOR U8054 ( .A(n6903), .B(n6904), .Z(n6897) );
  ANDN U8055 ( .A(n6905), .B(n4323), .Z(n6904) );
  XOR U8056 ( .A(n6906), .B(n6907), .Z(n4323) );
  IV U8057 ( .A(n6903), .Z(n6906) );
  XNOR U8058 ( .A(n4324), .B(n6903), .Z(n6905) );
  NAND U8059 ( .A(n6908), .B(nreg[899]), .Z(n4324) );
  NAND U8060 ( .A(n6107), .B(nreg[899]), .Z(n6908) );
  XOR U8061 ( .A(n6909), .B(n6910), .Z(n6903) );
  ANDN U8062 ( .A(n6911), .B(n4325), .Z(n6910) );
  XOR U8063 ( .A(n6912), .B(n6913), .Z(n4325) );
  IV U8064 ( .A(n6909), .Z(n6912) );
  XNOR U8065 ( .A(n4326), .B(n6909), .Z(n6911) );
  NAND U8066 ( .A(n6914), .B(nreg[898]), .Z(n4326) );
  NAND U8067 ( .A(n6107), .B(nreg[898]), .Z(n6914) );
  XOR U8068 ( .A(n6915), .B(n6916), .Z(n6909) );
  ANDN U8069 ( .A(n6917), .B(n4327), .Z(n6916) );
  XOR U8070 ( .A(n6918), .B(n6919), .Z(n4327) );
  IV U8071 ( .A(n6915), .Z(n6918) );
  XNOR U8072 ( .A(n4328), .B(n6915), .Z(n6917) );
  NAND U8073 ( .A(n6920), .B(nreg[897]), .Z(n4328) );
  NAND U8074 ( .A(n6107), .B(nreg[897]), .Z(n6920) );
  XOR U8075 ( .A(n6921), .B(n6922), .Z(n6915) );
  ANDN U8076 ( .A(n6923), .B(n4333), .Z(n6922) );
  XOR U8077 ( .A(n6924), .B(n6925), .Z(n4333) );
  IV U8078 ( .A(n6921), .Z(n6924) );
  XNOR U8079 ( .A(n4334), .B(n6921), .Z(n6923) );
  NAND U8080 ( .A(n6926), .B(nreg[896]), .Z(n4334) );
  NAND U8081 ( .A(n6107), .B(nreg[896]), .Z(n6926) );
  XOR U8082 ( .A(n6927), .B(n6928), .Z(n6921) );
  ANDN U8083 ( .A(n6929), .B(n4335), .Z(n6928) );
  XOR U8084 ( .A(n6930), .B(n6931), .Z(n4335) );
  IV U8085 ( .A(n6927), .Z(n6930) );
  XNOR U8086 ( .A(n4336), .B(n6927), .Z(n6929) );
  NAND U8087 ( .A(n6932), .B(nreg[895]), .Z(n4336) );
  NAND U8088 ( .A(n6107), .B(nreg[895]), .Z(n6932) );
  XOR U8089 ( .A(n6933), .B(n6934), .Z(n6927) );
  ANDN U8090 ( .A(n6935), .B(n4337), .Z(n6934) );
  XOR U8091 ( .A(n6936), .B(n6937), .Z(n4337) );
  IV U8092 ( .A(n6933), .Z(n6936) );
  XNOR U8093 ( .A(n4338), .B(n6933), .Z(n6935) );
  NAND U8094 ( .A(n6938), .B(nreg[894]), .Z(n4338) );
  NAND U8095 ( .A(n6107), .B(nreg[894]), .Z(n6938) );
  XOR U8096 ( .A(n6939), .B(n6940), .Z(n6933) );
  ANDN U8097 ( .A(n6941), .B(n4339), .Z(n6940) );
  XOR U8098 ( .A(n6942), .B(n6943), .Z(n4339) );
  IV U8099 ( .A(n6939), .Z(n6942) );
  XNOR U8100 ( .A(n4340), .B(n6939), .Z(n6941) );
  NAND U8101 ( .A(n6944), .B(nreg[893]), .Z(n4340) );
  NAND U8102 ( .A(n6107), .B(nreg[893]), .Z(n6944) );
  XOR U8103 ( .A(n6945), .B(n6946), .Z(n6939) );
  ANDN U8104 ( .A(n6947), .B(n4341), .Z(n6946) );
  XOR U8105 ( .A(n6948), .B(n6949), .Z(n4341) );
  IV U8106 ( .A(n6945), .Z(n6948) );
  XNOR U8107 ( .A(n4342), .B(n6945), .Z(n6947) );
  NAND U8108 ( .A(n6950), .B(nreg[892]), .Z(n4342) );
  NAND U8109 ( .A(n6107), .B(nreg[892]), .Z(n6950) );
  XOR U8110 ( .A(n6951), .B(n6952), .Z(n6945) );
  ANDN U8111 ( .A(n6953), .B(n4343), .Z(n6952) );
  XOR U8112 ( .A(n6954), .B(n6955), .Z(n4343) );
  IV U8113 ( .A(n6951), .Z(n6954) );
  XNOR U8114 ( .A(n4344), .B(n6951), .Z(n6953) );
  NAND U8115 ( .A(n6956), .B(nreg[891]), .Z(n4344) );
  NAND U8116 ( .A(n6107), .B(nreg[891]), .Z(n6956) );
  XOR U8117 ( .A(n6957), .B(n6958), .Z(n6951) );
  ANDN U8118 ( .A(n6959), .B(n4345), .Z(n6958) );
  XOR U8119 ( .A(n6960), .B(n6961), .Z(n4345) );
  IV U8120 ( .A(n6957), .Z(n6960) );
  XNOR U8121 ( .A(n4346), .B(n6957), .Z(n6959) );
  NAND U8122 ( .A(n6962), .B(nreg[890]), .Z(n4346) );
  NAND U8123 ( .A(n6107), .B(nreg[890]), .Z(n6962) );
  XOR U8124 ( .A(n6963), .B(n6964), .Z(n6957) );
  ANDN U8125 ( .A(n6965), .B(n4347), .Z(n6964) );
  XOR U8126 ( .A(n6966), .B(n6967), .Z(n4347) );
  IV U8127 ( .A(n6963), .Z(n6966) );
  XNOR U8128 ( .A(n4348), .B(n6963), .Z(n6965) );
  NAND U8129 ( .A(n6968), .B(nreg[889]), .Z(n4348) );
  NAND U8130 ( .A(n6107), .B(nreg[889]), .Z(n6968) );
  XOR U8131 ( .A(n6969), .B(n6970), .Z(n6963) );
  ANDN U8132 ( .A(n6971), .B(n4349), .Z(n6970) );
  XOR U8133 ( .A(n6972), .B(n6973), .Z(n4349) );
  IV U8134 ( .A(n6969), .Z(n6972) );
  XNOR U8135 ( .A(n4350), .B(n6969), .Z(n6971) );
  NAND U8136 ( .A(n6974), .B(nreg[888]), .Z(n4350) );
  NAND U8137 ( .A(n6107), .B(nreg[888]), .Z(n6974) );
  XOR U8138 ( .A(n6975), .B(n6976), .Z(n6969) );
  ANDN U8139 ( .A(n6977), .B(n4351), .Z(n6976) );
  XOR U8140 ( .A(n6978), .B(n6979), .Z(n4351) );
  IV U8141 ( .A(n6975), .Z(n6978) );
  XNOR U8142 ( .A(n4352), .B(n6975), .Z(n6977) );
  NAND U8143 ( .A(n6980), .B(nreg[887]), .Z(n4352) );
  NAND U8144 ( .A(n6107), .B(nreg[887]), .Z(n6980) );
  XOR U8145 ( .A(n6981), .B(n6982), .Z(n6975) );
  ANDN U8146 ( .A(n6983), .B(n4355), .Z(n6982) );
  XOR U8147 ( .A(n6984), .B(n6985), .Z(n4355) );
  IV U8148 ( .A(n6981), .Z(n6984) );
  XNOR U8149 ( .A(n4356), .B(n6981), .Z(n6983) );
  NAND U8150 ( .A(n6986), .B(nreg[886]), .Z(n4356) );
  NAND U8151 ( .A(n6107), .B(nreg[886]), .Z(n6986) );
  XOR U8152 ( .A(n6987), .B(n6988), .Z(n6981) );
  ANDN U8153 ( .A(n6989), .B(n4357), .Z(n6988) );
  XOR U8154 ( .A(n6990), .B(n6991), .Z(n4357) );
  IV U8155 ( .A(n6987), .Z(n6990) );
  XNOR U8156 ( .A(n4358), .B(n6987), .Z(n6989) );
  NAND U8157 ( .A(n6992), .B(nreg[885]), .Z(n4358) );
  NAND U8158 ( .A(n6107), .B(nreg[885]), .Z(n6992) );
  XOR U8159 ( .A(n6993), .B(n6994), .Z(n6987) );
  ANDN U8160 ( .A(n6995), .B(n4359), .Z(n6994) );
  XOR U8161 ( .A(n6996), .B(n6997), .Z(n4359) );
  IV U8162 ( .A(n6993), .Z(n6996) );
  XNOR U8163 ( .A(n4360), .B(n6993), .Z(n6995) );
  NAND U8164 ( .A(n6998), .B(nreg[884]), .Z(n4360) );
  NAND U8165 ( .A(n6107), .B(nreg[884]), .Z(n6998) );
  XOR U8166 ( .A(n6999), .B(n7000), .Z(n6993) );
  ANDN U8167 ( .A(n7001), .B(n4361), .Z(n7000) );
  XOR U8168 ( .A(n7002), .B(n7003), .Z(n4361) );
  IV U8169 ( .A(n6999), .Z(n7002) );
  XNOR U8170 ( .A(n4362), .B(n6999), .Z(n7001) );
  NAND U8171 ( .A(n7004), .B(nreg[883]), .Z(n4362) );
  NAND U8172 ( .A(n6107), .B(nreg[883]), .Z(n7004) );
  XOR U8173 ( .A(n7005), .B(n7006), .Z(n6999) );
  ANDN U8174 ( .A(n7007), .B(n4363), .Z(n7006) );
  XOR U8175 ( .A(n7008), .B(n7009), .Z(n4363) );
  IV U8176 ( .A(n7005), .Z(n7008) );
  XNOR U8177 ( .A(n4364), .B(n7005), .Z(n7007) );
  NAND U8178 ( .A(n7010), .B(nreg[882]), .Z(n4364) );
  NAND U8179 ( .A(n6107), .B(nreg[882]), .Z(n7010) );
  XOR U8180 ( .A(n7011), .B(n7012), .Z(n7005) );
  ANDN U8181 ( .A(n7013), .B(n4365), .Z(n7012) );
  XOR U8182 ( .A(n7014), .B(n7015), .Z(n4365) );
  IV U8183 ( .A(n7011), .Z(n7014) );
  XNOR U8184 ( .A(n4366), .B(n7011), .Z(n7013) );
  NAND U8185 ( .A(n7016), .B(nreg[881]), .Z(n4366) );
  NAND U8186 ( .A(n6107), .B(nreg[881]), .Z(n7016) );
  XOR U8187 ( .A(n7017), .B(n7018), .Z(n7011) );
  ANDN U8188 ( .A(n7019), .B(n4367), .Z(n7018) );
  XOR U8189 ( .A(n7020), .B(n7021), .Z(n4367) );
  IV U8190 ( .A(n7017), .Z(n7020) );
  XNOR U8191 ( .A(n4368), .B(n7017), .Z(n7019) );
  NAND U8192 ( .A(n7022), .B(nreg[880]), .Z(n4368) );
  NAND U8193 ( .A(n6107), .B(nreg[880]), .Z(n7022) );
  XOR U8194 ( .A(n7023), .B(n7024), .Z(n7017) );
  ANDN U8195 ( .A(n7025), .B(n4369), .Z(n7024) );
  XOR U8196 ( .A(n7026), .B(n7027), .Z(n4369) );
  IV U8197 ( .A(n7023), .Z(n7026) );
  XNOR U8198 ( .A(n4370), .B(n7023), .Z(n7025) );
  NAND U8199 ( .A(n7028), .B(nreg[879]), .Z(n4370) );
  NAND U8200 ( .A(n6107), .B(nreg[879]), .Z(n7028) );
  XOR U8201 ( .A(n7029), .B(n7030), .Z(n7023) );
  ANDN U8202 ( .A(n7031), .B(n4371), .Z(n7030) );
  XOR U8203 ( .A(n7032), .B(n7033), .Z(n4371) );
  IV U8204 ( .A(n7029), .Z(n7032) );
  XNOR U8205 ( .A(n4372), .B(n7029), .Z(n7031) );
  NAND U8206 ( .A(n7034), .B(nreg[878]), .Z(n4372) );
  NAND U8207 ( .A(n6107), .B(nreg[878]), .Z(n7034) );
  XOR U8208 ( .A(n7035), .B(n7036), .Z(n7029) );
  ANDN U8209 ( .A(n7037), .B(n4373), .Z(n7036) );
  XOR U8210 ( .A(n7038), .B(n7039), .Z(n4373) );
  IV U8211 ( .A(n7035), .Z(n7038) );
  XNOR U8212 ( .A(n4374), .B(n7035), .Z(n7037) );
  NAND U8213 ( .A(n7040), .B(nreg[877]), .Z(n4374) );
  NAND U8214 ( .A(n6107), .B(nreg[877]), .Z(n7040) );
  XOR U8215 ( .A(n7041), .B(n7042), .Z(n7035) );
  ANDN U8216 ( .A(n7043), .B(n4377), .Z(n7042) );
  XOR U8217 ( .A(n7044), .B(n7045), .Z(n4377) );
  IV U8218 ( .A(n7041), .Z(n7044) );
  XNOR U8219 ( .A(n4378), .B(n7041), .Z(n7043) );
  NAND U8220 ( .A(n7046), .B(nreg[876]), .Z(n4378) );
  NAND U8221 ( .A(n6107), .B(nreg[876]), .Z(n7046) );
  XOR U8222 ( .A(n7047), .B(n7048), .Z(n7041) );
  ANDN U8223 ( .A(n7049), .B(n4379), .Z(n7048) );
  XOR U8224 ( .A(n7050), .B(n7051), .Z(n4379) );
  IV U8225 ( .A(n7047), .Z(n7050) );
  XNOR U8226 ( .A(n4380), .B(n7047), .Z(n7049) );
  NAND U8227 ( .A(n7052), .B(nreg[875]), .Z(n4380) );
  NAND U8228 ( .A(n6107), .B(nreg[875]), .Z(n7052) );
  XOR U8229 ( .A(n7053), .B(n7054), .Z(n7047) );
  ANDN U8230 ( .A(n7055), .B(n4381), .Z(n7054) );
  XOR U8231 ( .A(n7056), .B(n7057), .Z(n4381) );
  IV U8232 ( .A(n7053), .Z(n7056) );
  XNOR U8233 ( .A(n4382), .B(n7053), .Z(n7055) );
  NAND U8234 ( .A(n7058), .B(nreg[874]), .Z(n4382) );
  NAND U8235 ( .A(n6107), .B(nreg[874]), .Z(n7058) );
  XOR U8236 ( .A(n7059), .B(n7060), .Z(n7053) );
  ANDN U8237 ( .A(n7061), .B(n4383), .Z(n7060) );
  XOR U8238 ( .A(n7062), .B(n7063), .Z(n4383) );
  IV U8239 ( .A(n7059), .Z(n7062) );
  XNOR U8240 ( .A(n4384), .B(n7059), .Z(n7061) );
  NAND U8241 ( .A(n7064), .B(nreg[873]), .Z(n4384) );
  NAND U8242 ( .A(n6107), .B(nreg[873]), .Z(n7064) );
  XOR U8243 ( .A(n7065), .B(n7066), .Z(n7059) );
  ANDN U8244 ( .A(n7067), .B(n4385), .Z(n7066) );
  XOR U8245 ( .A(n7068), .B(n7069), .Z(n4385) );
  IV U8246 ( .A(n7065), .Z(n7068) );
  XNOR U8247 ( .A(n4386), .B(n7065), .Z(n7067) );
  NAND U8248 ( .A(n7070), .B(nreg[872]), .Z(n4386) );
  NAND U8249 ( .A(n6107), .B(nreg[872]), .Z(n7070) );
  XOR U8250 ( .A(n7071), .B(n7072), .Z(n7065) );
  ANDN U8251 ( .A(n7073), .B(n4387), .Z(n7072) );
  XOR U8252 ( .A(n7074), .B(n7075), .Z(n4387) );
  IV U8253 ( .A(n7071), .Z(n7074) );
  XNOR U8254 ( .A(n4388), .B(n7071), .Z(n7073) );
  NAND U8255 ( .A(n7076), .B(nreg[871]), .Z(n4388) );
  NAND U8256 ( .A(n6107), .B(nreg[871]), .Z(n7076) );
  XOR U8257 ( .A(n7077), .B(n7078), .Z(n7071) );
  ANDN U8258 ( .A(n7079), .B(n4389), .Z(n7078) );
  XOR U8259 ( .A(n7080), .B(n7081), .Z(n4389) );
  IV U8260 ( .A(n7077), .Z(n7080) );
  XNOR U8261 ( .A(n4390), .B(n7077), .Z(n7079) );
  NAND U8262 ( .A(n7082), .B(nreg[870]), .Z(n4390) );
  NAND U8263 ( .A(n6107), .B(nreg[870]), .Z(n7082) );
  XOR U8264 ( .A(n7083), .B(n7084), .Z(n7077) );
  ANDN U8265 ( .A(n7085), .B(n4391), .Z(n7084) );
  XOR U8266 ( .A(n7086), .B(n7087), .Z(n4391) );
  IV U8267 ( .A(n7083), .Z(n7086) );
  XNOR U8268 ( .A(n4392), .B(n7083), .Z(n7085) );
  NAND U8269 ( .A(n7088), .B(nreg[869]), .Z(n4392) );
  NAND U8270 ( .A(n6107), .B(nreg[869]), .Z(n7088) );
  XOR U8271 ( .A(n7089), .B(n7090), .Z(n7083) );
  ANDN U8272 ( .A(n7091), .B(n4393), .Z(n7090) );
  XOR U8273 ( .A(n7092), .B(n7093), .Z(n4393) );
  IV U8274 ( .A(n7089), .Z(n7092) );
  XNOR U8275 ( .A(n4394), .B(n7089), .Z(n7091) );
  NAND U8276 ( .A(n7094), .B(nreg[868]), .Z(n4394) );
  NAND U8277 ( .A(n6107), .B(nreg[868]), .Z(n7094) );
  XOR U8278 ( .A(n7095), .B(n7096), .Z(n7089) );
  ANDN U8279 ( .A(n7097), .B(n4395), .Z(n7096) );
  XOR U8280 ( .A(n7098), .B(n7099), .Z(n4395) );
  IV U8281 ( .A(n7095), .Z(n7098) );
  XNOR U8282 ( .A(n4396), .B(n7095), .Z(n7097) );
  NAND U8283 ( .A(n7100), .B(nreg[867]), .Z(n4396) );
  NAND U8284 ( .A(n6107), .B(nreg[867]), .Z(n7100) );
  XOR U8285 ( .A(n7101), .B(n7102), .Z(n7095) );
  ANDN U8286 ( .A(n7103), .B(n4399), .Z(n7102) );
  XOR U8287 ( .A(n7104), .B(n7105), .Z(n4399) );
  IV U8288 ( .A(n7101), .Z(n7104) );
  XNOR U8289 ( .A(n4400), .B(n7101), .Z(n7103) );
  NAND U8290 ( .A(n7106), .B(nreg[866]), .Z(n4400) );
  NAND U8291 ( .A(n6107), .B(nreg[866]), .Z(n7106) );
  XOR U8292 ( .A(n7107), .B(n7108), .Z(n7101) );
  ANDN U8293 ( .A(n7109), .B(n4401), .Z(n7108) );
  XOR U8294 ( .A(n7110), .B(n7111), .Z(n4401) );
  IV U8295 ( .A(n7107), .Z(n7110) );
  XNOR U8296 ( .A(n4402), .B(n7107), .Z(n7109) );
  NAND U8297 ( .A(n7112), .B(nreg[865]), .Z(n4402) );
  NAND U8298 ( .A(n6107), .B(nreg[865]), .Z(n7112) );
  XOR U8299 ( .A(n7113), .B(n7114), .Z(n7107) );
  ANDN U8300 ( .A(n7115), .B(n4403), .Z(n7114) );
  XOR U8301 ( .A(n7116), .B(n7117), .Z(n4403) );
  IV U8302 ( .A(n7113), .Z(n7116) );
  XNOR U8303 ( .A(n4404), .B(n7113), .Z(n7115) );
  NAND U8304 ( .A(n7118), .B(nreg[864]), .Z(n4404) );
  NAND U8305 ( .A(n6107), .B(nreg[864]), .Z(n7118) );
  XOR U8306 ( .A(n7119), .B(n7120), .Z(n7113) );
  ANDN U8307 ( .A(n7121), .B(n4405), .Z(n7120) );
  XOR U8308 ( .A(n7122), .B(n7123), .Z(n4405) );
  IV U8309 ( .A(n7119), .Z(n7122) );
  XNOR U8310 ( .A(n4406), .B(n7119), .Z(n7121) );
  NAND U8311 ( .A(n7124), .B(nreg[863]), .Z(n4406) );
  NAND U8312 ( .A(n6107), .B(nreg[863]), .Z(n7124) );
  XOR U8313 ( .A(n7125), .B(n7126), .Z(n7119) );
  ANDN U8314 ( .A(n7127), .B(n4407), .Z(n7126) );
  XOR U8315 ( .A(n7128), .B(n7129), .Z(n4407) );
  IV U8316 ( .A(n7125), .Z(n7128) );
  XNOR U8317 ( .A(n4408), .B(n7125), .Z(n7127) );
  NAND U8318 ( .A(n7130), .B(nreg[862]), .Z(n4408) );
  NAND U8319 ( .A(n6107), .B(nreg[862]), .Z(n7130) );
  XOR U8320 ( .A(n7131), .B(n7132), .Z(n7125) );
  ANDN U8321 ( .A(n7133), .B(n4409), .Z(n7132) );
  XOR U8322 ( .A(n7134), .B(n7135), .Z(n4409) );
  IV U8323 ( .A(n7131), .Z(n7134) );
  XNOR U8324 ( .A(n4410), .B(n7131), .Z(n7133) );
  NAND U8325 ( .A(n7136), .B(nreg[861]), .Z(n4410) );
  NAND U8326 ( .A(n6107), .B(nreg[861]), .Z(n7136) );
  XOR U8327 ( .A(n7137), .B(n7138), .Z(n7131) );
  ANDN U8328 ( .A(n7139), .B(n4411), .Z(n7138) );
  XOR U8329 ( .A(n7140), .B(n7141), .Z(n4411) );
  IV U8330 ( .A(n7137), .Z(n7140) );
  XNOR U8331 ( .A(n4412), .B(n7137), .Z(n7139) );
  NAND U8332 ( .A(n7142), .B(nreg[860]), .Z(n4412) );
  NAND U8333 ( .A(n6107), .B(nreg[860]), .Z(n7142) );
  XOR U8334 ( .A(n7143), .B(n7144), .Z(n7137) );
  ANDN U8335 ( .A(n7145), .B(n4413), .Z(n7144) );
  XOR U8336 ( .A(n7146), .B(n7147), .Z(n4413) );
  IV U8337 ( .A(n7143), .Z(n7146) );
  XNOR U8338 ( .A(n4414), .B(n7143), .Z(n7145) );
  NAND U8339 ( .A(n7148), .B(nreg[859]), .Z(n4414) );
  NAND U8340 ( .A(n6107), .B(nreg[859]), .Z(n7148) );
  XOR U8341 ( .A(n7149), .B(n7150), .Z(n7143) );
  ANDN U8342 ( .A(n7151), .B(n4415), .Z(n7150) );
  XOR U8343 ( .A(n7152), .B(n7153), .Z(n4415) );
  IV U8344 ( .A(n7149), .Z(n7152) );
  XNOR U8345 ( .A(n4416), .B(n7149), .Z(n7151) );
  NAND U8346 ( .A(n7154), .B(nreg[858]), .Z(n4416) );
  NAND U8347 ( .A(n6107), .B(nreg[858]), .Z(n7154) );
  XOR U8348 ( .A(n7155), .B(n7156), .Z(n7149) );
  ANDN U8349 ( .A(n7157), .B(n4417), .Z(n7156) );
  XOR U8350 ( .A(n7158), .B(n7159), .Z(n4417) );
  IV U8351 ( .A(n7155), .Z(n7158) );
  XNOR U8352 ( .A(n4418), .B(n7155), .Z(n7157) );
  NAND U8353 ( .A(n7160), .B(nreg[857]), .Z(n4418) );
  NAND U8354 ( .A(n6107), .B(nreg[857]), .Z(n7160) );
  XOR U8355 ( .A(n7161), .B(n7162), .Z(n7155) );
  ANDN U8356 ( .A(n7163), .B(n4421), .Z(n7162) );
  XOR U8357 ( .A(n7164), .B(n7165), .Z(n4421) );
  IV U8358 ( .A(n7161), .Z(n7164) );
  XNOR U8359 ( .A(n4422), .B(n7161), .Z(n7163) );
  NAND U8360 ( .A(n7166), .B(nreg[856]), .Z(n4422) );
  NAND U8361 ( .A(n6107), .B(nreg[856]), .Z(n7166) );
  XOR U8362 ( .A(n7167), .B(n7168), .Z(n7161) );
  ANDN U8363 ( .A(n7169), .B(n4423), .Z(n7168) );
  XOR U8364 ( .A(n7170), .B(n7171), .Z(n4423) );
  IV U8365 ( .A(n7167), .Z(n7170) );
  XNOR U8366 ( .A(n4424), .B(n7167), .Z(n7169) );
  NAND U8367 ( .A(n7172), .B(nreg[855]), .Z(n4424) );
  NAND U8368 ( .A(n6107), .B(nreg[855]), .Z(n7172) );
  XOR U8369 ( .A(n7173), .B(n7174), .Z(n7167) );
  ANDN U8370 ( .A(n7175), .B(n4425), .Z(n7174) );
  XOR U8371 ( .A(n7176), .B(n7177), .Z(n4425) );
  IV U8372 ( .A(n7173), .Z(n7176) );
  XNOR U8373 ( .A(n4426), .B(n7173), .Z(n7175) );
  NAND U8374 ( .A(n7178), .B(nreg[854]), .Z(n4426) );
  NAND U8375 ( .A(n6107), .B(nreg[854]), .Z(n7178) );
  XOR U8376 ( .A(n7179), .B(n7180), .Z(n7173) );
  ANDN U8377 ( .A(n7181), .B(n4427), .Z(n7180) );
  XOR U8378 ( .A(n7182), .B(n7183), .Z(n4427) );
  IV U8379 ( .A(n7179), .Z(n7182) );
  XNOR U8380 ( .A(n4428), .B(n7179), .Z(n7181) );
  NAND U8381 ( .A(n7184), .B(nreg[853]), .Z(n4428) );
  NAND U8382 ( .A(n6107), .B(nreg[853]), .Z(n7184) );
  XOR U8383 ( .A(n7185), .B(n7186), .Z(n7179) );
  ANDN U8384 ( .A(n7187), .B(n4429), .Z(n7186) );
  XOR U8385 ( .A(n7188), .B(n7189), .Z(n4429) );
  IV U8386 ( .A(n7185), .Z(n7188) );
  XNOR U8387 ( .A(n4430), .B(n7185), .Z(n7187) );
  NAND U8388 ( .A(n7190), .B(nreg[852]), .Z(n4430) );
  NAND U8389 ( .A(n6107), .B(nreg[852]), .Z(n7190) );
  XOR U8390 ( .A(n7191), .B(n7192), .Z(n7185) );
  ANDN U8391 ( .A(n7193), .B(n4431), .Z(n7192) );
  XOR U8392 ( .A(n7194), .B(n7195), .Z(n4431) );
  IV U8393 ( .A(n7191), .Z(n7194) );
  XNOR U8394 ( .A(n4432), .B(n7191), .Z(n7193) );
  NAND U8395 ( .A(n7196), .B(nreg[851]), .Z(n4432) );
  NAND U8396 ( .A(n6107), .B(nreg[851]), .Z(n7196) );
  XOR U8397 ( .A(n7197), .B(n7198), .Z(n7191) );
  ANDN U8398 ( .A(n7199), .B(n4433), .Z(n7198) );
  XOR U8399 ( .A(n7200), .B(n7201), .Z(n4433) );
  IV U8400 ( .A(n7197), .Z(n7200) );
  XNOR U8401 ( .A(n4434), .B(n7197), .Z(n7199) );
  NAND U8402 ( .A(n7202), .B(nreg[850]), .Z(n4434) );
  NAND U8403 ( .A(n6107), .B(nreg[850]), .Z(n7202) );
  XOR U8404 ( .A(n7203), .B(n7204), .Z(n7197) );
  ANDN U8405 ( .A(n7205), .B(n4435), .Z(n7204) );
  XOR U8406 ( .A(n7206), .B(n7207), .Z(n4435) );
  IV U8407 ( .A(n7203), .Z(n7206) );
  XNOR U8408 ( .A(n4436), .B(n7203), .Z(n7205) );
  NAND U8409 ( .A(n7208), .B(nreg[849]), .Z(n4436) );
  NAND U8410 ( .A(n6107), .B(nreg[849]), .Z(n7208) );
  XOR U8411 ( .A(n7209), .B(n7210), .Z(n7203) );
  ANDN U8412 ( .A(n7211), .B(n4437), .Z(n7210) );
  XOR U8413 ( .A(n7212), .B(n7213), .Z(n4437) );
  IV U8414 ( .A(n7209), .Z(n7212) );
  XNOR U8415 ( .A(n4438), .B(n7209), .Z(n7211) );
  NAND U8416 ( .A(n7214), .B(nreg[848]), .Z(n4438) );
  NAND U8417 ( .A(n6107), .B(nreg[848]), .Z(n7214) );
  XOR U8418 ( .A(n7215), .B(n7216), .Z(n7209) );
  ANDN U8419 ( .A(n7217), .B(n4439), .Z(n7216) );
  XOR U8420 ( .A(n7218), .B(n7219), .Z(n4439) );
  IV U8421 ( .A(n7215), .Z(n7218) );
  XNOR U8422 ( .A(n4440), .B(n7215), .Z(n7217) );
  NAND U8423 ( .A(n7220), .B(nreg[847]), .Z(n4440) );
  NAND U8424 ( .A(n6107), .B(nreg[847]), .Z(n7220) );
  XOR U8425 ( .A(n7221), .B(n7222), .Z(n7215) );
  ANDN U8426 ( .A(n7223), .B(n4443), .Z(n7222) );
  XOR U8427 ( .A(n7224), .B(n7225), .Z(n4443) );
  IV U8428 ( .A(n7221), .Z(n7224) );
  XNOR U8429 ( .A(n4444), .B(n7221), .Z(n7223) );
  NAND U8430 ( .A(n7226), .B(nreg[846]), .Z(n4444) );
  NAND U8431 ( .A(n6107), .B(nreg[846]), .Z(n7226) );
  XOR U8432 ( .A(n7227), .B(n7228), .Z(n7221) );
  ANDN U8433 ( .A(n7229), .B(n4445), .Z(n7228) );
  XOR U8434 ( .A(n7230), .B(n7231), .Z(n4445) );
  IV U8435 ( .A(n7227), .Z(n7230) );
  XNOR U8436 ( .A(n4446), .B(n7227), .Z(n7229) );
  NAND U8437 ( .A(n7232), .B(nreg[845]), .Z(n4446) );
  NAND U8438 ( .A(n6107), .B(nreg[845]), .Z(n7232) );
  XOR U8439 ( .A(n7233), .B(n7234), .Z(n7227) );
  ANDN U8440 ( .A(n7235), .B(n4447), .Z(n7234) );
  XOR U8441 ( .A(n7236), .B(n7237), .Z(n4447) );
  IV U8442 ( .A(n7233), .Z(n7236) );
  XNOR U8443 ( .A(n4448), .B(n7233), .Z(n7235) );
  NAND U8444 ( .A(n7238), .B(nreg[844]), .Z(n4448) );
  NAND U8445 ( .A(n6107), .B(nreg[844]), .Z(n7238) );
  XOR U8446 ( .A(n7239), .B(n7240), .Z(n7233) );
  ANDN U8447 ( .A(n7241), .B(n4449), .Z(n7240) );
  XOR U8448 ( .A(n7242), .B(n7243), .Z(n4449) );
  IV U8449 ( .A(n7239), .Z(n7242) );
  XNOR U8450 ( .A(n4450), .B(n7239), .Z(n7241) );
  NAND U8451 ( .A(n7244), .B(nreg[843]), .Z(n4450) );
  NAND U8452 ( .A(n6107), .B(nreg[843]), .Z(n7244) );
  XOR U8453 ( .A(n7245), .B(n7246), .Z(n7239) );
  ANDN U8454 ( .A(n7247), .B(n4451), .Z(n7246) );
  XOR U8455 ( .A(n7248), .B(n7249), .Z(n4451) );
  IV U8456 ( .A(n7245), .Z(n7248) );
  XNOR U8457 ( .A(n4452), .B(n7245), .Z(n7247) );
  NAND U8458 ( .A(n7250), .B(nreg[842]), .Z(n4452) );
  NAND U8459 ( .A(n6107), .B(nreg[842]), .Z(n7250) );
  XOR U8460 ( .A(n7251), .B(n7252), .Z(n7245) );
  ANDN U8461 ( .A(n7253), .B(n4453), .Z(n7252) );
  XOR U8462 ( .A(n7254), .B(n7255), .Z(n4453) );
  IV U8463 ( .A(n7251), .Z(n7254) );
  XNOR U8464 ( .A(n4454), .B(n7251), .Z(n7253) );
  NAND U8465 ( .A(n7256), .B(nreg[841]), .Z(n4454) );
  NAND U8466 ( .A(n6107), .B(nreg[841]), .Z(n7256) );
  XOR U8467 ( .A(n7257), .B(n7258), .Z(n7251) );
  ANDN U8468 ( .A(n7259), .B(n4455), .Z(n7258) );
  XOR U8469 ( .A(n7260), .B(n7261), .Z(n4455) );
  IV U8470 ( .A(n7257), .Z(n7260) );
  XNOR U8471 ( .A(n4456), .B(n7257), .Z(n7259) );
  NAND U8472 ( .A(n7262), .B(nreg[840]), .Z(n4456) );
  NAND U8473 ( .A(n6107), .B(nreg[840]), .Z(n7262) );
  XOR U8474 ( .A(n7263), .B(n7264), .Z(n7257) );
  ANDN U8475 ( .A(n7265), .B(n4457), .Z(n7264) );
  XOR U8476 ( .A(n7266), .B(n7267), .Z(n4457) );
  IV U8477 ( .A(n7263), .Z(n7266) );
  XNOR U8478 ( .A(n4458), .B(n7263), .Z(n7265) );
  NAND U8479 ( .A(n7268), .B(nreg[839]), .Z(n4458) );
  NAND U8480 ( .A(n6107), .B(nreg[839]), .Z(n7268) );
  XOR U8481 ( .A(n7269), .B(n7270), .Z(n7263) );
  ANDN U8482 ( .A(n7271), .B(n4459), .Z(n7270) );
  XOR U8483 ( .A(n7272), .B(n7273), .Z(n4459) );
  IV U8484 ( .A(n7269), .Z(n7272) );
  XNOR U8485 ( .A(n4460), .B(n7269), .Z(n7271) );
  NAND U8486 ( .A(n7274), .B(nreg[838]), .Z(n4460) );
  NAND U8487 ( .A(n6107), .B(nreg[838]), .Z(n7274) );
  XOR U8488 ( .A(n7275), .B(n7276), .Z(n7269) );
  ANDN U8489 ( .A(n7277), .B(n4461), .Z(n7276) );
  XOR U8490 ( .A(n7278), .B(n7279), .Z(n4461) );
  IV U8491 ( .A(n7275), .Z(n7278) );
  XNOR U8492 ( .A(n4462), .B(n7275), .Z(n7277) );
  NAND U8493 ( .A(n7280), .B(nreg[837]), .Z(n4462) );
  NAND U8494 ( .A(n6107), .B(nreg[837]), .Z(n7280) );
  XOR U8495 ( .A(n7281), .B(n7282), .Z(n7275) );
  ANDN U8496 ( .A(n7283), .B(n4465), .Z(n7282) );
  XOR U8497 ( .A(n7284), .B(n7285), .Z(n4465) );
  IV U8498 ( .A(n7281), .Z(n7284) );
  XNOR U8499 ( .A(n4466), .B(n7281), .Z(n7283) );
  NAND U8500 ( .A(n7286), .B(nreg[836]), .Z(n4466) );
  NAND U8501 ( .A(n6107), .B(nreg[836]), .Z(n7286) );
  XOR U8502 ( .A(n7287), .B(n7288), .Z(n7281) );
  ANDN U8503 ( .A(n7289), .B(n4467), .Z(n7288) );
  XOR U8504 ( .A(n7290), .B(n7291), .Z(n4467) );
  IV U8505 ( .A(n7287), .Z(n7290) );
  XNOR U8506 ( .A(n4468), .B(n7287), .Z(n7289) );
  NAND U8507 ( .A(n7292), .B(nreg[835]), .Z(n4468) );
  NAND U8508 ( .A(n6107), .B(nreg[835]), .Z(n7292) );
  XOR U8509 ( .A(n7293), .B(n7294), .Z(n7287) );
  ANDN U8510 ( .A(n7295), .B(n4469), .Z(n7294) );
  XOR U8511 ( .A(n7296), .B(n7297), .Z(n4469) );
  IV U8512 ( .A(n7293), .Z(n7296) );
  XNOR U8513 ( .A(n4470), .B(n7293), .Z(n7295) );
  NAND U8514 ( .A(n7298), .B(nreg[834]), .Z(n4470) );
  NAND U8515 ( .A(n6107), .B(nreg[834]), .Z(n7298) );
  XOR U8516 ( .A(n7299), .B(n7300), .Z(n7293) );
  ANDN U8517 ( .A(n7301), .B(n4471), .Z(n7300) );
  XOR U8518 ( .A(n7302), .B(n7303), .Z(n4471) );
  IV U8519 ( .A(n7299), .Z(n7302) );
  XNOR U8520 ( .A(n4472), .B(n7299), .Z(n7301) );
  NAND U8521 ( .A(n7304), .B(nreg[833]), .Z(n4472) );
  NAND U8522 ( .A(n6107), .B(nreg[833]), .Z(n7304) );
  XOR U8523 ( .A(n7305), .B(n7306), .Z(n7299) );
  ANDN U8524 ( .A(n7307), .B(n4473), .Z(n7306) );
  XOR U8525 ( .A(n7308), .B(n7309), .Z(n4473) );
  IV U8526 ( .A(n7305), .Z(n7308) );
  XNOR U8527 ( .A(n4474), .B(n7305), .Z(n7307) );
  NAND U8528 ( .A(n7310), .B(nreg[832]), .Z(n4474) );
  NAND U8529 ( .A(n6107), .B(nreg[832]), .Z(n7310) );
  XOR U8530 ( .A(n7311), .B(n7312), .Z(n7305) );
  ANDN U8531 ( .A(n7313), .B(n4475), .Z(n7312) );
  XOR U8532 ( .A(n7314), .B(n7315), .Z(n4475) );
  IV U8533 ( .A(n7311), .Z(n7314) );
  XNOR U8534 ( .A(n4476), .B(n7311), .Z(n7313) );
  NAND U8535 ( .A(n7316), .B(nreg[831]), .Z(n4476) );
  NAND U8536 ( .A(n6107), .B(nreg[831]), .Z(n7316) );
  XOR U8537 ( .A(n7317), .B(n7318), .Z(n7311) );
  ANDN U8538 ( .A(n7319), .B(n4477), .Z(n7318) );
  XOR U8539 ( .A(n7320), .B(n7321), .Z(n4477) );
  IV U8540 ( .A(n7317), .Z(n7320) );
  XNOR U8541 ( .A(n4478), .B(n7317), .Z(n7319) );
  NAND U8542 ( .A(n7322), .B(nreg[830]), .Z(n4478) );
  NAND U8543 ( .A(n6107), .B(nreg[830]), .Z(n7322) );
  XOR U8544 ( .A(n7323), .B(n7324), .Z(n7317) );
  ANDN U8545 ( .A(n7325), .B(n4479), .Z(n7324) );
  XOR U8546 ( .A(n7326), .B(n7327), .Z(n4479) );
  IV U8547 ( .A(n7323), .Z(n7326) );
  XNOR U8548 ( .A(n4480), .B(n7323), .Z(n7325) );
  NAND U8549 ( .A(n7328), .B(nreg[829]), .Z(n4480) );
  NAND U8550 ( .A(n6107), .B(nreg[829]), .Z(n7328) );
  XOR U8551 ( .A(n7329), .B(n7330), .Z(n7323) );
  ANDN U8552 ( .A(n7331), .B(n4481), .Z(n7330) );
  XOR U8553 ( .A(n7332), .B(n7333), .Z(n4481) );
  IV U8554 ( .A(n7329), .Z(n7332) );
  XNOR U8555 ( .A(n4482), .B(n7329), .Z(n7331) );
  NAND U8556 ( .A(n7334), .B(nreg[828]), .Z(n4482) );
  NAND U8557 ( .A(n6107), .B(nreg[828]), .Z(n7334) );
  XOR U8558 ( .A(n7335), .B(n7336), .Z(n7329) );
  ANDN U8559 ( .A(n7337), .B(n4483), .Z(n7336) );
  XOR U8560 ( .A(n7338), .B(n7339), .Z(n4483) );
  IV U8561 ( .A(n7335), .Z(n7338) );
  XNOR U8562 ( .A(n4484), .B(n7335), .Z(n7337) );
  NAND U8563 ( .A(n7340), .B(nreg[827]), .Z(n4484) );
  NAND U8564 ( .A(n6107), .B(nreg[827]), .Z(n7340) );
  XOR U8565 ( .A(n7341), .B(n7342), .Z(n7335) );
  ANDN U8566 ( .A(n7343), .B(n4487), .Z(n7342) );
  XOR U8567 ( .A(n7344), .B(n7345), .Z(n4487) );
  IV U8568 ( .A(n7341), .Z(n7344) );
  XNOR U8569 ( .A(n4488), .B(n7341), .Z(n7343) );
  NAND U8570 ( .A(n7346), .B(nreg[826]), .Z(n4488) );
  NAND U8571 ( .A(n6107), .B(nreg[826]), .Z(n7346) );
  XOR U8572 ( .A(n7347), .B(n7348), .Z(n7341) );
  ANDN U8573 ( .A(n7349), .B(n4489), .Z(n7348) );
  XOR U8574 ( .A(n7350), .B(n7351), .Z(n4489) );
  IV U8575 ( .A(n7347), .Z(n7350) );
  XNOR U8576 ( .A(n4490), .B(n7347), .Z(n7349) );
  NAND U8577 ( .A(n7352), .B(nreg[825]), .Z(n4490) );
  NAND U8578 ( .A(n6107), .B(nreg[825]), .Z(n7352) );
  XOR U8579 ( .A(n7353), .B(n7354), .Z(n7347) );
  ANDN U8580 ( .A(n7355), .B(n4491), .Z(n7354) );
  XOR U8581 ( .A(n7356), .B(n7357), .Z(n4491) );
  IV U8582 ( .A(n7353), .Z(n7356) );
  XNOR U8583 ( .A(n4492), .B(n7353), .Z(n7355) );
  NAND U8584 ( .A(n7358), .B(nreg[824]), .Z(n4492) );
  NAND U8585 ( .A(n6107), .B(nreg[824]), .Z(n7358) );
  XOR U8586 ( .A(n7359), .B(n7360), .Z(n7353) );
  ANDN U8587 ( .A(n7361), .B(n4493), .Z(n7360) );
  XOR U8588 ( .A(n7362), .B(n7363), .Z(n4493) );
  IV U8589 ( .A(n7359), .Z(n7362) );
  XNOR U8590 ( .A(n4494), .B(n7359), .Z(n7361) );
  NAND U8591 ( .A(n7364), .B(nreg[823]), .Z(n4494) );
  NAND U8592 ( .A(n6107), .B(nreg[823]), .Z(n7364) );
  XOR U8593 ( .A(n7365), .B(n7366), .Z(n7359) );
  ANDN U8594 ( .A(n7367), .B(n4495), .Z(n7366) );
  XOR U8595 ( .A(n7368), .B(n7369), .Z(n4495) );
  IV U8596 ( .A(n7365), .Z(n7368) );
  XNOR U8597 ( .A(n4496), .B(n7365), .Z(n7367) );
  NAND U8598 ( .A(n7370), .B(nreg[822]), .Z(n4496) );
  NAND U8599 ( .A(n6107), .B(nreg[822]), .Z(n7370) );
  XOR U8600 ( .A(n7371), .B(n7372), .Z(n7365) );
  ANDN U8601 ( .A(n7373), .B(n4497), .Z(n7372) );
  XOR U8602 ( .A(n7374), .B(n7375), .Z(n4497) );
  IV U8603 ( .A(n7371), .Z(n7374) );
  XNOR U8604 ( .A(n4498), .B(n7371), .Z(n7373) );
  NAND U8605 ( .A(n7376), .B(nreg[821]), .Z(n4498) );
  NAND U8606 ( .A(n6107), .B(nreg[821]), .Z(n7376) );
  XOR U8607 ( .A(n7377), .B(n7378), .Z(n7371) );
  ANDN U8608 ( .A(n7379), .B(n4499), .Z(n7378) );
  XOR U8609 ( .A(n7380), .B(n7381), .Z(n4499) );
  IV U8610 ( .A(n7377), .Z(n7380) );
  XNOR U8611 ( .A(n4500), .B(n7377), .Z(n7379) );
  NAND U8612 ( .A(n7382), .B(nreg[820]), .Z(n4500) );
  NAND U8613 ( .A(n6107), .B(nreg[820]), .Z(n7382) );
  XOR U8614 ( .A(n7383), .B(n7384), .Z(n7377) );
  ANDN U8615 ( .A(n7385), .B(n4501), .Z(n7384) );
  XOR U8616 ( .A(n7386), .B(n7387), .Z(n4501) );
  IV U8617 ( .A(n7383), .Z(n7386) );
  XNOR U8618 ( .A(n4502), .B(n7383), .Z(n7385) );
  NAND U8619 ( .A(n7388), .B(nreg[819]), .Z(n4502) );
  NAND U8620 ( .A(n6107), .B(nreg[819]), .Z(n7388) );
  XOR U8621 ( .A(n7389), .B(n7390), .Z(n7383) );
  ANDN U8622 ( .A(n7391), .B(n4503), .Z(n7390) );
  XOR U8623 ( .A(n7392), .B(n7393), .Z(n4503) );
  IV U8624 ( .A(n7389), .Z(n7392) );
  XNOR U8625 ( .A(n4504), .B(n7389), .Z(n7391) );
  NAND U8626 ( .A(n7394), .B(nreg[818]), .Z(n4504) );
  NAND U8627 ( .A(n6107), .B(nreg[818]), .Z(n7394) );
  XOR U8628 ( .A(n7395), .B(n7396), .Z(n7389) );
  ANDN U8629 ( .A(n7397), .B(n4505), .Z(n7396) );
  XOR U8630 ( .A(n7398), .B(n7399), .Z(n4505) );
  IV U8631 ( .A(n7395), .Z(n7398) );
  XNOR U8632 ( .A(n4506), .B(n7395), .Z(n7397) );
  NAND U8633 ( .A(n7400), .B(nreg[817]), .Z(n4506) );
  NAND U8634 ( .A(n6107), .B(nreg[817]), .Z(n7400) );
  XOR U8635 ( .A(n7401), .B(n7402), .Z(n7395) );
  ANDN U8636 ( .A(n7403), .B(n4509), .Z(n7402) );
  XOR U8637 ( .A(n7404), .B(n7405), .Z(n4509) );
  IV U8638 ( .A(n7401), .Z(n7404) );
  XNOR U8639 ( .A(n4510), .B(n7401), .Z(n7403) );
  NAND U8640 ( .A(n7406), .B(nreg[816]), .Z(n4510) );
  NAND U8641 ( .A(n6107), .B(nreg[816]), .Z(n7406) );
  XOR U8642 ( .A(n7407), .B(n7408), .Z(n7401) );
  ANDN U8643 ( .A(n7409), .B(n4511), .Z(n7408) );
  XOR U8644 ( .A(n7410), .B(n7411), .Z(n4511) );
  IV U8645 ( .A(n7407), .Z(n7410) );
  XNOR U8646 ( .A(n4512), .B(n7407), .Z(n7409) );
  NAND U8647 ( .A(n7412), .B(nreg[815]), .Z(n4512) );
  NAND U8648 ( .A(n6107), .B(nreg[815]), .Z(n7412) );
  XOR U8649 ( .A(n7413), .B(n7414), .Z(n7407) );
  ANDN U8650 ( .A(n7415), .B(n4513), .Z(n7414) );
  XOR U8651 ( .A(n7416), .B(n7417), .Z(n4513) );
  IV U8652 ( .A(n7413), .Z(n7416) );
  XNOR U8653 ( .A(n4514), .B(n7413), .Z(n7415) );
  NAND U8654 ( .A(n7418), .B(nreg[814]), .Z(n4514) );
  NAND U8655 ( .A(n6107), .B(nreg[814]), .Z(n7418) );
  XOR U8656 ( .A(n7419), .B(n7420), .Z(n7413) );
  ANDN U8657 ( .A(n7421), .B(n4515), .Z(n7420) );
  XOR U8658 ( .A(n7422), .B(n7423), .Z(n4515) );
  IV U8659 ( .A(n7419), .Z(n7422) );
  XNOR U8660 ( .A(n4516), .B(n7419), .Z(n7421) );
  NAND U8661 ( .A(n7424), .B(nreg[813]), .Z(n4516) );
  NAND U8662 ( .A(n6107), .B(nreg[813]), .Z(n7424) );
  XOR U8663 ( .A(n7425), .B(n7426), .Z(n7419) );
  ANDN U8664 ( .A(n7427), .B(n4517), .Z(n7426) );
  XOR U8665 ( .A(n7428), .B(n7429), .Z(n4517) );
  IV U8666 ( .A(n7425), .Z(n7428) );
  XNOR U8667 ( .A(n4518), .B(n7425), .Z(n7427) );
  NAND U8668 ( .A(n7430), .B(nreg[812]), .Z(n4518) );
  NAND U8669 ( .A(n6107), .B(nreg[812]), .Z(n7430) );
  XOR U8670 ( .A(n7431), .B(n7432), .Z(n7425) );
  ANDN U8671 ( .A(n7433), .B(n4519), .Z(n7432) );
  XOR U8672 ( .A(n7434), .B(n7435), .Z(n4519) );
  IV U8673 ( .A(n7431), .Z(n7434) );
  XNOR U8674 ( .A(n4520), .B(n7431), .Z(n7433) );
  NAND U8675 ( .A(n7436), .B(nreg[811]), .Z(n4520) );
  NAND U8676 ( .A(n6107), .B(nreg[811]), .Z(n7436) );
  XOR U8677 ( .A(n7437), .B(n7438), .Z(n7431) );
  ANDN U8678 ( .A(n7439), .B(n4521), .Z(n7438) );
  XOR U8679 ( .A(n7440), .B(n7441), .Z(n4521) );
  IV U8680 ( .A(n7437), .Z(n7440) );
  XNOR U8681 ( .A(n4522), .B(n7437), .Z(n7439) );
  NAND U8682 ( .A(n7442), .B(nreg[810]), .Z(n4522) );
  NAND U8683 ( .A(n6107), .B(nreg[810]), .Z(n7442) );
  XOR U8684 ( .A(n7443), .B(n7444), .Z(n7437) );
  ANDN U8685 ( .A(n7445), .B(n4523), .Z(n7444) );
  XOR U8686 ( .A(n7446), .B(n7447), .Z(n4523) );
  IV U8687 ( .A(n7443), .Z(n7446) );
  XNOR U8688 ( .A(n4524), .B(n7443), .Z(n7445) );
  NAND U8689 ( .A(n7448), .B(nreg[809]), .Z(n4524) );
  NAND U8690 ( .A(n6107), .B(nreg[809]), .Z(n7448) );
  XOR U8691 ( .A(n7449), .B(n7450), .Z(n7443) );
  ANDN U8692 ( .A(n7451), .B(n4525), .Z(n7450) );
  XOR U8693 ( .A(n7452), .B(n7453), .Z(n4525) );
  IV U8694 ( .A(n7449), .Z(n7452) );
  XNOR U8695 ( .A(n4526), .B(n7449), .Z(n7451) );
  NAND U8696 ( .A(n7454), .B(nreg[808]), .Z(n4526) );
  NAND U8697 ( .A(n6107), .B(nreg[808]), .Z(n7454) );
  XOR U8698 ( .A(n7455), .B(n7456), .Z(n7449) );
  ANDN U8699 ( .A(n7457), .B(n4527), .Z(n7456) );
  XOR U8700 ( .A(n7458), .B(n7459), .Z(n4527) );
  IV U8701 ( .A(n7455), .Z(n7458) );
  XNOR U8702 ( .A(n4528), .B(n7455), .Z(n7457) );
  NAND U8703 ( .A(n7460), .B(nreg[807]), .Z(n4528) );
  NAND U8704 ( .A(n6107), .B(nreg[807]), .Z(n7460) );
  XOR U8705 ( .A(n7461), .B(n7462), .Z(n7455) );
  ANDN U8706 ( .A(n7463), .B(n4531), .Z(n7462) );
  XOR U8707 ( .A(n7464), .B(n7465), .Z(n4531) );
  IV U8708 ( .A(n7461), .Z(n7464) );
  XNOR U8709 ( .A(n4532), .B(n7461), .Z(n7463) );
  NAND U8710 ( .A(n7466), .B(nreg[806]), .Z(n4532) );
  NAND U8711 ( .A(n6107), .B(nreg[806]), .Z(n7466) );
  XOR U8712 ( .A(n7467), .B(n7468), .Z(n7461) );
  ANDN U8713 ( .A(n7469), .B(n4533), .Z(n7468) );
  XOR U8714 ( .A(n7470), .B(n7471), .Z(n4533) );
  IV U8715 ( .A(n7467), .Z(n7470) );
  XNOR U8716 ( .A(n4534), .B(n7467), .Z(n7469) );
  NAND U8717 ( .A(n7472), .B(nreg[805]), .Z(n4534) );
  NAND U8718 ( .A(n6107), .B(nreg[805]), .Z(n7472) );
  XOR U8719 ( .A(n7473), .B(n7474), .Z(n7467) );
  ANDN U8720 ( .A(n7475), .B(n4535), .Z(n7474) );
  XOR U8721 ( .A(n7476), .B(n7477), .Z(n4535) );
  IV U8722 ( .A(n7473), .Z(n7476) );
  XNOR U8723 ( .A(n4536), .B(n7473), .Z(n7475) );
  NAND U8724 ( .A(n7478), .B(nreg[804]), .Z(n4536) );
  NAND U8725 ( .A(n6107), .B(nreg[804]), .Z(n7478) );
  XOR U8726 ( .A(n7479), .B(n7480), .Z(n7473) );
  ANDN U8727 ( .A(n7481), .B(n4537), .Z(n7480) );
  XOR U8728 ( .A(n7482), .B(n7483), .Z(n4537) );
  IV U8729 ( .A(n7479), .Z(n7482) );
  XNOR U8730 ( .A(n4538), .B(n7479), .Z(n7481) );
  NAND U8731 ( .A(n7484), .B(nreg[803]), .Z(n4538) );
  NAND U8732 ( .A(n6107), .B(nreg[803]), .Z(n7484) );
  XOR U8733 ( .A(n7485), .B(n7486), .Z(n7479) );
  ANDN U8734 ( .A(n7487), .B(n4539), .Z(n7486) );
  XOR U8735 ( .A(n7488), .B(n7489), .Z(n4539) );
  IV U8736 ( .A(n7485), .Z(n7488) );
  XNOR U8737 ( .A(n4540), .B(n7485), .Z(n7487) );
  NAND U8738 ( .A(n7490), .B(nreg[802]), .Z(n4540) );
  NAND U8739 ( .A(n6107), .B(nreg[802]), .Z(n7490) );
  XOR U8740 ( .A(n7491), .B(n7492), .Z(n7485) );
  ANDN U8741 ( .A(n7493), .B(n4541), .Z(n7492) );
  XOR U8742 ( .A(n7494), .B(n7495), .Z(n4541) );
  IV U8743 ( .A(n7491), .Z(n7494) );
  XNOR U8744 ( .A(n4542), .B(n7491), .Z(n7493) );
  NAND U8745 ( .A(n7496), .B(nreg[801]), .Z(n4542) );
  NAND U8746 ( .A(n6107), .B(nreg[801]), .Z(n7496) );
  XOR U8747 ( .A(n7497), .B(n7498), .Z(n7491) );
  ANDN U8748 ( .A(n7499), .B(n4543), .Z(n7498) );
  XOR U8749 ( .A(n7500), .B(n7501), .Z(n4543) );
  IV U8750 ( .A(n7497), .Z(n7500) );
  XNOR U8751 ( .A(n4544), .B(n7497), .Z(n7499) );
  NAND U8752 ( .A(n7502), .B(nreg[800]), .Z(n4544) );
  NAND U8753 ( .A(n6107), .B(nreg[800]), .Z(n7502) );
  XOR U8754 ( .A(n7503), .B(n7504), .Z(n7497) );
  ANDN U8755 ( .A(n7505), .B(n4545), .Z(n7504) );
  XOR U8756 ( .A(n7506), .B(n7507), .Z(n4545) );
  IV U8757 ( .A(n7503), .Z(n7506) );
  XNOR U8758 ( .A(n4546), .B(n7503), .Z(n7505) );
  NAND U8759 ( .A(n7508), .B(nreg[799]), .Z(n4546) );
  NAND U8760 ( .A(n6107), .B(nreg[799]), .Z(n7508) );
  XOR U8761 ( .A(n7509), .B(n7510), .Z(n7503) );
  ANDN U8762 ( .A(n7511), .B(n4547), .Z(n7510) );
  XOR U8763 ( .A(n7512), .B(n7513), .Z(n4547) );
  IV U8764 ( .A(n7509), .Z(n7512) );
  XNOR U8765 ( .A(n4548), .B(n7509), .Z(n7511) );
  NAND U8766 ( .A(n7514), .B(nreg[798]), .Z(n4548) );
  NAND U8767 ( .A(n6107), .B(nreg[798]), .Z(n7514) );
  XOR U8768 ( .A(n7515), .B(n7516), .Z(n7509) );
  ANDN U8769 ( .A(n7517), .B(n4549), .Z(n7516) );
  XOR U8770 ( .A(n7518), .B(n7519), .Z(n4549) );
  IV U8771 ( .A(n7515), .Z(n7518) );
  XNOR U8772 ( .A(n4550), .B(n7515), .Z(n7517) );
  NAND U8773 ( .A(n7520), .B(nreg[797]), .Z(n4550) );
  NAND U8774 ( .A(n6107), .B(nreg[797]), .Z(n7520) );
  XOR U8775 ( .A(n7521), .B(n7522), .Z(n7515) );
  ANDN U8776 ( .A(n7523), .B(n4555), .Z(n7522) );
  XOR U8777 ( .A(n7524), .B(n7525), .Z(n4555) );
  IV U8778 ( .A(n7521), .Z(n7524) );
  XNOR U8779 ( .A(n4556), .B(n7521), .Z(n7523) );
  NAND U8780 ( .A(n7526), .B(nreg[796]), .Z(n4556) );
  NAND U8781 ( .A(n6107), .B(nreg[796]), .Z(n7526) );
  XOR U8782 ( .A(n7527), .B(n7528), .Z(n7521) );
  ANDN U8783 ( .A(n7529), .B(n4557), .Z(n7528) );
  XOR U8784 ( .A(n7530), .B(n7531), .Z(n4557) );
  IV U8785 ( .A(n7527), .Z(n7530) );
  XNOR U8786 ( .A(n4558), .B(n7527), .Z(n7529) );
  NAND U8787 ( .A(n7532), .B(nreg[795]), .Z(n4558) );
  NAND U8788 ( .A(n6107), .B(nreg[795]), .Z(n7532) );
  XOR U8789 ( .A(n7533), .B(n7534), .Z(n7527) );
  ANDN U8790 ( .A(n7535), .B(n4559), .Z(n7534) );
  XOR U8791 ( .A(n7536), .B(n7537), .Z(n4559) );
  IV U8792 ( .A(n7533), .Z(n7536) );
  XNOR U8793 ( .A(n4560), .B(n7533), .Z(n7535) );
  NAND U8794 ( .A(n7538), .B(nreg[794]), .Z(n4560) );
  NAND U8795 ( .A(n6107), .B(nreg[794]), .Z(n7538) );
  XOR U8796 ( .A(n7539), .B(n7540), .Z(n7533) );
  ANDN U8797 ( .A(n7541), .B(n4561), .Z(n7540) );
  XOR U8798 ( .A(n7542), .B(n7543), .Z(n4561) );
  IV U8799 ( .A(n7539), .Z(n7542) );
  XNOR U8800 ( .A(n4562), .B(n7539), .Z(n7541) );
  NAND U8801 ( .A(n7544), .B(nreg[793]), .Z(n4562) );
  NAND U8802 ( .A(n6107), .B(nreg[793]), .Z(n7544) );
  XOR U8803 ( .A(n7545), .B(n7546), .Z(n7539) );
  ANDN U8804 ( .A(n7547), .B(n4563), .Z(n7546) );
  XOR U8805 ( .A(n7548), .B(n7549), .Z(n4563) );
  IV U8806 ( .A(n7545), .Z(n7548) );
  XNOR U8807 ( .A(n4564), .B(n7545), .Z(n7547) );
  NAND U8808 ( .A(n7550), .B(nreg[792]), .Z(n4564) );
  NAND U8809 ( .A(n6107), .B(nreg[792]), .Z(n7550) );
  XOR U8810 ( .A(n7551), .B(n7552), .Z(n7545) );
  ANDN U8811 ( .A(n7553), .B(n4565), .Z(n7552) );
  XOR U8812 ( .A(n7554), .B(n7555), .Z(n4565) );
  IV U8813 ( .A(n7551), .Z(n7554) );
  XNOR U8814 ( .A(n4566), .B(n7551), .Z(n7553) );
  NAND U8815 ( .A(n7556), .B(nreg[791]), .Z(n4566) );
  NAND U8816 ( .A(n6107), .B(nreg[791]), .Z(n7556) );
  XOR U8817 ( .A(n7557), .B(n7558), .Z(n7551) );
  ANDN U8818 ( .A(n7559), .B(n4567), .Z(n7558) );
  XOR U8819 ( .A(n7560), .B(n7561), .Z(n4567) );
  IV U8820 ( .A(n7557), .Z(n7560) );
  XNOR U8821 ( .A(n4568), .B(n7557), .Z(n7559) );
  NAND U8822 ( .A(n7562), .B(nreg[790]), .Z(n4568) );
  NAND U8823 ( .A(n6107), .B(nreg[790]), .Z(n7562) );
  XOR U8824 ( .A(n7563), .B(n7564), .Z(n7557) );
  ANDN U8825 ( .A(n7565), .B(n4569), .Z(n7564) );
  XOR U8826 ( .A(n7566), .B(n7567), .Z(n4569) );
  IV U8827 ( .A(n7563), .Z(n7566) );
  XNOR U8828 ( .A(n4570), .B(n7563), .Z(n7565) );
  NAND U8829 ( .A(n7568), .B(nreg[789]), .Z(n4570) );
  NAND U8830 ( .A(n6107), .B(nreg[789]), .Z(n7568) );
  XOR U8831 ( .A(n7569), .B(n7570), .Z(n7563) );
  ANDN U8832 ( .A(n7571), .B(n4571), .Z(n7570) );
  XOR U8833 ( .A(n7572), .B(n7573), .Z(n4571) );
  IV U8834 ( .A(n7569), .Z(n7572) );
  XNOR U8835 ( .A(n4572), .B(n7569), .Z(n7571) );
  NAND U8836 ( .A(n7574), .B(nreg[788]), .Z(n4572) );
  NAND U8837 ( .A(n6107), .B(nreg[788]), .Z(n7574) );
  XOR U8838 ( .A(n7575), .B(n7576), .Z(n7569) );
  ANDN U8839 ( .A(n7577), .B(n4573), .Z(n7576) );
  XOR U8840 ( .A(n7578), .B(n7579), .Z(n4573) );
  IV U8841 ( .A(n7575), .Z(n7578) );
  XNOR U8842 ( .A(n4574), .B(n7575), .Z(n7577) );
  NAND U8843 ( .A(n7580), .B(nreg[787]), .Z(n4574) );
  NAND U8844 ( .A(n6107), .B(nreg[787]), .Z(n7580) );
  XOR U8845 ( .A(n7581), .B(n7582), .Z(n7575) );
  ANDN U8846 ( .A(n7583), .B(n4577), .Z(n7582) );
  XOR U8847 ( .A(n7584), .B(n7585), .Z(n4577) );
  IV U8848 ( .A(n7581), .Z(n7584) );
  XNOR U8849 ( .A(n4578), .B(n7581), .Z(n7583) );
  NAND U8850 ( .A(n7586), .B(nreg[786]), .Z(n4578) );
  NAND U8851 ( .A(n6107), .B(nreg[786]), .Z(n7586) );
  XOR U8852 ( .A(n7587), .B(n7588), .Z(n7581) );
  ANDN U8853 ( .A(n7589), .B(n4579), .Z(n7588) );
  XOR U8854 ( .A(n7590), .B(n7591), .Z(n4579) );
  IV U8855 ( .A(n7587), .Z(n7590) );
  XNOR U8856 ( .A(n4580), .B(n7587), .Z(n7589) );
  NAND U8857 ( .A(n7592), .B(nreg[785]), .Z(n4580) );
  NAND U8858 ( .A(n6107), .B(nreg[785]), .Z(n7592) );
  XOR U8859 ( .A(n7593), .B(n7594), .Z(n7587) );
  ANDN U8860 ( .A(n7595), .B(n4581), .Z(n7594) );
  XOR U8861 ( .A(n7596), .B(n7597), .Z(n4581) );
  IV U8862 ( .A(n7593), .Z(n7596) );
  XNOR U8863 ( .A(n4582), .B(n7593), .Z(n7595) );
  NAND U8864 ( .A(n7598), .B(nreg[784]), .Z(n4582) );
  NAND U8865 ( .A(n6107), .B(nreg[784]), .Z(n7598) );
  XOR U8866 ( .A(n7599), .B(n7600), .Z(n7593) );
  ANDN U8867 ( .A(n7601), .B(n4583), .Z(n7600) );
  XOR U8868 ( .A(n7602), .B(n7603), .Z(n4583) );
  IV U8869 ( .A(n7599), .Z(n7602) );
  XNOR U8870 ( .A(n4584), .B(n7599), .Z(n7601) );
  NAND U8871 ( .A(n7604), .B(nreg[783]), .Z(n4584) );
  NAND U8872 ( .A(n6107), .B(nreg[783]), .Z(n7604) );
  XOR U8873 ( .A(n7605), .B(n7606), .Z(n7599) );
  ANDN U8874 ( .A(n7607), .B(n4585), .Z(n7606) );
  XOR U8875 ( .A(n7608), .B(n7609), .Z(n4585) );
  IV U8876 ( .A(n7605), .Z(n7608) );
  XNOR U8877 ( .A(n4586), .B(n7605), .Z(n7607) );
  NAND U8878 ( .A(n7610), .B(nreg[782]), .Z(n4586) );
  NAND U8879 ( .A(n6107), .B(nreg[782]), .Z(n7610) );
  XOR U8880 ( .A(n7611), .B(n7612), .Z(n7605) );
  ANDN U8881 ( .A(n7613), .B(n4587), .Z(n7612) );
  XOR U8882 ( .A(n7614), .B(n7615), .Z(n4587) );
  IV U8883 ( .A(n7611), .Z(n7614) );
  XNOR U8884 ( .A(n4588), .B(n7611), .Z(n7613) );
  NAND U8885 ( .A(n7616), .B(nreg[781]), .Z(n4588) );
  NAND U8886 ( .A(n6107), .B(nreg[781]), .Z(n7616) );
  XOR U8887 ( .A(n7617), .B(n7618), .Z(n7611) );
  ANDN U8888 ( .A(n7619), .B(n4589), .Z(n7618) );
  XOR U8889 ( .A(n7620), .B(n7621), .Z(n4589) );
  IV U8890 ( .A(n7617), .Z(n7620) );
  XNOR U8891 ( .A(n4590), .B(n7617), .Z(n7619) );
  NAND U8892 ( .A(n7622), .B(nreg[780]), .Z(n4590) );
  NAND U8893 ( .A(n6107), .B(nreg[780]), .Z(n7622) );
  XOR U8894 ( .A(n7623), .B(n7624), .Z(n7617) );
  ANDN U8895 ( .A(n7625), .B(n4591), .Z(n7624) );
  XOR U8896 ( .A(n7626), .B(n7627), .Z(n4591) );
  IV U8897 ( .A(n7623), .Z(n7626) );
  XNOR U8898 ( .A(n4592), .B(n7623), .Z(n7625) );
  NAND U8899 ( .A(n7628), .B(nreg[779]), .Z(n4592) );
  NAND U8900 ( .A(n6107), .B(nreg[779]), .Z(n7628) );
  XOR U8901 ( .A(n7629), .B(n7630), .Z(n7623) );
  ANDN U8902 ( .A(n7631), .B(n4593), .Z(n7630) );
  XOR U8903 ( .A(n7632), .B(n7633), .Z(n4593) );
  IV U8904 ( .A(n7629), .Z(n7632) );
  XNOR U8905 ( .A(n4594), .B(n7629), .Z(n7631) );
  NAND U8906 ( .A(n7634), .B(nreg[778]), .Z(n4594) );
  NAND U8907 ( .A(n6107), .B(nreg[778]), .Z(n7634) );
  XOR U8908 ( .A(n7635), .B(n7636), .Z(n7629) );
  ANDN U8909 ( .A(n7637), .B(n4595), .Z(n7636) );
  XOR U8910 ( .A(n7638), .B(n7639), .Z(n4595) );
  IV U8911 ( .A(n7635), .Z(n7638) );
  XNOR U8912 ( .A(n4596), .B(n7635), .Z(n7637) );
  NAND U8913 ( .A(n7640), .B(nreg[777]), .Z(n4596) );
  NAND U8914 ( .A(n6107), .B(nreg[777]), .Z(n7640) );
  XOR U8915 ( .A(n7641), .B(n7642), .Z(n7635) );
  ANDN U8916 ( .A(n7643), .B(n4599), .Z(n7642) );
  XOR U8917 ( .A(n7644), .B(n7645), .Z(n4599) );
  IV U8918 ( .A(n7641), .Z(n7644) );
  XNOR U8919 ( .A(n4600), .B(n7641), .Z(n7643) );
  NAND U8920 ( .A(n7646), .B(nreg[776]), .Z(n4600) );
  NAND U8921 ( .A(n6107), .B(nreg[776]), .Z(n7646) );
  XOR U8922 ( .A(n7647), .B(n7648), .Z(n7641) );
  ANDN U8923 ( .A(n7649), .B(n4601), .Z(n7648) );
  XOR U8924 ( .A(n7650), .B(n7651), .Z(n4601) );
  IV U8925 ( .A(n7647), .Z(n7650) );
  XNOR U8926 ( .A(n4602), .B(n7647), .Z(n7649) );
  NAND U8927 ( .A(n7652), .B(nreg[775]), .Z(n4602) );
  NAND U8928 ( .A(n6107), .B(nreg[775]), .Z(n7652) );
  XOR U8929 ( .A(n7653), .B(n7654), .Z(n7647) );
  ANDN U8930 ( .A(n7655), .B(n4603), .Z(n7654) );
  XOR U8931 ( .A(n7656), .B(n7657), .Z(n4603) );
  IV U8932 ( .A(n7653), .Z(n7656) );
  XNOR U8933 ( .A(n4604), .B(n7653), .Z(n7655) );
  NAND U8934 ( .A(n7658), .B(nreg[774]), .Z(n4604) );
  NAND U8935 ( .A(n6107), .B(nreg[774]), .Z(n7658) );
  XOR U8936 ( .A(n7659), .B(n7660), .Z(n7653) );
  ANDN U8937 ( .A(n7661), .B(n4605), .Z(n7660) );
  XOR U8938 ( .A(n7662), .B(n7663), .Z(n4605) );
  IV U8939 ( .A(n7659), .Z(n7662) );
  XNOR U8940 ( .A(n4606), .B(n7659), .Z(n7661) );
  NAND U8941 ( .A(n7664), .B(nreg[773]), .Z(n4606) );
  NAND U8942 ( .A(n6107), .B(nreg[773]), .Z(n7664) );
  XOR U8943 ( .A(n7665), .B(n7666), .Z(n7659) );
  ANDN U8944 ( .A(n7667), .B(n4607), .Z(n7666) );
  XOR U8945 ( .A(n7668), .B(n7669), .Z(n4607) );
  IV U8946 ( .A(n7665), .Z(n7668) );
  XNOR U8947 ( .A(n4608), .B(n7665), .Z(n7667) );
  NAND U8948 ( .A(n7670), .B(nreg[772]), .Z(n4608) );
  NAND U8949 ( .A(n6107), .B(nreg[772]), .Z(n7670) );
  XOR U8950 ( .A(n7671), .B(n7672), .Z(n7665) );
  ANDN U8951 ( .A(n7673), .B(n4609), .Z(n7672) );
  XOR U8952 ( .A(n7674), .B(n7675), .Z(n4609) );
  IV U8953 ( .A(n7671), .Z(n7674) );
  XNOR U8954 ( .A(n4610), .B(n7671), .Z(n7673) );
  NAND U8955 ( .A(n7676), .B(nreg[771]), .Z(n4610) );
  NAND U8956 ( .A(n6107), .B(nreg[771]), .Z(n7676) );
  XOR U8957 ( .A(n7677), .B(n7678), .Z(n7671) );
  ANDN U8958 ( .A(n7679), .B(n4611), .Z(n7678) );
  XOR U8959 ( .A(n7680), .B(n7681), .Z(n4611) );
  IV U8960 ( .A(n7677), .Z(n7680) );
  XNOR U8961 ( .A(n4612), .B(n7677), .Z(n7679) );
  NAND U8962 ( .A(n7682), .B(nreg[770]), .Z(n4612) );
  NAND U8963 ( .A(n6107), .B(nreg[770]), .Z(n7682) );
  XOR U8964 ( .A(n7683), .B(n7684), .Z(n7677) );
  ANDN U8965 ( .A(n7685), .B(n4613), .Z(n7684) );
  XOR U8966 ( .A(n7686), .B(n7687), .Z(n4613) );
  IV U8967 ( .A(n7683), .Z(n7686) );
  XNOR U8968 ( .A(n4614), .B(n7683), .Z(n7685) );
  NAND U8969 ( .A(n7688), .B(nreg[769]), .Z(n4614) );
  NAND U8970 ( .A(n6107), .B(nreg[769]), .Z(n7688) );
  XOR U8971 ( .A(n7689), .B(n7690), .Z(n7683) );
  ANDN U8972 ( .A(n7691), .B(n4615), .Z(n7690) );
  XOR U8973 ( .A(n7692), .B(n7693), .Z(n4615) );
  IV U8974 ( .A(n7689), .Z(n7692) );
  XNOR U8975 ( .A(n4616), .B(n7689), .Z(n7691) );
  NAND U8976 ( .A(n7694), .B(nreg[768]), .Z(n4616) );
  NAND U8977 ( .A(n6107), .B(nreg[768]), .Z(n7694) );
  XOR U8978 ( .A(n7695), .B(n7696), .Z(n7689) );
  ANDN U8979 ( .A(n7697), .B(n4617), .Z(n7696) );
  XOR U8980 ( .A(n7698), .B(n7699), .Z(n4617) );
  IV U8981 ( .A(n7695), .Z(n7698) );
  XNOR U8982 ( .A(n4618), .B(n7695), .Z(n7697) );
  NAND U8983 ( .A(n7700), .B(nreg[767]), .Z(n4618) );
  NAND U8984 ( .A(n6107), .B(nreg[767]), .Z(n7700) );
  XOR U8985 ( .A(n7701), .B(n7702), .Z(n7695) );
  ANDN U8986 ( .A(n7703), .B(n4621), .Z(n7702) );
  XOR U8987 ( .A(n7704), .B(n7705), .Z(n4621) );
  IV U8988 ( .A(n7701), .Z(n7704) );
  XNOR U8989 ( .A(n4622), .B(n7701), .Z(n7703) );
  NAND U8990 ( .A(n7706), .B(nreg[766]), .Z(n4622) );
  NAND U8991 ( .A(n6107), .B(nreg[766]), .Z(n7706) );
  XOR U8992 ( .A(n7707), .B(n7708), .Z(n7701) );
  ANDN U8993 ( .A(n7709), .B(n4623), .Z(n7708) );
  XOR U8994 ( .A(n7710), .B(n7711), .Z(n4623) );
  IV U8995 ( .A(n7707), .Z(n7710) );
  XNOR U8996 ( .A(n4624), .B(n7707), .Z(n7709) );
  NAND U8997 ( .A(n7712), .B(nreg[765]), .Z(n4624) );
  NAND U8998 ( .A(n6107), .B(nreg[765]), .Z(n7712) );
  XOR U8999 ( .A(n7713), .B(n7714), .Z(n7707) );
  ANDN U9000 ( .A(n7715), .B(n4625), .Z(n7714) );
  XOR U9001 ( .A(n7716), .B(n7717), .Z(n4625) );
  IV U9002 ( .A(n7713), .Z(n7716) );
  XNOR U9003 ( .A(n4626), .B(n7713), .Z(n7715) );
  NAND U9004 ( .A(n7718), .B(nreg[764]), .Z(n4626) );
  NAND U9005 ( .A(n6107), .B(nreg[764]), .Z(n7718) );
  XOR U9006 ( .A(n7719), .B(n7720), .Z(n7713) );
  ANDN U9007 ( .A(n7721), .B(n4627), .Z(n7720) );
  XOR U9008 ( .A(n7722), .B(n7723), .Z(n4627) );
  IV U9009 ( .A(n7719), .Z(n7722) );
  XNOR U9010 ( .A(n4628), .B(n7719), .Z(n7721) );
  NAND U9011 ( .A(n7724), .B(nreg[763]), .Z(n4628) );
  NAND U9012 ( .A(n6107), .B(nreg[763]), .Z(n7724) );
  XOR U9013 ( .A(n7725), .B(n7726), .Z(n7719) );
  ANDN U9014 ( .A(n7727), .B(n4629), .Z(n7726) );
  XOR U9015 ( .A(n7728), .B(n7729), .Z(n4629) );
  IV U9016 ( .A(n7725), .Z(n7728) );
  XNOR U9017 ( .A(n4630), .B(n7725), .Z(n7727) );
  NAND U9018 ( .A(n7730), .B(nreg[762]), .Z(n4630) );
  NAND U9019 ( .A(n6107), .B(nreg[762]), .Z(n7730) );
  XOR U9020 ( .A(n7731), .B(n7732), .Z(n7725) );
  ANDN U9021 ( .A(n7733), .B(n4631), .Z(n7732) );
  XOR U9022 ( .A(n7734), .B(n7735), .Z(n4631) );
  IV U9023 ( .A(n7731), .Z(n7734) );
  XNOR U9024 ( .A(n4632), .B(n7731), .Z(n7733) );
  NAND U9025 ( .A(n7736), .B(nreg[761]), .Z(n4632) );
  NAND U9026 ( .A(n6107), .B(nreg[761]), .Z(n7736) );
  XOR U9027 ( .A(n7737), .B(n7738), .Z(n7731) );
  ANDN U9028 ( .A(n7739), .B(n4633), .Z(n7738) );
  XOR U9029 ( .A(n7740), .B(n7741), .Z(n4633) );
  IV U9030 ( .A(n7737), .Z(n7740) );
  XNOR U9031 ( .A(n4634), .B(n7737), .Z(n7739) );
  NAND U9032 ( .A(n7742), .B(nreg[760]), .Z(n4634) );
  NAND U9033 ( .A(n6107), .B(nreg[760]), .Z(n7742) );
  XOR U9034 ( .A(n7743), .B(n7744), .Z(n7737) );
  ANDN U9035 ( .A(n7745), .B(n4635), .Z(n7744) );
  XOR U9036 ( .A(n7746), .B(n7747), .Z(n4635) );
  IV U9037 ( .A(n7743), .Z(n7746) );
  XNOR U9038 ( .A(n4636), .B(n7743), .Z(n7745) );
  NAND U9039 ( .A(n7748), .B(nreg[759]), .Z(n4636) );
  NAND U9040 ( .A(n6107), .B(nreg[759]), .Z(n7748) );
  XOR U9041 ( .A(n7749), .B(n7750), .Z(n7743) );
  ANDN U9042 ( .A(n7751), .B(n4637), .Z(n7750) );
  XOR U9043 ( .A(n7752), .B(n7753), .Z(n4637) );
  IV U9044 ( .A(n7749), .Z(n7752) );
  XNOR U9045 ( .A(n4638), .B(n7749), .Z(n7751) );
  NAND U9046 ( .A(n7754), .B(nreg[758]), .Z(n4638) );
  NAND U9047 ( .A(n6107), .B(nreg[758]), .Z(n7754) );
  XOR U9048 ( .A(n7755), .B(n7756), .Z(n7749) );
  ANDN U9049 ( .A(n7757), .B(n4639), .Z(n7756) );
  XOR U9050 ( .A(n7758), .B(n7759), .Z(n4639) );
  IV U9051 ( .A(n7755), .Z(n7758) );
  XNOR U9052 ( .A(n4640), .B(n7755), .Z(n7757) );
  NAND U9053 ( .A(n7760), .B(nreg[757]), .Z(n4640) );
  NAND U9054 ( .A(n6107), .B(nreg[757]), .Z(n7760) );
  XOR U9055 ( .A(n7761), .B(n7762), .Z(n7755) );
  ANDN U9056 ( .A(n7763), .B(n4643), .Z(n7762) );
  XOR U9057 ( .A(n7764), .B(n7765), .Z(n4643) );
  IV U9058 ( .A(n7761), .Z(n7764) );
  XNOR U9059 ( .A(n4644), .B(n7761), .Z(n7763) );
  NAND U9060 ( .A(n7766), .B(nreg[756]), .Z(n4644) );
  NAND U9061 ( .A(n6107), .B(nreg[756]), .Z(n7766) );
  XOR U9062 ( .A(n7767), .B(n7768), .Z(n7761) );
  ANDN U9063 ( .A(n7769), .B(n4645), .Z(n7768) );
  XOR U9064 ( .A(n7770), .B(n7771), .Z(n4645) );
  IV U9065 ( .A(n7767), .Z(n7770) );
  XNOR U9066 ( .A(n4646), .B(n7767), .Z(n7769) );
  NAND U9067 ( .A(n7772), .B(nreg[755]), .Z(n4646) );
  NAND U9068 ( .A(n6107), .B(nreg[755]), .Z(n7772) );
  XOR U9069 ( .A(n7773), .B(n7774), .Z(n7767) );
  ANDN U9070 ( .A(n7775), .B(n4647), .Z(n7774) );
  XOR U9071 ( .A(n7776), .B(n7777), .Z(n4647) );
  IV U9072 ( .A(n7773), .Z(n7776) );
  XNOR U9073 ( .A(n4648), .B(n7773), .Z(n7775) );
  NAND U9074 ( .A(n7778), .B(nreg[754]), .Z(n4648) );
  NAND U9075 ( .A(n6107), .B(nreg[754]), .Z(n7778) );
  XOR U9076 ( .A(n7779), .B(n7780), .Z(n7773) );
  ANDN U9077 ( .A(n7781), .B(n4649), .Z(n7780) );
  XOR U9078 ( .A(n7782), .B(n7783), .Z(n4649) );
  IV U9079 ( .A(n7779), .Z(n7782) );
  XNOR U9080 ( .A(n4650), .B(n7779), .Z(n7781) );
  NAND U9081 ( .A(n7784), .B(nreg[753]), .Z(n4650) );
  NAND U9082 ( .A(n6107), .B(nreg[753]), .Z(n7784) );
  XOR U9083 ( .A(n7785), .B(n7786), .Z(n7779) );
  ANDN U9084 ( .A(n7787), .B(n4651), .Z(n7786) );
  XOR U9085 ( .A(n7788), .B(n7789), .Z(n4651) );
  IV U9086 ( .A(n7785), .Z(n7788) );
  XNOR U9087 ( .A(n4652), .B(n7785), .Z(n7787) );
  NAND U9088 ( .A(n7790), .B(nreg[752]), .Z(n4652) );
  NAND U9089 ( .A(n6107), .B(nreg[752]), .Z(n7790) );
  XOR U9090 ( .A(n7791), .B(n7792), .Z(n7785) );
  ANDN U9091 ( .A(n7793), .B(n4653), .Z(n7792) );
  XOR U9092 ( .A(n7794), .B(n7795), .Z(n4653) );
  IV U9093 ( .A(n7791), .Z(n7794) );
  XNOR U9094 ( .A(n4654), .B(n7791), .Z(n7793) );
  NAND U9095 ( .A(n7796), .B(nreg[751]), .Z(n4654) );
  NAND U9096 ( .A(n6107), .B(nreg[751]), .Z(n7796) );
  XOR U9097 ( .A(n7797), .B(n7798), .Z(n7791) );
  ANDN U9098 ( .A(n7799), .B(n4655), .Z(n7798) );
  XOR U9099 ( .A(n7800), .B(n7801), .Z(n4655) );
  IV U9100 ( .A(n7797), .Z(n7800) );
  XNOR U9101 ( .A(n4656), .B(n7797), .Z(n7799) );
  NAND U9102 ( .A(n7802), .B(nreg[750]), .Z(n4656) );
  NAND U9103 ( .A(n6107), .B(nreg[750]), .Z(n7802) );
  XOR U9104 ( .A(n7803), .B(n7804), .Z(n7797) );
  ANDN U9105 ( .A(n7805), .B(n4657), .Z(n7804) );
  XOR U9106 ( .A(n7806), .B(n7807), .Z(n4657) );
  IV U9107 ( .A(n7803), .Z(n7806) );
  XNOR U9108 ( .A(n4658), .B(n7803), .Z(n7805) );
  NAND U9109 ( .A(n7808), .B(nreg[749]), .Z(n4658) );
  NAND U9110 ( .A(n6107), .B(nreg[749]), .Z(n7808) );
  XOR U9111 ( .A(n7809), .B(n7810), .Z(n7803) );
  ANDN U9112 ( .A(n7811), .B(n4659), .Z(n7810) );
  XOR U9113 ( .A(n7812), .B(n7813), .Z(n4659) );
  IV U9114 ( .A(n7809), .Z(n7812) );
  XNOR U9115 ( .A(n4660), .B(n7809), .Z(n7811) );
  NAND U9116 ( .A(n7814), .B(nreg[748]), .Z(n4660) );
  NAND U9117 ( .A(n6107), .B(nreg[748]), .Z(n7814) );
  XOR U9118 ( .A(n7815), .B(n7816), .Z(n7809) );
  ANDN U9119 ( .A(n7817), .B(n4661), .Z(n7816) );
  XOR U9120 ( .A(n7818), .B(n7819), .Z(n4661) );
  IV U9121 ( .A(n7815), .Z(n7818) );
  XNOR U9122 ( .A(n4662), .B(n7815), .Z(n7817) );
  NAND U9123 ( .A(n7820), .B(nreg[747]), .Z(n4662) );
  NAND U9124 ( .A(n6107), .B(nreg[747]), .Z(n7820) );
  XOR U9125 ( .A(n7821), .B(n7822), .Z(n7815) );
  ANDN U9126 ( .A(n7823), .B(n4665), .Z(n7822) );
  XOR U9127 ( .A(n7824), .B(n7825), .Z(n4665) );
  IV U9128 ( .A(n7821), .Z(n7824) );
  XNOR U9129 ( .A(n4666), .B(n7821), .Z(n7823) );
  NAND U9130 ( .A(n7826), .B(nreg[746]), .Z(n4666) );
  NAND U9131 ( .A(n6107), .B(nreg[746]), .Z(n7826) );
  XOR U9132 ( .A(n7827), .B(n7828), .Z(n7821) );
  ANDN U9133 ( .A(n7829), .B(n4667), .Z(n7828) );
  XOR U9134 ( .A(n7830), .B(n7831), .Z(n4667) );
  IV U9135 ( .A(n7827), .Z(n7830) );
  XNOR U9136 ( .A(n4668), .B(n7827), .Z(n7829) );
  NAND U9137 ( .A(n7832), .B(nreg[745]), .Z(n4668) );
  NAND U9138 ( .A(n6107), .B(nreg[745]), .Z(n7832) );
  XOR U9139 ( .A(n7833), .B(n7834), .Z(n7827) );
  ANDN U9140 ( .A(n7835), .B(n4669), .Z(n7834) );
  XOR U9141 ( .A(n7836), .B(n7837), .Z(n4669) );
  IV U9142 ( .A(n7833), .Z(n7836) );
  XNOR U9143 ( .A(n4670), .B(n7833), .Z(n7835) );
  NAND U9144 ( .A(n7838), .B(nreg[744]), .Z(n4670) );
  NAND U9145 ( .A(n6107), .B(nreg[744]), .Z(n7838) );
  XOR U9146 ( .A(n7839), .B(n7840), .Z(n7833) );
  ANDN U9147 ( .A(n7841), .B(n4671), .Z(n7840) );
  XOR U9148 ( .A(n7842), .B(n7843), .Z(n4671) );
  IV U9149 ( .A(n7839), .Z(n7842) );
  XNOR U9150 ( .A(n4672), .B(n7839), .Z(n7841) );
  NAND U9151 ( .A(n7844), .B(nreg[743]), .Z(n4672) );
  NAND U9152 ( .A(n6107), .B(nreg[743]), .Z(n7844) );
  XOR U9153 ( .A(n7845), .B(n7846), .Z(n7839) );
  ANDN U9154 ( .A(n7847), .B(n4673), .Z(n7846) );
  XOR U9155 ( .A(n7848), .B(n7849), .Z(n4673) );
  IV U9156 ( .A(n7845), .Z(n7848) );
  XNOR U9157 ( .A(n4674), .B(n7845), .Z(n7847) );
  NAND U9158 ( .A(n7850), .B(nreg[742]), .Z(n4674) );
  NAND U9159 ( .A(n6107), .B(nreg[742]), .Z(n7850) );
  XOR U9160 ( .A(n7851), .B(n7852), .Z(n7845) );
  ANDN U9161 ( .A(n7853), .B(n4675), .Z(n7852) );
  XOR U9162 ( .A(n7854), .B(n7855), .Z(n4675) );
  IV U9163 ( .A(n7851), .Z(n7854) );
  XNOR U9164 ( .A(n4676), .B(n7851), .Z(n7853) );
  NAND U9165 ( .A(n7856), .B(nreg[741]), .Z(n4676) );
  NAND U9166 ( .A(n6107), .B(nreg[741]), .Z(n7856) );
  XOR U9167 ( .A(n7857), .B(n7858), .Z(n7851) );
  ANDN U9168 ( .A(n7859), .B(n4677), .Z(n7858) );
  XOR U9169 ( .A(n7860), .B(n7861), .Z(n4677) );
  IV U9170 ( .A(n7857), .Z(n7860) );
  XNOR U9171 ( .A(n4678), .B(n7857), .Z(n7859) );
  NAND U9172 ( .A(n7862), .B(nreg[740]), .Z(n4678) );
  NAND U9173 ( .A(n6107), .B(nreg[740]), .Z(n7862) );
  XOR U9174 ( .A(n7863), .B(n7864), .Z(n7857) );
  ANDN U9175 ( .A(n7865), .B(n4679), .Z(n7864) );
  XOR U9176 ( .A(n7866), .B(n7867), .Z(n4679) );
  IV U9177 ( .A(n7863), .Z(n7866) );
  XNOR U9178 ( .A(n4680), .B(n7863), .Z(n7865) );
  NAND U9179 ( .A(n7868), .B(nreg[739]), .Z(n4680) );
  NAND U9180 ( .A(n6107), .B(nreg[739]), .Z(n7868) );
  XOR U9181 ( .A(n7869), .B(n7870), .Z(n7863) );
  ANDN U9182 ( .A(n7871), .B(n4681), .Z(n7870) );
  XOR U9183 ( .A(n7872), .B(n7873), .Z(n4681) );
  IV U9184 ( .A(n7869), .Z(n7872) );
  XNOR U9185 ( .A(n4682), .B(n7869), .Z(n7871) );
  NAND U9186 ( .A(n7874), .B(nreg[738]), .Z(n4682) );
  NAND U9187 ( .A(n6107), .B(nreg[738]), .Z(n7874) );
  XOR U9188 ( .A(n7875), .B(n7876), .Z(n7869) );
  ANDN U9189 ( .A(n7877), .B(n4683), .Z(n7876) );
  XOR U9190 ( .A(n7878), .B(n7879), .Z(n4683) );
  IV U9191 ( .A(n7875), .Z(n7878) );
  XNOR U9192 ( .A(n4684), .B(n7875), .Z(n7877) );
  NAND U9193 ( .A(n7880), .B(nreg[737]), .Z(n4684) );
  NAND U9194 ( .A(n6107), .B(nreg[737]), .Z(n7880) );
  XOR U9195 ( .A(n7881), .B(n7882), .Z(n7875) );
  ANDN U9196 ( .A(n7883), .B(n4687), .Z(n7882) );
  XOR U9197 ( .A(n7884), .B(n7885), .Z(n4687) );
  IV U9198 ( .A(n7881), .Z(n7884) );
  XNOR U9199 ( .A(n4688), .B(n7881), .Z(n7883) );
  NAND U9200 ( .A(n7886), .B(nreg[736]), .Z(n4688) );
  NAND U9201 ( .A(n6107), .B(nreg[736]), .Z(n7886) );
  XOR U9202 ( .A(n7887), .B(n7888), .Z(n7881) );
  ANDN U9203 ( .A(n7889), .B(n4689), .Z(n7888) );
  XOR U9204 ( .A(n7890), .B(n7891), .Z(n4689) );
  IV U9205 ( .A(n7887), .Z(n7890) );
  XNOR U9206 ( .A(n4690), .B(n7887), .Z(n7889) );
  NAND U9207 ( .A(n7892), .B(nreg[735]), .Z(n4690) );
  NAND U9208 ( .A(n6107), .B(nreg[735]), .Z(n7892) );
  XOR U9209 ( .A(n7893), .B(n7894), .Z(n7887) );
  ANDN U9210 ( .A(n7895), .B(n4691), .Z(n7894) );
  XOR U9211 ( .A(n7896), .B(n7897), .Z(n4691) );
  IV U9212 ( .A(n7893), .Z(n7896) );
  XNOR U9213 ( .A(n4692), .B(n7893), .Z(n7895) );
  NAND U9214 ( .A(n7898), .B(nreg[734]), .Z(n4692) );
  NAND U9215 ( .A(n6107), .B(nreg[734]), .Z(n7898) );
  XOR U9216 ( .A(n7899), .B(n7900), .Z(n7893) );
  ANDN U9217 ( .A(n7901), .B(n4693), .Z(n7900) );
  XOR U9218 ( .A(n7902), .B(n7903), .Z(n4693) );
  IV U9219 ( .A(n7899), .Z(n7902) );
  XNOR U9220 ( .A(n4694), .B(n7899), .Z(n7901) );
  NAND U9221 ( .A(n7904), .B(nreg[733]), .Z(n4694) );
  NAND U9222 ( .A(n6107), .B(nreg[733]), .Z(n7904) );
  XOR U9223 ( .A(n7905), .B(n7906), .Z(n7899) );
  ANDN U9224 ( .A(n7907), .B(n4695), .Z(n7906) );
  XOR U9225 ( .A(n7908), .B(n7909), .Z(n4695) );
  IV U9226 ( .A(n7905), .Z(n7908) );
  XNOR U9227 ( .A(n4696), .B(n7905), .Z(n7907) );
  NAND U9228 ( .A(n7910), .B(nreg[732]), .Z(n4696) );
  NAND U9229 ( .A(n6107), .B(nreg[732]), .Z(n7910) );
  XOR U9230 ( .A(n7911), .B(n7912), .Z(n7905) );
  ANDN U9231 ( .A(n7913), .B(n4697), .Z(n7912) );
  XOR U9232 ( .A(n7914), .B(n7915), .Z(n4697) );
  IV U9233 ( .A(n7911), .Z(n7914) );
  XNOR U9234 ( .A(n4698), .B(n7911), .Z(n7913) );
  NAND U9235 ( .A(n7916), .B(nreg[731]), .Z(n4698) );
  NAND U9236 ( .A(n6107), .B(nreg[731]), .Z(n7916) );
  XOR U9237 ( .A(n7917), .B(n7918), .Z(n7911) );
  ANDN U9238 ( .A(n7919), .B(n4699), .Z(n7918) );
  XOR U9239 ( .A(n7920), .B(n7921), .Z(n4699) );
  IV U9240 ( .A(n7917), .Z(n7920) );
  XNOR U9241 ( .A(n4700), .B(n7917), .Z(n7919) );
  NAND U9242 ( .A(n7922), .B(nreg[730]), .Z(n4700) );
  NAND U9243 ( .A(n6107), .B(nreg[730]), .Z(n7922) );
  XOR U9244 ( .A(n7923), .B(n7924), .Z(n7917) );
  ANDN U9245 ( .A(n7925), .B(n4701), .Z(n7924) );
  XOR U9246 ( .A(n7926), .B(n7927), .Z(n4701) );
  IV U9247 ( .A(n7923), .Z(n7926) );
  XNOR U9248 ( .A(n4702), .B(n7923), .Z(n7925) );
  NAND U9249 ( .A(n7928), .B(nreg[729]), .Z(n4702) );
  NAND U9250 ( .A(n6107), .B(nreg[729]), .Z(n7928) );
  XOR U9251 ( .A(n7929), .B(n7930), .Z(n7923) );
  ANDN U9252 ( .A(n7931), .B(n4703), .Z(n7930) );
  XOR U9253 ( .A(n7932), .B(n7933), .Z(n4703) );
  IV U9254 ( .A(n7929), .Z(n7932) );
  XNOR U9255 ( .A(n4704), .B(n7929), .Z(n7931) );
  NAND U9256 ( .A(n7934), .B(nreg[728]), .Z(n4704) );
  NAND U9257 ( .A(n6107), .B(nreg[728]), .Z(n7934) );
  XOR U9258 ( .A(n7935), .B(n7936), .Z(n7929) );
  ANDN U9259 ( .A(n7937), .B(n4705), .Z(n7936) );
  XOR U9260 ( .A(n7938), .B(n7939), .Z(n4705) );
  IV U9261 ( .A(n7935), .Z(n7938) );
  XNOR U9262 ( .A(n4706), .B(n7935), .Z(n7937) );
  NAND U9263 ( .A(n7940), .B(nreg[727]), .Z(n4706) );
  NAND U9264 ( .A(n6107), .B(nreg[727]), .Z(n7940) );
  XOR U9265 ( .A(n7941), .B(n7942), .Z(n7935) );
  ANDN U9266 ( .A(n7943), .B(n4709), .Z(n7942) );
  XOR U9267 ( .A(n7944), .B(n7945), .Z(n4709) );
  IV U9268 ( .A(n7941), .Z(n7944) );
  XNOR U9269 ( .A(n4710), .B(n7941), .Z(n7943) );
  NAND U9270 ( .A(n7946), .B(nreg[726]), .Z(n4710) );
  NAND U9271 ( .A(n6107), .B(nreg[726]), .Z(n7946) );
  XOR U9272 ( .A(n7947), .B(n7948), .Z(n7941) );
  ANDN U9273 ( .A(n7949), .B(n4711), .Z(n7948) );
  XOR U9274 ( .A(n7950), .B(n7951), .Z(n4711) );
  IV U9275 ( .A(n7947), .Z(n7950) );
  XNOR U9276 ( .A(n4712), .B(n7947), .Z(n7949) );
  NAND U9277 ( .A(n7952), .B(nreg[725]), .Z(n4712) );
  NAND U9278 ( .A(n6107), .B(nreg[725]), .Z(n7952) );
  XOR U9279 ( .A(n7953), .B(n7954), .Z(n7947) );
  ANDN U9280 ( .A(n7955), .B(n4713), .Z(n7954) );
  XOR U9281 ( .A(n7956), .B(n7957), .Z(n4713) );
  IV U9282 ( .A(n7953), .Z(n7956) );
  XNOR U9283 ( .A(n4714), .B(n7953), .Z(n7955) );
  NAND U9284 ( .A(n7958), .B(nreg[724]), .Z(n4714) );
  NAND U9285 ( .A(n6107), .B(nreg[724]), .Z(n7958) );
  XOR U9286 ( .A(n7959), .B(n7960), .Z(n7953) );
  ANDN U9287 ( .A(n7961), .B(n4715), .Z(n7960) );
  XOR U9288 ( .A(n7962), .B(n7963), .Z(n4715) );
  IV U9289 ( .A(n7959), .Z(n7962) );
  XNOR U9290 ( .A(n4716), .B(n7959), .Z(n7961) );
  NAND U9291 ( .A(n7964), .B(nreg[723]), .Z(n4716) );
  NAND U9292 ( .A(n6107), .B(nreg[723]), .Z(n7964) );
  XOR U9293 ( .A(n7965), .B(n7966), .Z(n7959) );
  ANDN U9294 ( .A(n7967), .B(n4717), .Z(n7966) );
  XOR U9295 ( .A(n7968), .B(n7969), .Z(n4717) );
  IV U9296 ( .A(n7965), .Z(n7968) );
  XNOR U9297 ( .A(n4718), .B(n7965), .Z(n7967) );
  NAND U9298 ( .A(n7970), .B(nreg[722]), .Z(n4718) );
  NAND U9299 ( .A(n6107), .B(nreg[722]), .Z(n7970) );
  XOR U9300 ( .A(n7971), .B(n7972), .Z(n7965) );
  ANDN U9301 ( .A(n7973), .B(n4719), .Z(n7972) );
  XOR U9302 ( .A(n7974), .B(n7975), .Z(n4719) );
  IV U9303 ( .A(n7971), .Z(n7974) );
  XNOR U9304 ( .A(n4720), .B(n7971), .Z(n7973) );
  NAND U9305 ( .A(n7976), .B(nreg[721]), .Z(n4720) );
  NAND U9306 ( .A(n6107), .B(nreg[721]), .Z(n7976) );
  XOR U9307 ( .A(n7977), .B(n7978), .Z(n7971) );
  ANDN U9308 ( .A(n7979), .B(n4721), .Z(n7978) );
  XOR U9309 ( .A(n7980), .B(n7981), .Z(n4721) );
  IV U9310 ( .A(n7977), .Z(n7980) );
  XNOR U9311 ( .A(n4722), .B(n7977), .Z(n7979) );
  NAND U9312 ( .A(n7982), .B(nreg[720]), .Z(n4722) );
  NAND U9313 ( .A(n6107), .B(nreg[720]), .Z(n7982) );
  XOR U9314 ( .A(n7983), .B(n7984), .Z(n7977) );
  ANDN U9315 ( .A(n7985), .B(n4723), .Z(n7984) );
  XOR U9316 ( .A(n7986), .B(n7987), .Z(n4723) );
  IV U9317 ( .A(n7983), .Z(n7986) );
  XNOR U9318 ( .A(n4724), .B(n7983), .Z(n7985) );
  NAND U9319 ( .A(n7988), .B(nreg[719]), .Z(n4724) );
  NAND U9320 ( .A(n6107), .B(nreg[719]), .Z(n7988) );
  XOR U9321 ( .A(n7989), .B(n7990), .Z(n7983) );
  ANDN U9322 ( .A(n7991), .B(n4725), .Z(n7990) );
  XOR U9323 ( .A(n7992), .B(n7993), .Z(n4725) );
  IV U9324 ( .A(n7989), .Z(n7992) );
  XNOR U9325 ( .A(n4726), .B(n7989), .Z(n7991) );
  NAND U9326 ( .A(n7994), .B(nreg[718]), .Z(n4726) );
  NAND U9327 ( .A(n6107), .B(nreg[718]), .Z(n7994) );
  XOR U9328 ( .A(n7995), .B(n7996), .Z(n7989) );
  ANDN U9329 ( .A(n7997), .B(n4727), .Z(n7996) );
  XOR U9330 ( .A(n7998), .B(n7999), .Z(n4727) );
  IV U9331 ( .A(n7995), .Z(n7998) );
  XNOR U9332 ( .A(n4728), .B(n7995), .Z(n7997) );
  NAND U9333 ( .A(n8000), .B(nreg[717]), .Z(n4728) );
  NAND U9334 ( .A(n6107), .B(nreg[717]), .Z(n8000) );
  XOR U9335 ( .A(n8001), .B(n8002), .Z(n7995) );
  ANDN U9336 ( .A(n8003), .B(n4731), .Z(n8002) );
  XOR U9337 ( .A(n8004), .B(n8005), .Z(n4731) );
  IV U9338 ( .A(n8001), .Z(n8004) );
  XNOR U9339 ( .A(n4732), .B(n8001), .Z(n8003) );
  NAND U9340 ( .A(n8006), .B(nreg[716]), .Z(n4732) );
  NAND U9341 ( .A(n6107), .B(nreg[716]), .Z(n8006) );
  XOR U9342 ( .A(n8007), .B(n8008), .Z(n8001) );
  ANDN U9343 ( .A(n8009), .B(n4733), .Z(n8008) );
  XOR U9344 ( .A(n8010), .B(n8011), .Z(n4733) );
  IV U9345 ( .A(n8007), .Z(n8010) );
  XNOR U9346 ( .A(n4734), .B(n8007), .Z(n8009) );
  NAND U9347 ( .A(n8012), .B(nreg[715]), .Z(n4734) );
  NAND U9348 ( .A(n6107), .B(nreg[715]), .Z(n8012) );
  XOR U9349 ( .A(n8013), .B(n8014), .Z(n8007) );
  ANDN U9350 ( .A(n8015), .B(n4735), .Z(n8014) );
  XOR U9351 ( .A(n8016), .B(n8017), .Z(n4735) );
  IV U9352 ( .A(n8013), .Z(n8016) );
  XNOR U9353 ( .A(n4736), .B(n8013), .Z(n8015) );
  NAND U9354 ( .A(n8018), .B(nreg[714]), .Z(n4736) );
  NAND U9355 ( .A(n6107), .B(nreg[714]), .Z(n8018) );
  XOR U9356 ( .A(n8019), .B(n8020), .Z(n8013) );
  ANDN U9357 ( .A(n8021), .B(n4737), .Z(n8020) );
  XOR U9358 ( .A(n8022), .B(n8023), .Z(n4737) );
  IV U9359 ( .A(n8019), .Z(n8022) );
  XNOR U9360 ( .A(n4738), .B(n8019), .Z(n8021) );
  NAND U9361 ( .A(n8024), .B(nreg[713]), .Z(n4738) );
  NAND U9362 ( .A(n6107), .B(nreg[713]), .Z(n8024) );
  XOR U9363 ( .A(n8025), .B(n8026), .Z(n8019) );
  ANDN U9364 ( .A(n8027), .B(n4739), .Z(n8026) );
  XOR U9365 ( .A(n8028), .B(n8029), .Z(n4739) );
  IV U9366 ( .A(n8025), .Z(n8028) );
  XNOR U9367 ( .A(n4740), .B(n8025), .Z(n8027) );
  NAND U9368 ( .A(n8030), .B(nreg[712]), .Z(n4740) );
  NAND U9369 ( .A(n6107), .B(nreg[712]), .Z(n8030) );
  XOR U9370 ( .A(n8031), .B(n8032), .Z(n8025) );
  ANDN U9371 ( .A(n8033), .B(n4741), .Z(n8032) );
  XOR U9372 ( .A(n8034), .B(n8035), .Z(n4741) );
  IV U9373 ( .A(n8031), .Z(n8034) );
  XNOR U9374 ( .A(n4742), .B(n8031), .Z(n8033) );
  NAND U9375 ( .A(n8036), .B(nreg[711]), .Z(n4742) );
  NAND U9376 ( .A(n6107), .B(nreg[711]), .Z(n8036) );
  XOR U9377 ( .A(n8037), .B(n8038), .Z(n8031) );
  ANDN U9378 ( .A(n8039), .B(n4743), .Z(n8038) );
  XOR U9379 ( .A(n8040), .B(n8041), .Z(n4743) );
  IV U9380 ( .A(n8037), .Z(n8040) );
  XNOR U9381 ( .A(n4744), .B(n8037), .Z(n8039) );
  NAND U9382 ( .A(n8042), .B(nreg[710]), .Z(n4744) );
  NAND U9383 ( .A(n6107), .B(nreg[710]), .Z(n8042) );
  XOR U9384 ( .A(n8043), .B(n8044), .Z(n8037) );
  ANDN U9385 ( .A(n8045), .B(n4745), .Z(n8044) );
  XOR U9386 ( .A(n8046), .B(n8047), .Z(n4745) );
  IV U9387 ( .A(n8043), .Z(n8046) );
  XNOR U9388 ( .A(n4746), .B(n8043), .Z(n8045) );
  NAND U9389 ( .A(n8048), .B(nreg[709]), .Z(n4746) );
  NAND U9390 ( .A(n6107), .B(nreg[709]), .Z(n8048) );
  XOR U9391 ( .A(n8049), .B(n8050), .Z(n8043) );
  ANDN U9392 ( .A(n8051), .B(n4747), .Z(n8050) );
  XOR U9393 ( .A(n8052), .B(n8053), .Z(n4747) );
  IV U9394 ( .A(n8049), .Z(n8052) );
  XNOR U9395 ( .A(n4748), .B(n8049), .Z(n8051) );
  NAND U9396 ( .A(n8054), .B(nreg[708]), .Z(n4748) );
  NAND U9397 ( .A(n6107), .B(nreg[708]), .Z(n8054) );
  XOR U9398 ( .A(n8055), .B(n8056), .Z(n8049) );
  ANDN U9399 ( .A(n8057), .B(n4749), .Z(n8056) );
  XOR U9400 ( .A(n8058), .B(n8059), .Z(n4749) );
  IV U9401 ( .A(n8055), .Z(n8058) );
  XNOR U9402 ( .A(n4750), .B(n8055), .Z(n8057) );
  NAND U9403 ( .A(n8060), .B(nreg[707]), .Z(n4750) );
  NAND U9404 ( .A(n6107), .B(nreg[707]), .Z(n8060) );
  XOR U9405 ( .A(n8061), .B(n8062), .Z(n8055) );
  ANDN U9406 ( .A(n8063), .B(n4753), .Z(n8062) );
  XOR U9407 ( .A(n8064), .B(n8065), .Z(n4753) );
  IV U9408 ( .A(n8061), .Z(n8064) );
  XNOR U9409 ( .A(n4754), .B(n8061), .Z(n8063) );
  NAND U9410 ( .A(n8066), .B(nreg[706]), .Z(n4754) );
  NAND U9411 ( .A(n6107), .B(nreg[706]), .Z(n8066) );
  XOR U9412 ( .A(n8067), .B(n8068), .Z(n8061) );
  ANDN U9413 ( .A(n8069), .B(n4755), .Z(n8068) );
  XOR U9414 ( .A(n8070), .B(n8071), .Z(n4755) );
  IV U9415 ( .A(n8067), .Z(n8070) );
  XNOR U9416 ( .A(n4756), .B(n8067), .Z(n8069) );
  NAND U9417 ( .A(n8072), .B(nreg[705]), .Z(n4756) );
  NAND U9418 ( .A(n6107), .B(nreg[705]), .Z(n8072) );
  XOR U9419 ( .A(n8073), .B(n8074), .Z(n8067) );
  ANDN U9420 ( .A(n8075), .B(n4757), .Z(n8074) );
  XOR U9421 ( .A(n8076), .B(n8077), .Z(n4757) );
  IV U9422 ( .A(n8073), .Z(n8076) );
  XNOR U9423 ( .A(n4758), .B(n8073), .Z(n8075) );
  NAND U9424 ( .A(n8078), .B(nreg[704]), .Z(n4758) );
  NAND U9425 ( .A(n6107), .B(nreg[704]), .Z(n8078) );
  XOR U9426 ( .A(n8079), .B(n8080), .Z(n8073) );
  ANDN U9427 ( .A(n8081), .B(n4759), .Z(n8080) );
  XOR U9428 ( .A(n8082), .B(n8083), .Z(n4759) );
  IV U9429 ( .A(n8079), .Z(n8082) );
  XNOR U9430 ( .A(n4760), .B(n8079), .Z(n8081) );
  NAND U9431 ( .A(n8084), .B(nreg[703]), .Z(n4760) );
  NAND U9432 ( .A(n6107), .B(nreg[703]), .Z(n8084) );
  XOR U9433 ( .A(n8085), .B(n8086), .Z(n8079) );
  ANDN U9434 ( .A(n8087), .B(n4761), .Z(n8086) );
  XOR U9435 ( .A(n8088), .B(n8089), .Z(n4761) );
  IV U9436 ( .A(n8085), .Z(n8088) );
  XNOR U9437 ( .A(n4762), .B(n8085), .Z(n8087) );
  NAND U9438 ( .A(n8090), .B(nreg[702]), .Z(n4762) );
  NAND U9439 ( .A(n6107), .B(nreg[702]), .Z(n8090) );
  XOR U9440 ( .A(n8091), .B(n8092), .Z(n8085) );
  ANDN U9441 ( .A(n8093), .B(n4763), .Z(n8092) );
  XOR U9442 ( .A(n8094), .B(n8095), .Z(n4763) );
  IV U9443 ( .A(n8091), .Z(n8094) );
  XNOR U9444 ( .A(n4764), .B(n8091), .Z(n8093) );
  NAND U9445 ( .A(n8096), .B(nreg[701]), .Z(n4764) );
  NAND U9446 ( .A(n6107), .B(nreg[701]), .Z(n8096) );
  XOR U9447 ( .A(n8097), .B(n8098), .Z(n8091) );
  ANDN U9448 ( .A(n8099), .B(n4765), .Z(n8098) );
  XOR U9449 ( .A(n8100), .B(n8101), .Z(n4765) );
  IV U9450 ( .A(n8097), .Z(n8100) );
  XNOR U9451 ( .A(n4766), .B(n8097), .Z(n8099) );
  NAND U9452 ( .A(n8102), .B(nreg[700]), .Z(n4766) );
  NAND U9453 ( .A(n6107), .B(nreg[700]), .Z(n8102) );
  XOR U9454 ( .A(n8103), .B(n8104), .Z(n8097) );
  ANDN U9455 ( .A(n8105), .B(n4767), .Z(n8104) );
  XOR U9456 ( .A(n8106), .B(n8107), .Z(n4767) );
  IV U9457 ( .A(n8103), .Z(n8106) );
  XNOR U9458 ( .A(n4768), .B(n8103), .Z(n8105) );
  NAND U9459 ( .A(n8108), .B(nreg[699]), .Z(n4768) );
  NAND U9460 ( .A(n6107), .B(nreg[699]), .Z(n8108) );
  XOR U9461 ( .A(n8109), .B(n8110), .Z(n8103) );
  ANDN U9462 ( .A(n8111), .B(n4769), .Z(n8110) );
  XOR U9463 ( .A(n8112), .B(n8113), .Z(n4769) );
  IV U9464 ( .A(n8109), .Z(n8112) );
  XNOR U9465 ( .A(n4770), .B(n8109), .Z(n8111) );
  NAND U9466 ( .A(n8114), .B(nreg[698]), .Z(n4770) );
  NAND U9467 ( .A(n6107), .B(nreg[698]), .Z(n8114) );
  XOR U9468 ( .A(n8115), .B(n8116), .Z(n8109) );
  ANDN U9469 ( .A(n8117), .B(n4771), .Z(n8116) );
  XOR U9470 ( .A(n8118), .B(n8119), .Z(n4771) );
  IV U9471 ( .A(n8115), .Z(n8118) );
  XNOR U9472 ( .A(n4772), .B(n8115), .Z(n8117) );
  NAND U9473 ( .A(n8120), .B(nreg[697]), .Z(n4772) );
  NAND U9474 ( .A(n6107), .B(nreg[697]), .Z(n8120) );
  XOR U9475 ( .A(n8121), .B(n8122), .Z(n8115) );
  ANDN U9476 ( .A(n8123), .B(n4777), .Z(n8122) );
  XOR U9477 ( .A(n8124), .B(n8125), .Z(n4777) );
  IV U9478 ( .A(n8121), .Z(n8124) );
  XNOR U9479 ( .A(n4778), .B(n8121), .Z(n8123) );
  NAND U9480 ( .A(n8126), .B(nreg[696]), .Z(n4778) );
  NAND U9481 ( .A(n6107), .B(nreg[696]), .Z(n8126) );
  XOR U9482 ( .A(n8127), .B(n8128), .Z(n8121) );
  ANDN U9483 ( .A(n8129), .B(n4779), .Z(n8128) );
  XOR U9484 ( .A(n8130), .B(n8131), .Z(n4779) );
  IV U9485 ( .A(n8127), .Z(n8130) );
  XNOR U9486 ( .A(n4780), .B(n8127), .Z(n8129) );
  NAND U9487 ( .A(n8132), .B(nreg[695]), .Z(n4780) );
  NAND U9488 ( .A(n6107), .B(nreg[695]), .Z(n8132) );
  XOR U9489 ( .A(n8133), .B(n8134), .Z(n8127) );
  ANDN U9490 ( .A(n8135), .B(n4781), .Z(n8134) );
  XOR U9491 ( .A(n8136), .B(n8137), .Z(n4781) );
  IV U9492 ( .A(n8133), .Z(n8136) );
  XNOR U9493 ( .A(n4782), .B(n8133), .Z(n8135) );
  NAND U9494 ( .A(n8138), .B(nreg[694]), .Z(n4782) );
  NAND U9495 ( .A(n6107), .B(nreg[694]), .Z(n8138) );
  XOR U9496 ( .A(n8139), .B(n8140), .Z(n8133) );
  ANDN U9497 ( .A(n8141), .B(n4783), .Z(n8140) );
  XOR U9498 ( .A(n8142), .B(n8143), .Z(n4783) );
  IV U9499 ( .A(n8139), .Z(n8142) );
  XNOR U9500 ( .A(n4784), .B(n8139), .Z(n8141) );
  NAND U9501 ( .A(n8144), .B(nreg[693]), .Z(n4784) );
  NAND U9502 ( .A(n6107), .B(nreg[693]), .Z(n8144) );
  XOR U9503 ( .A(n8145), .B(n8146), .Z(n8139) );
  ANDN U9504 ( .A(n8147), .B(n4785), .Z(n8146) );
  XOR U9505 ( .A(n8148), .B(n8149), .Z(n4785) );
  IV U9506 ( .A(n8145), .Z(n8148) );
  XNOR U9507 ( .A(n4786), .B(n8145), .Z(n8147) );
  NAND U9508 ( .A(n8150), .B(nreg[692]), .Z(n4786) );
  NAND U9509 ( .A(n6107), .B(nreg[692]), .Z(n8150) );
  XOR U9510 ( .A(n8151), .B(n8152), .Z(n8145) );
  ANDN U9511 ( .A(n8153), .B(n4787), .Z(n8152) );
  XOR U9512 ( .A(n8154), .B(n8155), .Z(n4787) );
  IV U9513 ( .A(n8151), .Z(n8154) );
  XNOR U9514 ( .A(n4788), .B(n8151), .Z(n8153) );
  NAND U9515 ( .A(n8156), .B(nreg[691]), .Z(n4788) );
  NAND U9516 ( .A(n6107), .B(nreg[691]), .Z(n8156) );
  XOR U9517 ( .A(n8157), .B(n8158), .Z(n8151) );
  ANDN U9518 ( .A(n8159), .B(n4789), .Z(n8158) );
  XOR U9519 ( .A(n8160), .B(n8161), .Z(n4789) );
  IV U9520 ( .A(n8157), .Z(n8160) );
  XNOR U9521 ( .A(n4790), .B(n8157), .Z(n8159) );
  NAND U9522 ( .A(n8162), .B(nreg[690]), .Z(n4790) );
  NAND U9523 ( .A(n6107), .B(nreg[690]), .Z(n8162) );
  XOR U9524 ( .A(n8163), .B(n8164), .Z(n8157) );
  ANDN U9525 ( .A(n8165), .B(n4791), .Z(n8164) );
  XOR U9526 ( .A(n8166), .B(n8167), .Z(n4791) );
  IV U9527 ( .A(n8163), .Z(n8166) );
  XNOR U9528 ( .A(n4792), .B(n8163), .Z(n8165) );
  NAND U9529 ( .A(n8168), .B(nreg[689]), .Z(n4792) );
  NAND U9530 ( .A(n6107), .B(nreg[689]), .Z(n8168) );
  XOR U9531 ( .A(n8169), .B(n8170), .Z(n8163) );
  ANDN U9532 ( .A(n8171), .B(n4793), .Z(n8170) );
  XOR U9533 ( .A(n8172), .B(n8173), .Z(n4793) );
  IV U9534 ( .A(n8169), .Z(n8172) );
  XNOR U9535 ( .A(n4794), .B(n8169), .Z(n8171) );
  NAND U9536 ( .A(n8174), .B(nreg[688]), .Z(n4794) );
  NAND U9537 ( .A(n6107), .B(nreg[688]), .Z(n8174) );
  XOR U9538 ( .A(n8175), .B(n8176), .Z(n8169) );
  ANDN U9539 ( .A(n8177), .B(n4795), .Z(n8176) );
  XOR U9540 ( .A(n8178), .B(n8179), .Z(n4795) );
  IV U9541 ( .A(n8175), .Z(n8178) );
  XNOR U9542 ( .A(n4796), .B(n8175), .Z(n8177) );
  NAND U9543 ( .A(n8180), .B(nreg[687]), .Z(n4796) );
  NAND U9544 ( .A(n6107), .B(nreg[687]), .Z(n8180) );
  XOR U9545 ( .A(n8181), .B(n8182), .Z(n8175) );
  ANDN U9546 ( .A(n8183), .B(n4799), .Z(n8182) );
  XOR U9547 ( .A(n8184), .B(n8185), .Z(n4799) );
  IV U9548 ( .A(n8181), .Z(n8184) );
  XNOR U9549 ( .A(n4800), .B(n8181), .Z(n8183) );
  NAND U9550 ( .A(n8186), .B(nreg[686]), .Z(n4800) );
  NAND U9551 ( .A(n6107), .B(nreg[686]), .Z(n8186) );
  XOR U9552 ( .A(n8187), .B(n8188), .Z(n8181) );
  ANDN U9553 ( .A(n8189), .B(n4801), .Z(n8188) );
  XOR U9554 ( .A(n8190), .B(n8191), .Z(n4801) );
  IV U9555 ( .A(n8187), .Z(n8190) );
  XNOR U9556 ( .A(n4802), .B(n8187), .Z(n8189) );
  NAND U9557 ( .A(n8192), .B(nreg[685]), .Z(n4802) );
  NAND U9558 ( .A(n6107), .B(nreg[685]), .Z(n8192) );
  XOR U9559 ( .A(n8193), .B(n8194), .Z(n8187) );
  ANDN U9560 ( .A(n8195), .B(n4803), .Z(n8194) );
  XOR U9561 ( .A(n8196), .B(n8197), .Z(n4803) );
  IV U9562 ( .A(n8193), .Z(n8196) );
  XNOR U9563 ( .A(n4804), .B(n8193), .Z(n8195) );
  NAND U9564 ( .A(n8198), .B(nreg[684]), .Z(n4804) );
  NAND U9565 ( .A(n6107), .B(nreg[684]), .Z(n8198) );
  XOR U9566 ( .A(n8199), .B(n8200), .Z(n8193) );
  ANDN U9567 ( .A(n8201), .B(n4805), .Z(n8200) );
  XOR U9568 ( .A(n8202), .B(n8203), .Z(n4805) );
  IV U9569 ( .A(n8199), .Z(n8202) );
  XNOR U9570 ( .A(n4806), .B(n8199), .Z(n8201) );
  NAND U9571 ( .A(n8204), .B(nreg[683]), .Z(n4806) );
  NAND U9572 ( .A(n6107), .B(nreg[683]), .Z(n8204) );
  XOR U9573 ( .A(n8205), .B(n8206), .Z(n8199) );
  ANDN U9574 ( .A(n8207), .B(n4807), .Z(n8206) );
  XOR U9575 ( .A(n8208), .B(n8209), .Z(n4807) );
  IV U9576 ( .A(n8205), .Z(n8208) );
  XNOR U9577 ( .A(n4808), .B(n8205), .Z(n8207) );
  NAND U9578 ( .A(n8210), .B(nreg[682]), .Z(n4808) );
  NAND U9579 ( .A(n6107), .B(nreg[682]), .Z(n8210) );
  XOR U9580 ( .A(n8211), .B(n8212), .Z(n8205) );
  ANDN U9581 ( .A(n8213), .B(n4809), .Z(n8212) );
  XOR U9582 ( .A(n8214), .B(n8215), .Z(n4809) );
  IV U9583 ( .A(n8211), .Z(n8214) );
  XNOR U9584 ( .A(n4810), .B(n8211), .Z(n8213) );
  NAND U9585 ( .A(n8216), .B(nreg[681]), .Z(n4810) );
  NAND U9586 ( .A(n6107), .B(nreg[681]), .Z(n8216) );
  XOR U9587 ( .A(n8217), .B(n8218), .Z(n8211) );
  ANDN U9588 ( .A(n8219), .B(n4811), .Z(n8218) );
  XOR U9589 ( .A(n8220), .B(n8221), .Z(n4811) );
  IV U9590 ( .A(n8217), .Z(n8220) );
  XNOR U9591 ( .A(n4812), .B(n8217), .Z(n8219) );
  NAND U9592 ( .A(n8222), .B(nreg[680]), .Z(n4812) );
  NAND U9593 ( .A(n6107), .B(nreg[680]), .Z(n8222) );
  XOR U9594 ( .A(n8223), .B(n8224), .Z(n8217) );
  ANDN U9595 ( .A(n8225), .B(n4813), .Z(n8224) );
  XOR U9596 ( .A(n8226), .B(n8227), .Z(n4813) );
  IV U9597 ( .A(n8223), .Z(n8226) );
  XNOR U9598 ( .A(n4814), .B(n8223), .Z(n8225) );
  NAND U9599 ( .A(n8228), .B(nreg[679]), .Z(n4814) );
  NAND U9600 ( .A(n6107), .B(nreg[679]), .Z(n8228) );
  XOR U9601 ( .A(n8229), .B(n8230), .Z(n8223) );
  ANDN U9602 ( .A(n8231), .B(n4815), .Z(n8230) );
  XOR U9603 ( .A(n8232), .B(n8233), .Z(n4815) );
  IV U9604 ( .A(n8229), .Z(n8232) );
  XNOR U9605 ( .A(n4816), .B(n8229), .Z(n8231) );
  NAND U9606 ( .A(n8234), .B(nreg[678]), .Z(n4816) );
  NAND U9607 ( .A(n6107), .B(nreg[678]), .Z(n8234) );
  XOR U9608 ( .A(n8235), .B(n8236), .Z(n8229) );
  ANDN U9609 ( .A(n8237), .B(n4817), .Z(n8236) );
  XOR U9610 ( .A(n8238), .B(n8239), .Z(n4817) );
  IV U9611 ( .A(n8235), .Z(n8238) );
  XNOR U9612 ( .A(n4818), .B(n8235), .Z(n8237) );
  NAND U9613 ( .A(n8240), .B(nreg[677]), .Z(n4818) );
  NAND U9614 ( .A(n6107), .B(nreg[677]), .Z(n8240) );
  XOR U9615 ( .A(n8241), .B(n8242), .Z(n8235) );
  ANDN U9616 ( .A(n8243), .B(n4821), .Z(n8242) );
  XOR U9617 ( .A(n8244), .B(n8245), .Z(n4821) );
  IV U9618 ( .A(n8241), .Z(n8244) );
  XNOR U9619 ( .A(n4822), .B(n8241), .Z(n8243) );
  NAND U9620 ( .A(n8246), .B(nreg[676]), .Z(n4822) );
  NAND U9621 ( .A(n6107), .B(nreg[676]), .Z(n8246) );
  XOR U9622 ( .A(n8247), .B(n8248), .Z(n8241) );
  ANDN U9623 ( .A(n8249), .B(n4823), .Z(n8248) );
  XOR U9624 ( .A(n8250), .B(n8251), .Z(n4823) );
  IV U9625 ( .A(n8247), .Z(n8250) );
  XNOR U9626 ( .A(n4824), .B(n8247), .Z(n8249) );
  NAND U9627 ( .A(n8252), .B(nreg[675]), .Z(n4824) );
  NAND U9628 ( .A(n6107), .B(nreg[675]), .Z(n8252) );
  XOR U9629 ( .A(n8253), .B(n8254), .Z(n8247) );
  ANDN U9630 ( .A(n8255), .B(n4825), .Z(n8254) );
  XOR U9631 ( .A(n8256), .B(n8257), .Z(n4825) );
  IV U9632 ( .A(n8253), .Z(n8256) );
  XNOR U9633 ( .A(n4826), .B(n8253), .Z(n8255) );
  NAND U9634 ( .A(n8258), .B(nreg[674]), .Z(n4826) );
  NAND U9635 ( .A(n6107), .B(nreg[674]), .Z(n8258) );
  XOR U9636 ( .A(n8259), .B(n8260), .Z(n8253) );
  ANDN U9637 ( .A(n8261), .B(n4827), .Z(n8260) );
  XOR U9638 ( .A(n8262), .B(n8263), .Z(n4827) );
  IV U9639 ( .A(n8259), .Z(n8262) );
  XNOR U9640 ( .A(n4828), .B(n8259), .Z(n8261) );
  NAND U9641 ( .A(n8264), .B(nreg[673]), .Z(n4828) );
  NAND U9642 ( .A(n6107), .B(nreg[673]), .Z(n8264) );
  XOR U9643 ( .A(n8265), .B(n8266), .Z(n8259) );
  ANDN U9644 ( .A(n8267), .B(n4829), .Z(n8266) );
  XOR U9645 ( .A(n8268), .B(n8269), .Z(n4829) );
  IV U9646 ( .A(n8265), .Z(n8268) );
  XNOR U9647 ( .A(n4830), .B(n8265), .Z(n8267) );
  NAND U9648 ( .A(n8270), .B(nreg[672]), .Z(n4830) );
  NAND U9649 ( .A(n6107), .B(nreg[672]), .Z(n8270) );
  XOR U9650 ( .A(n8271), .B(n8272), .Z(n8265) );
  ANDN U9651 ( .A(n8273), .B(n4831), .Z(n8272) );
  XOR U9652 ( .A(n8274), .B(n8275), .Z(n4831) );
  IV U9653 ( .A(n8271), .Z(n8274) );
  XNOR U9654 ( .A(n4832), .B(n8271), .Z(n8273) );
  NAND U9655 ( .A(n8276), .B(nreg[671]), .Z(n4832) );
  NAND U9656 ( .A(n6107), .B(nreg[671]), .Z(n8276) );
  XOR U9657 ( .A(n8277), .B(n8278), .Z(n8271) );
  ANDN U9658 ( .A(n8279), .B(n4833), .Z(n8278) );
  XOR U9659 ( .A(n8280), .B(n8281), .Z(n4833) );
  IV U9660 ( .A(n8277), .Z(n8280) );
  XNOR U9661 ( .A(n4834), .B(n8277), .Z(n8279) );
  NAND U9662 ( .A(n8282), .B(nreg[670]), .Z(n4834) );
  NAND U9663 ( .A(n6107), .B(nreg[670]), .Z(n8282) );
  XOR U9664 ( .A(n8283), .B(n8284), .Z(n8277) );
  ANDN U9665 ( .A(n8285), .B(n4835), .Z(n8284) );
  XOR U9666 ( .A(n8286), .B(n8287), .Z(n4835) );
  IV U9667 ( .A(n8283), .Z(n8286) );
  XNOR U9668 ( .A(n4836), .B(n8283), .Z(n8285) );
  NAND U9669 ( .A(n8288), .B(nreg[669]), .Z(n4836) );
  NAND U9670 ( .A(n6107), .B(nreg[669]), .Z(n8288) );
  XOR U9671 ( .A(n8289), .B(n8290), .Z(n8283) );
  ANDN U9672 ( .A(n8291), .B(n4837), .Z(n8290) );
  XOR U9673 ( .A(n8292), .B(n8293), .Z(n4837) );
  IV U9674 ( .A(n8289), .Z(n8292) );
  XNOR U9675 ( .A(n4838), .B(n8289), .Z(n8291) );
  NAND U9676 ( .A(n8294), .B(nreg[668]), .Z(n4838) );
  NAND U9677 ( .A(n6107), .B(nreg[668]), .Z(n8294) );
  XOR U9678 ( .A(n8295), .B(n8296), .Z(n8289) );
  ANDN U9679 ( .A(n8297), .B(n4839), .Z(n8296) );
  XOR U9680 ( .A(n8298), .B(n8299), .Z(n4839) );
  IV U9681 ( .A(n8295), .Z(n8298) );
  XNOR U9682 ( .A(n4840), .B(n8295), .Z(n8297) );
  NAND U9683 ( .A(n8300), .B(nreg[667]), .Z(n4840) );
  NAND U9684 ( .A(n6107), .B(nreg[667]), .Z(n8300) );
  XOR U9685 ( .A(n8301), .B(n8302), .Z(n8295) );
  ANDN U9686 ( .A(n8303), .B(n4843), .Z(n8302) );
  XOR U9687 ( .A(n8304), .B(n8305), .Z(n4843) );
  IV U9688 ( .A(n8301), .Z(n8304) );
  XNOR U9689 ( .A(n4844), .B(n8301), .Z(n8303) );
  NAND U9690 ( .A(n8306), .B(nreg[666]), .Z(n4844) );
  NAND U9691 ( .A(n6107), .B(nreg[666]), .Z(n8306) );
  XOR U9692 ( .A(n8307), .B(n8308), .Z(n8301) );
  ANDN U9693 ( .A(n8309), .B(n4845), .Z(n8308) );
  XOR U9694 ( .A(n8310), .B(n8311), .Z(n4845) );
  IV U9695 ( .A(n8307), .Z(n8310) );
  XNOR U9696 ( .A(n4846), .B(n8307), .Z(n8309) );
  NAND U9697 ( .A(n8312), .B(nreg[665]), .Z(n4846) );
  NAND U9698 ( .A(n6107), .B(nreg[665]), .Z(n8312) );
  XOR U9699 ( .A(n8313), .B(n8314), .Z(n8307) );
  ANDN U9700 ( .A(n8315), .B(n4847), .Z(n8314) );
  XOR U9701 ( .A(n8316), .B(n8317), .Z(n4847) );
  IV U9702 ( .A(n8313), .Z(n8316) );
  XNOR U9703 ( .A(n4848), .B(n8313), .Z(n8315) );
  NAND U9704 ( .A(n8318), .B(nreg[664]), .Z(n4848) );
  NAND U9705 ( .A(n6107), .B(nreg[664]), .Z(n8318) );
  XOR U9706 ( .A(n8319), .B(n8320), .Z(n8313) );
  ANDN U9707 ( .A(n8321), .B(n4849), .Z(n8320) );
  XOR U9708 ( .A(n8322), .B(n8323), .Z(n4849) );
  IV U9709 ( .A(n8319), .Z(n8322) );
  XNOR U9710 ( .A(n4850), .B(n8319), .Z(n8321) );
  NAND U9711 ( .A(n8324), .B(nreg[663]), .Z(n4850) );
  NAND U9712 ( .A(n6107), .B(nreg[663]), .Z(n8324) );
  XOR U9713 ( .A(n8325), .B(n8326), .Z(n8319) );
  ANDN U9714 ( .A(n8327), .B(n4851), .Z(n8326) );
  XOR U9715 ( .A(n8328), .B(n8329), .Z(n4851) );
  IV U9716 ( .A(n8325), .Z(n8328) );
  XNOR U9717 ( .A(n4852), .B(n8325), .Z(n8327) );
  NAND U9718 ( .A(n8330), .B(nreg[662]), .Z(n4852) );
  NAND U9719 ( .A(n6107), .B(nreg[662]), .Z(n8330) );
  XOR U9720 ( .A(n8331), .B(n8332), .Z(n8325) );
  ANDN U9721 ( .A(n8333), .B(n4853), .Z(n8332) );
  XOR U9722 ( .A(n8334), .B(n8335), .Z(n4853) );
  IV U9723 ( .A(n8331), .Z(n8334) );
  XNOR U9724 ( .A(n4854), .B(n8331), .Z(n8333) );
  NAND U9725 ( .A(n8336), .B(nreg[661]), .Z(n4854) );
  NAND U9726 ( .A(n6107), .B(nreg[661]), .Z(n8336) );
  XOR U9727 ( .A(n8337), .B(n8338), .Z(n8331) );
  ANDN U9728 ( .A(n8339), .B(n4855), .Z(n8338) );
  XOR U9729 ( .A(n8340), .B(n8341), .Z(n4855) );
  IV U9730 ( .A(n8337), .Z(n8340) );
  XNOR U9731 ( .A(n4856), .B(n8337), .Z(n8339) );
  NAND U9732 ( .A(n8342), .B(nreg[660]), .Z(n4856) );
  NAND U9733 ( .A(n6107), .B(nreg[660]), .Z(n8342) );
  XOR U9734 ( .A(n8343), .B(n8344), .Z(n8337) );
  ANDN U9735 ( .A(n8345), .B(n4857), .Z(n8344) );
  XOR U9736 ( .A(n8346), .B(n8347), .Z(n4857) );
  IV U9737 ( .A(n8343), .Z(n8346) );
  XNOR U9738 ( .A(n4858), .B(n8343), .Z(n8345) );
  NAND U9739 ( .A(n8348), .B(nreg[659]), .Z(n4858) );
  NAND U9740 ( .A(n6107), .B(nreg[659]), .Z(n8348) );
  XOR U9741 ( .A(n8349), .B(n8350), .Z(n8343) );
  ANDN U9742 ( .A(n8351), .B(n4859), .Z(n8350) );
  XOR U9743 ( .A(n8352), .B(n8353), .Z(n4859) );
  IV U9744 ( .A(n8349), .Z(n8352) );
  XNOR U9745 ( .A(n4860), .B(n8349), .Z(n8351) );
  NAND U9746 ( .A(n8354), .B(nreg[658]), .Z(n4860) );
  NAND U9747 ( .A(n6107), .B(nreg[658]), .Z(n8354) );
  XOR U9748 ( .A(n8355), .B(n8356), .Z(n8349) );
  ANDN U9749 ( .A(n8357), .B(n4861), .Z(n8356) );
  XOR U9750 ( .A(n8358), .B(n8359), .Z(n4861) );
  IV U9751 ( .A(n8355), .Z(n8358) );
  XNOR U9752 ( .A(n4862), .B(n8355), .Z(n8357) );
  NAND U9753 ( .A(n8360), .B(nreg[657]), .Z(n4862) );
  NAND U9754 ( .A(n6107), .B(nreg[657]), .Z(n8360) );
  XOR U9755 ( .A(n8361), .B(n8362), .Z(n8355) );
  ANDN U9756 ( .A(n8363), .B(n4865), .Z(n8362) );
  XOR U9757 ( .A(n8364), .B(n8365), .Z(n4865) );
  IV U9758 ( .A(n8361), .Z(n8364) );
  XNOR U9759 ( .A(n4866), .B(n8361), .Z(n8363) );
  NAND U9760 ( .A(n8366), .B(nreg[656]), .Z(n4866) );
  NAND U9761 ( .A(n6107), .B(nreg[656]), .Z(n8366) );
  XOR U9762 ( .A(n8367), .B(n8368), .Z(n8361) );
  ANDN U9763 ( .A(n8369), .B(n4867), .Z(n8368) );
  XOR U9764 ( .A(n8370), .B(n8371), .Z(n4867) );
  IV U9765 ( .A(n8367), .Z(n8370) );
  XNOR U9766 ( .A(n4868), .B(n8367), .Z(n8369) );
  NAND U9767 ( .A(n8372), .B(nreg[655]), .Z(n4868) );
  NAND U9768 ( .A(n6107), .B(nreg[655]), .Z(n8372) );
  XOR U9769 ( .A(n8373), .B(n8374), .Z(n8367) );
  ANDN U9770 ( .A(n8375), .B(n4869), .Z(n8374) );
  XOR U9771 ( .A(n8376), .B(n8377), .Z(n4869) );
  IV U9772 ( .A(n8373), .Z(n8376) );
  XNOR U9773 ( .A(n4870), .B(n8373), .Z(n8375) );
  NAND U9774 ( .A(n8378), .B(nreg[654]), .Z(n4870) );
  NAND U9775 ( .A(n6107), .B(nreg[654]), .Z(n8378) );
  XOR U9776 ( .A(n8379), .B(n8380), .Z(n8373) );
  ANDN U9777 ( .A(n8381), .B(n4871), .Z(n8380) );
  XOR U9778 ( .A(n8382), .B(n8383), .Z(n4871) );
  IV U9779 ( .A(n8379), .Z(n8382) );
  XNOR U9780 ( .A(n4872), .B(n8379), .Z(n8381) );
  NAND U9781 ( .A(n8384), .B(nreg[653]), .Z(n4872) );
  NAND U9782 ( .A(n6107), .B(nreg[653]), .Z(n8384) );
  XOR U9783 ( .A(n8385), .B(n8386), .Z(n8379) );
  ANDN U9784 ( .A(n8387), .B(n4873), .Z(n8386) );
  XOR U9785 ( .A(n8388), .B(n8389), .Z(n4873) );
  IV U9786 ( .A(n8385), .Z(n8388) );
  XNOR U9787 ( .A(n4874), .B(n8385), .Z(n8387) );
  NAND U9788 ( .A(n8390), .B(nreg[652]), .Z(n4874) );
  NAND U9789 ( .A(n6107), .B(nreg[652]), .Z(n8390) );
  XOR U9790 ( .A(n8391), .B(n8392), .Z(n8385) );
  ANDN U9791 ( .A(n8393), .B(n4875), .Z(n8392) );
  XOR U9792 ( .A(n8394), .B(n8395), .Z(n4875) );
  IV U9793 ( .A(n8391), .Z(n8394) );
  XNOR U9794 ( .A(n4876), .B(n8391), .Z(n8393) );
  NAND U9795 ( .A(n8396), .B(nreg[651]), .Z(n4876) );
  NAND U9796 ( .A(n6107), .B(nreg[651]), .Z(n8396) );
  XOR U9797 ( .A(n8397), .B(n8398), .Z(n8391) );
  ANDN U9798 ( .A(n8399), .B(n4877), .Z(n8398) );
  XOR U9799 ( .A(n8400), .B(n8401), .Z(n4877) );
  IV U9800 ( .A(n8397), .Z(n8400) );
  XNOR U9801 ( .A(n4878), .B(n8397), .Z(n8399) );
  NAND U9802 ( .A(n8402), .B(nreg[650]), .Z(n4878) );
  NAND U9803 ( .A(n6107), .B(nreg[650]), .Z(n8402) );
  XOR U9804 ( .A(n8403), .B(n8404), .Z(n8397) );
  ANDN U9805 ( .A(n8405), .B(n4879), .Z(n8404) );
  XOR U9806 ( .A(n8406), .B(n8407), .Z(n4879) );
  IV U9807 ( .A(n8403), .Z(n8406) );
  XNOR U9808 ( .A(n4880), .B(n8403), .Z(n8405) );
  NAND U9809 ( .A(n8408), .B(nreg[649]), .Z(n4880) );
  NAND U9810 ( .A(n6107), .B(nreg[649]), .Z(n8408) );
  XOR U9811 ( .A(n8409), .B(n8410), .Z(n8403) );
  ANDN U9812 ( .A(n8411), .B(n4881), .Z(n8410) );
  XOR U9813 ( .A(n8412), .B(n8413), .Z(n4881) );
  IV U9814 ( .A(n8409), .Z(n8412) );
  XNOR U9815 ( .A(n4882), .B(n8409), .Z(n8411) );
  NAND U9816 ( .A(n8414), .B(nreg[648]), .Z(n4882) );
  NAND U9817 ( .A(n6107), .B(nreg[648]), .Z(n8414) );
  XOR U9818 ( .A(n8415), .B(n8416), .Z(n8409) );
  ANDN U9819 ( .A(n8417), .B(n4883), .Z(n8416) );
  XOR U9820 ( .A(n8418), .B(n8419), .Z(n4883) );
  IV U9821 ( .A(n8415), .Z(n8418) );
  XNOR U9822 ( .A(n4884), .B(n8415), .Z(n8417) );
  NAND U9823 ( .A(n8420), .B(nreg[647]), .Z(n4884) );
  NAND U9824 ( .A(n6107), .B(nreg[647]), .Z(n8420) );
  XOR U9825 ( .A(n8421), .B(n8422), .Z(n8415) );
  ANDN U9826 ( .A(n8423), .B(n4887), .Z(n8422) );
  XOR U9827 ( .A(n8424), .B(n8425), .Z(n4887) );
  IV U9828 ( .A(n8421), .Z(n8424) );
  XNOR U9829 ( .A(n4888), .B(n8421), .Z(n8423) );
  NAND U9830 ( .A(n8426), .B(nreg[646]), .Z(n4888) );
  NAND U9831 ( .A(n6107), .B(nreg[646]), .Z(n8426) );
  XOR U9832 ( .A(n8427), .B(n8428), .Z(n8421) );
  ANDN U9833 ( .A(n8429), .B(n4889), .Z(n8428) );
  XOR U9834 ( .A(n8430), .B(n8431), .Z(n4889) );
  IV U9835 ( .A(n8427), .Z(n8430) );
  XNOR U9836 ( .A(n4890), .B(n8427), .Z(n8429) );
  NAND U9837 ( .A(n8432), .B(nreg[645]), .Z(n4890) );
  NAND U9838 ( .A(n6107), .B(nreg[645]), .Z(n8432) );
  XOR U9839 ( .A(n8433), .B(n8434), .Z(n8427) );
  ANDN U9840 ( .A(n8435), .B(n4891), .Z(n8434) );
  XOR U9841 ( .A(n8436), .B(n8437), .Z(n4891) );
  IV U9842 ( .A(n8433), .Z(n8436) );
  XNOR U9843 ( .A(n4892), .B(n8433), .Z(n8435) );
  NAND U9844 ( .A(n8438), .B(nreg[644]), .Z(n4892) );
  NAND U9845 ( .A(n6107), .B(nreg[644]), .Z(n8438) );
  XOR U9846 ( .A(n8439), .B(n8440), .Z(n8433) );
  ANDN U9847 ( .A(n8441), .B(n4893), .Z(n8440) );
  XOR U9848 ( .A(n8442), .B(n8443), .Z(n4893) );
  IV U9849 ( .A(n8439), .Z(n8442) );
  XNOR U9850 ( .A(n4894), .B(n8439), .Z(n8441) );
  NAND U9851 ( .A(n8444), .B(nreg[643]), .Z(n4894) );
  NAND U9852 ( .A(n6107), .B(nreg[643]), .Z(n8444) );
  XOR U9853 ( .A(n8445), .B(n8446), .Z(n8439) );
  ANDN U9854 ( .A(n8447), .B(n4895), .Z(n8446) );
  XOR U9855 ( .A(n8448), .B(n8449), .Z(n4895) );
  IV U9856 ( .A(n8445), .Z(n8448) );
  XNOR U9857 ( .A(n4896), .B(n8445), .Z(n8447) );
  NAND U9858 ( .A(n8450), .B(nreg[642]), .Z(n4896) );
  NAND U9859 ( .A(n6107), .B(nreg[642]), .Z(n8450) );
  XOR U9860 ( .A(n8451), .B(n8452), .Z(n8445) );
  ANDN U9861 ( .A(n8453), .B(n4897), .Z(n8452) );
  XOR U9862 ( .A(n8454), .B(n8455), .Z(n4897) );
  IV U9863 ( .A(n8451), .Z(n8454) );
  XNOR U9864 ( .A(n4898), .B(n8451), .Z(n8453) );
  NAND U9865 ( .A(n8456), .B(nreg[641]), .Z(n4898) );
  NAND U9866 ( .A(n6107), .B(nreg[641]), .Z(n8456) );
  XOR U9867 ( .A(n8457), .B(n8458), .Z(n8451) );
  ANDN U9868 ( .A(n8459), .B(n4899), .Z(n8458) );
  XOR U9869 ( .A(n8460), .B(n8461), .Z(n4899) );
  IV U9870 ( .A(n8457), .Z(n8460) );
  XNOR U9871 ( .A(n4900), .B(n8457), .Z(n8459) );
  NAND U9872 ( .A(n8462), .B(nreg[640]), .Z(n4900) );
  NAND U9873 ( .A(n6107), .B(nreg[640]), .Z(n8462) );
  XOR U9874 ( .A(n8463), .B(n8464), .Z(n8457) );
  ANDN U9875 ( .A(n8465), .B(n4901), .Z(n8464) );
  XOR U9876 ( .A(n8466), .B(n8467), .Z(n4901) );
  IV U9877 ( .A(n8463), .Z(n8466) );
  XNOR U9878 ( .A(n4902), .B(n8463), .Z(n8465) );
  NAND U9879 ( .A(n8468), .B(nreg[639]), .Z(n4902) );
  NAND U9880 ( .A(n6107), .B(nreg[639]), .Z(n8468) );
  XOR U9881 ( .A(n8469), .B(n8470), .Z(n8463) );
  ANDN U9882 ( .A(n8471), .B(n4903), .Z(n8470) );
  XOR U9883 ( .A(n8472), .B(n8473), .Z(n4903) );
  IV U9884 ( .A(n8469), .Z(n8472) );
  XNOR U9885 ( .A(n4904), .B(n8469), .Z(n8471) );
  NAND U9886 ( .A(n8474), .B(nreg[638]), .Z(n4904) );
  NAND U9887 ( .A(n6107), .B(nreg[638]), .Z(n8474) );
  XOR U9888 ( .A(n8475), .B(n8476), .Z(n8469) );
  ANDN U9889 ( .A(n8477), .B(n4905), .Z(n8476) );
  XOR U9890 ( .A(n8478), .B(n8479), .Z(n4905) );
  IV U9891 ( .A(n8475), .Z(n8478) );
  XNOR U9892 ( .A(n4906), .B(n8475), .Z(n8477) );
  NAND U9893 ( .A(n8480), .B(nreg[637]), .Z(n4906) );
  NAND U9894 ( .A(n6107), .B(nreg[637]), .Z(n8480) );
  XOR U9895 ( .A(n8481), .B(n8482), .Z(n8475) );
  ANDN U9896 ( .A(n8483), .B(n4909), .Z(n8482) );
  XOR U9897 ( .A(n8484), .B(n8485), .Z(n4909) );
  IV U9898 ( .A(n8481), .Z(n8484) );
  XNOR U9899 ( .A(n4910), .B(n8481), .Z(n8483) );
  NAND U9900 ( .A(n8486), .B(nreg[636]), .Z(n4910) );
  NAND U9901 ( .A(n6107), .B(nreg[636]), .Z(n8486) );
  XOR U9902 ( .A(n8487), .B(n8488), .Z(n8481) );
  ANDN U9903 ( .A(n8489), .B(n4911), .Z(n8488) );
  XOR U9904 ( .A(n8490), .B(n8491), .Z(n4911) );
  IV U9905 ( .A(n8487), .Z(n8490) );
  XNOR U9906 ( .A(n4912), .B(n8487), .Z(n8489) );
  NAND U9907 ( .A(n8492), .B(nreg[635]), .Z(n4912) );
  NAND U9908 ( .A(n6107), .B(nreg[635]), .Z(n8492) );
  XOR U9909 ( .A(n8493), .B(n8494), .Z(n8487) );
  ANDN U9910 ( .A(n8495), .B(n4913), .Z(n8494) );
  XOR U9911 ( .A(n8496), .B(n8497), .Z(n4913) );
  IV U9912 ( .A(n8493), .Z(n8496) );
  XNOR U9913 ( .A(n4914), .B(n8493), .Z(n8495) );
  NAND U9914 ( .A(n8498), .B(nreg[634]), .Z(n4914) );
  NAND U9915 ( .A(n6107), .B(nreg[634]), .Z(n8498) );
  XOR U9916 ( .A(n8499), .B(n8500), .Z(n8493) );
  ANDN U9917 ( .A(n8501), .B(n4915), .Z(n8500) );
  XOR U9918 ( .A(n8502), .B(n8503), .Z(n4915) );
  IV U9919 ( .A(n8499), .Z(n8502) );
  XNOR U9920 ( .A(n4916), .B(n8499), .Z(n8501) );
  NAND U9921 ( .A(n8504), .B(nreg[633]), .Z(n4916) );
  NAND U9922 ( .A(n6107), .B(nreg[633]), .Z(n8504) );
  XOR U9923 ( .A(n8505), .B(n8506), .Z(n8499) );
  ANDN U9924 ( .A(n8507), .B(n4917), .Z(n8506) );
  XOR U9925 ( .A(n8508), .B(n8509), .Z(n4917) );
  IV U9926 ( .A(n8505), .Z(n8508) );
  XNOR U9927 ( .A(n4918), .B(n8505), .Z(n8507) );
  NAND U9928 ( .A(n8510), .B(nreg[632]), .Z(n4918) );
  NAND U9929 ( .A(n6107), .B(nreg[632]), .Z(n8510) );
  XOR U9930 ( .A(n8511), .B(n8512), .Z(n8505) );
  ANDN U9931 ( .A(n8513), .B(n4919), .Z(n8512) );
  XOR U9932 ( .A(n8514), .B(n8515), .Z(n4919) );
  IV U9933 ( .A(n8511), .Z(n8514) );
  XNOR U9934 ( .A(n4920), .B(n8511), .Z(n8513) );
  NAND U9935 ( .A(n8516), .B(nreg[631]), .Z(n4920) );
  NAND U9936 ( .A(n6107), .B(nreg[631]), .Z(n8516) );
  XOR U9937 ( .A(n8517), .B(n8518), .Z(n8511) );
  ANDN U9938 ( .A(n8519), .B(n4921), .Z(n8518) );
  XOR U9939 ( .A(n8520), .B(n8521), .Z(n4921) );
  IV U9940 ( .A(n8517), .Z(n8520) );
  XNOR U9941 ( .A(n4922), .B(n8517), .Z(n8519) );
  NAND U9942 ( .A(n8522), .B(nreg[630]), .Z(n4922) );
  NAND U9943 ( .A(n6107), .B(nreg[630]), .Z(n8522) );
  XOR U9944 ( .A(n8523), .B(n8524), .Z(n8517) );
  ANDN U9945 ( .A(n8525), .B(n4923), .Z(n8524) );
  XOR U9946 ( .A(n8526), .B(n8527), .Z(n4923) );
  IV U9947 ( .A(n8523), .Z(n8526) );
  XNOR U9948 ( .A(n4924), .B(n8523), .Z(n8525) );
  NAND U9949 ( .A(n8528), .B(nreg[629]), .Z(n4924) );
  NAND U9950 ( .A(n6107), .B(nreg[629]), .Z(n8528) );
  XOR U9951 ( .A(n8529), .B(n8530), .Z(n8523) );
  ANDN U9952 ( .A(n8531), .B(n4925), .Z(n8530) );
  XOR U9953 ( .A(n8532), .B(n8533), .Z(n4925) );
  IV U9954 ( .A(n8529), .Z(n8532) );
  XNOR U9955 ( .A(n4926), .B(n8529), .Z(n8531) );
  NAND U9956 ( .A(n8534), .B(nreg[628]), .Z(n4926) );
  NAND U9957 ( .A(n6107), .B(nreg[628]), .Z(n8534) );
  XOR U9958 ( .A(n8535), .B(n8536), .Z(n8529) );
  ANDN U9959 ( .A(n8537), .B(n4927), .Z(n8536) );
  XOR U9960 ( .A(n8538), .B(n8539), .Z(n4927) );
  IV U9961 ( .A(n8535), .Z(n8538) );
  XNOR U9962 ( .A(n4928), .B(n8535), .Z(n8537) );
  NAND U9963 ( .A(n8540), .B(nreg[627]), .Z(n4928) );
  NAND U9964 ( .A(n6107), .B(nreg[627]), .Z(n8540) );
  XOR U9965 ( .A(n8541), .B(n8542), .Z(n8535) );
  ANDN U9966 ( .A(n8543), .B(n4931), .Z(n8542) );
  XOR U9967 ( .A(n8544), .B(n8545), .Z(n4931) );
  IV U9968 ( .A(n8541), .Z(n8544) );
  XNOR U9969 ( .A(n4932), .B(n8541), .Z(n8543) );
  NAND U9970 ( .A(n8546), .B(nreg[626]), .Z(n4932) );
  NAND U9971 ( .A(n6107), .B(nreg[626]), .Z(n8546) );
  XOR U9972 ( .A(n8547), .B(n8548), .Z(n8541) );
  ANDN U9973 ( .A(n8549), .B(n4933), .Z(n8548) );
  XOR U9974 ( .A(n8550), .B(n8551), .Z(n4933) );
  IV U9975 ( .A(n8547), .Z(n8550) );
  XNOR U9976 ( .A(n4934), .B(n8547), .Z(n8549) );
  NAND U9977 ( .A(n8552), .B(nreg[625]), .Z(n4934) );
  NAND U9978 ( .A(n6107), .B(nreg[625]), .Z(n8552) );
  XOR U9979 ( .A(n8553), .B(n8554), .Z(n8547) );
  ANDN U9980 ( .A(n8555), .B(n4935), .Z(n8554) );
  XOR U9981 ( .A(n8556), .B(n8557), .Z(n4935) );
  IV U9982 ( .A(n8553), .Z(n8556) );
  XNOR U9983 ( .A(n4936), .B(n8553), .Z(n8555) );
  NAND U9984 ( .A(n8558), .B(nreg[624]), .Z(n4936) );
  NAND U9985 ( .A(n6107), .B(nreg[624]), .Z(n8558) );
  XOR U9986 ( .A(n8559), .B(n8560), .Z(n8553) );
  ANDN U9987 ( .A(n8561), .B(n4937), .Z(n8560) );
  XOR U9988 ( .A(n8562), .B(n8563), .Z(n4937) );
  IV U9989 ( .A(n8559), .Z(n8562) );
  XNOR U9990 ( .A(n4938), .B(n8559), .Z(n8561) );
  NAND U9991 ( .A(n8564), .B(nreg[623]), .Z(n4938) );
  NAND U9992 ( .A(n6107), .B(nreg[623]), .Z(n8564) );
  XOR U9993 ( .A(n8565), .B(n8566), .Z(n8559) );
  ANDN U9994 ( .A(n8567), .B(n4939), .Z(n8566) );
  XOR U9995 ( .A(n8568), .B(n8569), .Z(n4939) );
  IV U9996 ( .A(n8565), .Z(n8568) );
  XNOR U9997 ( .A(n4940), .B(n8565), .Z(n8567) );
  NAND U9998 ( .A(n8570), .B(nreg[622]), .Z(n4940) );
  NAND U9999 ( .A(n6107), .B(nreg[622]), .Z(n8570) );
  XOR U10000 ( .A(n8571), .B(n8572), .Z(n8565) );
  ANDN U10001 ( .A(n8573), .B(n4941), .Z(n8572) );
  XOR U10002 ( .A(n8574), .B(n8575), .Z(n4941) );
  IV U10003 ( .A(n8571), .Z(n8574) );
  XNOR U10004 ( .A(n4942), .B(n8571), .Z(n8573) );
  NAND U10005 ( .A(n8576), .B(nreg[621]), .Z(n4942) );
  NAND U10006 ( .A(n6107), .B(nreg[621]), .Z(n8576) );
  XOR U10007 ( .A(n8577), .B(n8578), .Z(n8571) );
  ANDN U10008 ( .A(n8579), .B(n4943), .Z(n8578) );
  XOR U10009 ( .A(n8580), .B(n8581), .Z(n4943) );
  IV U10010 ( .A(n8577), .Z(n8580) );
  XNOR U10011 ( .A(n4944), .B(n8577), .Z(n8579) );
  NAND U10012 ( .A(n8582), .B(nreg[620]), .Z(n4944) );
  NAND U10013 ( .A(n6107), .B(nreg[620]), .Z(n8582) );
  XOR U10014 ( .A(n8583), .B(n8584), .Z(n8577) );
  ANDN U10015 ( .A(n8585), .B(n4945), .Z(n8584) );
  XOR U10016 ( .A(n8586), .B(n8587), .Z(n4945) );
  IV U10017 ( .A(n8583), .Z(n8586) );
  XNOR U10018 ( .A(n4946), .B(n8583), .Z(n8585) );
  NAND U10019 ( .A(n8588), .B(nreg[619]), .Z(n4946) );
  NAND U10020 ( .A(n6107), .B(nreg[619]), .Z(n8588) );
  XOR U10021 ( .A(n8589), .B(n8590), .Z(n8583) );
  ANDN U10022 ( .A(n8591), .B(n4947), .Z(n8590) );
  XOR U10023 ( .A(n8592), .B(n8593), .Z(n4947) );
  IV U10024 ( .A(n8589), .Z(n8592) );
  XNOR U10025 ( .A(n4948), .B(n8589), .Z(n8591) );
  NAND U10026 ( .A(n8594), .B(nreg[618]), .Z(n4948) );
  NAND U10027 ( .A(n6107), .B(nreg[618]), .Z(n8594) );
  XOR U10028 ( .A(n8595), .B(n8596), .Z(n8589) );
  ANDN U10029 ( .A(n8597), .B(n4949), .Z(n8596) );
  XOR U10030 ( .A(n8598), .B(n8599), .Z(n4949) );
  IV U10031 ( .A(n8595), .Z(n8598) );
  XNOR U10032 ( .A(n4950), .B(n8595), .Z(n8597) );
  NAND U10033 ( .A(n8600), .B(nreg[617]), .Z(n4950) );
  NAND U10034 ( .A(n6107), .B(nreg[617]), .Z(n8600) );
  XOR U10035 ( .A(n8601), .B(n8602), .Z(n8595) );
  ANDN U10036 ( .A(n8603), .B(n4953), .Z(n8602) );
  XOR U10037 ( .A(n8604), .B(n8605), .Z(n4953) );
  IV U10038 ( .A(n8601), .Z(n8604) );
  XNOR U10039 ( .A(n4954), .B(n8601), .Z(n8603) );
  NAND U10040 ( .A(n8606), .B(nreg[616]), .Z(n4954) );
  NAND U10041 ( .A(n6107), .B(nreg[616]), .Z(n8606) );
  XOR U10042 ( .A(n8607), .B(n8608), .Z(n8601) );
  ANDN U10043 ( .A(n8609), .B(n4955), .Z(n8608) );
  XOR U10044 ( .A(n8610), .B(n8611), .Z(n4955) );
  IV U10045 ( .A(n8607), .Z(n8610) );
  XNOR U10046 ( .A(n4956), .B(n8607), .Z(n8609) );
  NAND U10047 ( .A(n8612), .B(nreg[615]), .Z(n4956) );
  NAND U10048 ( .A(n6107), .B(nreg[615]), .Z(n8612) );
  XOR U10049 ( .A(n8613), .B(n8614), .Z(n8607) );
  ANDN U10050 ( .A(n8615), .B(n4957), .Z(n8614) );
  XOR U10051 ( .A(n8616), .B(n8617), .Z(n4957) );
  IV U10052 ( .A(n8613), .Z(n8616) );
  XNOR U10053 ( .A(n4958), .B(n8613), .Z(n8615) );
  NAND U10054 ( .A(n8618), .B(nreg[614]), .Z(n4958) );
  NAND U10055 ( .A(n6107), .B(nreg[614]), .Z(n8618) );
  XOR U10056 ( .A(n8619), .B(n8620), .Z(n8613) );
  ANDN U10057 ( .A(n8621), .B(n4959), .Z(n8620) );
  XOR U10058 ( .A(n8622), .B(n8623), .Z(n4959) );
  IV U10059 ( .A(n8619), .Z(n8622) );
  XNOR U10060 ( .A(n4960), .B(n8619), .Z(n8621) );
  NAND U10061 ( .A(n8624), .B(nreg[613]), .Z(n4960) );
  NAND U10062 ( .A(n6107), .B(nreg[613]), .Z(n8624) );
  XOR U10063 ( .A(n8625), .B(n8626), .Z(n8619) );
  ANDN U10064 ( .A(n8627), .B(n4961), .Z(n8626) );
  XOR U10065 ( .A(n8628), .B(n8629), .Z(n4961) );
  IV U10066 ( .A(n8625), .Z(n8628) );
  XNOR U10067 ( .A(n4962), .B(n8625), .Z(n8627) );
  NAND U10068 ( .A(n8630), .B(nreg[612]), .Z(n4962) );
  NAND U10069 ( .A(n6107), .B(nreg[612]), .Z(n8630) );
  XOR U10070 ( .A(n8631), .B(n8632), .Z(n8625) );
  ANDN U10071 ( .A(n8633), .B(n4963), .Z(n8632) );
  XOR U10072 ( .A(n8634), .B(n8635), .Z(n4963) );
  IV U10073 ( .A(n8631), .Z(n8634) );
  XNOR U10074 ( .A(n4964), .B(n8631), .Z(n8633) );
  NAND U10075 ( .A(n8636), .B(nreg[611]), .Z(n4964) );
  NAND U10076 ( .A(n6107), .B(nreg[611]), .Z(n8636) );
  XOR U10077 ( .A(n8637), .B(n8638), .Z(n8631) );
  ANDN U10078 ( .A(n8639), .B(n4965), .Z(n8638) );
  XOR U10079 ( .A(n8640), .B(n8641), .Z(n4965) );
  IV U10080 ( .A(n8637), .Z(n8640) );
  XNOR U10081 ( .A(n4966), .B(n8637), .Z(n8639) );
  NAND U10082 ( .A(n8642), .B(nreg[610]), .Z(n4966) );
  NAND U10083 ( .A(n6107), .B(nreg[610]), .Z(n8642) );
  XOR U10084 ( .A(n8643), .B(n8644), .Z(n8637) );
  ANDN U10085 ( .A(n8645), .B(n4967), .Z(n8644) );
  XOR U10086 ( .A(n8646), .B(n8647), .Z(n4967) );
  IV U10087 ( .A(n8643), .Z(n8646) );
  XNOR U10088 ( .A(n4968), .B(n8643), .Z(n8645) );
  NAND U10089 ( .A(n8648), .B(nreg[609]), .Z(n4968) );
  NAND U10090 ( .A(n6107), .B(nreg[609]), .Z(n8648) );
  XOR U10091 ( .A(n8649), .B(n8650), .Z(n8643) );
  ANDN U10092 ( .A(n8651), .B(n4969), .Z(n8650) );
  XOR U10093 ( .A(n8652), .B(n8653), .Z(n4969) );
  IV U10094 ( .A(n8649), .Z(n8652) );
  XNOR U10095 ( .A(n4970), .B(n8649), .Z(n8651) );
  NAND U10096 ( .A(n8654), .B(nreg[608]), .Z(n4970) );
  NAND U10097 ( .A(n6107), .B(nreg[608]), .Z(n8654) );
  XOR U10098 ( .A(n8655), .B(n8656), .Z(n8649) );
  ANDN U10099 ( .A(n8657), .B(n4971), .Z(n8656) );
  XOR U10100 ( .A(n8658), .B(n8659), .Z(n4971) );
  IV U10101 ( .A(n8655), .Z(n8658) );
  XNOR U10102 ( .A(n4972), .B(n8655), .Z(n8657) );
  NAND U10103 ( .A(n8660), .B(nreg[607]), .Z(n4972) );
  NAND U10104 ( .A(n6107), .B(nreg[607]), .Z(n8660) );
  XOR U10105 ( .A(n8661), .B(n8662), .Z(n8655) );
  ANDN U10106 ( .A(n8663), .B(n4975), .Z(n8662) );
  XOR U10107 ( .A(n8664), .B(n8665), .Z(n4975) );
  IV U10108 ( .A(n8661), .Z(n8664) );
  XNOR U10109 ( .A(n4976), .B(n8661), .Z(n8663) );
  NAND U10110 ( .A(n8666), .B(nreg[606]), .Z(n4976) );
  NAND U10111 ( .A(n6107), .B(nreg[606]), .Z(n8666) );
  XOR U10112 ( .A(n8667), .B(n8668), .Z(n8661) );
  ANDN U10113 ( .A(n8669), .B(n4977), .Z(n8668) );
  XOR U10114 ( .A(n8670), .B(n8671), .Z(n4977) );
  IV U10115 ( .A(n8667), .Z(n8670) );
  XNOR U10116 ( .A(n4978), .B(n8667), .Z(n8669) );
  NAND U10117 ( .A(n8672), .B(nreg[605]), .Z(n4978) );
  NAND U10118 ( .A(n6107), .B(nreg[605]), .Z(n8672) );
  XOR U10119 ( .A(n8673), .B(n8674), .Z(n8667) );
  ANDN U10120 ( .A(n8675), .B(n4979), .Z(n8674) );
  XOR U10121 ( .A(n8676), .B(n8677), .Z(n4979) );
  IV U10122 ( .A(n8673), .Z(n8676) );
  XNOR U10123 ( .A(n4980), .B(n8673), .Z(n8675) );
  NAND U10124 ( .A(n8678), .B(nreg[604]), .Z(n4980) );
  NAND U10125 ( .A(n6107), .B(nreg[604]), .Z(n8678) );
  XOR U10126 ( .A(n8679), .B(n8680), .Z(n8673) );
  ANDN U10127 ( .A(n8681), .B(n4981), .Z(n8680) );
  XOR U10128 ( .A(n8682), .B(n8683), .Z(n4981) );
  IV U10129 ( .A(n8679), .Z(n8682) );
  XNOR U10130 ( .A(n4982), .B(n8679), .Z(n8681) );
  NAND U10131 ( .A(n8684), .B(nreg[603]), .Z(n4982) );
  NAND U10132 ( .A(n6107), .B(nreg[603]), .Z(n8684) );
  XOR U10133 ( .A(n8685), .B(n8686), .Z(n8679) );
  ANDN U10134 ( .A(n8687), .B(n4983), .Z(n8686) );
  XOR U10135 ( .A(n8688), .B(n8689), .Z(n4983) );
  IV U10136 ( .A(n8685), .Z(n8688) );
  XNOR U10137 ( .A(n4984), .B(n8685), .Z(n8687) );
  NAND U10138 ( .A(n8690), .B(nreg[602]), .Z(n4984) );
  NAND U10139 ( .A(n6107), .B(nreg[602]), .Z(n8690) );
  XOR U10140 ( .A(n8691), .B(n8692), .Z(n8685) );
  ANDN U10141 ( .A(n8693), .B(n4985), .Z(n8692) );
  XOR U10142 ( .A(n8694), .B(n8695), .Z(n4985) );
  IV U10143 ( .A(n8691), .Z(n8694) );
  XNOR U10144 ( .A(n4986), .B(n8691), .Z(n8693) );
  NAND U10145 ( .A(n8696), .B(nreg[601]), .Z(n4986) );
  NAND U10146 ( .A(n6107), .B(nreg[601]), .Z(n8696) );
  XOR U10147 ( .A(n8697), .B(n8698), .Z(n8691) );
  ANDN U10148 ( .A(n8699), .B(n4987), .Z(n8698) );
  XOR U10149 ( .A(n8700), .B(n8701), .Z(n4987) );
  IV U10150 ( .A(n8697), .Z(n8700) );
  XNOR U10151 ( .A(n4988), .B(n8697), .Z(n8699) );
  NAND U10152 ( .A(n8702), .B(nreg[600]), .Z(n4988) );
  NAND U10153 ( .A(n6107), .B(nreg[600]), .Z(n8702) );
  XOR U10154 ( .A(n8703), .B(n8704), .Z(n8697) );
  ANDN U10155 ( .A(n8705), .B(n4989), .Z(n8704) );
  XOR U10156 ( .A(n8706), .B(n8707), .Z(n4989) );
  IV U10157 ( .A(n8703), .Z(n8706) );
  XNOR U10158 ( .A(n4990), .B(n8703), .Z(n8705) );
  NAND U10159 ( .A(n8708), .B(nreg[599]), .Z(n4990) );
  NAND U10160 ( .A(n6107), .B(nreg[599]), .Z(n8708) );
  XOR U10161 ( .A(n8709), .B(n8710), .Z(n8703) );
  ANDN U10162 ( .A(n8711), .B(n4991), .Z(n8710) );
  XOR U10163 ( .A(n8712), .B(n8713), .Z(n4991) );
  IV U10164 ( .A(n8709), .Z(n8712) );
  XNOR U10165 ( .A(n4992), .B(n8709), .Z(n8711) );
  NAND U10166 ( .A(n8714), .B(nreg[598]), .Z(n4992) );
  NAND U10167 ( .A(n6107), .B(nreg[598]), .Z(n8714) );
  XOR U10168 ( .A(n8715), .B(n8716), .Z(n8709) );
  ANDN U10169 ( .A(n8717), .B(n4993), .Z(n8716) );
  XOR U10170 ( .A(n8718), .B(n8719), .Z(n4993) );
  IV U10171 ( .A(n8715), .Z(n8718) );
  XNOR U10172 ( .A(n4994), .B(n8715), .Z(n8717) );
  NAND U10173 ( .A(n8720), .B(nreg[597]), .Z(n4994) );
  NAND U10174 ( .A(n6107), .B(nreg[597]), .Z(n8720) );
  XOR U10175 ( .A(n8721), .B(n8722), .Z(n8715) );
  ANDN U10176 ( .A(n8723), .B(n4999), .Z(n8722) );
  XOR U10177 ( .A(n8724), .B(n8725), .Z(n4999) );
  IV U10178 ( .A(n8721), .Z(n8724) );
  XNOR U10179 ( .A(n5000), .B(n8721), .Z(n8723) );
  NAND U10180 ( .A(n8726), .B(nreg[596]), .Z(n5000) );
  NAND U10181 ( .A(n6107), .B(nreg[596]), .Z(n8726) );
  XOR U10182 ( .A(n8727), .B(n8728), .Z(n8721) );
  ANDN U10183 ( .A(n8729), .B(n5001), .Z(n8728) );
  XOR U10184 ( .A(n8730), .B(n8731), .Z(n5001) );
  IV U10185 ( .A(n8727), .Z(n8730) );
  XNOR U10186 ( .A(n5002), .B(n8727), .Z(n8729) );
  NAND U10187 ( .A(n8732), .B(nreg[595]), .Z(n5002) );
  NAND U10188 ( .A(n6107), .B(nreg[595]), .Z(n8732) );
  XOR U10189 ( .A(n8733), .B(n8734), .Z(n8727) );
  ANDN U10190 ( .A(n8735), .B(n5003), .Z(n8734) );
  XOR U10191 ( .A(n8736), .B(n8737), .Z(n5003) );
  IV U10192 ( .A(n8733), .Z(n8736) );
  XNOR U10193 ( .A(n5004), .B(n8733), .Z(n8735) );
  NAND U10194 ( .A(n8738), .B(nreg[594]), .Z(n5004) );
  NAND U10195 ( .A(n6107), .B(nreg[594]), .Z(n8738) );
  XOR U10196 ( .A(n8739), .B(n8740), .Z(n8733) );
  ANDN U10197 ( .A(n8741), .B(n5005), .Z(n8740) );
  XOR U10198 ( .A(n8742), .B(n8743), .Z(n5005) );
  IV U10199 ( .A(n8739), .Z(n8742) );
  XNOR U10200 ( .A(n5006), .B(n8739), .Z(n8741) );
  NAND U10201 ( .A(n8744), .B(nreg[593]), .Z(n5006) );
  NAND U10202 ( .A(n6107), .B(nreg[593]), .Z(n8744) );
  XOR U10203 ( .A(n8745), .B(n8746), .Z(n8739) );
  ANDN U10204 ( .A(n8747), .B(n5007), .Z(n8746) );
  XOR U10205 ( .A(n8748), .B(n8749), .Z(n5007) );
  IV U10206 ( .A(n8745), .Z(n8748) );
  XNOR U10207 ( .A(n5008), .B(n8745), .Z(n8747) );
  NAND U10208 ( .A(n8750), .B(nreg[592]), .Z(n5008) );
  NAND U10209 ( .A(n6107), .B(nreg[592]), .Z(n8750) );
  XOR U10210 ( .A(n8751), .B(n8752), .Z(n8745) );
  ANDN U10211 ( .A(n8753), .B(n5009), .Z(n8752) );
  XOR U10212 ( .A(n8754), .B(n8755), .Z(n5009) );
  IV U10213 ( .A(n8751), .Z(n8754) );
  XNOR U10214 ( .A(n5010), .B(n8751), .Z(n8753) );
  NAND U10215 ( .A(n8756), .B(nreg[591]), .Z(n5010) );
  NAND U10216 ( .A(n6107), .B(nreg[591]), .Z(n8756) );
  XOR U10217 ( .A(n8757), .B(n8758), .Z(n8751) );
  ANDN U10218 ( .A(n8759), .B(n5011), .Z(n8758) );
  XOR U10219 ( .A(n8760), .B(n8761), .Z(n5011) );
  IV U10220 ( .A(n8757), .Z(n8760) );
  XNOR U10221 ( .A(n5012), .B(n8757), .Z(n8759) );
  NAND U10222 ( .A(n8762), .B(nreg[590]), .Z(n5012) );
  NAND U10223 ( .A(n6107), .B(nreg[590]), .Z(n8762) );
  XOR U10224 ( .A(n8763), .B(n8764), .Z(n8757) );
  ANDN U10225 ( .A(n8765), .B(n5013), .Z(n8764) );
  XOR U10226 ( .A(n8766), .B(n8767), .Z(n5013) );
  IV U10227 ( .A(n8763), .Z(n8766) );
  XNOR U10228 ( .A(n5014), .B(n8763), .Z(n8765) );
  NAND U10229 ( .A(n8768), .B(nreg[589]), .Z(n5014) );
  NAND U10230 ( .A(n6107), .B(nreg[589]), .Z(n8768) );
  XOR U10231 ( .A(n8769), .B(n8770), .Z(n8763) );
  ANDN U10232 ( .A(n8771), .B(n5015), .Z(n8770) );
  XOR U10233 ( .A(n8772), .B(n8773), .Z(n5015) );
  IV U10234 ( .A(n8769), .Z(n8772) );
  XNOR U10235 ( .A(n5016), .B(n8769), .Z(n8771) );
  NAND U10236 ( .A(n8774), .B(nreg[588]), .Z(n5016) );
  NAND U10237 ( .A(n6107), .B(nreg[588]), .Z(n8774) );
  XOR U10238 ( .A(n8775), .B(n8776), .Z(n8769) );
  ANDN U10239 ( .A(n8777), .B(n5017), .Z(n8776) );
  XOR U10240 ( .A(n8778), .B(n8779), .Z(n5017) );
  IV U10241 ( .A(n8775), .Z(n8778) );
  XNOR U10242 ( .A(n5018), .B(n8775), .Z(n8777) );
  NAND U10243 ( .A(n8780), .B(nreg[587]), .Z(n5018) );
  NAND U10244 ( .A(n6107), .B(nreg[587]), .Z(n8780) );
  XOR U10245 ( .A(n8781), .B(n8782), .Z(n8775) );
  ANDN U10246 ( .A(n8783), .B(n5021), .Z(n8782) );
  XOR U10247 ( .A(n8784), .B(n8785), .Z(n5021) );
  IV U10248 ( .A(n8781), .Z(n8784) );
  XNOR U10249 ( .A(n5022), .B(n8781), .Z(n8783) );
  NAND U10250 ( .A(n8786), .B(nreg[586]), .Z(n5022) );
  NAND U10251 ( .A(n6107), .B(nreg[586]), .Z(n8786) );
  XOR U10252 ( .A(n8787), .B(n8788), .Z(n8781) );
  ANDN U10253 ( .A(n8789), .B(n5023), .Z(n8788) );
  XOR U10254 ( .A(n8790), .B(n8791), .Z(n5023) );
  IV U10255 ( .A(n8787), .Z(n8790) );
  XNOR U10256 ( .A(n5024), .B(n8787), .Z(n8789) );
  NAND U10257 ( .A(n8792), .B(nreg[585]), .Z(n5024) );
  NAND U10258 ( .A(n6107), .B(nreg[585]), .Z(n8792) );
  XOR U10259 ( .A(n8793), .B(n8794), .Z(n8787) );
  ANDN U10260 ( .A(n8795), .B(n5025), .Z(n8794) );
  XOR U10261 ( .A(n8796), .B(n8797), .Z(n5025) );
  IV U10262 ( .A(n8793), .Z(n8796) );
  XNOR U10263 ( .A(n5026), .B(n8793), .Z(n8795) );
  NAND U10264 ( .A(n8798), .B(nreg[584]), .Z(n5026) );
  NAND U10265 ( .A(n6107), .B(nreg[584]), .Z(n8798) );
  XOR U10266 ( .A(n8799), .B(n8800), .Z(n8793) );
  ANDN U10267 ( .A(n8801), .B(n5027), .Z(n8800) );
  XOR U10268 ( .A(n8802), .B(n8803), .Z(n5027) );
  IV U10269 ( .A(n8799), .Z(n8802) );
  XNOR U10270 ( .A(n5028), .B(n8799), .Z(n8801) );
  NAND U10271 ( .A(n8804), .B(nreg[583]), .Z(n5028) );
  NAND U10272 ( .A(n6107), .B(nreg[583]), .Z(n8804) );
  XOR U10273 ( .A(n8805), .B(n8806), .Z(n8799) );
  ANDN U10274 ( .A(n8807), .B(n5029), .Z(n8806) );
  XOR U10275 ( .A(n8808), .B(n8809), .Z(n5029) );
  IV U10276 ( .A(n8805), .Z(n8808) );
  XNOR U10277 ( .A(n5030), .B(n8805), .Z(n8807) );
  NAND U10278 ( .A(n8810), .B(nreg[582]), .Z(n5030) );
  NAND U10279 ( .A(n6107), .B(nreg[582]), .Z(n8810) );
  XOR U10280 ( .A(n8811), .B(n8812), .Z(n8805) );
  ANDN U10281 ( .A(n8813), .B(n5031), .Z(n8812) );
  XOR U10282 ( .A(n8814), .B(n8815), .Z(n5031) );
  IV U10283 ( .A(n8811), .Z(n8814) );
  XNOR U10284 ( .A(n5032), .B(n8811), .Z(n8813) );
  NAND U10285 ( .A(n8816), .B(nreg[581]), .Z(n5032) );
  NAND U10286 ( .A(n6107), .B(nreg[581]), .Z(n8816) );
  XOR U10287 ( .A(n8817), .B(n8818), .Z(n8811) );
  ANDN U10288 ( .A(n8819), .B(n5033), .Z(n8818) );
  XOR U10289 ( .A(n8820), .B(n8821), .Z(n5033) );
  IV U10290 ( .A(n8817), .Z(n8820) );
  XNOR U10291 ( .A(n5034), .B(n8817), .Z(n8819) );
  NAND U10292 ( .A(n8822), .B(nreg[580]), .Z(n5034) );
  NAND U10293 ( .A(n6107), .B(nreg[580]), .Z(n8822) );
  XOR U10294 ( .A(n8823), .B(n8824), .Z(n8817) );
  ANDN U10295 ( .A(n8825), .B(n5035), .Z(n8824) );
  XOR U10296 ( .A(n8826), .B(n8827), .Z(n5035) );
  IV U10297 ( .A(n8823), .Z(n8826) );
  XNOR U10298 ( .A(n5036), .B(n8823), .Z(n8825) );
  NAND U10299 ( .A(n8828), .B(nreg[579]), .Z(n5036) );
  NAND U10300 ( .A(n6107), .B(nreg[579]), .Z(n8828) );
  XOR U10301 ( .A(n8829), .B(n8830), .Z(n8823) );
  ANDN U10302 ( .A(n8831), .B(n5037), .Z(n8830) );
  XOR U10303 ( .A(n8832), .B(n8833), .Z(n5037) );
  IV U10304 ( .A(n8829), .Z(n8832) );
  XNOR U10305 ( .A(n5038), .B(n8829), .Z(n8831) );
  NAND U10306 ( .A(n8834), .B(nreg[578]), .Z(n5038) );
  NAND U10307 ( .A(n6107), .B(nreg[578]), .Z(n8834) );
  XOR U10308 ( .A(n8835), .B(n8836), .Z(n8829) );
  ANDN U10309 ( .A(n8837), .B(n5039), .Z(n8836) );
  XOR U10310 ( .A(n8838), .B(n8839), .Z(n5039) );
  IV U10311 ( .A(n8835), .Z(n8838) );
  XNOR U10312 ( .A(n5040), .B(n8835), .Z(n8837) );
  NAND U10313 ( .A(n8840), .B(nreg[577]), .Z(n5040) );
  NAND U10314 ( .A(n6107), .B(nreg[577]), .Z(n8840) );
  XOR U10315 ( .A(n8841), .B(n8842), .Z(n8835) );
  ANDN U10316 ( .A(n8843), .B(n5043), .Z(n8842) );
  XOR U10317 ( .A(n8844), .B(n8845), .Z(n5043) );
  IV U10318 ( .A(n8841), .Z(n8844) );
  XNOR U10319 ( .A(n5044), .B(n8841), .Z(n8843) );
  NAND U10320 ( .A(n8846), .B(nreg[576]), .Z(n5044) );
  NAND U10321 ( .A(n6107), .B(nreg[576]), .Z(n8846) );
  XOR U10322 ( .A(n8847), .B(n8848), .Z(n8841) );
  ANDN U10323 ( .A(n8849), .B(n5045), .Z(n8848) );
  XOR U10324 ( .A(n8850), .B(n8851), .Z(n5045) );
  IV U10325 ( .A(n8847), .Z(n8850) );
  XNOR U10326 ( .A(n5046), .B(n8847), .Z(n8849) );
  NAND U10327 ( .A(n8852), .B(nreg[575]), .Z(n5046) );
  NAND U10328 ( .A(n6107), .B(nreg[575]), .Z(n8852) );
  XOR U10329 ( .A(n8853), .B(n8854), .Z(n8847) );
  ANDN U10330 ( .A(n8855), .B(n5047), .Z(n8854) );
  XOR U10331 ( .A(n8856), .B(n8857), .Z(n5047) );
  IV U10332 ( .A(n8853), .Z(n8856) );
  XNOR U10333 ( .A(n5048), .B(n8853), .Z(n8855) );
  NAND U10334 ( .A(n8858), .B(nreg[574]), .Z(n5048) );
  NAND U10335 ( .A(n6107), .B(nreg[574]), .Z(n8858) );
  XOR U10336 ( .A(n8859), .B(n8860), .Z(n8853) );
  ANDN U10337 ( .A(n8861), .B(n5049), .Z(n8860) );
  XOR U10338 ( .A(n8862), .B(n8863), .Z(n5049) );
  IV U10339 ( .A(n8859), .Z(n8862) );
  XNOR U10340 ( .A(n5050), .B(n8859), .Z(n8861) );
  NAND U10341 ( .A(n8864), .B(nreg[573]), .Z(n5050) );
  NAND U10342 ( .A(n6107), .B(nreg[573]), .Z(n8864) );
  XOR U10343 ( .A(n8865), .B(n8866), .Z(n8859) );
  ANDN U10344 ( .A(n8867), .B(n5051), .Z(n8866) );
  XOR U10345 ( .A(n8868), .B(n8869), .Z(n5051) );
  IV U10346 ( .A(n8865), .Z(n8868) );
  XNOR U10347 ( .A(n5052), .B(n8865), .Z(n8867) );
  NAND U10348 ( .A(n8870), .B(nreg[572]), .Z(n5052) );
  NAND U10349 ( .A(n6107), .B(nreg[572]), .Z(n8870) );
  XOR U10350 ( .A(n8871), .B(n8872), .Z(n8865) );
  ANDN U10351 ( .A(n8873), .B(n5053), .Z(n8872) );
  XOR U10352 ( .A(n8874), .B(n8875), .Z(n5053) );
  IV U10353 ( .A(n8871), .Z(n8874) );
  XNOR U10354 ( .A(n5054), .B(n8871), .Z(n8873) );
  NAND U10355 ( .A(n8876), .B(nreg[571]), .Z(n5054) );
  NAND U10356 ( .A(n6107), .B(nreg[571]), .Z(n8876) );
  XOR U10357 ( .A(n8877), .B(n8878), .Z(n8871) );
  ANDN U10358 ( .A(n8879), .B(n5055), .Z(n8878) );
  XOR U10359 ( .A(n8880), .B(n8881), .Z(n5055) );
  IV U10360 ( .A(n8877), .Z(n8880) );
  XNOR U10361 ( .A(n5056), .B(n8877), .Z(n8879) );
  NAND U10362 ( .A(n8882), .B(nreg[570]), .Z(n5056) );
  NAND U10363 ( .A(n6107), .B(nreg[570]), .Z(n8882) );
  XOR U10364 ( .A(n8883), .B(n8884), .Z(n8877) );
  ANDN U10365 ( .A(n8885), .B(n5057), .Z(n8884) );
  XOR U10366 ( .A(n8886), .B(n8887), .Z(n5057) );
  IV U10367 ( .A(n8883), .Z(n8886) );
  XNOR U10368 ( .A(n5058), .B(n8883), .Z(n8885) );
  NAND U10369 ( .A(n8888), .B(nreg[569]), .Z(n5058) );
  NAND U10370 ( .A(n6107), .B(nreg[569]), .Z(n8888) );
  XOR U10371 ( .A(n8889), .B(n8890), .Z(n8883) );
  ANDN U10372 ( .A(n8891), .B(n5059), .Z(n8890) );
  XOR U10373 ( .A(n8892), .B(n8893), .Z(n5059) );
  IV U10374 ( .A(n8889), .Z(n8892) );
  XNOR U10375 ( .A(n5060), .B(n8889), .Z(n8891) );
  NAND U10376 ( .A(n8894), .B(nreg[568]), .Z(n5060) );
  NAND U10377 ( .A(n6107), .B(nreg[568]), .Z(n8894) );
  XOR U10378 ( .A(n8895), .B(n8896), .Z(n8889) );
  ANDN U10379 ( .A(n8897), .B(n5061), .Z(n8896) );
  XOR U10380 ( .A(n8898), .B(n8899), .Z(n5061) );
  IV U10381 ( .A(n8895), .Z(n8898) );
  XNOR U10382 ( .A(n5062), .B(n8895), .Z(n8897) );
  NAND U10383 ( .A(n8900), .B(nreg[567]), .Z(n5062) );
  NAND U10384 ( .A(n6107), .B(nreg[567]), .Z(n8900) );
  XOR U10385 ( .A(n8901), .B(n8902), .Z(n8895) );
  ANDN U10386 ( .A(n8903), .B(n5065), .Z(n8902) );
  XOR U10387 ( .A(n8904), .B(n8905), .Z(n5065) );
  IV U10388 ( .A(n8901), .Z(n8904) );
  XNOR U10389 ( .A(n5066), .B(n8901), .Z(n8903) );
  NAND U10390 ( .A(n8906), .B(nreg[566]), .Z(n5066) );
  NAND U10391 ( .A(n6107), .B(nreg[566]), .Z(n8906) );
  XOR U10392 ( .A(n8907), .B(n8908), .Z(n8901) );
  ANDN U10393 ( .A(n8909), .B(n5067), .Z(n8908) );
  XOR U10394 ( .A(n8910), .B(n8911), .Z(n5067) );
  IV U10395 ( .A(n8907), .Z(n8910) );
  XNOR U10396 ( .A(n5068), .B(n8907), .Z(n8909) );
  NAND U10397 ( .A(n8912), .B(nreg[565]), .Z(n5068) );
  NAND U10398 ( .A(n6107), .B(nreg[565]), .Z(n8912) );
  XOR U10399 ( .A(n8913), .B(n8914), .Z(n8907) );
  ANDN U10400 ( .A(n8915), .B(n5069), .Z(n8914) );
  XOR U10401 ( .A(n8916), .B(n8917), .Z(n5069) );
  IV U10402 ( .A(n8913), .Z(n8916) );
  XNOR U10403 ( .A(n5070), .B(n8913), .Z(n8915) );
  NAND U10404 ( .A(n8918), .B(nreg[564]), .Z(n5070) );
  NAND U10405 ( .A(n6107), .B(nreg[564]), .Z(n8918) );
  XOR U10406 ( .A(n8919), .B(n8920), .Z(n8913) );
  ANDN U10407 ( .A(n8921), .B(n5071), .Z(n8920) );
  XOR U10408 ( .A(n8922), .B(n8923), .Z(n5071) );
  IV U10409 ( .A(n8919), .Z(n8922) );
  XNOR U10410 ( .A(n5072), .B(n8919), .Z(n8921) );
  NAND U10411 ( .A(n8924), .B(nreg[563]), .Z(n5072) );
  NAND U10412 ( .A(n6107), .B(nreg[563]), .Z(n8924) );
  XOR U10413 ( .A(n8925), .B(n8926), .Z(n8919) );
  ANDN U10414 ( .A(n8927), .B(n5073), .Z(n8926) );
  XOR U10415 ( .A(n8928), .B(n8929), .Z(n5073) );
  IV U10416 ( .A(n8925), .Z(n8928) );
  XNOR U10417 ( .A(n5074), .B(n8925), .Z(n8927) );
  NAND U10418 ( .A(n8930), .B(nreg[562]), .Z(n5074) );
  NAND U10419 ( .A(n6107), .B(nreg[562]), .Z(n8930) );
  XOR U10420 ( .A(n8931), .B(n8932), .Z(n8925) );
  ANDN U10421 ( .A(n8933), .B(n5075), .Z(n8932) );
  XOR U10422 ( .A(n8934), .B(n8935), .Z(n5075) );
  IV U10423 ( .A(n8931), .Z(n8934) );
  XNOR U10424 ( .A(n5076), .B(n8931), .Z(n8933) );
  NAND U10425 ( .A(n8936), .B(nreg[561]), .Z(n5076) );
  NAND U10426 ( .A(n6107), .B(nreg[561]), .Z(n8936) );
  XOR U10427 ( .A(n8937), .B(n8938), .Z(n8931) );
  ANDN U10428 ( .A(n8939), .B(n5077), .Z(n8938) );
  XOR U10429 ( .A(n8940), .B(n8941), .Z(n5077) );
  IV U10430 ( .A(n8937), .Z(n8940) );
  XNOR U10431 ( .A(n5078), .B(n8937), .Z(n8939) );
  NAND U10432 ( .A(n8942), .B(nreg[560]), .Z(n5078) );
  NAND U10433 ( .A(n6107), .B(nreg[560]), .Z(n8942) );
  XOR U10434 ( .A(n8943), .B(n8944), .Z(n8937) );
  ANDN U10435 ( .A(n8945), .B(n5079), .Z(n8944) );
  XOR U10436 ( .A(n8946), .B(n8947), .Z(n5079) );
  IV U10437 ( .A(n8943), .Z(n8946) );
  XNOR U10438 ( .A(n5080), .B(n8943), .Z(n8945) );
  NAND U10439 ( .A(n8948), .B(nreg[559]), .Z(n5080) );
  NAND U10440 ( .A(n6107), .B(nreg[559]), .Z(n8948) );
  XOR U10441 ( .A(n8949), .B(n8950), .Z(n8943) );
  ANDN U10442 ( .A(n8951), .B(n5081), .Z(n8950) );
  XOR U10443 ( .A(n8952), .B(n8953), .Z(n5081) );
  IV U10444 ( .A(n8949), .Z(n8952) );
  XNOR U10445 ( .A(n5082), .B(n8949), .Z(n8951) );
  NAND U10446 ( .A(n8954), .B(nreg[558]), .Z(n5082) );
  NAND U10447 ( .A(n6107), .B(nreg[558]), .Z(n8954) );
  XOR U10448 ( .A(n8955), .B(n8956), .Z(n8949) );
  ANDN U10449 ( .A(n8957), .B(n5083), .Z(n8956) );
  XOR U10450 ( .A(n8958), .B(n8959), .Z(n5083) );
  IV U10451 ( .A(n8955), .Z(n8958) );
  XNOR U10452 ( .A(n5084), .B(n8955), .Z(n8957) );
  NAND U10453 ( .A(n8960), .B(nreg[557]), .Z(n5084) );
  NAND U10454 ( .A(n6107), .B(nreg[557]), .Z(n8960) );
  XOR U10455 ( .A(n8961), .B(n8962), .Z(n8955) );
  ANDN U10456 ( .A(n8963), .B(n5087), .Z(n8962) );
  XOR U10457 ( .A(n8964), .B(n8965), .Z(n5087) );
  IV U10458 ( .A(n8961), .Z(n8964) );
  XNOR U10459 ( .A(n5088), .B(n8961), .Z(n8963) );
  NAND U10460 ( .A(n8966), .B(nreg[556]), .Z(n5088) );
  NAND U10461 ( .A(n6107), .B(nreg[556]), .Z(n8966) );
  XOR U10462 ( .A(n8967), .B(n8968), .Z(n8961) );
  ANDN U10463 ( .A(n8969), .B(n5089), .Z(n8968) );
  XOR U10464 ( .A(n8970), .B(n8971), .Z(n5089) );
  IV U10465 ( .A(n8967), .Z(n8970) );
  XNOR U10466 ( .A(n5090), .B(n8967), .Z(n8969) );
  NAND U10467 ( .A(n8972), .B(nreg[555]), .Z(n5090) );
  NAND U10468 ( .A(n6107), .B(nreg[555]), .Z(n8972) );
  XOR U10469 ( .A(n8973), .B(n8974), .Z(n8967) );
  ANDN U10470 ( .A(n8975), .B(n5091), .Z(n8974) );
  XOR U10471 ( .A(n8976), .B(n8977), .Z(n5091) );
  IV U10472 ( .A(n8973), .Z(n8976) );
  XNOR U10473 ( .A(n5092), .B(n8973), .Z(n8975) );
  NAND U10474 ( .A(n8978), .B(nreg[554]), .Z(n5092) );
  NAND U10475 ( .A(n6107), .B(nreg[554]), .Z(n8978) );
  XOR U10476 ( .A(n8979), .B(n8980), .Z(n8973) );
  ANDN U10477 ( .A(n8981), .B(n5093), .Z(n8980) );
  XOR U10478 ( .A(n8982), .B(n8983), .Z(n5093) );
  IV U10479 ( .A(n8979), .Z(n8982) );
  XNOR U10480 ( .A(n5094), .B(n8979), .Z(n8981) );
  NAND U10481 ( .A(n8984), .B(nreg[553]), .Z(n5094) );
  NAND U10482 ( .A(n6107), .B(nreg[553]), .Z(n8984) );
  XOR U10483 ( .A(n8985), .B(n8986), .Z(n8979) );
  ANDN U10484 ( .A(n8987), .B(n5095), .Z(n8986) );
  XOR U10485 ( .A(n8988), .B(n8989), .Z(n5095) );
  IV U10486 ( .A(n8985), .Z(n8988) );
  XNOR U10487 ( .A(n5096), .B(n8985), .Z(n8987) );
  NAND U10488 ( .A(n8990), .B(nreg[552]), .Z(n5096) );
  NAND U10489 ( .A(n6107), .B(nreg[552]), .Z(n8990) );
  XOR U10490 ( .A(n8991), .B(n8992), .Z(n8985) );
  ANDN U10491 ( .A(n8993), .B(n5097), .Z(n8992) );
  XOR U10492 ( .A(n8994), .B(n8995), .Z(n5097) );
  IV U10493 ( .A(n8991), .Z(n8994) );
  XNOR U10494 ( .A(n5098), .B(n8991), .Z(n8993) );
  NAND U10495 ( .A(n8996), .B(nreg[551]), .Z(n5098) );
  NAND U10496 ( .A(n6107), .B(nreg[551]), .Z(n8996) );
  XOR U10497 ( .A(n8997), .B(n8998), .Z(n8991) );
  ANDN U10498 ( .A(n8999), .B(n5099), .Z(n8998) );
  XOR U10499 ( .A(n9000), .B(n9001), .Z(n5099) );
  IV U10500 ( .A(n8997), .Z(n9000) );
  XNOR U10501 ( .A(n5100), .B(n8997), .Z(n8999) );
  NAND U10502 ( .A(n9002), .B(nreg[550]), .Z(n5100) );
  NAND U10503 ( .A(n6107), .B(nreg[550]), .Z(n9002) );
  XOR U10504 ( .A(n9003), .B(n9004), .Z(n8997) );
  ANDN U10505 ( .A(n9005), .B(n5101), .Z(n9004) );
  XOR U10506 ( .A(n9006), .B(n9007), .Z(n5101) );
  IV U10507 ( .A(n9003), .Z(n9006) );
  XNOR U10508 ( .A(n5102), .B(n9003), .Z(n9005) );
  NAND U10509 ( .A(n9008), .B(nreg[549]), .Z(n5102) );
  NAND U10510 ( .A(n6107), .B(nreg[549]), .Z(n9008) );
  XOR U10511 ( .A(n9009), .B(n9010), .Z(n9003) );
  ANDN U10512 ( .A(n9011), .B(n5103), .Z(n9010) );
  XOR U10513 ( .A(n9012), .B(n9013), .Z(n5103) );
  IV U10514 ( .A(n9009), .Z(n9012) );
  XNOR U10515 ( .A(n5104), .B(n9009), .Z(n9011) );
  NAND U10516 ( .A(n9014), .B(nreg[548]), .Z(n5104) );
  NAND U10517 ( .A(n6107), .B(nreg[548]), .Z(n9014) );
  XOR U10518 ( .A(n9015), .B(n9016), .Z(n9009) );
  ANDN U10519 ( .A(n9017), .B(n5105), .Z(n9016) );
  XOR U10520 ( .A(n9018), .B(n9019), .Z(n5105) );
  IV U10521 ( .A(n9015), .Z(n9018) );
  XNOR U10522 ( .A(n5106), .B(n9015), .Z(n9017) );
  NAND U10523 ( .A(n9020), .B(nreg[547]), .Z(n5106) );
  NAND U10524 ( .A(n6107), .B(nreg[547]), .Z(n9020) );
  XOR U10525 ( .A(n9021), .B(n9022), .Z(n9015) );
  ANDN U10526 ( .A(n9023), .B(n5109), .Z(n9022) );
  XOR U10527 ( .A(n9024), .B(n9025), .Z(n5109) );
  IV U10528 ( .A(n9021), .Z(n9024) );
  XNOR U10529 ( .A(n5110), .B(n9021), .Z(n9023) );
  NAND U10530 ( .A(n9026), .B(nreg[546]), .Z(n5110) );
  NAND U10531 ( .A(n6107), .B(nreg[546]), .Z(n9026) );
  XOR U10532 ( .A(n9027), .B(n9028), .Z(n9021) );
  ANDN U10533 ( .A(n9029), .B(n5111), .Z(n9028) );
  XOR U10534 ( .A(n9030), .B(n9031), .Z(n5111) );
  IV U10535 ( .A(n9027), .Z(n9030) );
  XNOR U10536 ( .A(n5112), .B(n9027), .Z(n9029) );
  NAND U10537 ( .A(n9032), .B(nreg[545]), .Z(n5112) );
  NAND U10538 ( .A(n6107), .B(nreg[545]), .Z(n9032) );
  XOR U10539 ( .A(n9033), .B(n9034), .Z(n9027) );
  ANDN U10540 ( .A(n9035), .B(n5113), .Z(n9034) );
  XOR U10541 ( .A(n9036), .B(n9037), .Z(n5113) );
  IV U10542 ( .A(n9033), .Z(n9036) );
  XNOR U10543 ( .A(n5114), .B(n9033), .Z(n9035) );
  NAND U10544 ( .A(n9038), .B(nreg[544]), .Z(n5114) );
  NAND U10545 ( .A(n6107), .B(nreg[544]), .Z(n9038) );
  XOR U10546 ( .A(n9039), .B(n9040), .Z(n9033) );
  ANDN U10547 ( .A(n9041), .B(n5115), .Z(n9040) );
  XOR U10548 ( .A(n9042), .B(n9043), .Z(n5115) );
  IV U10549 ( .A(n9039), .Z(n9042) );
  XNOR U10550 ( .A(n5116), .B(n9039), .Z(n9041) );
  NAND U10551 ( .A(n9044), .B(nreg[543]), .Z(n5116) );
  NAND U10552 ( .A(n6107), .B(nreg[543]), .Z(n9044) );
  XOR U10553 ( .A(n9045), .B(n9046), .Z(n9039) );
  ANDN U10554 ( .A(n9047), .B(n5117), .Z(n9046) );
  XOR U10555 ( .A(n9048), .B(n9049), .Z(n5117) );
  IV U10556 ( .A(n9045), .Z(n9048) );
  XNOR U10557 ( .A(n5118), .B(n9045), .Z(n9047) );
  NAND U10558 ( .A(n9050), .B(nreg[542]), .Z(n5118) );
  NAND U10559 ( .A(n6107), .B(nreg[542]), .Z(n9050) );
  XOR U10560 ( .A(n9051), .B(n9052), .Z(n9045) );
  ANDN U10561 ( .A(n9053), .B(n5119), .Z(n9052) );
  XOR U10562 ( .A(n9054), .B(n9055), .Z(n5119) );
  IV U10563 ( .A(n9051), .Z(n9054) );
  XNOR U10564 ( .A(n5120), .B(n9051), .Z(n9053) );
  NAND U10565 ( .A(n9056), .B(nreg[541]), .Z(n5120) );
  NAND U10566 ( .A(n6107), .B(nreg[541]), .Z(n9056) );
  XOR U10567 ( .A(n9057), .B(n9058), .Z(n9051) );
  ANDN U10568 ( .A(n9059), .B(n5121), .Z(n9058) );
  XOR U10569 ( .A(n9060), .B(n9061), .Z(n5121) );
  IV U10570 ( .A(n9057), .Z(n9060) );
  XNOR U10571 ( .A(n5122), .B(n9057), .Z(n9059) );
  NAND U10572 ( .A(n9062), .B(nreg[540]), .Z(n5122) );
  NAND U10573 ( .A(n6107), .B(nreg[540]), .Z(n9062) );
  XOR U10574 ( .A(n9063), .B(n9064), .Z(n9057) );
  ANDN U10575 ( .A(n9065), .B(n5123), .Z(n9064) );
  XOR U10576 ( .A(n9066), .B(n9067), .Z(n5123) );
  IV U10577 ( .A(n9063), .Z(n9066) );
  XNOR U10578 ( .A(n5124), .B(n9063), .Z(n9065) );
  NAND U10579 ( .A(n9068), .B(nreg[539]), .Z(n5124) );
  NAND U10580 ( .A(n6107), .B(nreg[539]), .Z(n9068) );
  XOR U10581 ( .A(n9069), .B(n9070), .Z(n9063) );
  ANDN U10582 ( .A(n9071), .B(n5125), .Z(n9070) );
  XOR U10583 ( .A(n9072), .B(n9073), .Z(n5125) );
  IV U10584 ( .A(n9069), .Z(n9072) );
  XNOR U10585 ( .A(n5126), .B(n9069), .Z(n9071) );
  NAND U10586 ( .A(n9074), .B(nreg[538]), .Z(n5126) );
  NAND U10587 ( .A(n6107), .B(nreg[538]), .Z(n9074) );
  XOR U10588 ( .A(n9075), .B(n9076), .Z(n9069) );
  ANDN U10589 ( .A(n9077), .B(n5127), .Z(n9076) );
  XOR U10590 ( .A(n9078), .B(n9079), .Z(n5127) );
  IV U10591 ( .A(n9075), .Z(n9078) );
  XNOR U10592 ( .A(n5128), .B(n9075), .Z(n9077) );
  NAND U10593 ( .A(n9080), .B(nreg[537]), .Z(n5128) );
  NAND U10594 ( .A(n6107), .B(nreg[537]), .Z(n9080) );
  XOR U10595 ( .A(n9081), .B(n9082), .Z(n9075) );
  ANDN U10596 ( .A(n9083), .B(n5131), .Z(n9082) );
  XOR U10597 ( .A(n9084), .B(n9085), .Z(n5131) );
  IV U10598 ( .A(n9081), .Z(n9084) );
  XNOR U10599 ( .A(n5132), .B(n9081), .Z(n9083) );
  NAND U10600 ( .A(n9086), .B(nreg[536]), .Z(n5132) );
  NAND U10601 ( .A(n6107), .B(nreg[536]), .Z(n9086) );
  XOR U10602 ( .A(n9087), .B(n9088), .Z(n9081) );
  ANDN U10603 ( .A(n9089), .B(n5133), .Z(n9088) );
  XOR U10604 ( .A(n9090), .B(n9091), .Z(n5133) );
  IV U10605 ( .A(n9087), .Z(n9090) );
  XNOR U10606 ( .A(n5134), .B(n9087), .Z(n9089) );
  NAND U10607 ( .A(n9092), .B(nreg[535]), .Z(n5134) );
  NAND U10608 ( .A(n6107), .B(nreg[535]), .Z(n9092) );
  XOR U10609 ( .A(n9093), .B(n9094), .Z(n9087) );
  ANDN U10610 ( .A(n9095), .B(n5135), .Z(n9094) );
  XOR U10611 ( .A(n9096), .B(n9097), .Z(n5135) );
  IV U10612 ( .A(n9093), .Z(n9096) );
  XNOR U10613 ( .A(n5136), .B(n9093), .Z(n9095) );
  NAND U10614 ( .A(n9098), .B(nreg[534]), .Z(n5136) );
  NAND U10615 ( .A(n6107), .B(nreg[534]), .Z(n9098) );
  XOR U10616 ( .A(n9099), .B(n9100), .Z(n9093) );
  ANDN U10617 ( .A(n9101), .B(n5137), .Z(n9100) );
  XOR U10618 ( .A(n9102), .B(n9103), .Z(n5137) );
  IV U10619 ( .A(n9099), .Z(n9102) );
  XNOR U10620 ( .A(n5138), .B(n9099), .Z(n9101) );
  NAND U10621 ( .A(n9104), .B(nreg[533]), .Z(n5138) );
  NAND U10622 ( .A(n6107), .B(nreg[533]), .Z(n9104) );
  XOR U10623 ( .A(n9105), .B(n9106), .Z(n9099) );
  ANDN U10624 ( .A(n9107), .B(n5139), .Z(n9106) );
  XOR U10625 ( .A(n9108), .B(n9109), .Z(n5139) );
  IV U10626 ( .A(n9105), .Z(n9108) );
  XNOR U10627 ( .A(n5140), .B(n9105), .Z(n9107) );
  NAND U10628 ( .A(n9110), .B(nreg[532]), .Z(n5140) );
  NAND U10629 ( .A(n6107), .B(nreg[532]), .Z(n9110) );
  XOR U10630 ( .A(n9111), .B(n9112), .Z(n9105) );
  ANDN U10631 ( .A(n9113), .B(n5141), .Z(n9112) );
  XOR U10632 ( .A(n9114), .B(n9115), .Z(n5141) );
  IV U10633 ( .A(n9111), .Z(n9114) );
  XNOR U10634 ( .A(n5142), .B(n9111), .Z(n9113) );
  NAND U10635 ( .A(n9116), .B(nreg[531]), .Z(n5142) );
  NAND U10636 ( .A(n6107), .B(nreg[531]), .Z(n9116) );
  XOR U10637 ( .A(n9117), .B(n9118), .Z(n9111) );
  ANDN U10638 ( .A(n9119), .B(n5143), .Z(n9118) );
  XOR U10639 ( .A(n9120), .B(n9121), .Z(n5143) );
  IV U10640 ( .A(n9117), .Z(n9120) );
  XNOR U10641 ( .A(n5144), .B(n9117), .Z(n9119) );
  NAND U10642 ( .A(n9122), .B(nreg[530]), .Z(n5144) );
  NAND U10643 ( .A(n6107), .B(nreg[530]), .Z(n9122) );
  XOR U10644 ( .A(n9123), .B(n9124), .Z(n9117) );
  ANDN U10645 ( .A(n9125), .B(n5145), .Z(n9124) );
  XOR U10646 ( .A(n9126), .B(n9127), .Z(n5145) );
  IV U10647 ( .A(n9123), .Z(n9126) );
  XNOR U10648 ( .A(n5146), .B(n9123), .Z(n9125) );
  NAND U10649 ( .A(n9128), .B(nreg[529]), .Z(n5146) );
  NAND U10650 ( .A(n6107), .B(nreg[529]), .Z(n9128) );
  XOR U10651 ( .A(n9129), .B(n9130), .Z(n9123) );
  ANDN U10652 ( .A(n9131), .B(n5147), .Z(n9130) );
  XOR U10653 ( .A(n9132), .B(n9133), .Z(n5147) );
  IV U10654 ( .A(n9129), .Z(n9132) );
  XNOR U10655 ( .A(n5148), .B(n9129), .Z(n9131) );
  NAND U10656 ( .A(n9134), .B(nreg[528]), .Z(n5148) );
  NAND U10657 ( .A(n6107), .B(nreg[528]), .Z(n9134) );
  XOR U10658 ( .A(n9135), .B(n9136), .Z(n9129) );
  ANDN U10659 ( .A(n9137), .B(n5149), .Z(n9136) );
  XOR U10660 ( .A(n9138), .B(n9139), .Z(n5149) );
  IV U10661 ( .A(n9135), .Z(n9138) );
  XNOR U10662 ( .A(n5150), .B(n9135), .Z(n9137) );
  NAND U10663 ( .A(n9140), .B(nreg[527]), .Z(n5150) );
  NAND U10664 ( .A(n6107), .B(nreg[527]), .Z(n9140) );
  XOR U10665 ( .A(n9141), .B(n9142), .Z(n9135) );
  ANDN U10666 ( .A(n9143), .B(n5153), .Z(n9142) );
  XOR U10667 ( .A(n9144), .B(n9145), .Z(n5153) );
  IV U10668 ( .A(n9141), .Z(n9144) );
  XNOR U10669 ( .A(n5154), .B(n9141), .Z(n9143) );
  NAND U10670 ( .A(n9146), .B(nreg[526]), .Z(n5154) );
  NAND U10671 ( .A(n6107), .B(nreg[526]), .Z(n9146) );
  XOR U10672 ( .A(n9147), .B(n9148), .Z(n9141) );
  ANDN U10673 ( .A(n9149), .B(n5155), .Z(n9148) );
  XOR U10674 ( .A(n9150), .B(n9151), .Z(n5155) );
  IV U10675 ( .A(n9147), .Z(n9150) );
  XNOR U10676 ( .A(n5156), .B(n9147), .Z(n9149) );
  NAND U10677 ( .A(n9152), .B(nreg[525]), .Z(n5156) );
  NAND U10678 ( .A(n6107), .B(nreg[525]), .Z(n9152) );
  XOR U10679 ( .A(n9153), .B(n9154), .Z(n9147) );
  ANDN U10680 ( .A(n9155), .B(n5157), .Z(n9154) );
  XOR U10681 ( .A(n9156), .B(n9157), .Z(n5157) );
  IV U10682 ( .A(n9153), .Z(n9156) );
  XNOR U10683 ( .A(n5158), .B(n9153), .Z(n9155) );
  NAND U10684 ( .A(n9158), .B(nreg[524]), .Z(n5158) );
  NAND U10685 ( .A(n6107), .B(nreg[524]), .Z(n9158) );
  XOR U10686 ( .A(n9159), .B(n9160), .Z(n9153) );
  ANDN U10687 ( .A(n9161), .B(n5159), .Z(n9160) );
  XOR U10688 ( .A(n9162), .B(n9163), .Z(n5159) );
  IV U10689 ( .A(n9159), .Z(n9162) );
  XNOR U10690 ( .A(n5160), .B(n9159), .Z(n9161) );
  NAND U10691 ( .A(n9164), .B(nreg[523]), .Z(n5160) );
  NAND U10692 ( .A(n6107), .B(nreg[523]), .Z(n9164) );
  XOR U10693 ( .A(n9165), .B(n9166), .Z(n9159) );
  ANDN U10694 ( .A(n9167), .B(n5161), .Z(n9166) );
  XOR U10695 ( .A(n9168), .B(n9169), .Z(n5161) );
  IV U10696 ( .A(n9165), .Z(n9168) );
  XNOR U10697 ( .A(n5162), .B(n9165), .Z(n9167) );
  NAND U10698 ( .A(n9170), .B(nreg[522]), .Z(n5162) );
  NAND U10699 ( .A(n6107), .B(nreg[522]), .Z(n9170) );
  XOR U10700 ( .A(n9171), .B(n9172), .Z(n9165) );
  ANDN U10701 ( .A(n9173), .B(n5163), .Z(n9172) );
  XOR U10702 ( .A(n9174), .B(n9175), .Z(n5163) );
  IV U10703 ( .A(n9171), .Z(n9174) );
  XNOR U10704 ( .A(n5164), .B(n9171), .Z(n9173) );
  NAND U10705 ( .A(n9176), .B(nreg[521]), .Z(n5164) );
  NAND U10706 ( .A(n6107), .B(nreg[521]), .Z(n9176) );
  XOR U10707 ( .A(n9177), .B(n9178), .Z(n9171) );
  ANDN U10708 ( .A(n9179), .B(n5165), .Z(n9178) );
  XOR U10709 ( .A(n9180), .B(n9181), .Z(n5165) );
  IV U10710 ( .A(n9177), .Z(n9180) );
  XNOR U10711 ( .A(n5166), .B(n9177), .Z(n9179) );
  NAND U10712 ( .A(n9182), .B(nreg[520]), .Z(n5166) );
  NAND U10713 ( .A(n6107), .B(nreg[520]), .Z(n9182) );
  XOR U10714 ( .A(n9183), .B(n9184), .Z(n9177) );
  ANDN U10715 ( .A(n9185), .B(n5167), .Z(n9184) );
  XOR U10716 ( .A(n9186), .B(n9187), .Z(n5167) );
  IV U10717 ( .A(n9183), .Z(n9186) );
  XNOR U10718 ( .A(n5168), .B(n9183), .Z(n9185) );
  NAND U10719 ( .A(n9188), .B(nreg[519]), .Z(n5168) );
  NAND U10720 ( .A(n6107), .B(nreg[519]), .Z(n9188) );
  XOR U10721 ( .A(n9189), .B(n9190), .Z(n9183) );
  ANDN U10722 ( .A(n9191), .B(n5169), .Z(n9190) );
  XOR U10723 ( .A(n9192), .B(n9193), .Z(n5169) );
  IV U10724 ( .A(n9189), .Z(n9192) );
  XNOR U10725 ( .A(n5170), .B(n9189), .Z(n9191) );
  NAND U10726 ( .A(n9194), .B(nreg[518]), .Z(n5170) );
  NAND U10727 ( .A(n6107), .B(nreg[518]), .Z(n9194) );
  XOR U10728 ( .A(n9195), .B(n9196), .Z(n9189) );
  ANDN U10729 ( .A(n9197), .B(n5171), .Z(n9196) );
  XOR U10730 ( .A(n9198), .B(n9199), .Z(n5171) );
  IV U10731 ( .A(n9195), .Z(n9198) );
  XNOR U10732 ( .A(n5172), .B(n9195), .Z(n9197) );
  NAND U10733 ( .A(n9200), .B(nreg[517]), .Z(n5172) );
  NAND U10734 ( .A(n6107), .B(nreg[517]), .Z(n9200) );
  XOR U10735 ( .A(n9201), .B(n9202), .Z(n9195) );
  ANDN U10736 ( .A(n9203), .B(n5175), .Z(n9202) );
  XOR U10737 ( .A(n9204), .B(n9205), .Z(n5175) );
  IV U10738 ( .A(n9201), .Z(n9204) );
  XNOR U10739 ( .A(n5176), .B(n9201), .Z(n9203) );
  NAND U10740 ( .A(n9206), .B(nreg[516]), .Z(n5176) );
  NAND U10741 ( .A(n6107), .B(nreg[516]), .Z(n9206) );
  XOR U10742 ( .A(n9207), .B(n9208), .Z(n9201) );
  ANDN U10743 ( .A(n9209), .B(n5177), .Z(n9208) );
  XOR U10744 ( .A(n9210), .B(n9211), .Z(n5177) );
  IV U10745 ( .A(n9207), .Z(n9210) );
  XNOR U10746 ( .A(n5178), .B(n9207), .Z(n9209) );
  NAND U10747 ( .A(n9212), .B(nreg[515]), .Z(n5178) );
  NAND U10748 ( .A(n6107), .B(nreg[515]), .Z(n9212) );
  XOR U10749 ( .A(n9213), .B(n9214), .Z(n9207) );
  ANDN U10750 ( .A(n9215), .B(n5179), .Z(n9214) );
  XOR U10751 ( .A(n9216), .B(n9217), .Z(n5179) );
  IV U10752 ( .A(n9213), .Z(n9216) );
  XNOR U10753 ( .A(n5180), .B(n9213), .Z(n9215) );
  NAND U10754 ( .A(n9218), .B(nreg[514]), .Z(n5180) );
  NAND U10755 ( .A(n6107), .B(nreg[514]), .Z(n9218) );
  XOR U10756 ( .A(n9219), .B(n9220), .Z(n9213) );
  ANDN U10757 ( .A(n9221), .B(n5181), .Z(n9220) );
  XOR U10758 ( .A(n9222), .B(n9223), .Z(n5181) );
  IV U10759 ( .A(n9219), .Z(n9222) );
  XNOR U10760 ( .A(n5182), .B(n9219), .Z(n9221) );
  NAND U10761 ( .A(n9224), .B(nreg[513]), .Z(n5182) );
  NAND U10762 ( .A(n6107), .B(nreg[513]), .Z(n9224) );
  XOR U10763 ( .A(n9225), .B(n9226), .Z(n9219) );
  ANDN U10764 ( .A(n9227), .B(n5183), .Z(n9226) );
  XOR U10765 ( .A(n9228), .B(n9229), .Z(n5183) );
  IV U10766 ( .A(n9225), .Z(n9228) );
  XNOR U10767 ( .A(n5184), .B(n9225), .Z(n9227) );
  NAND U10768 ( .A(n9230), .B(nreg[512]), .Z(n5184) );
  NAND U10769 ( .A(n6107), .B(nreg[512]), .Z(n9230) );
  XOR U10770 ( .A(n9231), .B(n9232), .Z(n9225) );
  ANDN U10771 ( .A(n9233), .B(n5185), .Z(n9232) );
  XOR U10772 ( .A(n9234), .B(n9235), .Z(n5185) );
  IV U10773 ( .A(n9231), .Z(n9234) );
  XNOR U10774 ( .A(n5186), .B(n9231), .Z(n9233) );
  NAND U10775 ( .A(n9236), .B(nreg[511]), .Z(n5186) );
  NAND U10776 ( .A(n6107), .B(nreg[511]), .Z(n9236) );
  XOR U10777 ( .A(n9237), .B(n9238), .Z(n9231) );
  ANDN U10778 ( .A(n9239), .B(n5187), .Z(n9238) );
  XOR U10779 ( .A(n9240), .B(n9241), .Z(n5187) );
  IV U10780 ( .A(n9237), .Z(n9240) );
  XNOR U10781 ( .A(n5188), .B(n9237), .Z(n9239) );
  NAND U10782 ( .A(n9242), .B(nreg[510]), .Z(n5188) );
  NAND U10783 ( .A(n6107), .B(nreg[510]), .Z(n9242) );
  XOR U10784 ( .A(n9243), .B(n9244), .Z(n9237) );
  ANDN U10785 ( .A(n9245), .B(n5189), .Z(n9244) );
  XOR U10786 ( .A(n9246), .B(n9247), .Z(n5189) );
  IV U10787 ( .A(n9243), .Z(n9246) );
  XNOR U10788 ( .A(n5190), .B(n9243), .Z(n9245) );
  NAND U10789 ( .A(n9248), .B(nreg[509]), .Z(n5190) );
  NAND U10790 ( .A(n6107), .B(nreg[509]), .Z(n9248) );
  XOR U10791 ( .A(n9249), .B(n9250), .Z(n9243) );
  ANDN U10792 ( .A(n9251), .B(n5191), .Z(n9250) );
  XOR U10793 ( .A(n9252), .B(n9253), .Z(n5191) );
  IV U10794 ( .A(n9249), .Z(n9252) );
  XNOR U10795 ( .A(n5192), .B(n9249), .Z(n9251) );
  NAND U10796 ( .A(n9254), .B(nreg[508]), .Z(n5192) );
  NAND U10797 ( .A(n6107), .B(nreg[508]), .Z(n9254) );
  XOR U10798 ( .A(n9255), .B(n9256), .Z(n9249) );
  ANDN U10799 ( .A(n9257), .B(n5193), .Z(n9256) );
  XOR U10800 ( .A(n9258), .B(n9259), .Z(n5193) );
  IV U10801 ( .A(n9255), .Z(n9258) );
  XNOR U10802 ( .A(n5194), .B(n9255), .Z(n9257) );
  NAND U10803 ( .A(n9260), .B(nreg[507]), .Z(n5194) );
  NAND U10804 ( .A(n6107), .B(nreg[507]), .Z(n9260) );
  XOR U10805 ( .A(n9261), .B(n9262), .Z(n9255) );
  ANDN U10806 ( .A(n9263), .B(n5197), .Z(n9262) );
  XOR U10807 ( .A(n9264), .B(n9265), .Z(n5197) );
  IV U10808 ( .A(n9261), .Z(n9264) );
  XNOR U10809 ( .A(n5198), .B(n9261), .Z(n9263) );
  NAND U10810 ( .A(n9266), .B(nreg[506]), .Z(n5198) );
  NAND U10811 ( .A(n6107), .B(nreg[506]), .Z(n9266) );
  XOR U10812 ( .A(n9267), .B(n9268), .Z(n9261) );
  ANDN U10813 ( .A(n9269), .B(n5199), .Z(n9268) );
  XOR U10814 ( .A(n9270), .B(n9271), .Z(n5199) );
  IV U10815 ( .A(n9267), .Z(n9270) );
  XNOR U10816 ( .A(n5200), .B(n9267), .Z(n9269) );
  NAND U10817 ( .A(n9272), .B(nreg[505]), .Z(n5200) );
  NAND U10818 ( .A(n6107), .B(nreg[505]), .Z(n9272) );
  XOR U10819 ( .A(n9273), .B(n9274), .Z(n9267) );
  ANDN U10820 ( .A(n9275), .B(n5201), .Z(n9274) );
  XOR U10821 ( .A(n9276), .B(n9277), .Z(n5201) );
  IV U10822 ( .A(n9273), .Z(n9276) );
  XNOR U10823 ( .A(n5202), .B(n9273), .Z(n9275) );
  NAND U10824 ( .A(n9278), .B(nreg[504]), .Z(n5202) );
  NAND U10825 ( .A(n6107), .B(nreg[504]), .Z(n9278) );
  XOR U10826 ( .A(n9279), .B(n9280), .Z(n9273) );
  ANDN U10827 ( .A(n9281), .B(n5203), .Z(n9280) );
  XOR U10828 ( .A(n9282), .B(n9283), .Z(n5203) );
  IV U10829 ( .A(n9279), .Z(n9282) );
  XNOR U10830 ( .A(n5204), .B(n9279), .Z(n9281) );
  NAND U10831 ( .A(n9284), .B(nreg[503]), .Z(n5204) );
  NAND U10832 ( .A(n6107), .B(nreg[503]), .Z(n9284) );
  XOR U10833 ( .A(n9285), .B(n9286), .Z(n9279) );
  ANDN U10834 ( .A(n9287), .B(n5205), .Z(n9286) );
  XOR U10835 ( .A(n9288), .B(n9289), .Z(n5205) );
  IV U10836 ( .A(n9285), .Z(n9288) );
  XNOR U10837 ( .A(n5206), .B(n9285), .Z(n9287) );
  NAND U10838 ( .A(n9290), .B(nreg[502]), .Z(n5206) );
  NAND U10839 ( .A(n6107), .B(nreg[502]), .Z(n9290) );
  XOR U10840 ( .A(n9291), .B(n9292), .Z(n9285) );
  ANDN U10841 ( .A(n9293), .B(n5207), .Z(n9292) );
  XOR U10842 ( .A(n9294), .B(n9295), .Z(n5207) );
  IV U10843 ( .A(n9291), .Z(n9294) );
  XNOR U10844 ( .A(n5208), .B(n9291), .Z(n9293) );
  NAND U10845 ( .A(n9296), .B(nreg[501]), .Z(n5208) );
  NAND U10846 ( .A(n6107), .B(nreg[501]), .Z(n9296) );
  XOR U10847 ( .A(n9297), .B(n9298), .Z(n9291) );
  ANDN U10848 ( .A(n9299), .B(n5209), .Z(n9298) );
  XOR U10849 ( .A(n9300), .B(n9301), .Z(n5209) );
  IV U10850 ( .A(n9297), .Z(n9300) );
  XNOR U10851 ( .A(n5210), .B(n9297), .Z(n9299) );
  NAND U10852 ( .A(n9302), .B(nreg[500]), .Z(n5210) );
  NAND U10853 ( .A(n6107), .B(nreg[500]), .Z(n9302) );
  XOR U10854 ( .A(n9303), .B(n9304), .Z(n9297) );
  ANDN U10855 ( .A(n9305), .B(n5211), .Z(n9304) );
  XOR U10856 ( .A(n9306), .B(n9307), .Z(n5211) );
  IV U10857 ( .A(n9303), .Z(n9306) );
  XNOR U10858 ( .A(n5212), .B(n9303), .Z(n9305) );
  NAND U10859 ( .A(n9308), .B(nreg[499]), .Z(n5212) );
  NAND U10860 ( .A(n6107), .B(nreg[499]), .Z(n9308) );
  XOR U10861 ( .A(n9309), .B(n9310), .Z(n9303) );
  ANDN U10862 ( .A(n9311), .B(n5213), .Z(n9310) );
  XOR U10863 ( .A(n9312), .B(n9313), .Z(n5213) );
  IV U10864 ( .A(n9309), .Z(n9312) );
  XNOR U10865 ( .A(n5214), .B(n9309), .Z(n9311) );
  NAND U10866 ( .A(n9314), .B(nreg[498]), .Z(n5214) );
  NAND U10867 ( .A(n6107), .B(nreg[498]), .Z(n9314) );
  XOR U10868 ( .A(n9315), .B(n9316), .Z(n9309) );
  ANDN U10869 ( .A(n9317), .B(n5215), .Z(n9316) );
  XOR U10870 ( .A(n9318), .B(n9319), .Z(n5215) );
  IV U10871 ( .A(n9315), .Z(n9318) );
  XNOR U10872 ( .A(n5216), .B(n9315), .Z(n9317) );
  NAND U10873 ( .A(n9320), .B(nreg[497]), .Z(n5216) );
  NAND U10874 ( .A(n6107), .B(nreg[497]), .Z(n9320) );
  XOR U10875 ( .A(n9321), .B(n9322), .Z(n9315) );
  ANDN U10876 ( .A(n9323), .B(n5221), .Z(n9322) );
  XOR U10877 ( .A(n9324), .B(n9325), .Z(n5221) );
  IV U10878 ( .A(n9321), .Z(n9324) );
  XNOR U10879 ( .A(n5222), .B(n9321), .Z(n9323) );
  NAND U10880 ( .A(n9326), .B(nreg[496]), .Z(n5222) );
  NAND U10881 ( .A(n6107), .B(nreg[496]), .Z(n9326) );
  XOR U10882 ( .A(n9327), .B(n9328), .Z(n9321) );
  ANDN U10883 ( .A(n9329), .B(n5223), .Z(n9328) );
  XOR U10884 ( .A(n9330), .B(n9331), .Z(n5223) );
  IV U10885 ( .A(n9327), .Z(n9330) );
  XNOR U10886 ( .A(n5224), .B(n9327), .Z(n9329) );
  NAND U10887 ( .A(n9332), .B(nreg[495]), .Z(n5224) );
  NAND U10888 ( .A(n6107), .B(nreg[495]), .Z(n9332) );
  XOR U10889 ( .A(n9333), .B(n9334), .Z(n9327) );
  ANDN U10890 ( .A(n9335), .B(n5225), .Z(n9334) );
  XOR U10891 ( .A(n9336), .B(n9337), .Z(n5225) );
  IV U10892 ( .A(n9333), .Z(n9336) );
  XNOR U10893 ( .A(n5226), .B(n9333), .Z(n9335) );
  NAND U10894 ( .A(n9338), .B(nreg[494]), .Z(n5226) );
  NAND U10895 ( .A(n6107), .B(nreg[494]), .Z(n9338) );
  XOR U10896 ( .A(n9339), .B(n9340), .Z(n9333) );
  ANDN U10897 ( .A(n9341), .B(n5227), .Z(n9340) );
  XOR U10898 ( .A(n9342), .B(n9343), .Z(n5227) );
  IV U10899 ( .A(n9339), .Z(n9342) );
  XNOR U10900 ( .A(n5228), .B(n9339), .Z(n9341) );
  NAND U10901 ( .A(n9344), .B(nreg[493]), .Z(n5228) );
  NAND U10902 ( .A(n6107), .B(nreg[493]), .Z(n9344) );
  XOR U10903 ( .A(n9345), .B(n9346), .Z(n9339) );
  ANDN U10904 ( .A(n9347), .B(n5229), .Z(n9346) );
  XOR U10905 ( .A(n9348), .B(n9349), .Z(n5229) );
  IV U10906 ( .A(n9345), .Z(n9348) );
  XNOR U10907 ( .A(n5230), .B(n9345), .Z(n9347) );
  NAND U10908 ( .A(n9350), .B(nreg[492]), .Z(n5230) );
  NAND U10909 ( .A(n6107), .B(nreg[492]), .Z(n9350) );
  XOR U10910 ( .A(n9351), .B(n9352), .Z(n9345) );
  ANDN U10911 ( .A(n9353), .B(n5231), .Z(n9352) );
  XOR U10912 ( .A(n9354), .B(n9355), .Z(n5231) );
  IV U10913 ( .A(n9351), .Z(n9354) );
  XNOR U10914 ( .A(n5232), .B(n9351), .Z(n9353) );
  NAND U10915 ( .A(n9356), .B(nreg[491]), .Z(n5232) );
  NAND U10916 ( .A(n6107), .B(nreg[491]), .Z(n9356) );
  XOR U10917 ( .A(n9357), .B(n9358), .Z(n9351) );
  ANDN U10918 ( .A(n9359), .B(n5233), .Z(n9358) );
  XOR U10919 ( .A(n9360), .B(n9361), .Z(n5233) );
  IV U10920 ( .A(n9357), .Z(n9360) );
  XNOR U10921 ( .A(n5234), .B(n9357), .Z(n9359) );
  NAND U10922 ( .A(n9362), .B(nreg[490]), .Z(n5234) );
  NAND U10923 ( .A(n6107), .B(nreg[490]), .Z(n9362) );
  XOR U10924 ( .A(n9363), .B(n9364), .Z(n9357) );
  ANDN U10925 ( .A(n9365), .B(n5235), .Z(n9364) );
  XOR U10926 ( .A(n9366), .B(n9367), .Z(n5235) );
  IV U10927 ( .A(n9363), .Z(n9366) );
  XNOR U10928 ( .A(n5236), .B(n9363), .Z(n9365) );
  NAND U10929 ( .A(n9368), .B(nreg[489]), .Z(n5236) );
  NAND U10930 ( .A(n6107), .B(nreg[489]), .Z(n9368) );
  XOR U10931 ( .A(n9369), .B(n9370), .Z(n9363) );
  ANDN U10932 ( .A(n9371), .B(n5237), .Z(n9370) );
  XOR U10933 ( .A(n9372), .B(n9373), .Z(n5237) );
  IV U10934 ( .A(n9369), .Z(n9372) );
  XNOR U10935 ( .A(n5238), .B(n9369), .Z(n9371) );
  NAND U10936 ( .A(n9374), .B(nreg[488]), .Z(n5238) );
  NAND U10937 ( .A(n6107), .B(nreg[488]), .Z(n9374) );
  XOR U10938 ( .A(n9375), .B(n9376), .Z(n9369) );
  ANDN U10939 ( .A(n9377), .B(n5239), .Z(n9376) );
  XOR U10940 ( .A(n9378), .B(n9379), .Z(n5239) );
  IV U10941 ( .A(n9375), .Z(n9378) );
  XNOR U10942 ( .A(n5240), .B(n9375), .Z(n9377) );
  NAND U10943 ( .A(n9380), .B(nreg[487]), .Z(n5240) );
  NAND U10944 ( .A(n6107), .B(nreg[487]), .Z(n9380) );
  XOR U10945 ( .A(n9381), .B(n9382), .Z(n9375) );
  ANDN U10946 ( .A(n9383), .B(n5243), .Z(n9382) );
  XOR U10947 ( .A(n9384), .B(n9385), .Z(n5243) );
  IV U10948 ( .A(n9381), .Z(n9384) );
  XNOR U10949 ( .A(n5244), .B(n9381), .Z(n9383) );
  NAND U10950 ( .A(n9386), .B(nreg[486]), .Z(n5244) );
  NAND U10951 ( .A(n6107), .B(nreg[486]), .Z(n9386) );
  XOR U10952 ( .A(n9387), .B(n9388), .Z(n9381) );
  ANDN U10953 ( .A(n9389), .B(n5245), .Z(n9388) );
  XOR U10954 ( .A(n9390), .B(n9391), .Z(n5245) );
  IV U10955 ( .A(n9387), .Z(n9390) );
  XNOR U10956 ( .A(n5246), .B(n9387), .Z(n9389) );
  NAND U10957 ( .A(n9392), .B(nreg[485]), .Z(n5246) );
  NAND U10958 ( .A(n6107), .B(nreg[485]), .Z(n9392) );
  XOR U10959 ( .A(n9393), .B(n9394), .Z(n9387) );
  ANDN U10960 ( .A(n9395), .B(n5247), .Z(n9394) );
  XOR U10961 ( .A(n9396), .B(n9397), .Z(n5247) );
  IV U10962 ( .A(n9393), .Z(n9396) );
  XNOR U10963 ( .A(n5248), .B(n9393), .Z(n9395) );
  NAND U10964 ( .A(n9398), .B(nreg[484]), .Z(n5248) );
  NAND U10965 ( .A(n6107), .B(nreg[484]), .Z(n9398) );
  XOR U10966 ( .A(n9399), .B(n9400), .Z(n9393) );
  ANDN U10967 ( .A(n9401), .B(n5249), .Z(n9400) );
  XOR U10968 ( .A(n9402), .B(n9403), .Z(n5249) );
  IV U10969 ( .A(n9399), .Z(n9402) );
  XNOR U10970 ( .A(n5250), .B(n9399), .Z(n9401) );
  NAND U10971 ( .A(n9404), .B(nreg[483]), .Z(n5250) );
  NAND U10972 ( .A(n6107), .B(nreg[483]), .Z(n9404) );
  XOR U10973 ( .A(n9405), .B(n9406), .Z(n9399) );
  ANDN U10974 ( .A(n9407), .B(n5251), .Z(n9406) );
  XOR U10975 ( .A(n9408), .B(n9409), .Z(n5251) );
  IV U10976 ( .A(n9405), .Z(n9408) );
  XNOR U10977 ( .A(n5252), .B(n9405), .Z(n9407) );
  NAND U10978 ( .A(n9410), .B(nreg[482]), .Z(n5252) );
  NAND U10979 ( .A(n6107), .B(nreg[482]), .Z(n9410) );
  XOR U10980 ( .A(n9411), .B(n9412), .Z(n9405) );
  ANDN U10981 ( .A(n9413), .B(n5253), .Z(n9412) );
  XOR U10982 ( .A(n9414), .B(n9415), .Z(n5253) );
  IV U10983 ( .A(n9411), .Z(n9414) );
  XNOR U10984 ( .A(n5254), .B(n9411), .Z(n9413) );
  NAND U10985 ( .A(n9416), .B(nreg[481]), .Z(n5254) );
  NAND U10986 ( .A(n6107), .B(nreg[481]), .Z(n9416) );
  XOR U10987 ( .A(n9417), .B(n9418), .Z(n9411) );
  ANDN U10988 ( .A(n9419), .B(n5255), .Z(n9418) );
  XOR U10989 ( .A(n9420), .B(n9421), .Z(n5255) );
  IV U10990 ( .A(n9417), .Z(n9420) );
  XNOR U10991 ( .A(n5256), .B(n9417), .Z(n9419) );
  NAND U10992 ( .A(n9422), .B(nreg[480]), .Z(n5256) );
  NAND U10993 ( .A(n6107), .B(nreg[480]), .Z(n9422) );
  XOR U10994 ( .A(n9423), .B(n9424), .Z(n9417) );
  ANDN U10995 ( .A(n9425), .B(n5257), .Z(n9424) );
  XOR U10996 ( .A(n9426), .B(n9427), .Z(n5257) );
  IV U10997 ( .A(n9423), .Z(n9426) );
  XNOR U10998 ( .A(n5258), .B(n9423), .Z(n9425) );
  NAND U10999 ( .A(n9428), .B(nreg[479]), .Z(n5258) );
  NAND U11000 ( .A(n6107), .B(nreg[479]), .Z(n9428) );
  XOR U11001 ( .A(n9429), .B(n9430), .Z(n9423) );
  ANDN U11002 ( .A(n9431), .B(n5259), .Z(n9430) );
  XOR U11003 ( .A(n9432), .B(n9433), .Z(n5259) );
  IV U11004 ( .A(n9429), .Z(n9432) );
  XNOR U11005 ( .A(n5260), .B(n9429), .Z(n9431) );
  NAND U11006 ( .A(n9434), .B(nreg[478]), .Z(n5260) );
  NAND U11007 ( .A(n6107), .B(nreg[478]), .Z(n9434) );
  XOR U11008 ( .A(n9435), .B(n9436), .Z(n9429) );
  ANDN U11009 ( .A(n9437), .B(n5261), .Z(n9436) );
  XOR U11010 ( .A(n9438), .B(n9439), .Z(n5261) );
  IV U11011 ( .A(n9435), .Z(n9438) );
  XNOR U11012 ( .A(n5262), .B(n9435), .Z(n9437) );
  NAND U11013 ( .A(n9440), .B(nreg[477]), .Z(n5262) );
  NAND U11014 ( .A(n6107), .B(nreg[477]), .Z(n9440) );
  XOR U11015 ( .A(n9441), .B(n9442), .Z(n9435) );
  ANDN U11016 ( .A(n9443), .B(n5265), .Z(n9442) );
  XOR U11017 ( .A(n9444), .B(n9445), .Z(n5265) );
  IV U11018 ( .A(n9441), .Z(n9444) );
  XNOR U11019 ( .A(n5266), .B(n9441), .Z(n9443) );
  NAND U11020 ( .A(n9446), .B(nreg[476]), .Z(n5266) );
  NAND U11021 ( .A(n6107), .B(nreg[476]), .Z(n9446) );
  XOR U11022 ( .A(n9447), .B(n9448), .Z(n9441) );
  ANDN U11023 ( .A(n9449), .B(n5267), .Z(n9448) );
  XOR U11024 ( .A(n9450), .B(n9451), .Z(n5267) );
  IV U11025 ( .A(n9447), .Z(n9450) );
  XNOR U11026 ( .A(n5268), .B(n9447), .Z(n9449) );
  NAND U11027 ( .A(n9452), .B(nreg[475]), .Z(n5268) );
  NAND U11028 ( .A(n6107), .B(nreg[475]), .Z(n9452) );
  XOR U11029 ( .A(n9453), .B(n9454), .Z(n9447) );
  ANDN U11030 ( .A(n9455), .B(n5269), .Z(n9454) );
  XOR U11031 ( .A(n9456), .B(n9457), .Z(n5269) );
  IV U11032 ( .A(n9453), .Z(n9456) );
  XNOR U11033 ( .A(n5270), .B(n9453), .Z(n9455) );
  NAND U11034 ( .A(n9458), .B(nreg[474]), .Z(n5270) );
  NAND U11035 ( .A(n6107), .B(nreg[474]), .Z(n9458) );
  XOR U11036 ( .A(n9459), .B(n9460), .Z(n9453) );
  ANDN U11037 ( .A(n9461), .B(n5271), .Z(n9460) );
  XOR U11038 ( .A(n9462), .B(n9463), .Z(n5271) );
  IV U11039 ( .A(n9459), .Z(n9462) );
  XNOR U11040 ( .A(n5272), .B(n9459), .Z(n9461) );
  NAND U11041 ( .A(n9464), .B(nreg[473]), .Z(n5272) );
  NAND U11042 ( .A(n6107), .B(nreg[473]), .Z(n9464) );
  XOR U11043 ( .A(n9465), .B(n9466), .Z(n9459) );
  ANDN U11044 ( .A(n9467), .B(n5273), .Z(n9466) );
  XOR U11045 ( .A(n9468), .B(n9469), .Z(n5273) );
  IV U11046 ( .A(n9465), .Z(n9468) );
  XNOR U11047 ( .A(n5274), .B(n9465), .Z(n9467) );
  NAND U11048 ( .A(n9470), .B(nreg[472]), .Z(n5274) );
  NAND U11049 ( .A(n6107), .B(nreg[472]), .Z(n9470) );
  XOR U11050 ( .A(n9471), .B(n9472), .Z(n9465) );
  ANDN U11051 ( .A(n9473), .B(n5275), .Z(n9472) );
  XOR U11052 ( .A(n9474), .B(n9475), .Z(n5275) );
  IV U11053 ( .A(n9471), .Z(n9474) );
  XNOR U11054 ( .A(n5276), .B(n9471), .Z(n9473) );
  NAND U11055 ( .A(n9476), .B(nreg[471]), .Z(n5276) );
  NAND U11056 ( .A(n6107), .B(nreg[471]), .Z(n9476) );
  XOR U11057 ( .A(n9477), .B(n9478), .Z(n9471) );
  ANDN U11058 ( .A(n9479), .B(n5277), .Z(n9478) );
  XOR U11059 ( .A(n9480), .B(n9481), .Z(n5277) );
  IV U11060 ( .A(n9477), .Z(n9480) );
  XNOR U11061 ( .A(n5278), .B(n9477), .Z(n9479) );
  NAND U11062 ( .A(n9482), .B(nreg[470]), .Z(n5278) );
  NAND U11063 ( .A(n6107), .B(nreg[470]), .Z(n9482) );
  XOR U11064 ( .A(n9483), .B(n9484), .Z(n9477) );
  ANDN U11065 ( .A(n9485), .B(n5279), .Z(n9484) );
  XOR U11066 ( .A(n9486), .B(n9487), .Z(n5279) );
  IV U11067 ( .A(n9483), .Z(n9486) );
  XNOR U11068 ( .A(n5280), .B(n9483), .Z(n9485) );
  NAND U11069 ( .A(n9488), .B(nreg[469]), .Z(n5280) );
  NAND U11070 ( .A(n6107), .B(nreg[469]), .Z(n9488) );
  XOR U11071 ( .A(n9489), .B(n9490), .Z(n9483) );
  ANDN U11072 ( .A(n9491), .B(n5281), .Z(n9490) );
  XOR U11073 ( .A(n9492), .B(n9493), .Z(n5281) );
  IV U11074 ( .A(n9489), .Z(n9492) );
  XNOR U11075 ( .A(n5282), .B(n9489), .Z(n9491) );
  NAND U11076 ( .A(n9494), .B(nreg[468]), .Z(n5282) );
  NAND U11077 ( .A(n6107), .B(nreg[468]), .Z(n9494) );
  XOR U11078 ( .A(n9495), .B(n9496), .Z(n9489) );
  ANDN U11079 ( .A(n9497), .B(n5283), .Z(n9496) );
  XOR U11080 ( .A(n9498), .B(n9499), .Z(n5283) );
  IV U11081 ( .A(n9495), .Z(n9498) );
  XNOR U11082 ( .A(n5284), .B(n9495), .Z(n9497) );
  NAND U11083 ( .A(n9500), .B(nreg[467]), .Z(n5284) );
  NAND U11084 ( .A(n6107), .B(nreg[467]), .Z(n9500) );
  XOR U11085 ( .A(n9501), .B(n9502), .Z(n9495) );
  ANDN U11086 ( .A(n9503), .B(n5287), .Z(n9502) );
  XOR U11087 ( .A(n9504), .B(n9505), .Z(n5287) );
  IV U11088 ( .A(n9501), .Z(n9504) );
  XNOR U11089 ( .A(n5288), .B(n9501), .Z(n9503) );
  NAND U11090 ( .A(n9506), .B(nreg[466]), .Z(n5288) );
  NAND U11091 ( .A(n6107), .B(nreg[466]), .Z(n9506) );
  XOR U11092 ( .A(n9507), .B(n9508), .Z(n9501) );
  ANDN U11093 ( .A(n9509), .B(n5289), .Z(n9508) );
  XOR U11094 ( .A(n9510), .B(n9511), .Z(n5289) );
  IV U11095 ( .A(n9507), .Z(n9510) );
  XNOR U11096 ( .A(n5290), .B(n9507), .Z(n9509) );
  NAND U11097 ( .A(n9512), .B(nreg[465]), .Z(n5290) );
  NAND U11098 ( .A(n6107), .B(nreg[465]), .Z(n9512) );
  XOR U11099 ( .A(n9513), .B(n9514), .Z(n9507) );
  ANDN U11100 ( .A(n9515), .B(n5291), .Z(n9514) );
  XOR U11101 ( .A(n9516), .B(n9517), .Z(n5291) );
  IV U11102 ( .A(n9513), .Z(n9516) );
  XNOR U11103 ( .A(n5292), .B(n9513), .Z(n9515) );
  NAND U11104 ( .A(n9518), .B(nreg[464]), .Z(n5292) );
  NAND U11105 ( .A(n6107), .B(nreg[464]), .Z(n9518) );
  XOR U11106 ( .A(n9519), .B(n9520), .Z(n9513) );
  ANDN U11107 ( .A(n9521), .B(n5293), .Z(n9520) );
  XOR U11108 ( .A(n9522), .B(n9523), .Z(n5293) );
  IV U11109 ( .A(n9519), .Z(n9522) );
  XNOR U11110 ( .A(n5294), .B(n9519), .Z(n9521) );
  NAND U11111 ( .A(n9524), .B(nreg[463]), .Z(n5294) );
  NAND U11112 ( .A(n6107), .B(nreg[463]), .Z(n9524) );
  XOR U11113 ( .A(n9525), .B(n9526), .Z(n9519) );
  ANDN U11114 ( .A(n9527), .B(n5295), .Z(n9526) );
  XOR U11115 ( .A(n9528), .B(n9529), .Z(n5295) );
  IV U11116 ( .A(n9525), .Z(n9528) );
  XNOR U11117 ( .A(n5296), .B(n9525), .Z(n9527) );
  NAND U11118 ( .A(n9530), .B(nreg[462]), .Z(n5296) );
  NAND U11119 ( .A(n6107), .B(nreg[462]), .Z(n9530) );
  XOR U11120 ( .A(n9531), .B(n9532), .Z(n9525) );
  ANDN U11121 ( .A(n9533), .B(n5297), .Z(n9532) );
  XOR U11122 ( .A(n9534), .B(n9535), .Z(n5297) );
  IV U11123 ( .A(n9531), .Z(n9534) );
  XNOR U11124 ( .A(n5298), .B(n9531), .Z(n9533) );
  NAND U11125 ( .A(n9536), .B(nreg[461]), .Z(n5298) );
  NAND U11126 ( .A(n6107), .B(nreg[461]), .Z(n9536) );
  XOR U11127 ( .A(n9537), .B(n9538), .Z(n9531) );
  ANDN U11128 ( .A(n9539), .B(n5299), .Z(n9538) );
  XOR U11129 ( .A(n9540), .B(n9541), .Z(n5299) );
  IV U11130 ( .A(n9537), .Z(n9540) );
  XNOR U11131 ( .A(n5300), .B(n9537), .Z(n9539) );
  NAND U11132 ( .A(n9542), .B(nreg[460]), .Z(n5300) );
  NAND U11133 ( .A(n6107), .B(nreg[460]), .Z(n9542) );
  XOR U11134 ( .A(n9543), .B(n9544), .Z(n9537) );
  ANDN U11135 ( .A(n9545), .B(n5301), .Z(n9544) );
  XOR U11136 ( .A(n9546), .B(n9547), .Z(n5301) );
  IV U11137 ( .A(n9543), .Z(n9546) );
  XNOR U11138 ( .A(n5302), .B(n9543), .Z(n9545) );
  NAND U11139 ( .A(n9548), .B(nreg[459]), .Z(n5302) );
  NAND U11140 ( .A(n6107), .B(nreg[459]), .Z(n9548) );
  XOR U11141 ( .A(n9549), .B(n9550), .Z(n9543) );
  ANDN U11142 ( .A(n9551), .B(n5303), .Z(n9550) );
  XOR U11143 ( .A(n9552), .B(n9553), .Z(n5303) );
  IV U11144 ( .A(n9549), .Z(n9552) );
  XNOR U11145 ( .A(n5304), .B(n9549), .Z(n9551) );
  NAND U11146 ( .A(n9554), .B(nreg[458]), .Z(n5304) );
  NAND U11147 ( .A(n6107), .B(nreg[458]), .Z(n9554) );
  XOR U11148 ( .A(n9555), .B(n9556), .Z(n9549) );
  ANDN U11149 ( .A(n9557), .B(n5305), .Z(n9556) );
  XOR U11150 ( .A(n9558), .B(n9559), .Z(n5305) );
  IV U11151 ( .A(n9555), .Z(n9558) );
  XNOR U11152 ( .A(n5306), .B(n9555), .Z(n9557) );
  NAND U11153 ( .A(n9560), .B(nreg[457]), .Z(n5306) );
  NAND U11154 ( .A(n6107), .B(nreg[457]), .Z(n9560) );
  XOR U11155 ( .A(n9561), .B(n9562), .Z(n9555) );
  ANDN U11156 ( .A(n9563), .B(n5309), .Z(n9562) );
  XOR U11157 ( .A(n9564), .B(n9565), .Z(n5309) );
  IV U11158 ( .A(n9561), .Z(n9564) );
  XNOR U11159 ( .A(n5310), .B(n9561), .Z(n9563) );
  NAND U11160 ( .A(n9566), .B(nreg[456]), .Z(n5310) );
  NAND U11161 ( .A(n6107), .B(nreg[456]), .Z(n9566) );
  XOR U11162 ( .A(n9567), .B(n9568), .Z(n9561) );
  ANDN U11163 ( .A(n9569), .B(n5311), .Z(n9568) );
  XOR U11164 ( .A(n9570), .B(n9571), .Z(n5311) );
  IV U11165 ( .A(n9567), .Z(n9570) );
  XNOR U11166 ( .A(n5312), .B(n9567), .Z(n9569) );
  NAND U11167 ( .A(n9572), .B(nreg[455]), .Z(n5312) );
  NAND U11168 ( .A(n6107), .B(nreg[455]), .Z(n9572) );
  XOR U11169 ( .A(n9573), .B(n9574), .Z(n9567) );
  ANDN U11170 ( .A(n9575), .B(n5313), .Z(n9574) );
  XOR U11171 ( .A(n9576), .B(n9577), .Z(n5313) );
  IV U11172 ( .A(n9573), .Z(n9576) );
  XNOR U11173 ( .A(n5314), .B(n9573), .Z(n9575) );
  NAND U11174 ( .A(n9578), .B(nreg[454]), .Z(n5314) );
  NAND U11175 ( .A(n6107), .B(nreg[454]), .Z(n9578) );
  XOR U11176 ( .A(n9579), .B(n9580), .Z(n9573) );
  ANDN U11177 ( .A(n9581), .B(n5315), .Z(n9580) );
  XOR U11178 ( .A(n9582), .B(n9583), .Z(n5315) );
  IV U11179 ( .A(n9579), .Z(n9582) );
  XNOR U11180 ( .A(n5316), .B(n9579), .Z(n9581) );
  NAND U11181 ( .A(n9584), .B(nreg[453]), .Z(n5316) );
  NAND U11182 ( .A(n6107), .B(nreg[453]), .Z(n9584) );
  XOR U11183 ( .A(n9585), .B(n9586), .Z(n9579) );
  ANDN U11184 ( .A(n9587), .B(n5317), .Z(n9586) );
  XOR U11185 ( .A(n9588), .B(n9589), .Z(n5317) );
  IV U11186 ( .A(n9585), .Z(n9588) );
  XNOR U11187 ( .A(n5318), .B(n9585), .Z(n9587) );
  NAND U11188 ( .A(n9590), .B(nreg[452]), .Z(n5318) );
  NAND U11189 ( .A(n6107), .B(nreg[452]), .Z(n9590) );
  XOR U11190 ( .A(n9591), .B(n9592), .Z(n9585) );
  ANDN U11191 ( .A(n9593), .B(n5319), .Z(n9592) );
  XOR U11192 ( .A(n9594), .B(n9595), .Z(n5319) );
  IV U11193 ( .A(n9591), .Z(n9594) );
  XNOR U11194 ( .A(n5320), .B(n9591), .Z(n9593) );
  NAND U11195 ( .A(n9596), .B(nreg[451]), .Z(n5320) );
  NAND U11196 ( .A(n6107), .B(nreg[451]), .Z(n9596) );
  XOR U11197 ( .A(n9597), .B(n9598), .Z(n9591) );
  ANDN U11198 ( .A(n9599), .B(n5321), .Z(n9598) );
  XOR U11199 ( .A(n9600), .B(n9601), .Z(n5321) );
  IV U11200 ( .A(n9597), .Z(n9600) );
  XNOR U11201 ( .A(n5322), .B(n9597), .Z(n9599) );
  NAND U11202 ( .A(n9602), .B(nreg[450]), .Z(n5322) );
  NAND U11203 ( .A(n6107), .B(nreg[450]), .Z(n9602) );
  XOR U11204 ( .A(n9603), .B(n9604), .Z(n9597) );
  ANDN U11205 ( .A(n9605), .B(n5323), .Z(n9604) );
  XOR U11206 ( .A(n9606), .B(n9607), .Z(n5323) );
  IV U11207 ( .A(n9603), .Z(n9606) );
  XNOR U11208 ( .A(n5324), .B(n9603), .Z(n9605) );
  NAND U11209 ( .A(n9608), .B(nreg[449]), .Z(n5324) );
  NAND U11210 ( .A(n6107), .B(nreg[449]), .Z(n9608) );
  XOR U11211 ( .A(n9609), .B(n9610), .Z(n9603) );
  ANDN U11212 ( .A(n9611), .B(n5325), .Z(n9610) );
  XOR U11213 ( .A(n9612), .B(n9613), .Z(n5325) );
  IV U11214 ( .A(n9609), .Z(n9612) );
  XNOR U11215 ( .A(n5326), .B(n9609), .Z(n9611) );
  NAND U11216 ( .A(n9614), .B(nreg[448]), .Z(n5326) );
  NAND U11217 ( .A(n6107), .B(nreg[448]), .Z(n9614) );
  XOR U11218 ( .A(n9615), .B(n9616), .Z(n9609) );
  ANDN U11219 ( .A(n9617), .B(n5327), .Z(n9616) );
  XOR U11220 ( .A(n9618), .B(n9619), .Z(n5327) );
  IV U11221 ( .A(n9615), .Z(n9618) );
  XNOR U11222 ( .A(n5328), .B(n9615), .Z(n9617) );
  NAND U11223 ( .A(n9620), .B(nreg[447]), .Z(n5328) );
  NAND U11224 ( .A(n6107), .B(nreg[447]), .Z(n9620) );
  XOR U11225 ( .A(n9621), .B(n9622), .Z(n9615) );
  ANDN U11226 ( .A(n9623), .B(n5331), .Z(n9622) );
  XOR U11227 ( .A(n9624), .B(n9625), .Z(n5331) );
  IV U11228 ( .A(n9621), .Z(n9624) );
  XNOR U11229 ( .A(n5332), .B(n9621), .Z(n9623) );
  NAND U11230 ( .A(n9626), .B(nreg[446]), .Z(n5332) );
  NAND U11231 ( .A(n6107), .B(nreg[446]), .Z(n9626) );
  XOR U11232 ( .A(n9627), .B(n9628), .Z(n9621) );
  ANDN U11233 ( .A(n9629), .B(n5333), .Z(n9628) );
  XOR U11234 ( .A(n9630), .B(n9631), .Z(n5333) );
  IV U11235 ( .A(n9627), .Z(n9630) );
  XNOR U11236 ( .A(n5334), .B(n9627), .Z(n9629) );
  NAND U11237 ( .A(n9632), .B(nreg[445]), .Z(n5334) );
  NAND U11238 ( .A(n6107), .B(nreg[445]), .Z(n9632) );
  XOR U11239 ( .A(n9633), .B(n9634), .Z(n9627) );
  ANDN U11240 ( .A(n9635), .B(n5335), .Z(n9634) );
  XOR U11241 ( .A(n9636), .B(n9637), .Z(n5335) );
  IV U11242 ( .A(n9633), .Z(n9636) );
  XNOR U11243 ( .A(n5336), .B(n9633), .Z(n9635) );
  NAND U11244 ( .A(n9638), .B(nreg[444]), .Z(n5336) );
  NAND U11245 ( .A(n6107), .B(nreg[444]), .Z(n9638) );
  XOR U11246 ( .A(n9639), .B(n9640), .Z(n9633) );
  ANDN U11247 ( .A(n9641), .B(n5337), .Z(n9640) );
  XOR U11248 ( .A(n9642), .B(n9643), .Z(n5337) );
  IV U11249 ( .A(n9639), .Z(n9642) );
  XNOR U11250 ( .A(n5338), .B(n9639), .Z(n9641) );
  NAND U11251 ( .A(n9644), .B(nreg[443]), .Z(n5338) );
  NAND U11252 ( .A(n6107), .B(nreg[443]), .Z(n9644) );
  XOR U11253 ( .A(n9645), .B(n9646), .Z(n9639) );
  ANDN U11254 ( .A(n9647), .B(n5339), .Z(n9646) );
  XOR U11255 ( .A(n9648), .B(n9649), .Z(n5339) );
  IV U11256 ( .A(n9645), .Z(n9648) );
  XNOR U11257 ( .A(n5340), .B(n9645), .Z(n9647) );
  NAND U11258 ( .A(n9650), .B(nreg[442]), .Z(n5340) );
  NAND U11259 ( .A(n6107), .B(nreg[442]), .Z(n9650) );
  XOR U11260 ( .A(n9651), .B(n9652), .Z(n9645) );
  ANDN U11261 ( .A(n9653), .B(n5341), .Z(n9652) );
  XOR U11262 ( .A(n9654), .B(n9655), .Z(n5341) );
  IV U11263 ( .A(n9651), .Z(n9654) );
  XNOR U11264 ( .A(n5342), .B(n9651), .Z(n9653) );
  NAND U11265 ( .A(n9656), .B(nreg[441]), .Z(n5342) );
  NAND U11266 ( .A(n6107), .B(nreg[441]), .Z(n9656) );
  XOR U11267 ( .A(n9657), .B(n9658), .Z(n9651) );
  ANDN U11268 ( .A(n9659), .B(n5343), .Z(n9658) );
  XOR U11269 ( .A(n9660), .B(n9661), .Z(n5343) );
  IV U11270 ( .A(n9657), .Z(n9660) );
  XNOR U11271 ( .A(n5344), .B(n9657), .Z(n9659) );
  NAND U11272 ( .A(n9662), .B(nreg[440]), .Z(n5344) );
  NAND U11273 ( .A(n6107), .B(nreg[440]), .Z(n9662) );
  XOR U11274 ( .A(n9663), .B(n9664), .Z(n9657) );
  ANDN U11275 ( .A(n9665), .B(n5345), .Z(n9664) );
  XOR U11276 ( .A(n9666), .B(n9667), .Z(n5345) );
  IV U11277 ( .A(n9663), .Z(n9666) );
  XNOR U11278 ( .A(n5346), .B(n9663), .Z(n9665) );
  NAND U11279 ( .A(n9668), .B(nreg[439]), .Z(n5346) );
  NAND U11280 ( .A(n6107), .B(nreg[439]), .Z(n9668) );
  XOR U11281 ( .A(n9669), .B(n9670), .Z(n9663) );
  ANDN U11282 ( .A(n9671), .B(n5347), .Z(n9670) );
  XOR U11283 ( .A(n9672), .B(n9673), .Z(n5347) );
  IV U11284 ( .A(n9669), .Z(n9672) );
  XNOR U11285 ( .A(n5348), .B(n9669), .Z(n9671) );
  NAND U11286 ( .A(n9674), .B(nreg[438]), .Z(n5348) );
  NAND U11287 ( .A(n6107), .B(nreg[438]), .Z(n9674) );
  XOR U11288 ( .A(n9675), .B(n9676), .Z(n9669) );
  ANDN U11289 ( .A(n9677), .B(n5349), .Z(n9676) );
  XOR U11290 ( .A(n9678), .B(n9679), .Z(n5349) );
  IV U11291 ( .A(n9675), .Z(n9678) );
  XNOR U11292 ( .A(n5350), .B(n9675), .Z(n9677) );
  NAND U11293 ( .A(n9680), .B(nreg[437]), .Z(n5350) );
  NAND U11294 ( .A(n6107), .B(nreg[437]), .Z(n9680) );
  XOR U11295 ( .A(n9681), .B(n9682), .Z(n9675) );
  ANDN U11296 ( .A(n9683), .B(n5353), .Z(n9682) );
  XOR U11297 ( .A(n9684), .B(n9685), .Z(n5353) );
  IV U11298 ( .A(n9681), .Z(n9684) );
  XNOR U11299 ( .A(n5354), .B(n9681), .Z(n9683) );
  NAND U11300 ( .A(n9686), .B(nreg[436]), .Z(n5354) );
  NAND U11301 ( .A(n6107), .B(nreg[436]), .Z(n9686) );
  XOR U11302 ( .A(n9687), .B(n9688), .Z(n9681) );
  ANDN U11303 ( .A(n9689), .B(n5355), .Z(n9688) );
  XOR U11304 ( .A(n9690), .B(n9691), .Z(n5355) );
  IV U11305 ( .A(n9687), .Z(n9690) );
  XNOR U11306 ( .A(n5356), .B(n9687), .Z(n9689) );
  NAND U11307 ( .A(n9692), .B(nreg[435]), .Z(n5356) );
  NAND U11308 ( .A(n6107), .B(nreg[435]), .Z(n9692) );
  XOR U11309 ( .A(n9693), .B(n9694), .Z(n9687) );
  ANDN U11310 ( .A(n9695), .B(n5357), .Z(n9694) );
  XOR U11311 ( .A(n9696), .B(n9697), .Z(n5357) );
  IV U11312 ( .A(n9693), .Z(n9696) );
  XNOR U11313 ( .A(n5358), .B(n9693), .Z(n9695) );
  NAND U11314 ( .A(n9698), .B(nreg[434]), .Z(n5358) );
  NAND U11315 ( .A(n6107), .B(nreg[434]), .Z(n9698) );
  XOR U11316 ( .A(n9699), .B(n9700), .Z(n9693) );
  ANDN U11317 ( .A(n9701), .B(n5359), .Z(n9700) );
  XOR U11318 ( .A(n9702), .B(n9703), .Z(n5359) );
  IV U11319 ( .A(n9699), .Z(n9702) );
  XNOR U11320 ( .A(n5360), .B(n9699), .Z(n9701) );
  NAND U11321 ( .A(n9704), .B(nreg[433]), .Z(n5360) );
  NAND U11322 ( .A(n6107), .B(nreg[433]), .Z(n9704) );
  XOR U11323 ( .A(n9705), .B(n9706), .Z(n9699) );
  ANDN U11324 ( .A(n9707), .B(n5361), .Z(n9706) );
  XOR U11325 ( .A(n9708), .B(n9709), .Z(n5361) );
  IV U11326 ( .A(n9705), .Z(n9708) );
  XNOR U11327 ( .A(n5362), .B(n9705), .Z(n9707) );
  NAND U11328 ( .A(n9710), .B(nreg[432]), .Z(n5362) );
  NAND U11329 ( .A(n6107), .B(nreg[432]), .Z(n9710) );
  XOR U11330 ( .A(n9711), .B(n9712), .Z(n9705) );
  ANDN U11331 ( .A(n9713), .B(n5363), .Z(n9712) );
  XOR U11332 ( .A(n9714), .B(n9715), .Z(n5363) );
  IV U11333 ( .A(n9711), .Z(n9714) );
  XNOR U11334 ( .A(n5364), .B(n9711), .Z(n9713) );
  NAND U11335 ( .A(n9716), .B(nreg[431]), .Z(n5364) );
  NAND U11336 ( .A(n6107), .B(nreg[431]), .Z(n9716) );
  XOR U11337 ( .A(n9717), .B(n9718), .Z(n9711) );
  ANDN U11338 ( .A(n9719), .B(n5365), .Z(n9718) );
  XOR U11339 ( .A(n9720), .B(n9721), .Z(n5365) );
  IV U11340 ( .A(n9717), .Z(n9720) );
  XNOR U11341 ( .A(n5366), .B(n9717), .Z(n9719) );
  NAND U11342 ( .A(n9722), .B(nreg[430]), .Z(n5366) );
  NAND U11343 ( .A(n6107), .B(nreg[430]), .Z(n9722) );
  XOR U11344 ( .A(n9723), .B(n9724), .Z(n9717) );
  ANDN U11345 ( .A(n9725), .B(n5367), .Z(n9724) );
  XOR U11346 ( .A(n9726), .B(n9727), .Z(n5367) );
  IV U11347 ( .A(n9723), .Z(n9726) );
  XNOR U11348 ( .A(n5368), .B(n9723), .Z(n9725) );
  NAND U11349 ( .A(n9728), .B(nreg[429]), .Z(n5368) );
  NAND U11350 ( .A(n6107), .B(nreg[429]), .Z(n9728) );
  XOR U11351 ( .A(n9729), .B(n9730), .Z(n9723) );
  ANDN U11352 ( .A(n9731), .B(n5369), .Z(n9730) );
  XOR U11353 ( .A(n9732), .B(n9733), .Z(n5369) );
  IV U11354 ( .A(n9729), .Z(n9732) );
  XNOR U11355 ( .A(n5370), .B(n9729), .Z(n9731) );
  NAND U11356 ( .A(n9734), .B(nreg[428]), .Z(n5370) );
  NAND U11357 ( .A(n6107), .B(nreg[428]), .Z(n9734) );
  XOR U11358 ( .A(n9735), .B(n9736), .Z(n9729) );
  ANDN U11359 ( .A(n9737), .B(n5371), .Z(n9736) );
  XOR U11360 ( .A(n9738), .B(n9739), .Z(n5371) );
  IV U11361 ( .A(n9735), .Z(n9738) );
  XNOR U11362 ( .A(n5372), .B(n9735), .Z(n9737) );
  NAND U11363 ( .A(n9740), .B(nreg[427]), .Z(n5372) );
  NAND U11364 ( .A(n6107), .B(nreg[427]), .Z(n9740) );
  XOR U11365 ( .A(n9741), .B(n9742), .Z(n9735) );
  ANDN U11366 ( .A(n9743), .B(n5375), .Z(n9742) );
  XOR U11367 ( .A(n9744), .B(n9745), .Z(n5375) );
  IV U11368 ( .A(n9741), .Z(n9744) );
  XNOR U11369 ( .A(n5376), .B(n9741), .Z(n9743) );
  NAND U11370 ( .A(n9746), .B(nreg[426]), .Z(n5376) );
  NAND U11371 ( .A(n6107), .B(nreg[426]), .Z(n9746) );
  XOR U11372 ( .A(n9747), .B(n9748), .Z(n9741) );
  ANDN U11373 ( .A(n9749), .B(n5377), .Z(n9748) );
  XOR U11374 ( .A(n9750), .B(n9751), .Z(n5377) );
  IV U11375 ( .A(n9747), .Z(n9750) );
  XNOR U11376 ( .A(n5378), .B(n9747), .Z(n9749) );
  NAND U11377 ( .A(n9752), .B(nreg[425]), .Z(n5378) );
  NAND U11378 ( .A(n6107), .B(nreg[425]), .Z(n9752) );
  XOR U11379 ( .A(n9753), .B(n9754), .Z(n9747) );
  ANDN U11380 ( .A(n9755), .B(n5379), .Z(n9754) );
  XOR U11381 ( .A(n9756), .B(n9757), .Z(n5379) );
  IV U11382 ( .A(n9753), .Z(n9756) );
  XNOR U11383 ( .A(n5380), .B(n9753), .Z(n9755) );
  NAND U11384 ( .A(n9758), .B(nreg[424]), .Z(n5380) );
  NAND U11385 ( .A(n6107), .B(nreg[424]), .Z(n9758) );
  XOR U11386 ( .A(n9759), .B(n9760), .Z(n9753) );
  ANDN U11387 ( .A(n9761), .B(n5381), .Z(n9760) );
  XOR U11388 ( .A(n9762), .B(n9763), .Z(n5381) );
  IV U11389 ( .A(n9759), .Z(n9762) );
  XNOR U11390 ( .A(n5382), .B(n9759), .Z(n9761) );
  NAND U11391 ( .A(n9764), .B(nreg[423]), .Z(n5382) );
  NAND U11392 ( .A(n6107), .B(nreg[423]), .Z(n9764) );
  XOR U11393 ( .A(n9765), .B(n9766), .Z(n9759) );
  ANDN U11394 ( .A(n9767), .B(n5383), .Z(n9766) );
  XOR U11395 ( .A(n9768), .B(n9769), .Z(n5383) );
  IV U11396 ( .A(n9765), .Z(n9768) );
  XNOR U11397 ( .A(n5384), .B(n9765), .Z(n9767) );
  NAND U11398 ( .A(n9770), .B(nreg[422]), .Z(n5384) );
  NAND U11399 ( .A(n6107), .B(nreg[422]), .Z(n9770) );
  XOR U11400 ( .A(n9771), .B(n9772), .Z(n9765) );
  ANDN U11401 ( .A(n9773), .B(n5385), .Z(n9772) );
  XOR U11402 ( .A(n9774), .B(n9775), .Z(n5385) );
  IV U11403 ( .A(n9771), .Z(n9774) );
  XNOR U11404 ( .A(n5386), .B(n9771), .Z(n9773) );
  NAND U11405 ( .A(n9776), .B(nreg[421]), .Z(n5386) );
  NAND U11406 ( .A(n6107), .B(nreg[421]), .Z(n9776) );
  XOR U11407 ( .A(n9777), .B(n9778), .Z(n9771) );
  ANDN U11408 ( .A(n9779), .B(n5387), .Z(n9778) );
  XOR U11409 ( .A(n9780), .B(n9781), .Z(n5387) );
  IV U11410 ( .A(n9777), .Z(n9780) );
  XNOR U11411 ( .A(n5388), .B(n9777), .Z(n9779) );
  NAND U11412 ( .A(n9782), .B(nreg[420]), .Z(n5388) );
  NAND U11413 ( .A(n6107), .B(nreg[420]), .Z(n9782) );
  XOR U11414 ( .A(n9783), .B(n9784), .Z(n9777) );
  ANDN U11415 ( .A(n9785), .B(n5389), .Z(n9784) );
  XOR U11416 ( .A(n9786), .B(n9787), .Z(n5389) );
  IV U11417 ( .A(n9783), .Z(n9786) );
  XNOR U11418 ( .A(n5390), .B(n9783), .Z(n9785) );
  NAND U11419 ( .A(n9788), .B(nreg[419]), .Z(n5390) );
  NAND U11420 ( .A(n6107), .B(nreg[419]), .Z(n9788) );
  XOR U11421 ( .A(n9789), .B(n9790), .Z(n9783) );
  ANDN U11422 ( .A(n9791), .B(n5391), .Z(n9790) );
  XOR U11423 ( .A(n9792), .B(n9793), .Z(n5391) );
  IV U11424 ( .A(n9789), .Z(n9792) );
  XNOR U11425 ( .A(n5392), .B(n9789), .Z(n9791) );
  NAND U11426 ( .A(n9794), .B(nreg[418]), .Z(n5392) );
  NAND U11427 ( .A(n6107), .B(nreg[418]), .Z(n9794) );
  XOR U11428 ( .A(n9795), .B(n9796), .Z(n9789) );
  ANDN U11429 ( .A(n9797), .B(n5393), .Z(n9796) );
  XOR U11430 ( .A(n9798), .B(n9799), .Z(n5393) );
  IV U11431 ( .A(n9795), .Z(n9798) );
  XNOR U11432 ( .A(n5394), .B(n9795), .Z(n9797) );
  NAND U11433 ( .A(n9800), .B(nreg[417]), .Z(n5394) );
  NAND U11434 ( .A(n6107), .B(nreg[417]), .Z(n9800) );
  XOR U11435 ( .A(n9801), .B(n9802), .Z(n9795) );
  ANDN U11436 ( .A(n9803), .B(n5397), .Z(n9802) );
  XOR U11437 ( .A(n9804), .B(n9805), .Z(n5397) );
  IV U11438 ( .A(n9801), .Z(n9804) );
  XNOR U11439 ( .A(n5398), .B(n9801), .Z(n9803) );
  NAND U11440 ( .A(n9806), .B(nreg[416]), .Z(n5398) );
  NAND U11441 ( .A(n6107), .B(nreg[416]), .Z(n9806) );
  XOR U11442 ( .A(n9807), .B(n9808), .Z(n9801) );
  ANDN U11443 ( .A(n9809), .B(n5399), .Z(n9808) );
  XOR U11444 ( .A(n9810), .B(n9811), .Z(n5399) );
  IV U11445 ( .A(n9807), .Z(n9810) );
  XNOR U11446 ( .A(n5400), .B(n9807), .Z(n9809) );
  NAND U11447 ( .A(n9812), .B(nreg[415]), .Z(n5400) );
  NAND U11448 ( .A(n6107), .B(nreg[415]), .Z(n9812) );
  XOR U11449 ( .A(n9813), .B(n9814), .Z(n9807) );
  ANDN U11450 ( .A(n9815), .B(n5401), .Z(n9814) );
  XOR U11451 ( .A(n9816), .B(n9817), .Z(n5401) );
  IV U11452 ( .A(n9813), .Z(n9816) );
  XNOR U11453 ( .A(n5402), .B(n9813), .Z(n9815) );
  NAND U11454 ( .A(n9818), .B(nreg[414]), .Z(n5402) );
  NAND U11455 ( .A(n6107), .B(nreg[414]), .Z(n9818) );
  XOR U11456 ( .A(n9819), .B(n9820), .Z(n9813) );
  ANDN U11457 ( .A(n9821), .B(n5403), .Z(n9820) );
  XOR U11458 ( .A(n9822), .B(n9823), .Z(n5403) );
  IV U11459 ( .A(n9819), .Z(n9822) );
  XNOR U11460 ( .A(n5404), .B(n9819), .Z(n9821) );
  NAND U11461 ( .A(n9824), .B(nreg[413]), .Z(n5404) );
  NAND U11462 ( .A(n6107), .B(nreg[413]), .Z(n9824) );
  XOR U11463 ( .A(n9825), .B(n9826), .Z(n9819) );
  ANDN U11464 ( .A(n9827), .B(n5405), .Z(n9826) );
  XOR U11465 ( .A(n9828), .B(n9829), .Z(n5405) );
  IV U11466 ( .A(n9825), .Z(n9828) );
  XNOR U11467 ( .A(n5406), .B(n9825), .Z(n9827) );
  NAND U11468 ( .A(n9830), .B(nreg[412]), .Z(n5406) );
  NAND U11469 ( .A(n6107), .B(nreg[412]), .Z(n9830) );
  XOR U11470 ( .A(n9831), .B(n9832), .Z(n9825) );
  ANDN U11471 ( .A(n9833), .B(n5407), .Z(n9832) );
  XOR U11472 ( .A(n9834), .B(n9835), .Z(n5407) );
  IV U11473 ( .A(n9831), .Z(n9834) );
  XNOR U11474 ( .A(n5408), .B(n9831), .Z(n9833) );
  NAND U11475 ( .A(n9836), .B(nreg[411]), .Z(n5408) );
  NAND U11476 ( .A(n6107), .B(nreg[411]), .Z(n9836) );
  XOR U11477 ( .A(n9837), .B(n9838), .Z(n9831) );
  ANDN U11478 ( .A(n9839), .B(n5409), .Z(n9838) );
  XOR U11479 ( .A(n9840), .B(n9841), .Z(n5409) );
  IV U11480 ( .A(n9837), .Z(n9840) );
  XNOR U11481 ( .A(n5410), .B(n9837), .Z(n9839) );
  NAND U11482 ( .A(n9842), .B(nreg[410]), .Z(n5410) );
  NAND U11483 ( .A(n6107), .B(nreg[410]), .Z(n9842) );
  XOR U11484 ( .A(n9843), .B(n9844), .Z(n9837) );
  ANDN U11485 ( .A(n9845), .B(n5411), .Z(n9844) );
  XOR U11486 ( .A(n9846), .B(n9847), .Z(n5411) );
  IV U11487 ( .A(n9843), .Z(n9846) );
  XNOR U11488 ( .A(n5412), .B(n9843), .Z(n9845) );
  NAND U11489 ( .A(n9848), .B(nreg[409]), .Z(n5412) );
  NAND U11490 ( .A(n6107), .B(nreg[409]), .Z(n9848) );
  XOR U11491 ( .A(n9849), .B(n9850), .Z(n9843) );
  ANDN U11492 ( .A(n9851), .B(n5413), .Z(n9850) );
  XOR U11493 ( .A(n9852), .B(n9853), .Z(n5413) );
  IV U11494 ( .A(n9849), .Z(n9852) );
  XNOR U11495 ( .A(n5414), .B(n9849), .Z(n9851) );
  NAND U11496 ( .A(n9854), .B(nreg[408]), .Z(n5414) );
  NAND U11497 ( .A(n6107), .B(nreg[408]), .Z(n9854) );
  XOR U11498 ( .A(n9855), .B(n9856), .Z(n9849) );
  ANDN U11499 ( .A(n9857), .B(n5415), .Z(n9856) );
  XOR U11500 ( .A(n9858), .B(n9859), .Z(n5415) );
  IV U11501 ( .A(n9855), .Z(n9858) );
  XNOR U11502 ( .A(n5416), .B(n9855), .Z(n9857) );
  NAND U11503 ( .A(n9860), .B(nreg[407]), .Z(n5416) );
  NAND U11504 ( .A(n6107), .B(nreg[407]), .Z(n9860) );
  XOR U11505 ( .A(n9861), .B(n9862), .Z(n9855) );
  ANDN U11506 ( .A(n9863), .B(n5419), .Z(n9862) );
  XOR U11507 ( .A(n9864), .B(n9865), .Z(n5419) );
  IV U11508 ( .A(n9861), .Z(n9864) );
  XNOR U11509 ( .A(n5420), .B(n9861), .Z(n9863) );
  NAND U11510 ( .A(n9866), .B(nreg[406]), .Z(n5420) );
  NAND U11511 ( .A(n6107), .B(nreg[406]), .Z(n9866) );
  XOR U11512 ( .A(n9867), .B(n9868), .Z(n9861) );
  ANDN U11513 ( .A(n9869), .B(n5421), .Z(n9868) );
  XOR U11514 ( .A(n9870), .B(n9871), .Z(n5421) );
  IV U11515 ( .A(n9867), .Z(n9870) );
  XNOR U11516 ( .A(n5422), .B(n9867), .Z(n9869) );
  NAND U11517 ( .A(n9872), .B(nreg[405]), .Z(n5422) );
  NAND U11518 ( .A(n6107), .B(nreg[405]), .Z(n9872) );
  XOR U11519 ( .A(n9873), .B(n9874), .Z(n9867) );
  ANDN U11520 ( .A(n9875), .B(n5423), .Z(n9874) );
  XOR U11521 ( .A(n9876), .B(n9877), .Z(n5423) );
  IV U11522 ( .A(n9873), .Z(n9876) );
  XNOR U11523 ( .A(n5424), .B(n9873), .Z(n9875) );
  NAND U11524 ( .A(n9878), .B(nreg[404]), .Z(n5424) );
  NAND U11525 ( .A(n6107), .B(nreg[404]), .Z(n9878) );
  XOR U11526 ( .A(n9879), .B(n9880), .Z(n9873) );
  ANDN U11527 ( .A(n9881), .B(n5425), .Z(n9880) );
  XOR U11528 ( .A(n9882), .B(n9883), .Z(n5425) );
  IV U11529 ( .A(n9879), .Z(n9882) );
  XNOR U11530 ( .A(n5426), .B(n9879), .Z(n9881) );
  NAND U11531 ( .A(n9884), .B(nreg[403]), .Z(n5426) );
  NAND U11532 ( .A(n6107), .B(nreg[403]), .Z(n9884) );
  XOR U11533 ( .A(n9885), .B(n9886), .Z(n9879) );
  ANDN U11534 ( .A(n9887), .B(n5427), .Z(n9886) );
  XOR U11535 ( .A(n9888), .B(n9889), .Z(n5427) );
  IV U11536 ( .A(n9885), .Z(n9888) );
  XNOR U11537 ( .A(n5428), .B(n9885), .Z(n9887) );
  NAND U11538 ( .A(n9890), .B(nreg[402]), .Z(n5428) );
  NAND U11539 ( .A(n6107), .B(nreg[402]), .Z(n9890) );
  XOR U11540 ( .A(n9891), .B(n9892), .Z(n9885) );
  ANDN U11541 ( .A(n9893), .B(n5429), .Z(n9892) );
  XOR U11542 ( .A(n9894), .B(n9895), .Z(n5429) );
  IV U11543 ( .A(n9891), .Z(n9894) );
  XNOR U11544 ( .A(n5430), .B(n9891), .Z(n9893) );
  NAND U11545 ( .A(n9896), .B(nreg[401]), .Z(n5430) );
  NAND U11546 ( .A(n6107), .B(nreg[401]), .Z(n9896) );
  XOR U11547 ( .A(n9897), .B(n9898), .Z(n9891) );
  ANDN U11548 ( .A(n9899), .B(n5431), .Z(n9898) );
  XOR U11549 ( .A(n9900), .B(n9901), .Z(n5431) );
  IV U11550 ( .A(n9897), .Z(n9900) );
  XNOR U11551 ( .A(n5432), .B(n9897), .Z(n9899) );
  NAND U11552 ( .A(n9902), .B(nreg[400]), .Z(n5432) );
  NAND U11553 ( .A(n6107), .B(nreg[400]), .Z(n9902) );
  XOR U11554 ( .A(n9903), .B(n9904), .Z(n9897) );
  ANDN U11555 ( .A(n9905), .B(n5433), .Z(n9904) );
  XOR U11556 ( .A(n9906), .B(n9907), .Z(n5433) );
  IV U11557 ( .A(n9903), .Z(n9906) );
  XNOR U11558 ( .A(n5434), .B(n9903), .Z(n9905) );
  NAND U11559 ( .A(n9908), .B(nreg[399]), .Z(n5434) );
  NAND U11560 ( .A(n6107), .B(nreg[399]), .Z(n9908) );
  XOR U11561 ( .A(n9909), .B(n9910), .Z(n9903) );
  ANDN U11562 ( .A(n9911), .B(n5435), .Z(n9910) );
  XOR U11563 ( .A(n9912), .B(n9913), .Z(n5435) );
  IV U11564 ( .A(n9909), .Z(n9912) );
  XNOR U11565 ( .A(n5436), .B(n9909), .Z(n9911) );
  NAND U11566 ( .A(n9914), .B(nreg[398]), .Z(n5436) );
  NAND U11567 ( .A(n6107), .B(nreg[398]), .Z(n9914) );
  XOR U11568 ( .A(n9915), .B(n9916), .Z(n9909) );
  ANDN U11569 ( .A(n9917), .B(n5437), .Z(n9916) );
  XOR U11570 ( .A(n9918), .B(n9919), .Z(n5437) );
  IV U11571 ( .A(n9915), .Z(n9918) );
  XNOR U11572 ( .A(n5438), .B(n9915), .Z(n9917) );
  NAND U11573 ( .A(n9920), .B(nreg[397]), .Z(n5438) );
  NAND U11574 ( .A(n6107), .B(nreg[397]), .Z(n9920) );
  XOR U11575 ( .A(n9921), .B(n9922), .Z(n9915) );
  ANDN U11576 ( .A(n9923), .B(n5443), .Z(n9922) );
  XOR U11577 ( .A(n9924), .B(n9925), .Z(n5443) );
  IV U11578 ( .A(n9921), .Z(n9924) );
  XNOR U11579 ( .A(n5444), .B(n9921), .Z(n9923) );
  NAND U11580 ( .A(n9926), .B(nreg[396]), .Z(n5444) );
  NAND U11581 ( .A(n6107), .B(nreg[396]), .Z(n9926) );
  XOR U11582 ( .A(n9927), .B(n9928), .Z(n9921) );
  ANDN U11583 ( .A(n9929), .B(n5445), .Z(n9928) );
  XOR U11584 ( .A(n9930), .B(n9931), .Z(n5445) );
  IV U11585 ( .A(n9927), .Z(n9930) );
  XNOR U11586 ( .A(n5446), .B(n9927), .Z(n9929) );
  NAND U11587 ( .A(n9932), .B(nreg[395]), .Z(n5446) );
  NAND U11588 ( .A(n6107), .B(nreg[395]), .Z(n9932) );
  XOR U11589 ( .A(n9933), .B(n9934), .Z(n9927) );
  ANDN U11590 ( .A(n9935), .B(n5447), .Z(n9934) );
  XOR U11591 ( .A(n9936), .B(n9937), .Z(n5447) );
  IV U11592 ( .A(n9933), .Z(n9936) );
  XNOR U11593 ( .A(n5448), .B(n9933), .Z(n9935) );
  NAND U11594 ( .A(n9938), .B(nreg[394]), .Z(n5448) );
  NAND U11595 ( .A(n6107), .B(nreg[394]), .Z(n9938) );
  XOR U11596 ( .A(n9939), .B(n9940), .Z(n9933) );
  ANDN U11597 ( .A(n9941), .B(n5449), .Z(n9940) );
  XOR U11598 ( .A(n9942), .B(n9943), .Z(n5449) );
  IV U11599 ( .A(n9939), .Z(n9942) );
  XNOR U11600 ( .A(n5450), .B(n9939), .Z(n9941) );
  NAND U11601 ( .A(n9944), .B(nreg[393]), .Z(n5450) );
  NAND U11602 ( .A(n6107), .B(nreg[393]), .Z(n9944) );
  XOR U11603 ( .A(n9945), .B(n9946), .Z(n9939) );
  ANDN U11604 ( .A(n9947), .B(n5451), .Z(n9946) );
  XOR U11605 ( .A(n9948), .B(n9949), .Z(n5451) );
  IV U11606 ( .A(n9945), .Z(n9948) );
  XNOR U11607 ( .A(n5452), .B(n9945), .Z(n9947) );
  NAND U11608 ( .A(n9950), .B(nreg[392]), .Z(n5452) );
  NAND U11609 ( .A(n6107), .B(nreg[392]), .Z(n9950) );
  XOR U11610 ( .A(n9951), .B(n9952), .Z(n9945) );
  ANDN U11611 ( .A(n9953), .B(n5453), .Z(n9952) );
  XOR U11612 ( .A(n9954), .B(n9955), .Z(n5453) );
  IV U11613 ( .A(n9951), .Z(n9954) );
  XNOR U11614 ( .A(n5454), .B(n9951), .Z(n9953) );
  NAND U11615 ( .A(n9956), .B(nreg[391]), .Z(n5454) );
  NAND U11616 ( .A(n6107), .B(nreg[391]), .Z(n9956) );
  XOR U11617 ( .A(n9957), .B(n9958), .Z(n9951) );
  ANDN U11618 ( .A(n9959), .B(n5455), .Z(n9958) );
  XOR U11619 ( .A(n9960), .B(n9961), .Z(n5455) );
  IV U11620 ( .A(n9957), .Z(n9960) );
  XNOR U11621 ( .A(n5456), .B(n9957), .Z(n9959) );
  NAND U11622 ( .A(n9962), .B(nreg[390]), .Z(n5456) );
  NAND U11623 ( .A(n6107), .B(nreg[390]), .Z(n9962) );
  XOR U11624 ( .A(n9963), .B(n9964), .Z(n9957) );
  ANDN U11625 ( .A(n9965), .B(n5457), .Z(n9964) );
  XOR U11626 ( .A(n9966), .B(n9967), .Z(n5457) );
  IV U11627 ( .A(n9963), .Z(n9966) );
  XNOR U11628 ( .A(n5458), .B(n9963), .Z(n9965) );
  NAND U11629 ( .A(n9968), .B(nreg[389]), .Z(n5458) );
  NAND U11630 ( .A(n6107), .B(nreg[389]), .Z(n9968) );
  XOR U11631 ( .A(n9969), .B(n9970), .Z(n9963) );
  ANDN U11632 ( .A(n9971), .B(n5459), .Z(n9970) );
  XOR U11633 ( .A(n9972), .B(n9973), .Z(n5459) );
  IV U11634 ( .A(n9969), .Z(n9972) );
  XNOR U11635 ( .A(n5460), .B(n9969), .Z(n9971) );
  NAND U11636 ( .A(n9974), .B(nreg[388]), .Z(n5460) );
  NAND U11637 ( .A(n6107), .B(nreg[388]), .Z(n9974) );
  XOR U11638 ( .A(n9975), .B(n9976), .Z(n9969) );
  ANDN U11639 ( .A(n9977), .B(n5461), .Z(n9976) );
  XOR U11640 ( .A(n9978), .B(n9979), .Z(n5461) );
  IV U11641 ( .A(n9975), .Z(n9978) );
  XNOR U11642 ( .A(n5462), .B(n9975), .Z(n9977) );
  NAND U11643 ( .A(n9980), .B(nreg[387]), .Z(n5462) );
  NAND U11644 ( .A(n6107), .B(nreg[387]), .Z(n9980) );
  XOR U11645 ( .A(n9981), .B(n9982), .Z(n9975) );
  ANDN U11646 ( .A(n9983), .B(n5465), .Z(n9982) );
  XOR U11647 ( .A(n9984), .B(n9985), .Z(n5465) );
  IV U11648 ( .A(n9981), .Z(n9984) );
  XNOR U11649 ( .A(n5466), .B(n9981), .Z(n9983) );
  NAND U11650 ( .A(n9986), .B(nreg[386]), .Z(n5466) );
  NAND U11651 ( .A(n6107), .B(nreg[386]), .Z(n9986) );
  XOR U11652 ( .A(n9987), .B(n9988), .Z(n9981) );
  ANDN U11653 ( .A(n9989), .B(n5467), .Z(n9988) );
  XOR U11654 ( .A(n9990), .B(n9991), .Z(n5467) );
  IV U11655 ( .A(n9987), .Z(n9990) );
  XNOR U11656 ( .A(n5468), .B(n9987), .Z(n9989) );
  NAND U11657 ( .A(n9992), .B(nreg[385]), .Z(n5468) );
  NAND U11658 ( .A(n6107), .B(nreg[385]), .Z(n9992) );
  XOR U11659 ( .A(n9993), .B(n9994), .Z(n9987) );
  ANDN U11660 ( .A(n9995), .B(n5469), .Z(n9994) );
  XOR U11661 ( .A(n9996), .B(n9997), .Z(n5469) );
  IV U11662 ( .A(n9993), .Z(n9996) );
  XNOR U11663 ( .A(n5470), .B(n9993), .Z(n9995) );
  NAND U11664 ( .A(n9998), .B(nreg[384]), .Z(n5470) );
  NAND U11665 ( .A(n6107), .B(nreg[384]), .Z(n9998) );
  XOR U11666 ( .A(n9999), .B(n10000), .Z(n9993) );
  ANDN U11667 ( .A(n10001), .B(n5471), .Z(n10000) );
  XOR U11668 ( .A(n10002), .B(n10003), .Z(n5471) );
  IV U11669 ( .A(n9999), .Z(n10002) );
  XNOR U11670 ( .A(n5472), .B(n9999), .Z(n10001) );
  NAND U11671 ( .A(n10004), .B(nreg[383]), .Z(n5472) );
  NAND U11672 ( .A(n6107), .B(nreg[383]), .Z(n10004) );
  XOR U11673 ( .A(n10005), .B(n10006), .Z(n9999) );
  ANDN U11674 ( .A(n10007), .B(n5473), .Z(n10006) );
  XOR U11675 ( .A(n10008), .B(n10009), .Z(n5473) );
  IV U11676 ( .A(n10005), .Z(n10008) );
  XNOR U11677 ( .A(n5474), .B(n10005), .Z(n10007) );
  NAND U11678 ( .A(n10010), .B(nreg[382]), .Z(n5474) );
  NAND U11679 ( .A(n6107), .B(nreg[382]), .Z(n10010) );
  XOR U11680 ( .A(n10011), .B(n10012), .Z(n10005) );
  ANDN U11681 ( .A(n10013), .B(n5475), .Z(n10012) );
  XOR U11682 ( .A(n10014), .B(n10015), .Z(n5475) );
  IV U11683 ( .A(n10011), .Z(n10014) );
  XNOR U11684 ( .A(n5476), .B(n10011), .Z(n10013) );
  NAND U11685 ( .A(n10016), .B(nreg[381]), .Z(n5476) );
  NAND U11686 ( .A(n6107), .B(nreg[381]), .Z(n10016) );
  XOR U11687 ( .A(n10017), .B(n10018), .Z(n10011) );
  ANDN U11688 ( .A(n10019), .B(n5477), .Z(n10018) );
  XOR U11689 ( .A(n10020), .B(n10021), .Z(n5477) );
  IV U11690 ( .A(n10017), .Z(n10020) );
  XNOR U11691 ( .A(n5478), .B(n10017), .Z(n10019) );
  NAND U11692 ( .A(n10022), .B(nreg[380]), .Z(n5478) );
  NAND U11693 ( .A(n6107), .B(nreg[380]), .Z(n10022) );
  XOR U11694 ( .A(n10023), .B(n10024), .Z(n10017) );
  ANDN U11695 ( .A(n10025), .B(n5479), .Z(n10024) );
  XOR U11696 ( .A(n10026), .B(n10027), .Z(n5479) );
  IV U11697 ( .A(n10023), .Z(n10026) );
  XNOR U11698 ( .A(n5480), .B(n10023), .Z(n10025) );
  NAND U11699 ( .A(n10028), .B(nreg[379]), .Z(n5480) );
  NAND U11700 ( .A(n6107), .B(nreg[379]), .Z(n10028) );
  XOR U11701 ( .A(n10029), .B(n10030), .Z(n10023) );
  ANDN U11702 ( .A(n10031), .B(n5481), .Z(n10030) );
  XOR U11703 ( .A(n10032), .B(n10033), .Z(n5481) );
  IV U11704 ( .A(n10029), .Z(n10032) );
  XNOR U11705 ( .A(n5482), .B(n10029), .Z(n10031) );
  NAND U11706 ( .A(n10034), .B(nreg[378]), .Z(n5482) );
  NAND U11707 ( .A(n6107), .B(nreg[378]), .Z(n10034) );
  XOR U11708 ( .A(n10035), .B(n10036), .Z(n10029) );
  ANDN U11709 ( .A(n10037), .B(n5483), .Z(n10036) );
  XOR U11710 ( .A(n10038), .B(n10039), .Z(n5483) );
  IV U11711 ( .A(n10035), .Z(n10038) );
  XNOR U11712 ( .A(n5484), .B(n10035), .Z(n10037) );
  NAND U11713 ( .A(n10040), .B(nreg[377]), .Z(n5484) );
  NAND U11714 ( .A(n6107), .B(nreg[377]), .Z(n10040) );
  XOR U11715 ( .A(n10041), .B(n10042), .Z(n10035) );
  ANDN U11716 ( .A(n10043), .B(n5487), .Z(n10042) );
  XOR U11717 ( .A(n10044), .B(n10045), .Z(n5487) );
  IV U11718 ( .A(n10041), .Z(n10044) );
  XNOR U11719 ( .A(n5488), .B(n10041), .Z(n10043) );
  NAND U11720 ( .A(n10046), .B(nreg[376]), .Z(n5488) );
  NAND U11721 ( .A(n6107), .B(nreg[376]), .Z(n10046) );
  XOR U11722 ( .A(n10047), .B(n10048), .Z(n10041) );
  ANDN U11723 ( .A(n10049), .B(n5489), .Z(n10048) );
  XOR U11724 ( .A(n10050), .B(n10051), .Z(n5489) );
  IV U11725 ( .A(n10047), .Z(n10050) );
  XNOR U11726 ( .A(n5490), .B(n10047), .Z(n10049) );
  NAND U11727 ( .A(n10052), .B(nreg[375]), .Z(n5490) );
  NAND U11728 ( .A(n6107), .B(nreg[375]), .Z(n10052) );
  XOR U11729 ( .A(n10053), .B(n10054), .Z(n10047) );
  ANDN U11730 ( .A(n10055), .B(n5491), .Z(n10054) );
  XOR U11731 ( .A(n10056), .B(n10057), .Z(n5491) );
  IV U11732 ( .A(n10053), .Z(n10056) );
  XNOR U11733 ( .A(n5492), .B(n10053), .Z(n10055) );
  NAND U11734 ( .A(n10058), .B(nreg[374]), .Z(n5492) );
  NAND U11735 ( .A(n6107), .B(nreg[374]), .Z(n10058) );
  XOR U11736 ( .A(n10059), .B(n10060), .Z(n10053) );
  ANDN U11737 ( .A(n10061), .B(n5493), .Z(n10060) );
  XOR U11738 ( .A(n10062), .B(n10063), .Z(n5493) );
  IV U11739 ( .A(n10059), .Z(n10062) );
  XNOR U11740 ( .A(n5494), .B(n10059), .Z(n10061) );
  NAND U11741 ( .A(n10064), .B(nreg[373]), .Z(n5494) );
  NAND U11742 ( .A(n6107), .B(nreg[373]), .Z(n10064) );
  XOR U11743 ( .A(n10065), .B(n10066), .Z(n10059) );
  ANDN U11744 ( .A(n10067), .B(n5495), .Z(n10066) );
  XOR U11745 ( .A(n10068), .B(n10069), .Z(n5495) );
  IV U11746 ( .A(n10065), .Z(n10068) );
  XNOR U11747 ( .A(n5496), .B(n10065), .Z(n10067) );
  NAND U11748 ( .A(n10070), .B(nreg[372]), .Z(n5496) );
  NAND U11749 ( .A(n6107), .B(nreg[372]), .Z(n10070) );
  XOR U11750 ( .A(n10071), .B(n10072), .Z(n10065) );
  ANDN U11751 ( .A(n10073), .B(n5497), .Z(n10072) );
  XOR U11752 ( .A(n10074), .B(n10075), .Z(n5497) );
  IV U11753 ( .A(n10071), .Z(n10074) );
  XNOR U11754 ( .A(n5498), .B(n10071), .Z(n10073) );
  NAND U11755 ( .A(n10076), .B(nreg[371]), .Z(n5498) );
  NAND U11756 ( .A(n6107), .B(nreg[371]), .Z(n10076) );
  XOR U11757 ( .A(n10077), .B(n10078), .Z(n10071) );
  ANDN U11758 ( .A(n10079), .B(n5499), .Z(n10078) );
  XOR U11759 ( .A(n10080), .B(n10081), .Z(n5499) );
  IV U11760 ( .A(n10077), .Z(n10080) );
  XNOR U11761 ( .A(n5500), .B(n10077), .Z(n10079) );
  NAND U11762 ( .A(n10082), .B(nreg[370]), .Z(n5500) );
  NAND U11763 ( .A(n6107), .B(nreg[370]), .Z(n10082) );
  XOR U11764 ( .A(n10083), .B(n10084), .Z(n10077) );
  ANDN U11765 ( .A(n10085), .B(n5501), .Z(n10084) );
  XOR U11766 ( .A(n10086), .B(n10087), .Z(n5501) );
  IV U11767 ( .A(n10083), .Z(n10086) );
  XNOR U11768 ( .A(n5502), .B(n10083), .Z(n10085) );
  NAND U11769 ( .A(n10088), .B(nreg[369]), .Z(n5502) );
  NAND U11770 ( .A(n6107), .B(nreg[369]), .Z(n10088) );
  XOR U11771 ( .A(n10089), .B(n10090), .Z(n10083) );
  ANDN U11772 ( .A(n10091), .B(n5503), .Z(n10090) );
  XOR U11773 ( .A(n10092), .B(n10093), .Z(n5503) );
  IV U11774 ( .A(n10089), .Z(n10092) );
  XNOR U11775 ( .A(n5504), .B(n10089), .Z(n10091) );
  NAND U11776 ( .A(n10094), .B(nreg[368]), .Z(n5504) );
  NAND U11777 ( .A(n6107), .B(nreg[368]), .Z(n10094) );
  XOR U11778 ( .A(n10095), .B(n10096), .Z(n10089) );
  ANDN U11779 ( .A(n10097), .B(n5505), .Z(n10096) );
  XOR U11780 ( .A(n10098), .B(n10099), .Z(n5505) );
  IV U11781 ( .A(n10095), .Z(n10098) );
  XNOR U11782 ( .A(n5506), .B(n10095), .Z(n10097) );
  NAND U11783 ( .A(n10100), .B(nreg[367]), .Z(n5506) );
  NAND U11784 ( .A(n6107), .B(nreg[367]), .Z(n10100) );
  XOR U11785 ( .A(n10101), .B(n10102), .Z(n10095) );
  ANDN U11786 ( .A(n10103), .B(n5509), .Z(n10102) );
  XOR U11787 ( .A(n10104), .B(n10105), .Z(n5509) );
  IV U11788 ( .A(n10101), .Z(n10104) );
  XNOR U11789 ( .A(n5510), .B(n10101), .Z(n10103) );
  NAND U11790 ( .A(n10106), .B(nreg[366]), .Z(n5510) );
  NAND U11791 ( .A(n6107), .B(nreg[366]), .Z(n10106) );
  XOR U11792 ( .A(n10107), .B(n10108), .Z(n10101) );
  ANDN U11793 ( .A(n10109), .B(n5511), .Z(n10108) );
  XOR U11794 ( .A(n10110), .B(n10111), .Z(n5511) );
  IV U11795 ( .A(n10107), .Z(n10110) );
  XNOR U11796 ( .A(n5512), .B(n10107), .Z(n10109) );
  NAND U11797 ( .A(n10112), .B(nreg[365]), .Z(n5512) );
  NAND U11798 ( .A(n6107), .B(nreg[365]), .Z(n10112) );
  XOR U11799 ( .A(n10113), .B(n10114), .Z(n10107) );
  ANDN U11800 ( .A(n10115), .B(n5513), .Z(n10114) );
  XOR U11801 ( .A(n10116), .B(n10117), .Z(n5513) );
  IV U11802 ( .A(n10113), .Z(n10116) );
  XNOR U11803 ( .A(n5514), .B(n10113), .Z(n10115) );
  NAND U11804 ( .A(n10118), .B(nreg[364]), .Z(n5514) );
  NAND U11805 ( .A(n6107), .B(nreg[364]), .Z(n10118) );
  XOR U11806 ( .A(n10119), .B(n10120), .Z(n10113) );
  ANDN U11807 ( .A(n10121), .B(n5515), .Z(n10120) );
  XOR U11808 ( .A(n10122), .B(n10123), .Z(n5515) );
  IV U11809 ( .A(n10119), .Z(n10122) );
  XNOR U11810 ( .A(n5516), .B(n10119), .Z(n10121) );
  NAND U11811 ( .A(n10124), .B(nreg[363]), .Z(n5516) );
  NAND U11812 ( .A(n6107), .B(nreg[363]), .Z(n10124) );
  XOR U11813 ( .A(n10125), .B(n10126), .Z(n10119) );
  ANDN U11814 ( .A(n10127), .B(n5517), .Z(n10126) );
  XOR U11815 ( .A(n10128), .B(n10129), .Z(n5517) );
  IV U11816 ( .A(n10125), .Z(n10128) );
  XNOR U11817 ( .A(n5518), .B(n10125), .Z(n10127) );
  NAND U11818 ( .A(n10130), .B(nreg[362]), .Z(n5518) );
  NAND U11819 ( .A(n6107), .B(nreg[362]), .Z(n10130) );
  XOR U11820 ( .A(n10131), .B(n10132), .Z(n10125) );
  ANDN U11821 ( .A(n10133), .B(n5519), .Z(n10132) );
  XOR U11822 ( .A(n10134), .B(n10135), .Z(n5519) );
  IV U11823 ( .A(n10131), .Z(n10134) );
  XNOR U11824 ( .A(n5520), .B(n10131), .Z(n10133) );
  NAND U11825 ( .A(n10136), .B(nreg[361]), .Z(n5520) );
  NAND U11826 ( .A(n6107), .B(nreg[361]), .Z(n10136) );
  XOR U11827 ( .A(n10137), .B(n10138), .Z(n10131) );
  ANDN U11828 ( .A(n10139), .B(n5521), .Z(n10138) );
  XOR U11829 ( .A(n10140), .B(n10141), .Z(n5521) );
  IV U11830 ( .A(n10137), .Z(n10140) );
  XNOR U11831 ( .A(n5522), .B(n10137), .Z(n10139) );
  NAND U11832 ( .A(n10142), .B(nreg[360]), .Z(n5522) );
  NAND U11833 ( .A(n6107), .B(nreg[360]), .Z(n10142) );
  XOR U11834 ( .A(n10143), .B(n10144), .Z(n10137) );
  ANDN U11835 ( .A(n10145), .B(n5523), .Z(n10144) );
  XOR U11836 ( .A(n10146), .B(n10147), .Z(n5523) );
  IV U11837 ( .A(n10143), .Z(n10146) );
  XNOR U11838 ( .A(n5524), .B(n10143), .Z(n10145) );
  NAND U11839 ( .A(n10148), .B(nreg[359]), .Z(n5524) );
  NAND U11840 ( .A(n6107), .B(nreg[359]), .Z(n10148) );
  XOR U11841 ( .A(n10149), .B(n10150), .Z(n10143) );
  ANDN U11842 ( .A(n10151), .B(n5525), .Z(n10150) );
  XOR U11843 ( .A(n10152), .B(n10153), .Z(n5525) );
  IV U11844 ( .A(n10149), .Z(n10152) );
  XNOR U11845 ( .A(n5526), .B(n10149), .Z(n10151) );
  NAND U11846 ( .A(n10154), .B(nreg[358]), .Z(n5526) );
  NAND U11847 ( .A(n6107), .B(nreg[358]), .Z(n10154) );
  XOR U11848 ( .A(n10155), .B(n10156), .Z(n10149) );
  ANDN U11849 ( .A(n10157), .B(n5527), .Z(n10156) );
  XOR U11850 ( .A(n10158), .B(n10159), .Z(n5527) );
  IV U11851 ( .A(n10155), .Z(n10158) );
  XNOR U11852 ( .A(n5528), .B(n10155), .Z(n10157) );
  NAND U11853 ( .A(n10160), .B(nreg[357]), .Z(n5528) );
  NAND U11854 ( .A(n6107), .B(nreg[357]), .Z(n10160) );
  XOR U11855 ( .A(n10161), .B(n10162), .Z(n10155) );
  ANDN U11856 ( .A(n10163), .B(n5531), .Z(n10162) );
  XOR U11857 ( .A(n10164), .B(n10165), .Z(n5531) );
  IV U11858 ( .A(n10161), .Z(n10164) );
  XNOR U11859 ( .A(n5532), .B(n10161), .Z(n10163) );
  NAND U11860 ( .A(n10166), .B(nreg[356]), .Z(n5532) );
  NAND U11861 ( .A(n6107), .B(nreg[356]), .Z(n10166) );
  XOR U11862 ( .A(n10167), .B(n10168), .Z(n10161) );
  ANDN U11863 ( .A(n10169), .B(n5533), .Z(n10168) );
  XOR U11864 ( .A(n10170), .B(n10171), .Z(n5533) );
  IV U11865 ( .A(n10167), .Z(n10170) );
  XNOR U11866 ( .A(n5534), .B(n10167), .Z(n10169) );
  NAND U11867 ( .A(n10172), .B(nreg[355]), .Z(n5534) );
  NAND U11868 ( .A(n6107), .B(nreg[355]), .Z(n10172) );
  XOR U11869 ( .A(n10173), .B(n10174), .Z(n10167) );
  ANDN U11870 ( .A(n10175), .B(n5535), .Z(n10174) );
  XOR U11871 ( .A(n10176), .B(n10177), .Z(n5535) );
  IV U11872 ( .A(n10173), .Z(n10176) );
  XNOR U11873 ( .A(n5536), .B(n10173), .Z(n10175) );
  NAND U11874 ( .A(n10178), .B(nreg[354]), .Z(n5536) );
  NAND U11875 ( .A(n6107), .B(nreg[354]), .Z(n10178) );
  XOR U11876 ( .A(n10179), .B(n10180), .Z(n10173) );
  ANDN U11877 ( .A(n10181), .B(n5537), .Z(n10180) );
  XOR U11878 ( .A(n10182), .B(n10183), .Z(n5537) );
  IV U11879 ( .A(n10179), .Z(n10182) );
  XNOR U11880 ( .A(n5538), .B(n10179), .Z(n10181) );
  NAND U11881 ( .A(n10184), .B(nreg[353]), .Z(n5538) );
  NAND U11882 ( .A(n6107), .B(nreg[353]), .Z(n10184) );
  XOR U11883 ( .A(n10185), .B(n10186), .Z(n10179) );
  ANDN U11884 ( .A(n10187), .B(n5539), .Z(n10186) );
  XOR U11885 ( .A(n10188), .B(n10189), .Z(n5539) );
  IV U11886 ( .A(n10185), .Z(n10188) );
  XNOR U11887 ( .A(n5540), .B(n10185), .Z(n10187) );
  NAND U11888 ( .A(n10190), .B(nreg[352]), .Z(n5540) );
  NAND U11889 ( .A(n6107), .B(nreg[352]), .Z(n10190) );
  XOR U11890 ( .A(n10191), .B(n10192), .Z(n10185) );
  ANDN U11891 ( .A(n10193), .B(n5541), .Z(n10192) );
  XOR U11892 ( .A(n10194), .B(n10195), .Z(n5541) );
  IV U11893 ( .A(n10191), .Z(n10194) );
  XNOR U11894 ( .A(n5542), .B(n10191), .Z(n10193) );
  NAND U11895 ( .A(n10196), .B(nreg[351]), .Z(n5542) );
  NAND U11896 ( .A(n6107), .B(nreg[351]), .Z(n10196) );
  XOR U11897 ( .A(n10197), .B(n10198), .Z(n10191) );
  ANDN U11898 ( .A(n10199), .B(n5543), .Z(n10198) );
  XOR U11899 ( .A(n10200), .B(n10201), .Z(n5543) );
  IV U11900 ( .A(n10197), .Z(n10200) );
  XNOR U11901 ( .A(n5544), .B(n10197), .Z(n10199) );
  NAND U11902 ( .A(n10202), .B(nreg[350]), .Z(n5544) );
  NAND U11903 ( .A(n6107), .B(nreg[350]), .Z(n10202) );
  XOR U11904 ( .A(n10203), .B(n10204), .Z(n10197) );
  ANDN U11905 ( .A(n10205), .B(n5545), .Z(n10204) );
  XOR U11906 ( .A(n10206), .B(n10207), .Z(n5545) );
  IV U11907 ( .A(n10203), .Z(n10206) );
  XNOR U11908 ( .A(n5546), .B(n10203), .Z(n10205) );
  NAND U11909 ( .A(n10208), .B(nreg[349]), .Z(n5546) );
  NAND U11910 ( .A(n6107), .B(nreg[349]), .Z(n10208) );
  XOR U11911 ( .A(n10209), .B(n10210), .Z(n10203) );
  ANDN U11912 ( .A(n10211), .B(n5547), .Z(n10210) );
  XOR U11913 ( .A(n10212), .B(n10213), .Z(n5547) );
  IV U11914 ( .A(n10209), .Z(n10212) );
  XNOR U11915 ( .A(n5548), .B(n10209), .Z(n10211) );
  NAND U11916 ( .A(n10214), .B(nreg[348]), .Z(n5548) );
  NAND U11917 ( .A(n6107), .B(nreg[348]), .Z(n10214) );
  XOR U11918 ( .A(n10215), .B(n10216), .Z(n10209) );
  ANDN U11919 ( .A(n10217), .B(n5549), .Z(n10216) );
  XOR U11920 ( .A(n10218), .B(n10219), .Z(n5549) );
  IV U11921 ( .A(n10215), .Z(n10218) );
  XNOR U11922 ( .A(n5550), .B(n10215), .Z(n10217) );
  NAND U11923 ( .A(n10220), .B(nreg[347]), .Z(n5550) );
  NAND U11924 ( .A(n6107), .B(nreg[347]), .Z(n10220) );
  XOR U11925 ( .A(n10221), .B(n10222), .Z(n10215) );
  ANDN U11926 ( .A(n10223), .B(n5553), .Z(n10222) );
  XOR U11927 ( .A(n10224), .B(n10225), .Z(n5553) );
  IV U11928 ( .A(n10221), .Z(n10224) );
  XNOR U11929 ( .A(n5554), .B(n10221), .Z(n10223) );
  NAND U11930 ( .A(n10226), .B(nreg[346]), .Z(n5554) );
  NAND U11931 ( .A(n6107), .B(nreg[346]), .Z(n10226) );
  XOR U11932 ( .A(n10227), .B(n10228), .Z(n10221) );
  ANDN U11933 ( .A(n10229), .B(n5555), .Z(n10228) );
  XOR U11934 ( .A(n10230), .B(n10231), .Z(n5555) );
  IV U11935 ( .A(n10227), .Z(n10230) );
  XNOR U11936 ( .A(n5556), .B(n10227), .Z(n10229) );
  NAND U11937 ( .A(n10232), .B(nreg[345]), .Z(n5556) );
  NAND U11938 ( .A(n6107), .B(nreg[345]), .Z(n10232) );
  XOR U11939 ( .A(n10233), .B(n10234), .Z(n10227) );
  ANDN U11940 ( .A(n10235), .B(n5557), .Z(n10234) );
  XOR U11941 ( .A(n10236), .B(n10237), .Z(n5557) );
  IV U11942 ( .A(n10233), .Z(n10236) );
  XNOR U11943 ( .A(n5558), .B(n10233), .Z(n10235) );
  NAND U11944 ( .A(n10238), .B(nreg[344]), .Z(n5558) );
  NAND U11945 ( .A(n6107), .B(nreg[344]), .Z(n10238) );
  XOR U11946 ( .A(n10239), .B(n10240), .Z(n10233) );
  ANDN U11947 ( .A(n10241), .B(n5559), .Z(n10240) );
  XOR U11948 ( .A(n10242), .B(n10243), .Z(n5559) );
  IV U11949 ( .A(n10239), .Z(n10242) );
  XNOR U11950 ( .A(n5560), .B(n10239), .Z(n10241) );
  NAND U11951 ( .A(n10244), .B(nreg[343]), .Z(n5560) );
  NAND U11952 ( .A(n6107), .B(nreg[343]), .Z(n10244) );
  XOR U11953 ( .A(n10245), .B(n10246), .Z(n10239) );
  ANDN U11954 ( .A(n10247), .B(n5561), .Z(n10246) );
  XOR U11955 ( .A(n10248), .B(n10249), .Z(n5561) );
  IV U11956 ( .A(n10245), .Z(n10248) );
  XNOR U11957 ( .A(n5562), .B(n10245), .Z(n10247) );
  NAND U11958 ( .A(n10250), .B(nreg[342]), .Z(n5562) );
  NAND U11959 ( .A(n6107), .B(nreg[342]), .Z(n10250) );
  XOR U11960 ( .A(n10251), .B(n10252), .Z(n10245) );
  ANDN U11961 ( .A(n10253), .B(n5563), .Z(n10252) );
  XOR U11962 ( .A(n10254), .B(n10255), .Z(n5563) );
  IV U11963 ( .A(n10251), .Z(n10254) );
  XNOR U11964 ( .A(n5564), .B(n10251), .Z(n10253) );
  NAND U11965 ( .A(n10256), .B(nreg[341]), .Z(n5564) );
  NAND U11966 ( .A(n6107), .B(nreg[341]), .Z(n10256) );
  XOR U11967 ( .A(n10257), .B(n10258), .Z(n10251) );
  ANDN U11968 ( .A(n10259), .B(n5565), .Z(n10258) );
  XOR U11969 ( .A(n10260), .B(n10261), .Z(n5565) );
  IV U11970 ( .A(n10257), .Z(n10260) );
  XNOR U11971 ( .A(n5566), .B(n10257), .Z(n10259) );
  NAND U11972 ( .A(n10262), .B(nreg[340]), .Z(n5566) );
  NAND U11973 ( .A(n6107), .B(nreg[340]), .Z(n10262) );
  XOR U11974 ( .A(n10263), .B(n10264), .Z(n10257) );
  ANDN U11975 ( .A(n10265), .B(n5567), .Z(n10264) );
  XOR U11976 ( .A(n10266), .B(n10267), .Z(n5567) );
  IV U11977 ( .A(n10263), .Z(n10266) );
  XNOR U11978 ( .A(n5568), .B(n10263), .Z(n10265) );
  NAND U11979 ( .A(n10268), .B(nreg[339]), .Z(n5568) );
  NAND U11980 ( .A(n6107), .B(nreg[339]), .Z(n10268) );
  XOR U11981 ( .A(n10269), .B(n10270), .Z(n10263) );
  ANDN U11982 ( .A(n10271), .B(n5569), .Z(n10270) );
  XOR U11983 ( .A(n10272), .B(n10273), .Z(n5569) );
  IV U11984 ( .A(n10269), .Z(n10272) );
  XNOR U11985 ( .A(n5570), .B(n10269), .Z(n10271) );
  NAND U11986 ( .A(n10274), .B(nreg[338]), .Z(n5570) );
  NAND U11987 ( .A(n6107), .B(nreg[338]), .Z(n10274) );
  XOR U11988 ( .A(n10275), .B(n10276), .Z(n10269) );
  ANDN U11989 ( .A(n10277), .B(n5571), .Z(n10276) );
  XOR U11990 ( .A(n10278), .B(n10279), .Z(n5571) );
  IV U11991 ( .A(n10275), .Z(n10278) );
  XNOR U11992 ( .A(n5572), .B(n10275), .Z(n10277) );
  NAND U11993 ( .A(n10280), .B(nreg[337]), .Z(n5572) );
  NAND U11994 ( .A(n6107), .B(nreg[337]), .Z(n10280) );
  XOR U11995 ( .A(n10281), .B(n10282), .Z(n10275) );
  ANDN U11996 ( .A(n10283), .B(n5575), .Z(n10282) );
  XOR U11997 ( .A(n10284), .B(n10285), .Z(n5575) );
  IV U11998 ( .A(n10281), .Z(n10284) );
  XNOR U11999 ( .A(n5576), .B(n10281), .Z(n10283) );
  NAND U12000 ( .A(n10286), .B(nreg[336]), .Z(n5576) );
  NAND U12001 ( .A(n6107), .B(nreg[336]), .Z(n10286) );
  XOR U12002 ( .A(n10287), .B(n10288), .Z(n10281) );
  ANDN U12003 ( .A(n10289), .B(n5577), .Z(n10288) );
  XOR U12004 ( .A(n10290), .B(n10291), .Z(n5577) );
  IV U12005 ( .A(n10287), .Z(n10290) );
  XNOR U12006 ( .A(n5578), .B(n10287), .Z(n10289) );
  NAND U12007 ( .A(n10292), .B(nreg[335]), .Z(n5578) );
  NAND U12008 ( .A(n6107), .B(nreg[335]), .Z(n10292) );
  XOR U12009 ( .A(n10293), .B(n10294), .Z(n10287) );
  ANDN U12010 ( .A(n10295), .B(n5579), .Z(n10294) );
  XOR U12011 ( .A(n10296), .B(n10297), .Z(n5579) );
  IV U12012 ( .A(n10293), .Z(n10296) );
  XNOR U12013 ( .A(n5580), .B(n10293), .Z(n10295) );
  NAND U12014 ( .A(n10298), .B(nreg[334]), .Z(n5580) );
  NAND U12015 ( .A(n6107), .B(nreg[334]), .Z(n10298) );
  XOR U12016 ( .A(n10299), .B(n10300), .Z(n10293) );
  ANDN U12017 ( .A(n10301), .B(n5581), .Z(n10300) );
  XOR U12018 ( .A(n10302), .B(n10303), .Z(n5581) );
  IV U12019 ( .A(n10299), .Z(n10302) );
  XNOR U12020 ( .A(n5582), .B(n10299), .Z(n10301) );
  NAND U12021 ( .A(n10304), .B(nreg[333]), .Z(n5582) );
  NAND U12022 ( .A(n6107), .B(nreg[333]), .Z(n10304) );
  XOR U12023 ( .A(n10305), .B(n10306), .Z(n10299) );
  ANDN U12024 ( .A(n10307), .B(n5583), .Z(n10306) );
  XOR U12025 ( .A(n10308), .B(n10309), .Z(n5583) );
  IV U12026 ( .A(n10305), .Z(n10308) );
  XNOR U12027 ( .A(n5584), .B(n10305), .Z(n10307) );
  NAND U12028 ( .A(n10310), .B(nreg[332]), .Z(n5584) );
  NAND U12029 ( .A(n6107), .B(nreg[332]), .Z(n10310) );
  XOR U12030 ( .A(n10311), .B(n10312), .Z(n10305) );
  ANDN U12031 ( .A(n10313), .B(n5585), .Z(n10312) );
  XOR U12032 ( .A(n10314), .B(n10315), .Z(n5585) );
  IV U12033 ( .A(n10311), .Z(n10314) );
  XNOR U12034 ( .A(n5586), .B(n10311), .Z(n10313) );
  NAND U12035 ( .A(n10316), .B(nreg[331]), .Z(n5586) );
  NAND U12036 ( .A(n6107), .B(nreg[331]), .Z(n10316) );
  XOR U12037 ( .A(n10317), .B(n10318), .Z(n10311) );
  ANDN U12038 ( .A(n10319), .B(n5587), .Z(n10318) );
  XOR U12039 ( .A(n10320), .B(n10321), .Z(n5587) );
  IV U12040 ( .A(n10317), .Z(n10320) );
  XNOR U12041 ( .A(n5588), .B(n10317), .Z(n10319) );
  NAND U12042 ( .A(n10322), .B(nreg[330]), .Z(n5588) );
  NAND U12043 ( .A(n6107), .B(nreg[330]), .Z(n10322) );
  XOR U12044 ( .A(n10323), .B(n10324), .Z(n10317) );
  ANDN U12045 ( .A(n10325), .B(n5589), .Z(n10324) );
  XOR U12046 ( .A(n10326), .B(n10327), .Z(n5589) );
  IV U12047 ( .A(n10323), .Z(n10326) );
  XNOR U12048 ( .A(n5590), .B(n10323), .Z(n10325) );
  NAND U12049 ( .A(n10328), .B(nreg[329]), .Z(n5590) );
  NAND U12050 ( .A(n6107), .B(nreg[329]), .Z(n10328) );
  XOR U12051 ( .A(n10329), .B(n10330), .Z(n10323) );
  ANDN U12052 ( .A(n10331), .B(n5591), .Z(n10330) );
  XOR U12053 ( .A(n10332), .B(n10333), .Z(n5591) );
  IV U12054 ( .A(n10329), .Z(n10332) );
  XNOR U12055 ( .A(n5592), .B(n10329), .Z(n10331) );
  NAND U12056 ( .A(n10334), .B(nreg[328]), .Z(n5592) );
  NAND U12057 ( .A(n6107), .B(nreg[328]), .Z(n10334) );
  XOR U12058 ( .A(n10335), .B(n10336), .Z(n10329) );
  ANDN U12059 ( .A(n10337), .B(n5593), .Z(n10336) );
  XOR U12060 ( .A(n10338), .B(n10339), .Z(n5593) );
  IV U12061 ( .A(n10335), .Z(n10338) );
  XNOR U12062 ( .A(n5594), .B(n10335), .Z(n10337) );
  NAND U12063 ( .A(n10340), .B(nreg[327]), .Z(n5594) );
  NAND U12064 ( .A(n6107), .B(nreg[327]), .Z(n10340) );
  XOR U12065 ( .A(n10341), .B(n10342), .Z(n10335) );
  ANDN U12066 ( .A(n10343), .B(n5597), .Z(n10342) );
  XOR U12067 ( .A(n10344), .B(n10345), .Z(n5597) );
  IV U12068 ( .A(n10341), .Z(n10344) );
  XNOR U12069 ( .A(n5598), .B(n10341), .Z(n10343) );
  NAND U12070 ( .A(n10346), .B(nreg[326]), .Z(n5598) );
  NAND U12071 ( .A(n6107), .B(nreg[326]), .Z(n10346) );
  XOR U12072 ( .A(n10347), .B(n10348), .Z(n10341) );
  ANDN U12073 ( .A(n10349), .B(n5599), .Z(n10348) );
  XOR U12074 ( .A(n10350), .B(n10351), .Z(n5599) );
  IV U12075 ( .A(n10347), .Z(n10350) );
  XNOR U12076 ( .A(n5600), .B(n10347), .Z(n10349) );
  NAND U12077 ( .A(n10352), .B(nreg[325]), .Z(n5600) );
  NAND U12078 ( .A(n6107), .B(nreg[325]), .Z(n10352) );
  XOR U12079 ( .A(n10353), .B(n10354), .Z(n10347) );
  ANDN U12080 ( .A(n10355), .B(n5601), .Z(n10354) );
  XOR U12081 ( .A(n10356), .B(n10357), .Z(n5601) );
  IV U12082 ( .A(n10353), .Z(n10356) );
  XNOR U12083 ( .A(n5602), .B(n10353), .Z(n10355) );
  NAND U12084 ( .A(n10358), .B(nreg[324]), .Z(n5602) );
  NAND U12085 ( .A(n6107), .B(nreg[324]), .Z(n10358) );
  XOR U12086 ( .A(n10359), .B(n10360), .Z(n10353) );
  ANDN U12087 ( .A(n10361), .B(n5603), .Z(n10360) );
  XOR U12088 ( .A(n10362), .B(n10363), .Z(n5603) );
  IV U12089 ( .A(n10359), .Z(n10362) );
  XNOR U12090 ( .A(n5604), .B(n10359), .Z(n10361) );
  NAND U12091 ( .A(n10364), .B(nreg[323]), .Z(n5604) );
  NAND U12092 ( .A(n6107), .B(nreg[323]), .Z(n10364) );
  XOR U12093 ( .A(n10365), .B(n10366), .Z(n10359) );
  ANDN U12094 ( .A(n10367), .B(n5605), .Z(n10366) );
  XOR U12095 ( .A(n10368), .B(n10369), .Z(n5605) );
  IV U12096 ( .A(n10365), .Z(n10368) );
  XNOR U12097 ( .A(n5606), .B(n10365), .Z(n10367) );
  NAND U12098 ( .A(n10370), .B(nreg[322]), .Z(n5606) );
  NAND U12099 ( .A(n6107), .B(nreg[322]), .Z(n10370) );
  XOR U12100 ( .A(n10371), .B(n10372), .Z(n10365) );
  ANDN U12101 ( .A(n10373), .B(n5607), .Z(n10372) );
  XOR U12102 ( .A(n10374), .B(n10375), .Z(n5607) );
  IV U12103 ( .A(n10371), .Z(n10374) );
  XNOR U12104 ( .A(n5608), .B(n10371), .Z(n10373) );
  NAND U12105 ( .A(n10376), .B(nreg[321]), .Z(n5608) );
  NAND U12106 ( .A(n6107), .B(nreg[321]), .Z(n10376) );
  XOR U12107 ( .A(n10377), .B(n10378), .Z(n10371) );
  ANDN U12108 ( .A(n10379), .B(n5609), .Z(n10378) );
  XOR U12109 ( .A(n10380), .B(n10381), .Z(n5609) );
  IV U12110 ( .A(n10377), .Z(n10380) );
  XNOR U12111 ( .A(n5610), .B(n10377), .Z(n10379) );
  NAND U12112 ( .A(n10382), .B(nreg[320]), .Z(n5610) );
  NAND U12113 ( .A(n6107), .B(nreg[320]), .Z(n10382) );
  XOR U12114 ( .A(n10383), .B(n10384), .Z(n10377) );
  ANDN U12115 ( .A(n10385), .B(n5611), .Z(n10384) );
  XOR U12116 ( .A(n10386), .B(n10387), .Z(n5611) );
  IV U12117 ( .A(n10383), .Z(n10386) );
  XNOR U12118 ( .A(n5612), .B(n10383), .Z(n10385) );
  NAND U12119 ( .A(n10388), .B(nreg[319]), .Z(n5612) );
  NAND U12120 ( .A(n6107), .B(nreg[319]), .Z(n10388) );
  XOR U12121 ( .A(n10389), .B(n10390), .Z(n10383) );
  ANDN U12122 ( .A(n10391), .B(n5613), .Z(n10390) );
  XOR U12123 ( .A(n10392), .B(n10393), .Z(n5613) );
  IV U12124 ( .A(n10389), .Z(n10392) );
  XNOR U12125 ( .A(n5614), .B(n10389), .Z(n10391) );
  NAND U12126 ( .A(n10394), .B(nreg[318]), .Z(n5614) );
  NAND U12127 ( .A(n6107), .B(nreg[318]), .Z(n10394) );
  XOR U12128 ( .A(n10395), .B(n10396), .Z(n10389) );
  ANDN U12129 ( .A(n10397), .B(n5615), .Z(n10396) );
  XOR U12130 ( .A(n10398), .B(n10399), .Z(n5615) );
  IV U12131 ( .A(n10395), .Z(n10398) );
  XNOR U12132 ( .A(n5616), .B(n10395), .Z(n10397) );
  NAND U12133 ( .A(n10400), .B(nreg[317]), .Z(n5616) );
  NAND U12134 ( .A(n6107), .B(nreg[317]), .Z(n10400) );
  XOR U12135 ( .A(n10401), .B(n10402), .Z(n10395) );
  ANDN U12136 ( .A(n10403), .B(n5619), .Z(n10402) );
  XOR U12137 ( .A(n10404), .B(n10405), .Z(n5619) );
  IV U12138 ( .A(n10401), .Z(n10404) );
  XNOR U12139 ( .A(n5620), .B(n10401), .Z(n10403) );
  NAND U12140 ( .A(n10406), .B(nreg[316]), .Z(n5620) );
  NAND U12141 ( .A(n6107), .B(nreg[316]), .Z(n10406) );
  XOR U12142 ( .A(n10407), .B(n10408), .Z(n10401) );
  ANDN U12143 ( .A(n10409), .B(n5621), .Z(n10408) );
  XOR U12144 ( .A(n10410), .B(n10411), .Z(n5621) );
  IV U12145 ( .A(n10407), .Z(n10410) );
  XNOR U12146 ( .A(n5622), .B(n10407), .Z(n10409) );
  NAND U12147 ( .A(n10412), .B(nreg[315]), .Z(n5622) );
  NAND U12148 ( .A(n6107), .B(nreg[315]), .Z(n10412) );
  XOR U12149 ( .A(n10413), .B(n10414), .Z(n10407) );
  ANDN U12150 ( .A(n10415), .B(n5623), .Z(n10414) );
  XOR U12151 ( .A(n10416), .B(n10417), .Z(n5623) );
  IV U12152 ( .A(n10413), .Z(n10416) );
  XNOR U12153 ( .A(n5624), .B(n10413), .Z(n10415) );
  NAND U12154 ( .A(n10418), .B(nreg[314]), .Z(n5624) );
  NAND U12155 ( .A(n6107), .B(nreg[314]), .Z(n10418) );
  XOR U12156 ( .A(n10419), .B(n10420), .Z(n10413) );
  ANDN U12157 ( .A(n10421), .B(n5625), .Z(n10420) );
  XOR U12158 ( .A(n10422), .B(n10423), .Z(n5625) );
  IV U12159 ( .A(n10419), .Z(n10422) );
  XNOR U12160 ( .A(n5626), .B(n10419), .Z(n10421) );
  NAND U12161 ( .A(n10424), .B(nreg[313]), .Z(n5626) );
  NAND U12162 ( .A(n6107), .B(nreg[313]), .Z(n10424) );
  XOR U12163 ( .A(n10425), .B(n10426), .Z(n10419) );
  ANDN U12164 ( .A(n10427), .B(n5627), .Z(n10426) );
  XOR U12165 ( .A(n10428), .B(n10429), .Z(n5627) );
  IV U12166 ( .A(n10425), .Z(n10428) );
  XNOR U12167 ( .A(n5628), .B(n10425), .Z(n10427) );
  NAND U12168 ( .A(n10430), .B(nreg[312]), .Z(n5628) );
  NAND U12169 ( .A(n6107), .B(nreg[312]), .Z(n10430) );
  XOR U12170 ( .A(n10431), .B(n10432), .Z(n10425) );
  ANDN U12171 ( .A(n10433), .B(n5629), .Z(n10432) );
  XOR U12172 ( .A(n10434), .B(n10435), .Z(n5629) );
  IV U12173 ( .A(n10431), .Z(n10434) );
  XNOR U12174 ( .A(n5630), .B(n10431), .Z(n10433) );
  NAND U12175 ( .A(n10436), .B(nreg[311]), .Z(n5630) );
  NAND U12176 ( .A(n6107), .B(nreg[311]), .Z(n10436) );
  XOR U12177 ( .A(n10437), .B(n10438), .Z(n10431) );
  ANDN U12178 ( .A(n10439), .B(n5631), .Z(n10438) );
  XOR U12179 ( .A(n10440), .B(n10441), .Z(n5631) );
  IV U12180 ( .A(n10437), .Z(n10440) );
  XNOR U12181 ( .A(n5632), .B(n10437), .Z(n10439) );
  NAND U12182 ( .A(n10442), .B(nreg[310]), .Z(n5632) );
  NAND U12183 ( .A(n6107), .B(nreg[310]), .Z(n10442) );
  XOR U12184 ( .A(n10443), .B(n10444), .Z(n10437) );
  ANDN U12185 ( .A(n10445), .B(n5633), .Z(n10444) );
  XOR U12186 ( .A(n10446), .B(n10447), .Z(n5633) );
  IV U12187 ( .A(n10443), .Z(n10446) );
  XNOR U12188 ( .A(n5634), .B(n10443), .Z(n10445) );
  NAND U12189 ( .A(n10448), .B(nreg[309]), .Z(n5634) );
  NAND U12190 ( .A(n6107), .B(nreg[309]), .Z(n10448) );
  XOR U12191 ( .A(n10449), .B(n10450), .Z(n10443) );
  ANDN U12192 ( .A(n10451), .B(n5635), .Z(n10450) );
  XOR U12193 ( .A(n10452), .B(n10453), .Z(n5635) );
  IV U12194 ( .A(n10449), .Z(n10452) );
  XNOR U12195 ( .A(n5636), .B(n10449), .Z(n10451) );
  NAND U12196 ( .A(n10454), .B(nreg[308]), .Z(n5636) );
  NAND U12197 ( .A(n6107), .B(nreg[308]), .Z(n10454) );
  XOR U12198 ( .A(n10455), .B(n10456), .Z(n10449) );
  ANDN U12199 ( .A(n10457), .B(n5637), .Z(n10456) );
  XOR U12200 ( .A(n10458), .B(n10459), .Z(n5637) );
  IV U12201 ( .A(n10455), .Z(n10458) );
  XNOR U12202 ( .A(n5638), .B(n10455), .Z(n10457) );
  NAND U12203 ( .A(n10460), .B(nreg[307]), .Z(n5638) );
  NAND U12204 ( .A(n6107), .B(nreg[307]), .Z(n10460) );
  XOR U12205 ( .A(n10461), .B(n10462), .Z(n10455) );
  ANDN U12206 ( .A(n10463), .B(n5641), .Z(n10462) );
  XOR U12207 ( .A(n10464), .B(n10465), .Z(n5641) );
  IV U12208 ( .A(n10461), .Z(n10464) );
  XNOR U12209 ( .A(n5642), .B(n10461), .Z(n10463) );
  NAND U12210 ( .A(n10466), .B(nreg[306]), .Z(n5642) );
  NAND U12211 ( .A(n6107), .B(nreg[306]), .Z(n10466) );
  XOR U12212 ( .A(n10467), .B(n10468), .Z(n10461) );
  ANDN U12213 ( .A(n10469), .B(n5643), .Z(n10468) );
  XOR U12214 ( .A(n10470), .B(n10471), .Z(n5643) );
  IV U12215 ( .A(n10467), .Z(n10470) );
  XNOR U12216 ( .A(n5644), .B(n10467), .Z(n10469) );
  NAND U12217 ( .A(n10472), .B(nreg[305]), .Z(n5644) );
  NAND U12218 ( .A(n6107), .B(nreg[305]), .Z(n10472) );
  XOR U12219 ( .A(n10473), .B(n10474), .Z(n10467) );
  ANDN U12220 ( .A(n10475), .B(n5645), .Z(n10474) );
  XOR U12221 ( .A(n10476), .B(n10477), .Z(n5645) );
  IV U12222 ( .A(n10473), .Z(n10476) );
  XNOR U12223 ( .A(n5646), .B(n10473), .Z(n10475) );
  NAND U12224 ( .A(n10478), .B(nreg[304]), .Z(n5646) );
  NAND U12225 ( .A(n6107), .B(nreg[304]), .Z(n10478) );
  XOR U12226 ( .A(n10479), .B(n10480), .Z(n10473) );
  ANDN U12227 ( .A(n10481), .B(n5647), .Z(n10480) );
  XOR U12228 ( .A(n10482), .B(n10483), .Z(n5647) );
  IV U12229 ( .A(n10479), .Z(n10482) );
  XNOR U12230 ( .A(n5648), .B(n10479), .Z(n10481) );
  NAND U12231 ( .A(n10484), .B(nreg[303]), .Z(n5648) );
  NAND U12232 ( .A(n6107), .B(nreg[303]), .Z(n10484) );
  XOR U12233 ( .A(n10485), .B(n10486), .Z(n10479) );
  ANDN U12234 ( .A(n10487), .B(n5649), .Z(n10486) );
  XOR U12235 ( .A(n10488), .B(n10489), .Z(n5649) );
  IV U12236 ( .A(n10485), .Z(n10488) );
  XNOR U12237 ( .A(n5650), .B(n10485), .Z(n10487) );
  NAND U12238 ( .A(n10490), .B(nreg[302]), .Z(n5650) );
  NAND U12239 ( .A(n6107), .B(nreg[302]), .Z(n10490) );
  XOR U12240 ( .A(n10491), .B(n10492), .Z(n10485) );
  ANDN U12241 ( .A(n10493), .B(n5651), .Z(n10492) );
  XOR U12242 ( .A(n10494), .B(n10495), .Z(n5651) );
  IV U12243 ( .A(n10491), .Z(n10494) );
  XNOR U12244 ( .A(n5652), .B(n10491), .Z(n10493) );
  NAND U12245 ( .A(n10496), .B(nreg[301]), .Z(n5652) );
  NAND U12246 ( .A(n6107), .B(nreg[301]), .Z(n10496) );
  XOR U12247 ( .A(n10497), .B(n10498), .Z(n10491) );
  ANDN U12248 ( .A(n10499), .B(n5653), .Z(n10498) );
  XOR U12249 ( .A(n10500), .B(n10501), .Z(n5653) );
  IV U12250 ( .A(n10497), .Z(n10500) );
  XNOR U12251 ( .A(n5654), .B(n10497), .Z(n10499) );
  NAND U12252 ( .A(n10502), .B(nreg[300]), .Z(n5654) );
  NAND U12253 ( .A(n6107), .B(nreg[300]), .Z(n10502) );
  XOR U12254 ( .A(n10503), .B(n10504), .Z(n10497) );
  ANDN U12255 ( .A(n10505), .B(n5655), .Z(n10504) );
  XOR U12256 ( .A(n10506), .B(n10507), .Z(n5655) );
  IV U12257 ( .A(n10503), .Z(n10506) );
  XNOR U12258 ( .A(n5656), .B(n10503), .Z(n10505) );
  NAND U12259 ( .A(n10508), .B(nreg[299]), .Z(n5656) );
  NAND U12260 ( .A(n6107), .B(nreg[299]), .Z(n10508) );
  XOR U12261 ( .A(n10509), .B(n10510), .Z(n10503) );
  ANDN U12262 ( .A(n10511), .B(n5657), .Z(n10510) );
  XOR U12263 ( .A(n10512), .B(n10513), .Z(n5657) );
  IV U12264 ( .A(n10509), .Z(n10512) );
  XNOR U12265 ( .A(n5658), .B(n10509), .Z(n10511) );
  NAND U12266 ( .A(n10514), .B(nreg[298]), .Z(n5658) );
  NAND U12267 ( .A(n6107), .B(nreg[298]), .Z(n10514) );
  XOR U12268 ( .A(n10515), .B(n10516), .Z(n10509) );
  ANDN U12269 ( .A(n10517), .B(n5659), .Z(n10516) );
  XOR U12270 ( .A(n10518), .B(n10519), .Z(n5659) );
  IV U12271 ( .A(n10515), .Z(n10518) );
  XNOR U12272 ( .A(n5660), .B(n10515), .Z(n10517) );
  NAND U12273 ( .A(n10520), .B(nreg[297]), .Z(n5660) );
  NAND U12274 ( .A(n6107), .B(nreg[297]), .Z(n10520) );
  XOR U12275 ( .A(n10521), .B(n10522), .Z(n10515) );
  ANDN U12276 ( .A(n10523), .B(n5665), .Z(n10522) );
  XOR U12277 ( .A(n10524), .B(n10525), .Z(n5665) );
  IV U12278 ( .A(n10521), .Z(n10524) );
  XNOR U12279 ( .A(n5666), .B(n10521), .Z(n10523) );
  NAND U12280 ( .A(n10526), .B(nreg[296]), .Z(n5666) );
  NAND U12281 ( .A(n6107), .B(nreg[296]), .Z(n10526) );
  XOR U12282 ( .A(n10527), .B(n10528), .Z(n10521) );
  ANDN U12283 ( .A(n10529), .B(n5667), .Z(n10528) );
  XOR U12284 ( .A(n10530), .B(n10531), .Z(n5667) );
  IV U12285 ( .A(n10527), .Z(n10530) );
  XNOR U12286 ( .A(n5668), .B(n10527), .Z(n10529) );
  NAND U12287 ( .A(n10532), .B(nreg[295]), .Z(n5668) );
  NAND U12288 ( .A(n6107), .B(nreg[295]), .Z(n10532) );
  XOR U12289 ( .A(n10533), .B(n10534), .Z(n10527) );
  ANDN U12290 ( .A(n10535), .B(n5669), .Z(n10534) );
  XOR U12291 ( .A(n10536), .B(n10537), .Z(n5669) );
  IV U12292 ( .A(n10533), .Z(n10536) );
  XNOR U12293 ( .A(n5670), .B(n10533), .Z(n10535) );
  NAND U12294 ( .A(n10538), .B(nreg[294]), .Z(n5670) );
  NAND U12295 ( .A(n6107), .B(nreg[294]), .Z(n10538) );
  XOR U12296 ( .A(n10539), .B(n10540), .Z(n10533) );
  ANDN U12297 ( .A(n10541), .B(n5671), .Z(n10540) );
  XOR U12298 ( .A(n10542), .B(n10543), .Z(n5671) );
  IV U12299 ( .A(n10539), .Z(n10542) );
  XNOR U12300 ( .A(n5672), .B(n10539), .Z(n10541) );
  NAND U12301 ( .A(n10544), .B(nreg[293]), .Z(n5672) );
  NAND U12302 ( .A(n6107), .B(nreg[293]), .Z(n10544) );
  XOR U12303 ( .A(n10545), .B(n10546), .Z(n10539) );
  ANDN U12304 ( .A(n10547), .B(n5673), .Z(n10546) );
  XOR U12305 ( .A(n10548), .B(n10549), .Z(n5673) );
  IV U12306 ( .A(n10545), .Z(n10548) );
  XNOR U12307 ( .A(n5674), .B(n10545), .Z(n10547) );
  NAND U12308 ( .A(n10550), .B(nreg[292]), .Z(n5674) );
  NAND U12309 ( .A(n6107), .B(nreg[292]), .Z(n10550) );
  XOR U12310 ( .A(n10551), .B(n10552), .Z(n10545) );
  ANDN U12311 ( .A(n10553), .B(n5675), .Z(n10552) );
  XOR U12312 ( .A(n10554), .B(n10555), .Z(n5675) );
  IV U12313 ( .A(n10551), .Z(n10554) );
  XNOR U12314 ( .A(n5676), .B(n10551), .Z(n10553) );
  NAND U12315 ( .A(n10556), .B(nreg[291]), .Z(n5676) );
  NAND U12316 ( .A(n6107), .B(nreg[291]), .Z(n10556) );
  XOR U12317 ( .A(n10557), .B(n10558), .Z(n10551) );
  ANDN U12318 ( .A(n10559), .B(n5677), .Z(n10558) );
  XOR U12319 ( .A(n10560), .B(n10561), .Z(n5677) );
  IV U12320 ( .A(n10557), .Z(n10560) );
  XNOR U12321 ( .A(n5678), .B(n10557), .Z(n10559) );
  NAND U12322 ( .A(n10562), .B(nreg[290]), .Z(n5678) );
  NAND U12323 ( .A(n6107), .B(nreg[290]), .Z(n10562) );
  XOR U12324 ( .A(n10563), .B(n10564), .Z(n10557) );
  ANDN U12325 ( .A(n10565), .B(n5679), .Z(n10564) );
  XOR U12326 ( .A(n10566), .B(n10567), .Z(n5679) );
  IV U12327 ( .A(n10563), .Z(n10566) );
  XNOR U12328 ( .A(n5680), .B(n10563), .Z(n10565) );
  NAND U12329 ( .A(n10568), .B(nreg[289]), .Z(n5680) );
  NAND U12330 ( .A(n6107), .B(nreg[289]), .Z(n10568) );
  XOR U12331 ( .A(n10569), .B(n10570), .Z(n10563) );
  ANDN U12332 ( .A(n10571), .B(n5681), .Z(n10570) );
  XOR U12333 ( .A(n10572), .B(n10573), .Z(n5681) );
  IV U12334 ( .A(n10569), .Z(n10572) );
  XNOR U12335 ( .A(n5682), .B(n10569), .Z(n10571) );
  NAND U12336 ( .A(n10574), .B(nreg[288]), .Z(n5682) );
  NAND U12337 ( .A(n6107), .B(nreg[288]), .Z(n10574) );
  XOR U12338 ( .A(n10575), .B(n10576), .Z(n10569) );
  ANDN U12339 ( .A(n10577), .B(n5683), .Z(n10576) );
  XOR U12340 ( .A(n10578), .B(n10579), .Z(n5683) );
  IV U12341 ( .A(n10575), .Z(n10578) );
  XNOR U12342 ( .A(n5684), .B(n10575), .Z(n10577) );
  NAND U12343 ( .A(n10580), .B(nreg[287]), .Z(n5684) );
  NAND U12344 ( .A(n6107), .B(nreg[287]), .Z(n10580) );
  XOR U12345 ( .A(n10581), .B(n10582), .Z(n10575) );
  ANDN U12346 ( .A(n10583), .B(n5687), .Z(n10582) );
  XOR U12347 ( .A(n10584), .B(n10585), .Z(n5687) );
  IV U12348 ( .A(n10581), .Z(n10584) );
  XNOR U12349 ( .A(n5688), .B(n10581), .Z(n10583) );
  NAND U12350 ( .A(n10586), .B(nreg[286]), .Z(n5688) );
  NAND U12351 ( .A(n6107), .B(nreg[286]), .Z(n10586) );
  XOR U12352 ( .A(n10587), .B(n10588), .Z(n10581) );
  ANDN U12353 ( .A(n10589), .B(n5689), .Z(n10588) );
  XOR U12354 ( .A(n10590), .B(n10591), .Z(n5689) );
  IV U12355 ( .A(n10587), .Z(n10590) );
  XNOR U12356 ( .A(n5690), .B(n10587), .Z(n10589) );
  NAND U12357 ( .A(n10592), .B(nreg[285]), .Z(n5690) );
  NAND U12358 ( .A(n6107), .B(nreg[285]), .Z(n10592) );
  XOR U12359 ( .A(n10593), .B(n10594), .Z(n10587) );
  ANDN U12360 ( .A(n10595), .B(n5691), .Z(n10594) );
  XOR U12361 ( .A(n10596), .B(n10597), .Z(n5691) );
  IV U12362 ( .A(n10593), .Z(n10596) );
  XNOR U12363 ( .A(n5692), .B(n10593), .Z(n10595) );
  NAND U12364 ( .A(n10598), .B(nreg[284]), .Z(n5692) );
  NAND U12365 ( .A(n6107), .B(nreg[284]), .Z(n10598) );
  XOR U12366 ( .A(n10599), .B(n10600), .Z(n10593) );
  ANDN U12367 ( .A(n10601), .B(n5693), .Z(n10600) );
  XOR U12368 ( .A(n10602), .B(n10603), .Z(n5693) );
  IV U12369 ( .A(n10599), .Z(n10602) );
  XNOR U12370 ( .A(n5694), .B(n10599), .Z(n10601) );
  NAND U12371 ( .A(n10604), .B(nreg[283]), .Z(n5694) );
  NAND U12372 ( .A(n6107), .B(nreg[283]), .Z(n10604) );
  XOR U12373 ( .A(n10605), .B(n10606), .Z(n10599) );
  ANDN U12374 ( .A(n10607), .B(n5695), .Z(n10606) );
  XOR U12375 ( .A(n10608), .B(n10609), .Z(n5695) );
  IV U12376 ( .A(n10605), .Z(n10608) );
  XNOR U12377 ( .A(n5696), .B(n10605), .Z(n10607) );
  NAND U12378 ( .A(n10610), .B(nreg[282]), .Z(n5696) );
  NAND U12379 ( .A(n6107), .B(nreg[282]), .Z(n10610) );
  XOR U12380 ( .A(n10611), .B(n10612), .Z(n10605) );
  ANDN U12381 ( .A(n10613), .B(n5697), .Z(n10612) );
  XOR U12382 ( .A(n10614), .B(n10615), .Z(n5697) );
  IV U12383 ( .A(n10611), .Z(n10614) );
  XNOR U12384 ( .A(n5698), .B(n10611), .Z(n10613) );
  NAND U12385 ( .A(n10616), .B(nreg[281]), .Z(n5698) );
  NAND U12386 ( .A(n6107), .B(nreg[281]), .Z(n10616) );
  XOR U12387 ( .A(n10617), .B(n10618), .Z(n10611) );
  ANDN U12388 ( .A(n10619), .B(n5699), .Z(n10618) );
  XOR U12389 ( .A(n10620), .B(n10621), .Z(n5699) );
  IV U12390 ( .A(n10617), .Z(n10620) );
  XNOR U12391 ( .A(n5700), .B(n10617), .Z(n10619) );
  NAND U12392 ( .A(n10622), .B(nreg[280]), .Z(n5700) );
  NAND U12393 ( .A(n6107), .B(nreg[280]), .Z(n10622) );
  XOR U12394 ( .A(n10623), .B(n10624), .Z(n10617) );
  ANDN U12395 ( .A(n10625), .B(n5701), .Z(n10624) );
  XOR U12396 ( .A(n10626), .B(n10627), .Z(n5701) );
  IV U12397 ( .A(n10623), .Z(n10626) );
  XNOR U12398 ( .A(n5702), .B(n10623), .Z(n10625) );
  NAND U12399 ( .A(n10628), .B(nreg[279]), .Z(n5702) );
  NAND U12400 ( .A(n6107), .B(nreg[279]), .Z(n10628) );
  XOR U12401 ( .A(n10629), .B(n10630), .Z(n10623) );
  ANDN U12402 ( .A(n10631), .B(n5703), .Z(n10630) );
  XOR U12403 ( .A(n10632), .B(n10633), .Z(n5703) );
  IV U12404 ( .A(n10629), .Z(n10632) );
  XNOR U12405 ( .A(n5704), .B(n10629), .Z(n10631) );
  NAND U12406 ( .A(n10634), .B(nreg[278]), .Z(n5704) );
  NAND U12407 ( .A(n6107), .B(nreg[278]), .Z(n10634) );
  XOR U12408 ( .A(n10635), .B(n10636), .Z(n10629) );
  ANDN U12409 ( .A(n10637), .B(n5705), .Z(n10636) );
  XOR U12410 ( .A(n10638), .B(n10639), .Z(n5705) );
  IV U12411 ( .A(n10635), .Z(n10638) );
  XNOR U12412 ( .A(n5706), .B(n10635), .Z(n10637) );
  NAND U12413 ( .A(n10640), .B(nreg[277]), .Z(n5706) );
  NAND U12414 ( .A(n6107), .B(nreg[277]), .Z(n10640) );
  XOR U12415 ( .A(n10641), .B(n10642), .Z(n10635) );
  ANDN U12416 ( .A(n10643), .B(n5709), .Z(n10642) );
  XOR U12417 ( .A(n10644), .B(n10645), .Z(n5709) );
  IV U12418 ( .A(n10641), .Z(n10644) );
  XNOR U12419 ( .A(n5710), .B(n10641), .Z(n10643) );
  NAND U12420 ( .A(n10646), .B(nreg[276]), .Z(n5710) );
  NAND U12421 ( .A(n6107), .B(nreg[276]), .Z(n10646) );
  XOR U12422 ( .A(n10647), .B(n10648), .Z(n10641) );
  ANDN U12423 ( .A(n10649), .B(n5711), .Z(n10648) );
  XOR U12424 ( .A(n10650), .B(n10651), .Z(n5711) );
  IV U12425 ( .A(n10647), .Z(n10650) );
  XNOR U12426 ( .A(n5712), .B(n10647), .Z(n10649) );
  NAND U12427 ( .A(n10652), .B(nreg[275]), .Z(n5712) );
  NAND U12428 ( .A(n6107), .B(nreg[275]), .Z(n10652) );
  XOR U12429 ( .A(n10653), .B(n10654), .Z(n10647) );
  ANDN U12430 ( .A(n10655), .B(n5713), .Z(n10654) );
  XOR U12431 ( .A(n10656), .B(n10657), .Z(n5713) );
  IV U12432 ( .A(n10653), .Z(n10656) );
  XNOR U12433 ( .A(n5714), .B(n10653), .Z(n10655) );
  NAND U12434 ( .A(n10658), .B(nreg[274]), .Z(n5714) );
  NAND U12435 ( .A(n6107), .B(nreg[274]), .Z(n10658) );
  XOR U12436 ( .A(n10659), .B(n10660), .Z(n10653) );
  ANDN U12437 ( .A(n10661), .B(n5715), .Z(n10660) );
  XOR U12438 ( .A(n10662), .B(n10663), .Z(n5715) );
  IV U12439 ( .A(n10659), .Z(n10662) );
  XNOR U12440 ( .A(n5716), .B(n10659), .Z(n10661) );
  NAND U12441 ( .A(n10664), .B(nreg[273]), .Z(n5716) );
  NAND U12442 ( .A(n6107), .B(nreg[273]), .Z(n10664) );
  XOR U12443 ( .A(n10665), .B(n10666), .Z(n10659) );
  ANDN U12444 ( .A(n10667), .B(n5717), .Z(n10666) );
  XOR U12445 ( .A(n10668), .B(n10669), .Z(n5717) );
  IV U12446 ( .A(n10665), .Z(n10668) );
  XNOR U12447 ( .A(n5718), .B(n10665), .Z(n10667) );
  NAND U12448 ( .A(n10670), .B(nreg[272]), .Z(n5718) );
  NAND U12449 ( .A(n6107), .B(nreg[272]), .Z(n10670) );
  XOR U12450 ( .A(n10671), .B(n10672), .Z(n10665) );
  ANDN U12451 ( .A(n10673), .B(n5719), .Z(n10672) );
  XOR U12452 ( .A(n10674), .B(n10675), .Z(n5719) );
  IV U12453 ( .A(n10671), .Z(n10674) );
  XNOR U12454 ( .A(n5720), .B(n10671), .Z(n10673) );
  NAND U12455 ( .A(n10676), .B(nreg[271]), .Z(n5720) );
  NAND U12456 ( .A(n6107), .B(nreg[271]), .Z(n10676) );
  XOR U12457 ( .A(n10677), .B(n10678), .Z(n10671) );
  ANDN U12458 ( .A(n10679), .B(n5721), .Z(n10678) );
  XOR U12459 ( .A(n10680), .B(n10681), .Z(n5721) );
  IV U12460 ( .A(n10677), .Z(n10680) );
  XNOR U12461 ( .A(n5722), .B(n10677), .Z(n10679) );
  NAND U12462 ( .A(n10682), .B(nreg[270]), .Z(n5722) );
  NAND U12463 ( .A(n6107), .B(nreg[270]), .Z(n10682) );
  XOR U12464 ( .A(n10683), .B(n10684), .Z(n10677) );
  ANDN U12465 ( .A(n10685), .B(n5723), .Z(n10684) );
  XOR U12466 ( .A(n10686), .B(n10687), .Z(n5723) );
  IV U12467 ( .A(n10683), .Z(n10686) );
  XNOR U12468 ( .A(n5724), .B(n10683), .Z(n10685) );
  NAND U12469 ( .A(n10688), .B(nreg[269]), .Z(n5724) );
  NAND U12470 ( .A(n6107), .B(nreg[269]), .Z(n10688) );
  XOR U12471 ( .A(n10689), .B(n10690), .Z(n10683) );
  ANDN U12472 ( .A(n10691), .B(n5725), .Z(n10690) );
  XOR U12473 ( .A(n10692), .B(n10693), .Z(n5725) );
  IV U12474 ( .A(n10689), .Z(n10692) );
  XNOR U12475 ( .A(n5726), .B(n10689), .Z(n10691) );
  NAND U12476 ( .A(n10694), .B(nreg[268]), .Z(n5726) );
  NAND U12477 ( .A(n6107), .B(nreg[268]), .Z(n10694) );
  XOR U12478 ( .A(n10695), .B(n10696), .Z(n10689) );
  ANDN U12479 ( .A(n10697), .B(n5727), .Z(n10696) );
  XOR U12480 ( .A(n10698), .B(n10699), .Z(n5727) );
  IV U12481 ( .A(n10695), .Z(n10698) );
  XNOR U12482 ( .A(n5728), .B(n10695), .Z(n10697) );
  NAND U12483 ( .A(n10700), .B(nreg[267]), .Z(n5728) );
  NAND U12484 ( .A(n6107), .B(nreg[267]), .Z(n10700) );
  XOR U12485 ( .A(n10701), .B(n10702), .Z(n10695) );
  ANDN U12486 ( .A(n10703), .B(n5731), .Z(n10702) );
  XOR U12487 ( .A(n10704), .B(n10705), .Z(n5731) );
  IV U12488 ( .A(n10701), .Z(n10704) );
  XNOR U12489 ( .A(n5732), .B(n10701), .Z(n10703) );
  NAND U12490 ( .A(n10706), .B(nreg[266]), .Z(n5732) );
  NAND U12491 ( .A(n6107), .B(nreg[266]), .Z(n10706) );
  XOR U12492 ( .A(n10707), .B(n10708), .Z(n10701) );
  ANDN U12493 ( .A(n10709), .B(n5733), .Z(n10708) );
  XOR U12494 ( .A(n10710), .B(n10711), .Z(n5733) );
  IV U12495 ( .A(n10707), .Z(n10710) );
  XNOR U12496 ( .A(n5734), .B(n10707), .Z(n10709) );
  NAND U12497 ( .A(n10712), .B(nreg[265]), .Z(n5734) );
  NAND U12498 ( .A(n6107), .B(nreg[265]), .Z(n10712) );
  XOR U12499 ( .A(n10713), .B(n10714), .Z(n10707) );
  ANDN U12500 ( .A(n10715), .B(n5735), .Z(n10714) );
  XOR U12501 ( .A(n10716), .B(n10717), .Z(n5735) );
  IV U12502 ( .A(n10713), .Z(n10716) );
  XNOR U12503 ( .A(n5736), .B(n10713), .Z(n10715) );
  NAND U12504 ( .A(n10718), .B(nreg[264]), .Z(n5736) );
  NAND U12505 ( .A(n6107), .B(nreg[264]), .Z(n10718) );
  XOR U12506 ( .A(n10719), .B(n10720), .Z(n10713) );
  ANDN U12507 ( .A(n10721), .B(n5737), .Z(n10720) );
  XOR U12508 ( .A(n10722), .B(n10723), .Z(n5737) );
  IV U12509 ( .A(n10719), .Z(n10722) );
  XNOR U12510 ( .A(n5738), .B(n10719), .Z(n10721) );
  NAND U12511 ( .A(n10724), .B(nreg[263]), .Z(n5738) );
  NAND U12512 ( .A(n6107), .B(nreg[263]), .Z(n10724) );
  XOR U12513 ( .A(n10725), .B(n10726), .Z(n10719) );
  ANDN U12514 ( .A(n10727), .B(n5739), .Z(n10726) );
  XOR U12515 ( .A(n10728), .B(n10729), .Z(n5739) );
  IV U12516 ( .A(n10725), .Z(n10728) );
  XNOR U12517 ( .A(n5740), .B(n10725), .Z(n10727) );
  NAND U12518 ( .A(n10730), .B(nreg[262]), .Z(n5740) );
  NAND U12519 ( .A(n6107), .B(nreg[262]), .Z(n10730) );
  XOR U12520 ( .A(n10731), .B(n10732), .Z(n10725) );
  ANDN U12521 ( .A(n10733), .B(n5741), .Z(n10732) );
  XOR U12522 ( .A(n10734), .B(n10735), .Z(n5741) );
  IV U12523 ( .A(n10731), .Z(n10734) );
  XNOR U12524 ( .A(n5742), .B(n10731), .Z(n10733) );
  NAND U12525 ( .A(n10736), .B(nreg[261]), .Z(n5742) );
  NAND U12526 ( .A(n6107), .B(nreg[261]), .Z(n10736) );
  XOR U12527 ( .A(n10737), .B(n10738), .Z(n10731) );
  ANDN U12528 ( .A(n10739), .B(n5743), .Z(n10738) );
  XOR U12529 ( .A(n10740), .B(n10741), .Z(n5743) );
  IV U12530 ( .A(n10737), .Z(n10740) );
  XNOR U12531 ( .A(n5744), .B(n10737), .Z(n10739) );
  NAND U12532 ( .A(n10742), .B(nreg[260]), .Z(n5744) );
  NAND U12533 ( .A(n6107), .B(nreg[260]), .Z(n10742) );
  XOR U12534 ( .A(n10743), .B(n10744), .Z(n10737) );
  ANDN U12535 ( .A(n10745), .B(n5745), .Z(n10744) );
  XOR U12536 ( .A(n10746), .B(n10747), .Z(n5745) );
  IV U12537 ( .A(n10743), .Z(n10746) );
  XNOR U12538 ( .A(n5746), .B(n10743), .Z(n10745) );
  NAND U12539 ( .A(n10748), .B(nreg[259]), .Z(n5746) );
  NAND U12540 ( .A(n6107), .B(nreg[259]), .Z(n10748) );
  XOR U12541 ( .A(n10749), .B(n10750), .Z(n10743) );
  ANDN U12542 ( .A(n10751), .B(n5747), .Z(n10750) );
  XOR U12543 ( .A(n10752), .B(n10753), .Z(n5747) );
  IV U12544 ( .A(n10749), .Z(n10752) );
  XNOR U12545 ( .A(n5748), .B(n10749), .Z(n10751) );
  NAND U12546 ( .A(n10754), .B(nreg[258]), .Z(n5748) );
  NAND U12547 ( .A(n6107), .B(nreg[258]), .Z(n10754) );
  XOR U12548 ( .A(n10755), .B(n10756), .Z(n10749) );
  ANDN U12549 ( .A(n10757), .B(n5749), .Z(n10756) );
  XOR U12550 ( .A(n10758), .B(n10759), .Z(n5749) );
  IV U12551 ( .A(n10755), .Z(n10758) );
  XNOR U12552 ( .A(n5750), .B(n10755), .Z(n10757) );
  NAND U12553 ( .A(n10760), .B(nreg[257]), .Z(n5750) );
  NAND U12554 ( .A(n6107), .B(nreg[257]), .Z(n10760) );
  XOR U12555 ( .A(n10761), .B(n10762), .Z(n10755) );
  ANDN U12556 ( .A(n10763), .B(n5753), .Z(n10762) );
  XOR U12557 ( .A(n10764), .B(n10765), .Z(n5753) );
  IV U12558 ( .A(n10761), .Z(n10764) );
  XNOR U12559 ( .A(n5754), .B(n10761), .Z(n10763) );
  NAND U12560 ( .A(n10766), .B(nreg[256]), .Z(n5754) );
  NAND U12561 ( .A(n6107), .B(nreg[256]), .Z(n10766) );
  XOR U12562 ( .A(n10767), .B(n10768), .Z(n10761) );
  ANDN U12563 ( .A(n10769), .B(n5755), .Z(n10768) );
  XOR U12564 ( .A(n10770), .B(n10771), .Z(n5755) );
  IV U12565 ( .A(n10767), .Z(n10770) );
  XNOR U12566 ( .A(n5756), .B(n10767), .Z(n10769) );
  NAND U12567 ( .A(n10772), .B(nreg[255]), .Z(n5756) );
  NAND U12568 ( .A(n6107), .B(nreg[255]), .Z(n10772) );
  XOR U12569 ( .A(n10773), .B(n10774), .Z(n10767) );
  ANDN U12570 ( .A(n10775), .B(n5757), .Z(n10774) );
  XOR U12571 ( .A(n10776), .B(n10777), .Z(n5757) );
  IV U12572 ( .A(n10773), .Z(n10776) );
  XNOR U12573 ( .A(n5758), .B(n10773), .Z(n10775) );
  NAND U12574 ( .A(n10778), .B(nreg[254]), .Z(n5758) );
  NAND U12575 ( .A(n6107), .B(nreg[254]), .Z(n10778) );
  XOR U12576 ( .A(n10779), .B(n10780), .Z(n10773) );
  ANDN U12577 ( .A(n10781), .B(n5759), .Z(n10780) );
  XOR U12578 ( .A(n10782), .B(n10783), .Z(n5759) );
  IV U12579 ( .A(n10779), .Z(n10782) );
  XNOR U12580 ( .A(n5760), .B(n10779), .Z(n10781) );
  NAND U12581 ( .A(n10784), .B(nreg[253]), .Z(n5760) );
  NAND U12582 ( .A(n6107), .B(nreg[253]), .Z(n10784) );
  XOR U12583 ( .A(n10785), .B(n10786), .Z(n10779) );
  ANDN U12584 ( .A(n10787), .B(n5761), .Z(n10786) );
  XOR U12585 ( .A(n10788), .B(n10789), .Z(n5761) );
  IV U12586 ( .A(n10785), .Z(n10788) );
  XNOR U12587 ( .A(n5762), .B(n10785), .Z(n10787) );
  NAND U12588 ( .A(n10790), .B(nreg[252]), .Z(n5762) );
  NAND U12589 ( .A(n6107), .B(nreg[252]), .Z(n10790) );
  XOR U12590 ( .A(n10791), .B(n10792), .Z(n10785) );
  ANDN U12591 ( .A(n10793), .B(n5763), .Z(n10792) );
  XOR U12592 ( .A(n10794), .B(n10795), .Z(n5763) );
  IV U12593 ( .A(n10791), .Z(n10794) );
  XNOR U12594 ( .A(n5764), .B(n10791), .Z(n10793) );
  NAND U12595 ( .A(n10796), .B(nreg[251]), .Z(n5764) );
  NAND U12596 ( .A(n6107), .B(nreg[251]), .Z(n10796) );
  XOR U12597 ( .A(n10797), .B(n10798), .Z(n10791) );
  ANDN U12598 ( .A(n10799), .B(n5765), .Z(n10798) );
  XOR U12599 ( .A(n10800), .B(n10801), .Z(n5765) );
  IV U12600 ( .A(n10797), .Z(n10800) );
  XNOR U12601 ( .A(n5766), .B(n10797), .Z(n10799) );
  NAND U12602 ( .A(n10802), .B(nreg[250]), .Z(n5766) );
  NAND U12603 ( .A(n6107), .B(nreg[250]), .Z(n10802) );
  XOR U12604 ( .A(n10803), .B(n10804), .Z(n10797) );
  ANDN U12605 ( .A(n10805), .B(n5767), .Z(n10804) );
  XOR U12606 ( .A(n10806), .B(n10807), .Z(n5767) );
  IV U12607 ( .A(n10803), .Z(n10806) );
  XNOR U12608 ( .A(n5768), .B(n10803), .Z(n10805) );
  NAND U12609 ( .A(n10808), .B(nreg[249]), .Z(n5768) );
  NAND U12610 ( .A(n6107), .B(nreg[249]), .Z(n10808) );
  XOR U12611 ( .A(n10809), .B(n10810), .Z(n10803) );
  ANDN U12612 ( .A(n10811), .B(n5769), .Z(n10810) );
  XOR U12613 ( .A(n10812), .B(n10813), .Z(n5769) );
  IV U12614 ( .A(n10809), .Z(n10812) );
  XNOR U12615 ( .A(n5770), .B(n10809), .Z(n10811) );
  NAND U12616 ( .A(n10814), .B(nreg[248]), .Z(n5770) );
  NAND U12617 ( .A(n6107), .B(nreg[248]), .Z(n10814) );
  XOR U12618 ( .A(n10815), .B(n10816), .Z(n10809) );
  ANDN U12619 ( .A(n10817), .B(n5771), .Z(n10816) );
  XOR U12620 ( .A(n10818), .B(n10819), .Z(n5771) );
  IV U12621 ( .A(n10815), .Z(n10818) );
  XNOR U12622 ( .A(n5772), .B(n10815), .Z(n10817) );
  NAND U12623 ( .A(n10820), .B(nreg[247]), .Z(n5772) );
  NAND U12624 ( .A(n6107), .B(nreg[247]), .Z(n10820) );
  XOR U12625 ( .A(n10821), .B(n10822), .Z(n10815) );
  ANDN U12626 ( .A(n10823), .B(n5775), .Z(n10822) );
  XOR U12627 ( .A(n10824), .B(n10825), .Z(n5775) );
  IV U12628 ( .A(n10821), .Z(n10824) );
  XNOR U12629 ( .A(n5776), .B(n10821), .Z(n10823) );
  NAND U12630 ( .A(n10826), .B(nreg[246]), .Z(n5776) );
  NAND U12631 ( .A(n6107), .B(nreg[246]), .Z(n10826) );
  XOR U12632 ( .A(n10827), .B(n10828), .Z(n10821) );
  ANDN U12633 ( .A(n10829), .B(n5777), .Z(n10828) );
  XOR U12634 ( .A(n10830), .B(n10831), .Z(n5777) );
  IV U12635 ( .A(n10827), .Z(n10830) );
  XNOR U12636 ( .A(n5778), .B(n10827), .Z(n10829) );
  NAND U12637 ( .A(n10832), .B(nreg[245]), .Z(n5778) );
  NAND U12638 ( .A(n6107), .B(nreg[245]), .Z(n10832) );
  XOR U12639 ( .A(n10833), .B(n10834), .Z(n10827) );
  ANDN U12640 ( .A(n10835), .B(n5779), .Z(n10834) );
  XOR U12641 ( .A(n10836), .B(n10837), .Z(n5779) );
  IV U12642 ( .A(n10833), .Z(n10836) );
  XNOR U12643 ( .A(n5780), .B(n10833), .Z(n10835) );
  NAND U12644 ( .A(n10838), .B(nreg[244]), .Z(n5780) );
  NAND U12645 ( .A(n6107), .B(nreg[244]), .Z(n10838) );
  XOR U12646 ( .A(n10839), .B(n10840), .Z(n10833) );
  ANDN U12647 ( .A(n10841), .B(n5781), .Z(n10840) );
  XOR U12648 ( .A(n10842), .B(n10843), .Z(n5781) );
  IV U12649 ( .A(n10839), .Z(n10842) );
  XNOR U12650 ( .A(n5782), .B(n10839), .Z(n10841) );
  NAND U12651 ( .A(n10844), .B(nreg[243]), .Z(n5782) );
  NAND U12652 ( .A(n6107), .B(nreg[243]), .Z(n10844) );
  XOR U12653 ( .A(n10845), .B(n10846), .Z(n10839) );
  ANDN U12654 ( .A(n10847), .B(n5783), .Z(n10846) );
  XOR U12655 ( .A(n10848), .B(n10849), .Z(n5783) );
  IV U12656 ( .A(n10845), .Z(n10848) );
  XNOR U12657 ( .A(n5784), .B(n10845), .Z(n10847) );
  NAND U12658 ( .A(n10850), .B(nreg[242]), .Z(n5784) );
  NAND U12659 ( .A(n6107), .B(nreg[242]), .Z(n10850) );
  XOR U12660 ( .A(n10851), .B(n10852), .Z(n10845) );
  ANDN U12661 ( .A(n10853), .B(n5785), .Z(n10852) );
  XOR U12662 ( .A(n10854), .B(n10855), .Z(n5785) );
  IV U12663 ( .A(n10851), .Z(n10854) );
  XNOR U12664 ( .A(n5786), .B(n10851), .Z(n10853) );
  NAND U12665 ( .A(n10856), .B(nreg[241]), .Z(n5786) );
  NAND U12666 ( .A(n6107), .B(nreg[241]), .Z(n10856) );
  XOR U12667 ( .A(n10857), .B(n10858), .Z(n10851) );
  ANDN U12668 ( .A(n10859), .B(n5787), .Z(n10858) );
  XOR U12669 ( .A(n10860), .B(n10861), .Z(n5787) );
  IV U12670 ( .A(n10857), .Z(n10860) );
  XNOR U12671 ( .A(n5788), .B(n10857), .Z(n10859) );
  NAND U12672 ( .A(n10862), .B(nreg[240]), .Z(n5788) );
  NAND U12673 ( .A(n6107), .B(nreg[240]), .Z(n10862) );
  XOR U12674 ( .A(n10863), .B(n10864), .Z(n10857) );
  ANDN U12675 ( .A(n10865), .B(n5789), .Z(n10864) );
  XOR U12676 ( .A(n10866), .B(n10867), .Z(n5789) );
  IV U12677 ( .A(n10863), .Z(n10866) );
  XNOR U12678 ( .A(n5790), .B(n10863), .Z(n10865) );
  NAND U12679 ( .A(n10868), .B(nreg[239]), .Z(n5790) );
  NAND U12680 ( .A(n6107), .B(nreg[239]), .Z(n10868) );
  XOR U12681 ( .A(n10869), .B(n10870), .Z(n10863) );
  ANDN U12682 ( .A(n10871), .B(n5791), .Z(n10870) );
  XOR U12683 ( .A(n10872), .B(n10873), .Z(n5791) );
  IV U12684 ( .A(n10869), .Z(n10872) );
  XNOR U12685 ( .A(n5792), .B(n10869), .Z(n10871) );
  NAND U12686 ( .A(n10874), .B(nreg[238]), .Z(n5792) );
  NAND U12687 ( .A(n6107), .B(nreg[238]), .Z(n10874) );
  XOR U12688 ( .A(n10875), .B(n10876), .Z(n10869) );
  ANDN U12689 ( .A(n10877), .B(n5793), .Z(n10876) );
  XOR U12690 ( .A(n10878), .B(n10879), .Z(n5793) );
  IV U12691 ( .A(n10875), .Z(n10878) );
  XNOR U12692 ( .A(n5794), .B(n10875), .Z(n10877) );
  NAND U12693 ( .A(n10880), .B(nreg[237]), .Z(n5794) );
  NAND U12694 ( .A(n6107), .B(nreg[237]), .Z(n10880) );
  XOR U12695 ( .A(n10881), .B(n10882), .Z(n10875) );
  ANDN U12696 ( .A(n10883), .B(n5797), .Z(n10882) );
  XOR U12697 ( .A(n10884), .B(n10885), .Z(n5797) );
  IV U12698 ( .A(n10881), .Z(n10884) );
  XNOR U12699 ( .A(n5798), .B(n10881), .Z(n10883) );
  NAND U12700 ( .A(n10886), .B(nreg[236]), .Z(n5798) );
  NAND U12701 ( .A(n6107), .B(nreg[236]), .Z(n10886) );
  XOR U12702 ( .A(n10887), .B(n10888), .Z(n10881) );
  ANDN U12703 ( .A(n10889), .B(n5799), .Z(n10888) );
  XOR U12704 ( .A(n10890), .B(n10891), .Z(n5799) );
  IV U12705 ( .A(n10887), .Z(n10890) );
  XNOR U12706 ( .A(n5800), .B(n10887), .Z(n10889) );
  NAND U12707 ( .A(n10892), .B(nreg[235]), .Z(n5800) );
  NAND U12708 ( .A(n6107), .B(nreg[235]), .Z(n10892) );
  XOR U12709 ( .A(n10893), .B(n10894), .Z(n10887) );
  ANDN U12710 ( .A(n10895), .B(n5801), .Z(n10894) );
  XOR U12711 ( .A(n10896), .B(n10897), .Z(n5801) );
  IV U12712 ( .A(n10893), .Z(n10896) );
  XNOR U12713 ( .A(n5802), .B(n10893), .Z(n10895) );
  NAND U12714 ( .A(n10898), .B(nreg[234]), .Z(n5802) );
  NAND U12715 ( .A(n6107), .B(nreg[234]), .Z(n10898) );
  XOR U12716 ( .A(n10899), .B(n10900), .Z(n10893) );
  ANDN U12717 ( .A(n10901), .B(n5803), .Z(n10900) );
  XOR U12718 ( .A(n10902), .B(n10903), .Z(n5803) );
  IV U12719 ( .A(n10899), .Z(n10902) );
  XNOR U12720 ( .A(n5804), .B(n10899), .Z(n10901) );
  NAND U12721 ( .A(n10904), .B(nreg[233]), .Z(n5804) );
  NAND U12722 ( .A(n6107), .B(nreg[233]), .Z(n10904) );
  XOR U12723 ( .A(n10905), .B(n10906), .Z(n10899) );
  ANDN U12724 ( .A(n10907), .B(n5805), .Z(n10906) );
  XOR U12725 ( .A(n10908), .B(n10909), .Z(n5805) );
  IV U12726 ( .A(n10905), .Z(n10908) );
  XNOR U12727 ( .A(n5806), .B(n10905), .Z(n10907) );
  NAND U12728 ( .A(n10910), .B(nreg[232]), .Z(n5806) );
  NAND U12729 ( .A(n6107), .B(nreg[232]), .Z(n10910) );
  XOR U12730 ( .A(n10911), .B(n10912), .Z(n10905) );
  ANDN U12731 ( .A(n10913), .B(n5807), .Z(n10912) );
  XOR U12732 ( .A(n10914), .B(n10915), .Z(n5807) );
  IV U12733 ( .A(n10911), .Z(n10914) );
  XNOR U12734 ( .A(n5808), .B(n10911), .Z(n10913) );
  NAND U12735 ( .A(n10916), .B(nreg[231]), .Z(n5808) );
  NAND U12736 ( .A(n6107), .B(nreg[231]), .Z(n10916) );
  XOR U12737 ( .A(n10917), .B(n10918), .Z(n10911) );
  ANDN U12738 ( .A(n10919), .B(n5809), .Z(n10918) );
  XOR U12739 ( .A(n10920), .B(n10921), .Z(n5809) );
  IV U12740 ( .A(n10917), .Z(n10920) );
  XNOR U12741 ( .A(n5810), .B(n10917), .Z(n10919) );
  NAND U12742 ( .A(n10922), .B(nreg[230]), .Z(n5810) );
  NAND U12743 ( .A(n6107), .B(nreg[230]), .Z(n10922) );
  XOR U12744 ( .A(n10923), .B(n10924), .Z(n10917) );
  ANDN U12745 ( .A(n10925), .B(n5811), .Z(n10924) );
  XOR U12746 ( .A(n10926), .B(n10927), .Z(n5811) );
  IV U12747 ( .A(n10923), .Z(n10926) );
  XNOR U12748 ( .A(n5812), .B(n10923), .Z(n10925) );
  NAND U12749 ( .A(n10928), .B(nreg[229]), .Z(n5812) );
  NAND U12750 ( .A(n6107), .B(nreg[229]), .Z(n10928) );
  XOR U12751 ( .A(n10929), .B(n10930), .Z(n10923) );
  ANDN U12752 ( .A(n10931), .B(n5813), .Z(n10930) );
  XOR U12753 ( .A(n10932), .B(n10933), .Z(n5813) );
  IV U12754 ( .A(n10929), .Z(n10932) );
  XNOR U12755 ( .A(n5814), .B(n10929), .Z(n10931) );
  NAND U12756 ( .A(n10934), .B(nreg[228]), .Z(n5814) );
  NAND U12757 ( .A(n6107), .B(nreg[228]), .Z(n10934) );
  XOR U12758 ( .A(n10935), .B(n10936), .Z(n10929) );
  ANDN U12759 ( .A(n10937), .B(n5815), .Z(n10936) );
  XOR U12760 ( .A(n10938), .B(n10939), .Z(n5815) );
  IV U12761 ( .A(n10935), .Z(n10938) );
  XNOR U12762 ( .A(n5816), .B(n10935), .Z(n10937) );
  NAND U12763 ( .A(n10940), .B(nreg[227]), .Z(n5816) );
  NAND U12764 ( .A(n6107), .B(nreg[227]), .Z(n10940) );
  XOR U12765 ( .A(n10941), .B(n10942), .Z(n10935) );
  ANDN U12766 ( .A(n10943), .B(n5819), .Z(n10942) );
  XOR U12767 ( .A(n10944), .B(n10945), .Z(n5819) );
  IV U12768 ( .A(n10941), .Z(n10944) );
  XNOR U12769 ( .A(n5820), .B(n10941), .Z(n10943) );
  NAND U12770 ( .A(n10946), .B(nreg[226]), .Z(n5820) );
  NAND U12771 ( .A(n6107), .B(nreg[226]), .Z(n10946) );
  XOR U12772 ( .A(n10947), .B(n10948), .Z(n10941) );
  ANDN U12773 ( .A(n10949), .B(n5821), .Z(n10948) );
  XOR U12774 ( .A(n10950), .B(n10951), .Z(n5821) );
  IV U12775 ( .A(n10947), .Z(n10950) );
  XNOR U12776 ( .A(n5822), .B(n10947), .Z(n10949) );
  NAND U12777 ( .A(n10952), .B(nreg[225]), .Z(n5822) );
  NAND U12778 ( .A(n6107), .B(nreg[225]), .Z(n10952) );
  XOR U12779 ( .A(n10953), .B(n10954), .Z(n10947) );
  ANDN U12780 ( .A(n10955), .B(n5823), .Z(n10954) );
  XOR U12781 ( .A(n10956), .B(n10957), .Z(n5823) );
  IV U12782 ( .A(n10953), .Z(n10956) );
  XNOR U12783 ( .A(n5824), .B(n10953), .Z(n10955) );
  NAND U12784 ( .A(n10958), .B(nreg[224]), .Z(n5824) );
  NAND U12785 ( .A(n6107), .B(nreg[224]), .Z(n10958) );
  XOR U12786 ( .A(n10959), .B(n10960), .Z(n10953) );
  ANDN U12787 ( .A(n10961), .B(n5825), .Z(n10960) );
  XOR U12788 ( .A(n10962), .B(n10963), .Z(n5825) );
  IV U12789 ( .A(n10959), .Z(n10962) );
  XNOR U12790 ( .A(n5826), .B(n10959), .Z(n10961) );
  NAND U12791 ( .A(n10964), .B(nreg[223]), .Z(n5826) );
  NAND U12792 ( .A(n6107), .B(nreg[223]), .Z(n10964) );
  XOR U12793 ( .A(n10965), .B(n10966), .Z(n10959) );
  ANDN U12794 ( .A(n10967), .B(n5827), .Z(n10966) );
  XOR U12795 ( .A(n10968), .B(n10969), .Z(n5827) );
  IV U12796 ( .A(n10965), .Z(n10968) );
  XNOR U12797 ( .A(n5828), .B(n10965), .Z(n10967) );
  NAND U12798 ( .A(n10970), .B(nreg[222]), .Z(n5828) );
  NAND U12799 ( .A(n6107), .B(nreg[222]), .Z(n10970) );
  XOR U12800 ( .A(n10971), .B(n10972), .Z(n10965) );
  ANDN U12801 ( .A(n10973), .B(n5829), .Z(n10972) );
  XOR U12802 ( .A(n10974), .B(n10975), .Z(n5829) );
  IV U12803 ( .A(n10971), .Z(n10974) );
  XNOR U12804 ( .A(n5830), .B(n10971), .Z(n10973) );
  NAND U12805 ( .A(n10976), .B(nreg[221]), .Z(n5830) );
  NAND U12806 ( .A(n6107), .B(nreg[221]), .Z(n10976) );
  XOR U12807 ( .A(n10977), .B(n10978), .Z(n10971) );
  ANDN U12808 ( .A(n10979), .B(n5831), .Z(n10978) );
  XOR U12809 ( .A(n10980), .B(n10981), .Z(n5831) );
  IV U12810 ( .A(n10977), .Z(n10980) );
  XNOR U12811 ( .A(n5832), .B(n10977), .Z(n10979) );
  NAND U12812 ( .A(n10982), .B(nreg[220]), .Z(n5832) );
  NAND U12813 ( .A(n6107), .B(nreg[220]), .Z(n10982) );
  XOR U12814 ( .A(n10983), .B(n10984), .Z(n10977) );
  ANDN U12815 ( .A(n10985), .B(n5833), .Z(n10984) );
  XOR U12816 ( .A(n10986), .B(n10987), .Z(n5833) );
  IV U12817 ( .A(n10983), .Z(n10986) );
  XNOR U12818 ( .A(n5834), .B(n10983), .Z(n10985) );
  NAND U12819 ( .A(n10988), .B(nreg[219]), .Z(n5834) );
  NAND U12820 ( .A(n6107), .B(nreg[219]), .Z(n10988) );
  XOR U12821 ( .A(n10989), .B(n10990), .Z(n10983) );
  ANDN U12822 ( .A(n10991), .B(n5835), .Z(n10990) );
  XOR U12823 ( .A(n10992), .B(n10993), .Z(n5835) );
  IV U12824 ( .A(n10989), .Z(n10992) );
  XNOR U12825 ( .A(n5836), .B(n10989), .Z(n10991) );
  NAND U12826 ( .A(n10994), .B(nreg[218]), .Z(n5836) );
  NAND U12827 ( .A(n6107), .B(nreg[218]), .Z(n10994) );
  XOR U12828 ( .A(n10995), .B(n10996), .Z(n10989) );
  ANDN U12829 ( .A(n10997), .B(n5837), .Z(n10996) );
  XOR U12830 ( .A(n10998), .B(n10999), .Z(n5837) );
  IV U12831 ( .A(n10995), .Z(n10998) );
  XNOR U12832 ( .A(n5838), .B(n10995), .Z(n10997) );
  NAND U12833 ( .A(n11000), .B(nreg[217]), .Z(n5838) );
  NAND U12834 ( .A(n6107), .B(nreg[217]), .Z(n11000) );
  XOR U12835 ( .A(n11001), .B(n11002), .Z(n10995) );
  ANDN U12836 ( .A(n11003), .B(n5841), .Z(n11002) );
  XOR U12837 ( .A(n11004), .B(n11005), .Z(n5841) );
  IV U12838 ( .A(n11001), .Z(n11004) );
  XNOR U12839 ( .A(n5842), .B(n11001), .Z(n11003) );
  NAND U12840 ( .A(n11006), .B(nreg[216]), .Z(n5842) );
  NAND U12841 ( .A(n6107), .B(nreg[216]), .Z(n11006) );
  XOR U12842 ( .A(n11007), .B(n11008), .Z(n11001) );
  ANDN U12843 ( .A(n11009), .B(n5843), .Z(n11008) );
  XOR U12844 ( .A(n11010), .B(n11011), .Z(n5843) );
  IV U12845 ( .A(n11007), .Z(n11010) );
  XNOR U12846 ( .A(n5844), .B(n11007), .Z(n11009) );
  NAND U12847 ( .A(n11012), .B(nreg[215]), .Z(n5844) );
  NAND U12848 ( .A(n6107), .B(nreg[215]), .Z(n11012) );
  XOR U12849 ( .A(n11013), .B(n11014), .Z(n11007) );
  ANDN U12850 ( .A(n11015), .B(n5845), .Z(n11014) );
  XOR U12851 ( .A(n11016), .B(n11017), .Z(n5845) );
  IV U12852 ( .A(n11013), .Z(n11016) );
  XNOR U12853 ( .A(n5846), .B(n11013), .Z(n11015) );
  NAND U12854 ( .A(n11018), .B(nreg[214]), .Z(n5846) );
  NAND U12855 ( .A(n6107), .B(nreg[214]), .Z(n11018) );
  XOR U12856 ( .A(n11019), .B(n11020), .Z(n11013) );
  ANDN U12857 ( .A(n11021), .B(n5847), .Z(n11020) );
  XOR U12858 ( .A(n11022), .B(n11023), .Z(n5847) );
  IV U12859 ( .A(n11019), .Z(n11022) );
  XNOR U12860 ( .A(n5848), .B(n11019), .Z(n11021) );
  NAND U12861 ( .A(n11024), .B(nreg[213]), .Z(n5848) );
  NAND U12862 ( .A(n6107), .B(nreg[213]), .Z(n11024) );
  XOR U12863 ( .A(n11025), .B(n11026), .Z(n11019) );
  ANDN U12864 ( .A(n11027), .B(n5849), .Z(n11026) );
  XOR U12865 ( .A(n11028), .B(n11029), .Z(n5849) );
  IV U12866 ( .A(n11025), .Z(n11028) );
  XNOR U12867 ( .A(n5850), .B(n11025), .Z(n11027) );
  NAND U12868 ( .A(n11030), .B(nreg[212]), .Z(n5850) );
  NAND U12869 ( .A(n6107), .B(nreg[212]), .Z(n11030) );
  XOR U12870 ( .A(n11031), .B(n11032), .Z(n11025) );
  ANDN U12871 ( .A(n11033), .B(n5851), .Z(n11032) );
  XOR U12872 ( .A(n11034), .B(n11035), .Z(n5851) );
  IV U12873 ( .A(n11031), .Z(n11034) );
  XNOR U12874 ( .A(n5852), .B(n11031), .Z(n11033) );
  NAND U12875 ( .A(n11036), .B(nreg[211]), .Z(n5852) );
  NAND U12876 ( .A(n6107), .B(nreg[211]), .Z(n11036) );
  XOR U12877 ( .A(n11037), .B(n11038), .Z(n11031) );
  ANDN U12878 ( .A(n11039), .B(n5853), .Z(n11038) );
  XOR U12879 ( .A(n11040), .B(n11041), .Z(n5853) );
  IV U12880 ( .A(n11037), .Z(n11040) );
  XNOR U12881 ( .A(n5854), .B(n11037), .Z(n11039) );
  NAND U12882 ( .A(n11042), .B(nreg[210]), .Z(n5854) );
  NAND U12883 ( .A(n6107), .B(nreg[210]), .Z(n11042) );
  XOR U12884 ( .A(n11043), .B(n11044), .Z(n11037) );
  ANDN U12885 ( .A(n11045), .B(n5855), .Z(n11044) );
  XOR U12886 ( .A(n11046), .B(n11047), .Z(n5855) );
  IV U12887 ( .A(n11043), .Z(n11046) );
  XNOR U12888 ( .A(n5856), .B(n11043), .Z(n11045) );
  NAND U12889 ( .A(n11048), .B(nreg[209]), .Z(n5856) );
  NAND U12890 ( .A(n6107), .B(nreg[209]), .Z(n11048) );
  XOR U12891 ( .A(n11049), .B(n11050), .Z(n11043) );
  ANDN U12892 ( .A(n11051), .B(n5857), .Z(n11050) );
  XOR U12893 ( .A(n11052), .B(n11053), .Z(n5857) );
  IV U12894 ( .A(n11049), .Z(n11052) );
  XNOR U12895 ( .A(n5858), .B(n11049), .Z(n11051) );
  NAND U12896 ( .A(n11054), .B(nreg[208]), .Z(n5858) );
  NAND U12897 ( .A(n6107), .B(nreg[208]), .Z(n11054) );
  XOR U12898 ( .A(n11055), .B(n11056), .Z(n11049) );
  ANDN U12899 ( .A(n11057), .B(n5859), .Z(n11056) );
  XOR U12900 ( .A(n11058), .B(n11059), .Z(n5859) );
  IV U12901 ( .A(n11055), .Z(n11058) );
  XNOR U12902 ( .A(n5860), .B(n11055), .Z(n11057) );
  NAND U12903 ( .A(n11060), .B(nreg[207]), .Z(n5860) );
  NAND U12904 ( .A(n6107), .B(nreg[207]), .Z(n11060) );
  XOR U12905 ( .A(n11061), .B(n11062), .Z(n11055) );
  ANDN U12906 ( .A(n11063), .B(n5863), .Z(n11062) );
  XOR U12907 ( .A(n11064), .B(n11065), .Z(n5863) );
  IV U12908 ( .A(n11061), .Z(n11064) );
  XNOR U12909 ( .A(n5864), .B(n11061), .Z(n11063) );
  NAND U12910 ( .A(n11066), .B(nreg[206]), .Z(n5864) );
  NAND U12911 ( .A(n6107), .B(nreg[206]), .Z(n11066) );
  XOR U12912 ( .A(n11067), .B(n11068), .Z(n11061) );
  ANDN U12913 ( .A(n11069), .B(n5865), .Z(n11068) );
  XOR U12914 ( .A(n11070), .B(n11071), .Z(n5865) );
  IV U12915 ( .A(n11067), .Z(n11070) );
  XNOR U12916 ( .A(n5866), .B(n11067), .Z(n11069) );
  NAND U12917 ( .A(n11072), .B(nreg[205]), .Z(n5866) );
  NAND U12918 ( .A(n6107), .B(nreg[205]), .Z(n11072) );
  XOR U12919 ( .A(n11073), .B(n11074), .Z(n11067) );
  ANDN U12920 ( .A(n11075), .B(n5867), .Z(n11074) );
  XOR U12921 ( .A(n11076), .B(n11077), .Z(n5867) );
  IV U12922 ( .A(n11073), .Z(n11076) );
  XNOR U12923 ( .A(n5868), .B(n11073), .Z(n11075) );
  NAND U12924 ( .A(n11078), .B(nreg[204]), .Z(n5868) );
  NAND U12925 ( .A(n6107), .B(nreg[204]), .Z(n11078) );
  XOR U12926 ( .A(n11079), .B(n11080), .Z(n11073) );
  ANDN U12927 ( .A(n11081), .B(n5869), .Z(n11080) );
  XOR U12928 ( .A(n11082), .B(n11083), .Z(n5869) );
  IV U12929 ( .A(n11079), .Z(n11082) );
  XNOR U12930 ( .A(n5870), .B(n11079), .Z(n11081) );
  NAND U12931 ( .A(n11084), .B(nreg[203]), .Z(n5870) );
  NAND U12932 ( .A(n6107), .B(nreg[203]), .Z(n11084) );
  XOR U12933 ( .A(n11085), .B(n11086), .Z(n11079) );
  ANDN U12934 ( .A(n11087), .B(n5871), .Z(n11086) );
  XOR U12935 ( .A(n11088), .B(n11089), .Z(n5871) );
  IV U12936 ( .A(n11085), .Z(n11088) );
  XNOR U12937 ( .A(n5872), .B(n11085), .Z(n11087) );
  NAND U12938 ( .A(n11090), .B(nreg[202]), .Z(n5872) );
  NAND U12939 ( .A(n6107), .B(nreg[202]), .Z(n11090) );
  XOR U12940 ( .A(n11091), .B(n11092), .Z(n11085) );
  ANDN U12941 ( .A(n11093), .B(n5873), .Z(n11092) );
  XOR U12942 ( .A(n11094), .B(n11095), .Z(n5873) );
  IV U12943 ( .A(n11091), .Z(n11094) );
  XNOR U12944 ( .A(n5874), .B(n11091), .Z(n11093) );
  NAND U12945 ( .A(n11096), .B(nreg[201]), .Z(n5874) );
  NAND U12946 ( .A(n6107), .B(nreg[201]), .Z(n11096) );
  XOR U12947 ( .A(n11097), .B(n11098), .Z(n11091) );
  ANDN U12948 ( .A(n11099), .B(n5875), .Z(n11098) );
  XOR U12949 ( .A(n11100), .B(n11101), .Z(n5875) );
  IV U12950 ( .A(n11097), .Z(n11100) );
  XNOR U12951 ( .A(n5876), .B(n11097), .Z(n11099) );
  NAND U12952 ( .A(n11102), .B(nreg[200]), .Z(n5876) );
  NAND U12953 ( .A(n6107), .B(nreg[200]), .Z(n11102) );
  XOR U12954 ( .A(n11103), .B(n11104), .Z(n11097) );
  ANDN U12955 ( .A(n11105), .B(n5877), .Z(n11104) );
  XOR U12956 ( .A(n11106), .B(n11107), .Z(n5877) );
  IV U12957 ( .A(n11103), .Z(n11106) );
  XNOR U12958 ( .A(n5878), .B(n11103), .Z(n11105) );
  NAND U12959 ( .A(n11108), .B(nreg[199]), .Z(n5878) );
  NAND U12960 ( .A(n6107), .B(nreg[199]), .Z(n11108) );
  XOR U12961 ( .A(n11109), .B(n11110), .Z(n11103) );
  ANDN U12962 ( .A(n11111), .B(n5879), .Z(n11110) );
  XOR U12963 ( .A(n11112), .B(n11113), .Z(n5879) );
  IV U12964 ( .A(n11109), .Z(n11112) );
  XNOR U12965 ( .A(n5880), .B(n11109), .Z(n11111) );
  NAND U12966 ( .A(n11114), .B(nreg[198]), .Z(n5880) );
  NAND U12967 ( .A(n6107), .B(nreg[198]), .Z(n11114) );
  XOR U12968 ( .A(n11115), .B(n11116), .Z(n11109) );
  ANDN U12969 ( .A(n11117), .B(n5881), .Z(n11116) );
  XOR U12970 ( .A(n11118), .B(n11119), .Z(n5881) );
  IV U12971 ( .A(n11115), .Z(n11118) );
  XNOR U12972 ( .A(n5882), .B(n11115), .Z(n11117) );
  NAND U12973 ( .A(n11120), .B(nreg[197]), .Z(n5882) );
  NAND U12974 ( .A(n6107), .B(nreg[197]), .Z(n11120) );
  XOR U12975 ( .A(n11121), .B(n11122), .Z(n11115) );
  ANDN U12976 ( .A(n11123), .B(n5885), .Z(n11122) );
  XOR U12977 ( .A(n11124), .B(n11125), .Z(n5885) );
  IV U12978 ( .A(n11121), .Z(n11124) );
  XNOR U12979 ( .A(n5886), .B(n11121), .Z(n11123) );
  NAND U12980 ( .A(n11126), .B(nreg[196]), .Z(n5886) );
  NAND U12981 ( .A(n6107), .B(nreg[196]), .Z(n11126) );
  XOR U12982 ( .A(n11127), .B(n11128), .Z(n11121) );
  ANDN U12983 ( .A(n11129), .B(n5887), .Z(n11128) );
  XOR U12984 ( .A(n11130), .B(n11131), .Z(n5887) );
  IV U12985 ( .A(n11127), .Z(n11130) );
  XNOR U12986 ( .A(n5888), .B(n11127), .Z(n11129) );
  NAND U12987 ( .A(n11132), .B(nreg[195]), .Z(n5888) );
  NAND U12988 ( .A(n6107), .B(nreg[195]), .Z(n11132) );
  XOR U12989 ( .A(n11133), .B(n11134), .Z(n11127) );
  ANDN U12990 ( .A(n11135), .B(n5889), .Z(n11134) );
  XOR U12991 ( .A(n11136), .B(n11137), .Z(n5889) );
  IV U12992 ( .A(n11133), .Z(n11136) );
  XNOR U12993 ( .A(n5890), .B(n11133), .Z(n11135) );
  NAND U12994 ( .A(n11138), .B(nreg[194]), .Z(n5890) );
  NAND U12995 ( .A(n6107), .B(nreg[194]), .Z(n11138) );
  XOR U12996 ( .A(n11139), .B(n11140), .Z(n11133) );
  ANDN U12997 ( .A(n11141), .B(n5891), .Z(n11140) );
  XOR U12998 ( .A(n11142), .B(n11143), .Z(n5891) );
  IV U12999 ( .A(n11139), .Z(n11142) );
  XNOR U13000 ( .A(n5892), .B(n11139), .Z(n11141) );
  NAND U13001 ( .A(n11144), .B(nreg[193]), .Z(n5892) );
  NAND U13002 ( .A(n6107), .B(nreg[193]), .Z(n11144) );
  XOR U13003 ( .A(n11145), .B(n11146), .Z(n11139) );
  ANDN U13004 ( .A(n11147), .B(n5893), .Z(n11146) );
  XOR U13005 ( .A(n11148), .B(n11149), .Z(n5893) );
  IV U13006 ( .A(n11145), .Z(n11148) );
  XNOR U13007 ( .A(n5894), .B(n11145), .Z(n11147) );
  NAND U13008 ( .A(n11150), .B(nreg[192]), .Z(n5894) );
  NAND U13009 ( .A(n6107), .B(nreg[192]), .Z(n11150) );
  XOR U13010 ( .A(n11151), .B(n11152), .Z(n11145) );
  ANDN U13011 ( .A(n11153), .B(n5895), .Z(n11152) );
  XOR U13012 ( .A(n11154), .B(n11155), .Z(n5895) );
  IV U13013 ( .A(n11151), .Z(n11154) );
  XNOR U13014 ( .A(n5896), .B(n11151), .Z(n11153) );
  NAND U13015 ( .A(n11156), .B(nreg[191]), .Z(n5896) );
  NAND U13016 ( .A(n6107), .B(nreg[191]), .Z(n11156) );
  XOR U13017 ( .A(n11157), .B(n11158), .Z(n11151) );
  ANDN U13018 ( .A(n11159), .B(n5897), .Z(n11158) );
  XOR U13019 ( .A(n11160), .B(n11161), .Z(n5897) );
  IV U13020 ( .A(n11157), .Z(n11160) );
  XNOR U13021 ( .A(n5898), .B(n11157), .Z(n11159) );
  NAND U13022 ( .A(n11162), .B(nreg[190]), .Z(n5898) );
  NAND U13023 ( .A(n6107), .B(nreg[190]), .Z(n11162) );
  XOR U13024 ( .A(n11163), .B(n11164), .Z(n11157) );
  ANDN U13025 ( .A(n11165), .B(n5899), .Z(n11164) );
  XOR U13026 ( .A(n11166), .B(n11167), .Z(n5899) );
  IV U13027 ( .A(n11163), .Z(n11166) );
  XNOR U13028 ( .A(n5900), .B(n11163), .Z(n11165) );
  NAND U13029 ( .A(n11168), .B(nreg[189]), .Z(n5900) );
  NAND U13030 ( .A(n6107), .B(nreg[189]), .Z(n11168) );
  XOR U13031 ( .A(n11169), .B(n11170), .Z(n11163) );
  ANDN U13032 ( .A(n11171), .B(n5901), .Z(n11170) );
  XOR U13033 ( .A(n11172), .B(n11173), .Z(n5901) );
  IV U13034 ( .A(n11169), .Z(n11172) );
  XNOR U13035 ( .A(n5902), .B(n11169), .Z(n11171) );
  NAND U13036 ( .A(n11174), .B(nreg[188]), .Z(n5902) );
  NAND U13037 ( .A(n6107), .B(nreg[188]), .Z(n11174) );
  XOR U13038 ( .A(n11175), .B(n11176), .Z(n11169) );
  ANDN U13039 ( .A(n11177), .B(n5903), .Z(n11176) );
  XOR U13040 ( .A(n11178), .B(n11179), .Z(n5903) );
  IV U13041 ( .A(n11175), .Z(n11178) );
  XNOR U13042 ( .A(n5904), .B(n11175), .Z(n11177) );
  NAND U13043 ( .A(n11180), .B(nreg[187]), .Z(n5904) );
  NAND U13044 ( .A(n6107), .B(nreg[187]), .Z(n11180) );
  XOR U13045 ( .A(n11181), .B(n11182), .Z(n11175) );
  ANDN U13046 ( .A(n11183), .B(n5907), .Z(n11182) );
  XOR U13047 ( .A(n11184), .B(n11185), .Z(n5907) );
  IV U13048 ( .A(n11181), .Z(n11184) );
  XNOR U13049 ( .A(n5908), .B(n11181), .Z(n11183) );
  NAND U13050 ( .A(n11186), .B(nreg[186]), .Z(n5908) );
  NAND U13051 ( .A(n6107), .B(nreg[186]), .Z(n11186) );
  XOR U13052 ( .A(n11187), .B(n11188), .Z(n11181) );
  ANDN U13053 ( .A(n11189), .B(n5909), .Z(n11188) );
  XOR U13054 ( .A(n11190), .B(n11191), .Z(n5909) );
  IV U13055 ( .A(n11187), .Z(n11190) );
  XNOR U13056 ( .A(n5910), .B(n11187), .Z(n11189) );
  NAND U13057 ( .A(n11192), .B(nreg[185]), .Z(n5910) );
  NAND U13058 ( .A(n6107), .B(nreg[185]), .Z(n11192) );
  XOR U13059 ( .A(n11193), .B(n11194), .Z(n11187) );
  ANDN U13060 ( .A(n11195), .B(n5911), .Z(n11194) );
  XOR U13061 ( .A(n11196), .B(n11197), .Z(n5911) );
  IV U13062 ( .A(n11193), .Z(n11196) );
  XNOR U13063 ( .A(n5912), .B(n11193), .Z(n11195) );
  NAND U13064 ( .A(n11198), .B(nreg[184]), .Z(n5912) );
  NAND U13065 ( .A(n6107), .B(nreg[184]), .Z(n11198) );
  XOR U13066 ( .A(n11199), .B(n11200), .Z(n11193) );
  ANDN U13067 ( .A(n11201), .B(n5913), .Z(n11200) );
  XOR U13068 ( .A(n11202), .B(n11203), .Z(n5913) );
  IV U13069 ( .A(n11199), .Z(n11202) );
  XNOR U13070 ( .A(n5914), .B(n11199), .Z(n11201) );
  NAND U13071 ( .A(n11204), .B(nreg[183]), .Z(n5914) );
  NAND U13072 ( .A(n6107), .B(nreg[183]), .Z(n11204) );
  XOR U13073 ( .A(n11205), .B(n11206), .Z(n11199) );
  ANDN U13074 ( .A(n11207), .B(n5915), .Z(n11206) );
  XOR U13075 ( .A(n11208), .B(n11209), .Z(n5915) );
  IV U13076 ( .A(n11205), .Z(n11208) );
  XNOR U13077 ( .A(n5916), .B(n11205), .Z(n11207) );
  NAND U13078 ( .A(n11210), .B(nreg[182]), .Z(n5916) );
  NAND U13079 ( .A(n6107), .B(nreg[182]), .Z(n11210) );
  XOR U13080 ( .A(n11211), .B(n11212), .Z(n11205) );
  ANDN U13081 ( .A(n11213), .B(n5917), .Z(n11212) );
  XOR U13082 ( .A(n11214), .B(n11215), .Z(n5917) );
  IV U13083 ( .A(n11211), .Z(n11214) );
  XNOR U13084 ( .A(n5918), .B(n11211), .Z(n11213) );
  NAND U13085 ( .A(n11216), .B(nreg[181]), .Z(n5918) );
  NAND U13086 ( .A(n6107), .B(nreg[181]), .Z(n11216) );
  XOR U13087 ( .A(n11217), .B(n11218), .Z(n11211) );
  ANDN U13088 ( .A(n11219), .B(n5919), .Z(n11218) );
  XOR U13089 ( .A(n11220), .B(n11221), .Z(n5919) );
  IV U13090 ( .A(n11217), .Z(n11220) );
  XNOR U13091 ( .A(n5920), .B(n11217), .Z(n11219) );
  NAND U13092 ( .A(n11222), .B(nreg[180]), .Z(n5920) );
  NAND U13093 ( .A(n6107), .B(nreg[180]), .Z(n11222) );
  XOR U13094 ( .A(n11223), .B(n11224), .Z(n11217) );
  ANDN U13095 ( .A(n11225), .B(n5921), .Z(n11224) );
  XOR U13096 ( .A(n11226), .B(n11227), .Z(n5921) );
  IV U13097 ( .A(n11223), .Z(n11226) );
  XNOR U13098 ( .A(n5922), .B(n11223), .Z(n11225) );
  NAND U13099 ( .A(n11228), .B(nreg[179]), .Z(n5922) );
  NAND U13100 ( .A(n6107), .B(nreg[179]), .Z(n11228) );
  XOR U13101 ( .A(n11229), .B(n11230), .Z(n11223) );
  ANDN U13102 ( .A(n11231), .B(n5923), .Z(n11230) );
  XOR U13103 ( .A(n11232), .B(n11233), .Z(n5923) );
  IV U13104 ( .A(n11229), .Z(n11232) );
  XNOR U13105 ( .A(n5924), .B(n11229), .Z(n11231) );
  NAND U13106 ( .A(n11234), .B(nreg[178]), .Z(n5924) );
  NAND U13107 ( .A(n6107), .B(nreg[178]), .Z(n11234) );
  XOR U13108 ( .A(n11235), .B(n11236), .Z(n11229) );
  ANDN U13109 ( .A(n11237), .B(n5925), .Z(n11236) );
  XOR U13110 ( .A(n11238), .B(n11239), .Z(n5925) );
  IV U13111 ( .A(n11235), .Z(n11238) );
  XNOR U13112 ( .A(n5926), .B(n11235), .Z(n11237) );
  NAND U13113 ( .A(n11240), .B(nreg[177]), .Z(n5926) );
  NAND U13114 ( .A(n6107), .B(nreg[177]), .Z(n11240) );
  XOR U13115 ( .A(n11241), .B(n11242), .Z(n11235) );
  ANDN U13116 ( .A(n11243), .B(n5929), .Z(n11242) );
  XOR U13117 ( .A(n11244), .B(n11245), .Z(n5929) );
  IV U13118 ( .A(n11241), .Z(n11244) );
  XNOR U13119 ( .A(n5930), .B(n11241), .Z(n11243) );
  NAND U13120 ( .A(n11246), .B(nreg[176]), .Z(n5930) );
  NAND U13121 ( .A(n6107), .B(nreg[176]), .Z(n11246) );
  XOR U13122 ( .A(n11247), .B(n11248), .Z(n11241) );
  ANDN U13123 ( .A(n11249), .B(n5931), .Z(n11248) );
  XOR U13124 ( .A(n11250), .B(n11251), .Z(n5931) );
  IV U13125 ( .A(n11247), .Z(n11250) );
  XNOR U13126 ( .A(n5932), .B(n11247), .Z(n11249) );
  NAND U13127 ( .A(n11252), .B(nreg[175]), .Z(n5932) );
  NAND U13128 ( .A(n6107), .B(nreg[175]), .Z(n11252) );
  XOR U13129 ( .A(n11253), .B(n11254), .Z(n11247) );
  ANDN U13130 ( .A(n11255), .B(n5933), .Z(n11254) );
  XOR U13131 ( .A(n11256), .B(n11257), .Z(n5933) );
  IV U13132 ( .A(n11253), .Z(n11256) );
  XNOR U13133 ( .A(n5934), .B(n11253), .Z(n11255) );
  NAND U13134 ( .A(n11258), .B(nreg[174]), .Z(n5934) );
  NAND U13135 ( .A(n6107), .B(nreg[174]), .Z(n11258) );
  XOR U13136 ( .A(n11259), .B(n11260), .Z(n11253) );
  ANDN U13137 ( .A(n11261), .B(n5935), .Z(n11260) );
  XOR U13138 ( .A(n11262), .B(n11263), .Z(n5935) );
  IV U13139 ( .A(n11259), .Z(n11262) );
  XNOR U13140 ( .A(n5936), .B(n11259), .Z(n11261) );
  NAND U13141 ( .A(n11264), .B(nreg[173]), .Z(n5936) );
  NAND U13142 ( .A(n6107), .B(nreg[173]), .Z(n11264) );
  XOR U13143 ( .A(n11265), .B(n11266), .Z(n11259) );
  ANDN U13144 ( .A(n11267), .B(n5937), .Z(n11266) );
  XOR U13145 ( .A(n11268), .B(n11269), .Z(n5937) );
  IV U13146 ( .A(n11265), .Z(n11268) );
  XNOR U13147 ( .A(n5938), .B(n11265), .Z(n11267) );
  NAND U13148 ( .A(n11270), .B(nreg[172]), .Z(n5938) );
  NAND U13149 ( .A(n6107), .B(nreg[172]), .Z(n11270) );
  XOR U13150 ( .A(n11271), .B(n11272), .Z(n11265) );
  ANDN U13151 ( .A(n11273), .B(n5939), .Z(n11272) );
  XOR U13152 ( .A(n11274), .B(n11275), .Z(n5939) );
  IV U13153 ( .A(n11271), .Z(n11274) );
  XNOR U13154 ( .A(n5940), .B(n11271), .Z(n11273) );
  NAND U13155 ( .A(n11276), .B(nreg[171]), .Z(n5940) );
  NAND U13156 ( .A(n6107), .B(nreg[171]), .Z(n11276) );
  XOR U13157 ( .A(n11277), .B(n11278), .Z(n11271) );
  ANDN U13158 ( .A(n11279), .B(n5941), .Z(n11278) );
  XOR U13159 ( .A(n11280), .B(n11281), .Z(n5941) );
  IV U13160 ( .A(n11277), .Z(n11280) );
  XNOR U13161 ( .A(n5942), .B(n11277), .Z(n11279) );
  NAND U13162 ( .A(n11282), .B(nreg[170]), .Z(n5942) );
  NAND U13163 ( .A(n6107), .B(nreg[170]), .Z(n11282) );
  XOR U13164 ( .A(n11283), .B(n11284), .Z(n11277) );
  ANDN U13165 ( .A(n11285), .B(n5943), .Z(n11284) );
  XOR U13166 ( .A(n11286), .B(n11287), .Z(n5943) );
  IV U13167 ( .A(n11283), .Z(n11286) );
  XNOR U13168 ( .A(n5944), .B(n11283), .Z(n11285) );
  NAND U13169 ( .A(n11288), .B(nreg[169]), .Z(n5944) );
  NAND U13170 ( .A(n6107), .B(nreg[169]), .Z(n11288) );
  XOR U13171 ( .A(n11289), .B(n11290), .Z(n11283) );
  ANDN U13172 ( .A(n11291), .B(n5945), .Z(n11290) );
  XOR U13173 ( .A(n11292), .B(n11293), .Z(n5945) );
  IV U13174 ( .A(n11289), .Z(n11292) );
  XNOR U13175 ( .A(n5946), .B(n11289), .Z(n11291) );
  NAND U13176 ( .A(n11294), .B(nreg[168]), .Z(n5946) );
  NAND U13177 ( .A(n6107), .B(nreg[168]), .Z(n11294) );
  XOR U13178 ( .A(n11295), .B(n11296), .Z(n11289) );
  ANDN U13179 ( .A(n11297), .B(n5947), .Z(n11296) );
  XOR U13180 ( .A(n11298), .B(n11299), .Z(n5947) );
  IV U13181 ( .A(n11295), .Z(n11298) );
  XNOR U13182 ( .A(n5948), .B(n11295), .Z(n11297) );
  NAND U13183 ( .A(n11300), .B(nreg[167]), .Z(n5948) );
  NAND U13184 ( .A(n6107), .B(nreg[167]), .Z(n11300) );
  XOR U13185 ( .A(n11301), .B(n11302), .Z(n11295) );
  ANDN U13186 ( .A(n11303), .B(n5951), .Z(n11302) );
  XOR U13187 ( .A(n11304), .B(n11305), .Z(n5951) );
  IV U13188 ( .A(n11301), .Z(n11304) );
  XNOR U13189 ( .A(n5952), .B(n11301), .Z(n11303) );
  NAND U13190 ( .A(n11306), .B(nreg[166]), .Z(n5952) );
  NAND U13191 ( .A(n6107), .B(nreg[166]), .Z(n11306) );
  XOR U13192 ( .A(n11307), .B(n11308), .Z(n11301) );
  ANDN U13193 ( .A(n11309), .B(n5953), .Z(n11308) );
  XOR U13194 ( .A(n11310), .B(n11311), .Z(n5953) );
  IV U13195 ( .A(n11307), .Z(n11310) );
  XNOR U13196 ( .A(n5954), .B(n11307), .Z(n11309) );
  NAND U13197 ( .A(n11312), .B(nreg[165]), .Z(n5954) );
  NAND U13198 ( .A(n6107), .B(nreg[165]), .Z(n11312) );
  XOR U13199 ( .A(n11313), .B(n11314), .Z(n11307) );
  ANDN U13200 ( .A(n11315), .B(n5955), .Z(n11314) );
  XOR U13201 ( .A(n11316), .B(n11317), .Z(n5955) );
  IV U13202 ( .A(n11313), .Z(n11316) );
  XNOR U13203 ( .A(n5956), .B(n11313), .Z(n11315) );
  NAND U13204 ( .A(n11318), .B(nreg[164]), .Z(n5956) );
  NAND U13205 ( .A(n6107), .B(nreg[164]), .Z(n11318) );
  XOR U13206 ( .A(n11319), .B(n11320), .Z(n11313) );
  ANDN U13207 ( .A(n11321), .B(n5957), .Z(n11320) );
  XOR U13208 ( .A(n11322), .B(n11323), .Z(n5957) );
  IV U13209 ( .A(n11319), .Z(n11322) );
  XNOR U13210 ( .A(n5958), .B(n11319), .Z(n11321) );
  NAND U13211 ( .A(n11324), .B(nreg[163]), .Z(n5958) );
  NAND U13212 ( .A(n6107), .B(nreg[163]), .Z(n11324) );
  XOR U13213 ( .A(n11325), .B(n11326), .Z(n11319) );
  ANDN U13214 ( .A(n11327), .B(n5959), .Z(n11326) );
  XOR U13215 ( .A(n11328), .B(n11329), .Z(n5959) );
  IV U13216 ( .A(n11325), .Z(n11328) );
  XNOR U13217 ( .A(n5960), .B(n11325), .Z(n11327) );
  NAND U13218 ( .A(n11330), .B(nreg[162]), .Z(n5960) );
  NAND U13219 ( .A(n6107), .B(nreg[162]), .Z(n11330) );
  XOR U13220 ( .A(n11331), .B(n11332), .Z(n11325) );
  ANDN U13221 ( .A(n11333), .B(n5961), .Z(n11332) );
  XOR U13222 ( .A(n11334), .B(n11335), .Z(n5961) );
  IV U13223 ( .A(n11331), .Z(n11334) );
  XNOR U13224 ( .A(n5962), .B(n11331), .Z(n11333) );
  NAND U13225 ( .A(n11336), .B(nreg[161]), .Z(n5962) );
  NAND U13226 ( .A(n6107), .B(nreg[161]), .Z(n11336) );
  XOR U13227 ( .A(n11337), .B(n11338), .Z(n11331) );
  ANDN U13228 ( .A(n11339), .B(n5963), .Z(n11338) );
  XOR U13229 ( .A(n11340), .B(n11341), .Z(n5963) );
  IV U13230 ( .A(n11337), .Z(n11340) );
  XNOR U13231 ( .A(n5964), .B(n11337), .Z(n11339) );
  NAND U13232 ( .A(n11342), .B(nreg[160]), .Z(n5964) );
  NAND U13233 ( .A(n6107), .B(nreg[160]), .Z(n11342) );
  XOR U13234 ( .A(n11343), .B(n11344), .Z(n11337) );
  ANDN U13235 ( .A(n11345), .B(n5965), .Z(n11344) );
  XOR U13236 ( .A(n11346), .B(n11347), .Z(n5965) );
  IV U13237 ( .A(n11343), .Z(n11346) );
  XNOR U13238 ( .A(n5966), .B(n11343), .Z(n11345) );
  NAND U13239 ( .A(n11348), .B(nreg[159]), .Z(n5966) );
  NAND U13240 ( .A(n6107), .B(nreg[159]), .Z(n11348) );
  XOR U13241 ( .A(n11349), .B(n11350), .Z(n11343) );
  ANDN U13242 ( .A(n11351), .B(n5967), .Z(n11350) );
  XOR U13243 ( .A(n11352), .B(n11353), .Z(n5967) );
  IV U13244 ( .A(n11349), .Z(n11352) );
  XNOR U13245 ( .A(n5968), .B(n11349), .Z(n11351) );
  NAND U13246 ( .A(n11354), .B(nreg[158]), .Z(n5968) );
  NAND U13247 ( .A(n6107), .B(nreg[158]), .Z(n11354) );
  XOR U13248 ( .A(n11355), .B(n11356), .Z(n11349) );
  ANDN U13249 ( .A(n11357), .B(n5969), .Z(n11356) );
  XOR U13250 ( .A(n11358), .B(n11359), .Z(n5969) );
  IV U13251 ( .A(n11355), .Z(n11358) );
  XNOR U13252 ( .A(n5970), .B(n11355), .Z(n11357) );
  NAND U13253 ( .A(n11360), .B(nreg[157]), .Z(n5970) );
  NAND U13254 ( .A(n6107), .B(nreg[157]), .Z(n11360) );
  XOR U13255 ( .A(n11361), .B(n11362), .Z(n11355) );
  ANDN U13256 ( .A(n11363), .B(n5973), .Z(n11362) );
  XOR U13257 ( .A(n11364), .B(n11365), .Z(n5973) );
  IV U13258 ( .A(n11361), .Z(n11364) );
  XNOR U13259 ( .A(n5974), .B(n11361), .Z(n11363) );
  NAND U13260 ( .A(n11366), .B(nreg[156]), .Z(n5974) );
  NAND U13261 ( .A(n6107), .B(nreg[156]), .Z(n11366) );
  XOR U13262 ( .A(n11367), .B(n11368), .Z(n11361) );
  ANDN U13263 ( .A(n11369), .B(n5975), .Z(n11368) );
  XOR U13264 ( .A(n11370), .B(n11371), .Z(n5975) );
  IV U13265 ( .A(n11367), .Z(n11370) );
  XNOR U13266 ( .A(n5976), .B(n11367), .Z(n11369) );
  NAND U13267 ( .A(n11372), .B(nreg[155]), .Z(n5976) );
  NAND U13268 ( .A(n6107), .B(nreg[155]), .Z(n11372) );
  XOR U13269 ( .A(n11373), .B(n11374), .Z(n11367) );
  ANDN U13270 ( .A(n11375), .B(n5977), .Z(n11374) );
  XOR U13271 ( .A(n11376), .B(n11377), .Z(n5977) );
  IV U13272 ( .A(n11373), .Z(n11376) );
  XNOR U13273 ( .A(n5978), .B(n11373), .Z(n11375) );
  NAND U13274 ( .A(n11378), .B(nreg[154]), .Z(n5978) );
  NAND U13275 ( .A(n6107), .B(nreg[154]), .Z(n11378) );
  XOR U13276 ( .A(n11379), .B(n11380), .Z(n11373) );
  ANDN U13277 ( .A(n11381), .B(n5979), .Z(n11380) );
  XOR U13278 ( .A(n11382), .B(n11383), .Z(n5979) );
  IV U13279 ( .A(n11379), .Z(n11382) );
  XNOR U13280 ( .A(n5980), .B(n11379), .Z(n11381) );
  NAND U13281 ( .A(n11384), .B(nreg[153]), .Z(n5980) );
  NAND U13282 ( .A(n6107), .B(nreg[153]), .Z(n11384) );
  XOR U13283 ( .A(n11385), .B(n11386), .Z(n11379) );
  ANDN U13284 ( .A(n11387), .B(n5981), .Z(n11386) );
  XOR U13285 ( .A(n11388), .B(n11389), .Z(n5981) );
  IV U13286 ( .A(n11385), .Z(n11388) );
  XNOR U13287 ( .A(n5982), .B(n11385), .Z(n11387) );
  NAND U13288 ( .A(n11390), .B(nreg[152]), .Z(n5982) );
  NAND U13289 ( .A(n6107), .B(nreg[152]), .Z(n11390) );
  XOR U13290 ( .A(n11391), .B(n11392), .Z(n11385) );
  ANDN U13291 ( .A(n11393), .B(n5983), .Z(n11392) );
  XOR U13292 ( .A(n11394), .B(n11395), .Z(n5983) );
  IV U13293 ( .A(n11391), .Z(n11394) );
  XNOR U13294 ( .A(n5984), .B(n11391), .Z(n11393) );
  NAND U13295 ( .A(n11396), .B(nreg[151]), .Z(n5984) );
  NAND U13296 ( .A(n6107), .B(nreg[151]), .Z(n11396) );
  XOR U13297 ( .A(n11397), .B(n11398), .Z(n11391) );
  ANDN U13298 ( .A(n11399), .B(n5985), .Z(n11398) );
  XOR U13299 ( .A(n11400), .B(n11401), .Z(n5985) );
  IV U13300 ( .A(n11397), .Z(n11400) );
  XNOR U13301 ( .A(n5986), .B(n11397), .Z(n11399) );
  NAND U13302 ( .A(n11402), .B(nreg[150]), .Z(n5986) );
  NAND U13303 ( .A(n6107), .B(nreg[150]), .Z(n11402) );
  XOR U13304 ( .A(n11403), .B(n11404), .Z(n11397) );
  ANDN U13305 ( .A(n11405), .B(n5987), .Z(n11404) );
  XOR U13306 ( .A(n11406), .B(n11407), .Z(n5987) );
  IV U13307 ( .A(n11403), .Z(n11406) );
  XNOR U13308 ( .A(n5988), .B(n11403), .Z(n11405) );
  NAND U13309 ( .A(n11408), .B(nreg[149]), .Z(n5988) );
  NAND U13310 ( .A(n6107), .B(nreg[149]), .Z(n11408) );
  XOR U13311 ( .A(n11409), .B(n11410), .Z(n11403) );
  ANDN U13312 ( .A(n11411), .B(n5989), .Z(n11410) );
  XOR U13313 ( .A(n11412), .B(n11413), .Z(n5989) );
  IV U13314 ( .A(n11409), .Z(n11412) );
  XNOR U13315 ( .A(n5990), .B(n11409), .Z(n11411) );
  NAND U13316 ( .A(n11414), .B(nreg[148]), .Z(n5990) );
  NAND U13317 ( .A(n6107), .B(nreg[148]), .Z(n11414) );
  XOR U13318 ( .A(n11415), .B(n11416), .Z(n11409) );
  ANDN U13319 ( .A(n11417), .B(n5991), .Z(n11416) );
  XOR U13320 ( .A(n11418), .B(n11419), .Z(n5991) );
  IV U13321 ( .A(n11415), .Z(n11418) );
  XNOR U13322 ( .A(n5992), .B(n11415), .Z(n11417) );
  NAND U13323 ( .A(n11420), .B(nreg[147]), .Z(n5992) );
  NAND U13324 ( .A(n6107), .B(nreg[147]), .Z(n11420) );
  XOR U13325 ( .A(n11421), .B(n11422), .Z(n11415) );
  ANDN U13326 ( .A(n11423), .B(n5995), .Z(n11422) );
  XOR U13327 ( .A(n11424), .B(n11425), .Z(n5995) );
  IV U13328 ( .A(n11421), .Z(n11424) );
  XNOR U13329 ( .A(n5996), .B(n11421), .Z(n11423) );
  NAND U13330 ( .A(n11426), .B(nreg[146]), .Z(n5996) );
  NAND U13331 ( .A(n6107), .B(nreg[146]), .Z(n11426) );
  XOR U13332 ( .A(n11427), .B(n11428), .Z(n11421) );
  ANDN U13333 ( .A(n11429), .B(n5997), .Z(n11428) );
  XOR U13334 ( .A(n11430), .B(n11431), .Z(n5997) );
  IV U13335 ( .A(n11427), .Z(n11430) );
  XNOR U13336 ( .A(n5998), .B(n11427), .Z(n11429) );
  NAND U13337 ( .A(n11432), .B(nreg[145]), .Z(n5998) );
  NAND U13338 ( .A(n6107), .B(nreg[145]), .Z(n11432) );
  XOR U13339 ( .A(n11433), .B(n11434), .Z(n11427) );
  ANDN U13340 ( .A(n11435), .B(n5999), .Z(n11434) );
  XOR U13341 ( .A(n11436), .B(n11437), .Z(n5999) );
  IV U13342 ( .A(n11433), .Z(n11436) );
  XNOR U13343 ( .A(n6000), .B(n11433), .Z(n11435) );
  NAND U13344 ( .A(n11438), .B(nreg[144]), .Z(n6000) );
  NAND U13345 ( .A(n6107), .B(nreg[144]), .Z(n11438) );
  XOR U13346 ( .A(n11439), .B(n11440), .Z(n11433) );
  ANDN U13347 ( .A(n11441), .B(n6001), .Z(n11440) );
  XOR U13348 ( .A(n11442), .B(n11443), .Z(n6001) );
  IV U13349 ( .A(n11439), .Z(n11442) );
  XNOR U13350 ( .A(n6002), .B(n11439), .Z(n11441) );
  NAND U13351 ( .A(n11444), .B(nreg[143]), .Z(n6002) );
  NAND U13352 ( .A(n6107), .B(nreg[143]), .Z(n11444) );
  XOR U13353 ( .A(n11445), .B(n11446), .Z(n11439) );
  ANDN U13354 ( .A(n11447), .B(n6003), .Z(n11446) );
  XOR U13355 ( .A(n11448), .B(n11449), .Z(n6003) );
  IV U13356 ( .A(n11445), .Z(n11448) );
  XNOR U13357 ( .A(n6004), .B(n11445), .Z(n11447) );
  NAND U13358 ( .A(n11450), .B(nreg[142]), .Z(n6004) );
  NAND U13359 ( .A(n6107), .B(nreg[142]), .Z(n11450) );
  XOR U13360 ( .A(n11451), .B(n11452), .Z(n11445) );
  ANDN U13361 ( .A(n11453), .B(n6005), .Z(n11452) );
  XOR U13362 ( .A(n11454), .B(n11455), .Z(n6005) );
  IV U13363 ( .A(n11451), .Z(n11454) );
  XNOR U13364 ( .A(n6006), .B(n11451), .Z(n11453) );
  NAND U13365 ( .A(n11456), .B(nreg[141]), .Z(n6006) );
  NAND U13366 ( .A(n6107), .B(nreg[141]), .Z(n11456) );
  XOR U13367 ( .A(n11457), .B(n11458), .Z(n11451) );
  ANDN U13368 ( .A(n11459), .B(n6007), .Z(n11458) );
  XOR U13369 ( .A(n11460), .B(n11461), .Z(n6007) );
  IV U13370 ( .A(n11457), .Z(n11460) );
  XNOR U13371 ( .A(n6008), .B(n11457), .Z(n11459) );
  NAND U13372 ( .A(n11462), .B(nreg[140]), .Z(n6008) );
  NAND U13373 ( .A(n6107), .B(nreg[140]), .Z(n11462) );
  XOR U13374 ( .A(n11463), .B(n11464), .Z(n11457) );
  ANDN U13375 ( .A(n11465), .B(n6009), .Z(n11464) );
  XOR U13376 ( .A(n11466), .B(n11467), .Z(n6009) );
  IV U13377 ( .A(n11463), .Z(n11466) );
  XNOR U13378 ( .A(n6010), .B(n11463), .Z(n11465) );
  NAND U13379 ( .A(n11468), .B(nreg[139]), .Z(n6010) );
  NAND U13380 ( .A(n6107), .B(nreg[139]), .Z(n11468) );
  XOR U13381 ( .A(n11469), .B(n11470), .Z(n11463) );
  ANDN U13382 ( .A(n11471), .B(n6011), .Z(n11470) );
  XOR U13383 ( .A(n11472), .B(n11473), .Z(n6011) );
  IV U13384 ( .A(n11469), .Z(n11472) );
  XNOR U13385 ( .A(n6012), .B(n11469), .Z(n11471) );
  NAND U13386 ( .A(n11474), .B(nreg[138]), .Z(n6012) );
  NAND U13387 ( .A(n6107), .B(nreg[138]), .Z(n11474) );
  XOR U13388 ( .A(n11475), .B(n11476), .Z(n11469) );
  ANDN U13389 ( .A(n11477), .B(n6013), .Z(n11476) );
  XOR U13390 ( .A(n11478), .B(n11479), .Z(n6013) );
  IV U13391 ( .A(n11475), .Z(n11478) );
  XNOR U13392 ( .A(n6014), .B(n11475), .Z(n11477) );
  NAND U13393 ( .A(n11480), .B(nreg[137]), .Z(n6014) );
  NAND U13394 ( .A(n6107), .B(nreg[137]), .Z(n11480) );
  XOR U13395 ( .A(n11481), .B(n11482), .Z(n11475) );
  ANDN U13396 ( .A(n11483), .B(n6017), .Z(n11482) );
  XOR U13397 ( .A(n11484), .B(n11485), .Z(n6017) );
  IV U13398 ( .A(n11481), .Z(n11484) );
  XNOR U13399 ( .A(n6018), .B(n11481), .Z(n11483) );
  NAND U13400 ( .A(n11486), .B(nreg[136]), .Z(n6018) );
  NAND U13401 ( .A(n6107), .B(nreg[136]), .Z(n11486) );
  XOR U13402 ( .A(n11487), .B(n11488), .Z(n11481) );
  ANDN U13403 ( .A(n11489), .B(n6019), .Z(n11488) );
  XOR U13404 ( .A(n11490), .B(n11491), .Z(n6019) );
  IV U13405 ( .A(n11487), .Z(n11490) );
  XNOR U13406 ( .A(n6020), .B(n11487), .Z(n11489) );
  NAND U13407 ( .A(n11492), .B(nreg[135]), .Z(n6020) );
  NAND U13408 ( .A(n6107), .B(nreg[135]), .Z(n11492) );
  XOR U13409 ( .A(n11493), .B(n11494), .Z(n11487) );
  ANDN U13410 ( .A(n11495), .B(n6021), .Z(n11494) );
  XOR U13411 ( .A(n11496), .B(n11497), .Z(n6021) );
  IV U13412 ( .A(n11493), .Z(n11496) );
  XNOR U13413 ( .A(n6022), .B(n11493), .Z(n11495) );
  NAND U13414 ( .A(n11498), .B(nreg[134]), .Z(n6022) );
  NAND U13415 ( .A(n6107), .B(nreg[134]), .Z(n11498) );
  XOR U13416 ( .A(n11499), .B(n11500), .Z(n11493) );
  ANDN U13417 ( .A(n11501), .B(n6023), .Z(n11500) );
  XOR U13418 ( .A(n11502), .B(n11503), .Z(n6023) );
  IV U13419 ( .A(n11499), .Z(n11502) );
  XNOR U13420 ( .A(n6024), .B(n11499), .Z(n11501) );
  NAND U13421 ( .A(n11504), .B(nreg[133]), .Z(n6024) );
  NAND U13422 ( .A(n6107), .B(nreg[133]), .Z(n11504) );
  XOR U13423 ( .A(n11505), .B(n11506), .Z(n11499) );
  ANDN U13424 ( .A(n11507), .B(n6025), .Z(n11506) );
  XOR U13425 ( .A(n11508), .B(n11509), .Z(n6025) );
  IV U13426 ( .A(n11505), .Z(n11508) );
  XNOR U13427 ( .A(n6026), .B(n11505), .Z(n11507) );
  NAND U13428 ( .A(n11510), .B(nreg[132]), .Z(n6026) );
  NAND U13429 ( .A(n6107), .B(nreg[132]), .Z(n11510) );
  XOR U13430 ( .A(n11511), .B(n11512), .Z(n11505) );
  ANDN U13431 ( .A(n11513), .B(n6027), .Z(n11512) );
  XOR U13432 ( .A(n11514), .B(n11515), .Z(n6027) );
  IV U13433 ( .A(n11511), .Z(n11514) );
  XNOR U13434 ( .A(n6028), .B(n11511), .Z(n11513) );
  NAND U13435 ( .A(n11516), .B(nreg[131]), .Z(n6028) );
  NAND U13436 ( .A(n6107), .B(nreg[131]), .Z(n11516) );
  XOR U13437 ( .A(n11517), .B(n11518), .Z(n11511) );
  ANDN U13438 ( .A(n11519), .B(n6029), .Z(n11518) );
  XOR U13439 ( .A(n11520), .B(n11521), .Z(n6029) );
  IV U13440 ( .A(n11517), .Z(n11520) );
  XNOR U13441 ( .A(n6030), .B(n11517), .Z(n11519) );
  NAND U13442 ( .A(n11522), .B(nreg[130]), .Z(n6030) );
  NAND U13443 ( .A(n6107), .B(nreg[130]), .Z(n11522) );
  XOR U13444 ( .A(n11523), .B(n11524), .Z(n11517) );
  ANDN U13445 ( .A(n11525), .B(n6031), .Z(n11524) );
  XOR U13446 ( .A(n11526), .B(n11527), .Z(n6031) );
  IV U13447 ( .A(n11523), .Z(n11526) );
  XNOR U13448 ( .A(n6032), .B(n11523), .Z(n11525) );
  NAND U13449 ( .A(n11528), .B(nreg[129]), .Z(n6032) );
  NAND U13450 ( .A(n6107), .B(nreg[129]), .Z(n11528) );
  XOR U13451 ( .A(n11529), .B(n11530), .Z(n11523) );
  ANDN U13452 ( .A(n11531), .B(n6033), .Z(n11530) );
  XOR U13453 ( .A(n11532), .B(n11533), .Z(n6033) );
  IV U13454 ( .A(n11529), .Z(n11532) );
  XNOR U13455 ( .A(n6034), .B(n11529), .Z(n11531) );
  NAND U13456 ( .A(n11534), .B(nreg[128]), .Z(n6034) );
  NAND U13457 ( .A(n6107), .B(nreg[128]), .Z(n11534) );
  XOR U13458 ( .A(n11535), .B(n11536), .Z(n11529) );
  ANDN U13459 ( .A(n11537), .B(n6035), .Z(n11536) );
  XOR U13460 ( .A(n11538), .B(n11539), .Z(n6035) );
  IV U13461 ( .A(n11535), .Z(n11538) );
  XNOR U13462 ( .A(n6036), .B(n11535), .Z(n11537) );
  NAND U13463 ( .A(n11540), .B(nreg[127]), .Z(n6036) );
  NAND U13464 ( .A(n6107), .B(nreg[127]), .Z(n11540) );
  XOR U13465 ( .A(n11541), .B(n11542), .Z(n11535) );
  ANDN U13466 ( .A(n11543), .B(n6039), .Z(n11542) );
  XOR U13467 ( .A(n11544), .B(n11545), .Z(n6039) );
  IV U13468 ( .A(n11541), .Z(n11544) );
  XNOR U13469 ( .A(n6040), .B(n11541), .Z(n11543) );
  NAND U13470 ( .A(n11546), .B(nreg[126]), .Z(n6040) );
  NAND U13471 ( .A(n6107), .B(nreg[126]), .Z(n11546) );
  XOR U13472 ( .A(n11547), .B(n11548), .Z(n11541) );
  ANDN U13473 ( .A(n11549), .B(n6041), .Z(n11548) );
  XOR U13474 ( .A(n11550), .B(n11551), .Z(n6041) );
  IV U13475 ( .A(n11547), .Z(n11550) );
  XNOR U13476 ( .A(n6042), .B(n11547), .Z(n11549) );
  NAND U13477 ( .A(n11552), .B(nreg[125]), .Z(n6042) );
  NAND U13478 ( .A(n6107), .B(nreg[125]), .Z(n11552) );
  XOR U13479 ( .A(n11553), .B(n11554), .Z(n11547) );
  ANDN U13480 ( .A(n11555), .B(n6043), .Z(n11554) );
  XOR U13481 ( .A(n11556), .B(n11557), .Z(n6043) );
  IV U13482 ( .A(n11553), .Z(n11556) );
  XNOR U13483 ( .A(n6044), .B(n11553), .Z(n11555) );
  NAND U13484 ( .A(n11558), .B(nreg[124]), .Z(n6044) );
  NAND U13485 ( .A(n6107), .B(nreg[124]), .Z(n11558) );
  XOR U13486 ( .A(n11559), .B(n11560), .Z(n11553) );
  ANDN U13487 ( .A(n11561), .B(n6045), .Z(n11560) );
  XOR U13488 ( .A(n11562), .B(n11563), .Z(n6045) );
  IV U13489 ( .A(n11559), .Z(n11562) );
  XNOR U13490 ( .A(n6046), .B(n11559), .Z(n11561) );
  NAND U13491 ( .A(n11564), .B(nreg[123]), .Z(n6046) );
  NAND U13492 ( .A(n6107), .B(nreg[123]), .Z(n11564) );
  XOR U13493 ( .A(n11565), .B(n11566), .Z(n11559) );
  ANDN U13494 ( .A(n11567), .B(n6047), .Z(n11566) );
  XOR U13495 ( .A(n11568), .B(n11569), .Z(n6047) );
  IV U13496 ( .A(n11565), .Z(n11568) );
  XNOR U13497 ( .A(n6048), .B(n11565), .Z(n11567) );
  NAND U13498 ( .A(n11570), .B(nreg[122]), .Z(n6048) );
  NAND U13499 ( .A(n6107), .B(nreg[122]), .Z(n11570) );
  XOR U13500 ( .A(n11571), .B(n11572), .Z(n11565) );
  ANDN U13501 ( .A(n11573), .B(n6049), .Z(n11572) );
  XOR U13502 ( .A(n11574), .B(n11575), .Z(n6049) );
  IV U13503 ( .A(n11571), .Z(n11574) );
  XNOR U13504 ( .A(n6050), .B(n11571), .Z(n11573) );
  NAND U13505 ( .A(n11576), .B(nreg[121]), .Z(n6050) );
  NAND U13506 ( .A(n6107), .B(nreg[121]), .Z(n11576) );
  XOR U13507 ( .A(n11577), .B(n11578), .Z(n11571) );
  ANDN U13508 ( .A(n11579), .B(n6051), .Z(n11578) );
  XOR U13509 ( .A(n11580), .B(n11581), .Z(n6051) );
  IV U13510 ( .A(n11577), .Z(n11580) );
  XNOR U13511 ( .A(n6052), .B(n11577), .Z(n11579) );
  NAND U13512 ( .A(n11582), .B(nreg[120]), .Z(n6052) );
  NAND U13513 ( .A(n6107), .B(nreg[120]), .Z(n11582) );
  XOR U13514 ( .A(n11583), .B(n11584), .Z(n11577) );
  ANDN U13515 ( .A(n11585), .B(n6053), .Z(n11584) );
  XOR U13516 ( .A(n11586), .B(n11587), .Z(n6053) );
  IV U13517 ( .A(n11583), .Z(n11586) );
  XNOR U13518 ( .A(n6054), .B(n11583), .Z(n11585) );
  NAND U13519 ( .A(n11588), .B(nreg[119]), .Z(n6054) );
  NAND U13520 ( .A(n6107), .B(nreg[119]), .Z(n11588) );
  XOR U13521 ( .A(n11589), .B(n11590), .Z(n11583) );
  ANDN U13522 ( .A(n11591), .B(n6055), .Z(n11590) );
  XOR U13523 ( .A(n11592), .B(n11593), .Z(n6055) );
  IV U13524 ( .A(n11589), .Z(n11592) );
  XNOR U13525 ( .A(n6056), .B(n11589), .Z(n11591) );
  NAND U13526 ( .A(n11594), .B(nreg[118]), .Z(n6056) );
  NAND U13527 ( .A(n6107), .B(nreg[118]), .Z(n11594) );
  XOR U13528 ( .A(n11595), .B(n11596), .Z(n11589) );
  ANDN U13529 ( .A(n11597), .B(n6057), .Z(n11596) );
  XOR U13530 ( .A(n11598), .B(n11599), .Z(n6057) );
  IV U13531 ( .A(n11595), .Z(n11598) );
  XNOR U13532 ( .A(n6058), .B(n11595), .Z(n11597) );
  NAND U13533 ( .A(n11600), .B(nreg[117]), .Z(n6058) );
  NAND U13534 ( .A(n6107), .B(nreg[117]), .Z(n11600) );
  XOR U13535 ( .A(n11601), .B(n11602), .Z(n11595) );
  ANDN U13536 ( .A(n11603), .B(n6061), .Z(n11602) );
  XOR U13537 ( .A(n11604), .B(n11605), .Z(n6061) );
  IV U13538 ( .A(n11601), .Z(n11604) );
  XNOR U13539 ( .A(n6062), .B(n11601), .Z(n11603) );
  NAND U13540 ( .A(n11606), .B(nreg[116]), .Z(n6062) );
  NAND U13541 ( .A(n6107), .B(nreg[116]), .Z(n11606) );
  XOR U13542 ( .A(n11607), .B(n11608), .Z(n11601) );
  ANDN U13543 ( .A(n11609), .B(n6063), .Z(n11608) );
  XOR U13544 ( .A(n11610), .B(n11611), .Z(n6063) );
  IV U13545 ( .A(n11607), .Z(n11610) );
  XNOR U13546 ( .A(n6064), .B(n11607), .Z(n11609) );
  NAND U13547 ( .A(n11612), .B(nreg[115]), .Z(n6064) );
  NAND U13548 ( .A(n6107), .B(nreg[115]), .Z(n11612) );
  XOR U13549 ( .A(n11613), .B(n11614), .Z(n11607) );
  ANDN U13550 ( .A(n11615), .B(n6065), .Z(n11614) );
  XOR U13551 ( .A(n11616), .B(n11617), .Z(n6065) );
  IV U13552 ( .A(n11613), .Z(n11616) );
  XNOR U13553 ( .A(n6066), .B(n11613), .Z(n11615) );
  NAND U13554 ( .A(n11618), .B(nreg[114]), .Z(n6066) );
  NAND U13555 ( .A(n6107), .B(nreg[114]), .Z(n11618) );
  XOR U13556 ( .A(n11619), .B(n11620), .Z(n11613) );
  ANDN U13557 ( .A(n11621), .B(n6067), .Z(n11620) );
  XOR U13558 ( .A(n11622), .B(n11623), .Z(n6067) );
  IV U13559 ( .A(n11619), .Z(n11622) );
  XNOR U13560 ( .A(n6068), .B(n11619), .Z(n11621) );
  NAND U13561 ( .A(n11624), .B(nreg[113]), .Z(n6068) );
  NAND U13562 ( .A(n6107), .B(nreg[113]), .Z(n11624) );
  XOR U13563 ( .A(n11625), .B(n11626), .Z(n11619) );
  ANDN U13564 ( .A(n11627), .B(n6069), .Z(n11626) );
  XOR U13565 ( .A(n11628), .B(n11629), .Z(n6069) );
  IV U13566 ( .A(n11625), .Z(n11628) );
  XNOR U13567 ( .A(n6070), .B(n11625), .Z(n11627) );
  NAND U13568 ( .A(n11630), .B(nreg[112]), .Z(n6070) );
  NAND U13569 ( .A(n6107), .B(nreg[112]), .Z(n11630) );
  XOR U13570 ( .A(n11631), .B(n11632), .Z(n11625) );
  ANDN U13571 ( .A(n11633), .B(n6071), .Z(n11632) );
  XOR U13572 ( .A(n11634), .B(n11635), .Z(n6071) );
  IV U13573 ( .A(n11631), .Z(n11634) );
  XNOR U13574 ( .A(n6072), .B(n11631), .Z(n11633) );
  NAND U13575 ( .A(n11636), .B(nreg[111]), .Z(n6072) );
  NAND U13576 ( .A(n6107), .B(nreg[111]), .Z(n11636) );
  XOR U13577 ( .A(n11637), .B(n11638), .Z(n11631) );
  ANDN U13578 ( .A(n11639), .B(n6073), .Z(n11638) );
  XOR U13579 ( .A(n11640), .B(n11641), .Z(n6073) );
  IV U13580 ( .A(n11637), .Z(n11640) );
  XNOR U13581 ( .A(n6074), .B(n11637), .Z(n11639) );
  NAND U13582 ( .A(n11642), .B(nreg[110]), .Z(n6074) );
  NAND U13583 ( .A(n6107), .B(nreg[110]), .Z(n11642) );
  XOR U13584 ( .A(n11643), .B(n11644), .Z(n11637) );
  ANDN U13585 ( .A(n11645), .B(n6075), .Z(n11644) );
  XOR U13586 ( .A(n11646), .B(n11647), .Z(n6075) );
  IV U13587 ( .A(n11643), .Z(n11646) );
  XNOR U13588 ( .A(n6076), .B(n11643), .Z(n11645) );
  NAND U13589 ( .A(n11648), .B(nreg[109]), .Z(n6076) );
  NAND U13590 ( .A(n6107), .B(nreg[109]), .Z(n11648) );
  XOR U13591 ( .A(n11649), .B(n11650), .Z(n11643) );
  ANDN U13592 ( .A(n11651), .B(n6077), .Z(n11650) );
  XOR U13593 ( .A(n11652), .B(n11653), .Z(n6077) );
  IV U13594 ( .A(n11649), .Z(n11652) );
  XNOR U13595 ( .A(n6078), .B(n11649), .Z(n11651) );
  NAND U13596 ( .A(n11654), .B(nreg[108]), .Z(n6078) );
  NAND U13597 ( .A(n6107), .B(nreg[108]), .Z(n11654) );
  XOR U13598 ( .A(n11655), .B(n11656), .Z(n11649) );
  ANDN U13599 ( .A(n11657), .B(n6079), .Z(n11656) );
  XOR U13600 ( .A(n11658), .B(n11659), .Z(n6079) );
  IV U13601 ( .A(n11655), .Z(n11658) );
  XNOR U13602 ( .A(n6080), .B(n11655), .Z(n11657) );
  NAND U13603 ( .A(n11660), .B(nreg[107]), .Z(n6080) );
  NAND U13604 ( .A(n6107), .B(nreg[107]), .Z(n11660) );
  XOR U13605 ( .A(n11661), .B(n11662), .Z(n11655) );
  ANDN U13606 ( .A(n11663), .B(n6083), .Z(n11662) );
  XOR U13607 ( .A(n11664), .B(n11665), .Z(n6083) );
  IV U13608 ( .A(n11661), .Z(n11664) );
  XNOR U13609 ( .A(n6084), .B(n11661), .Z(n11663) );
  NAND U13610 ( .A(n11666), .B(nreg[106]), .Z(n6084) );
  NAND U13611 ( .A(n6107), .B(nreg[106]), .Z(n11666) );
  XOR U13612 ( .A(n11667), .B(n11668), .Z(n11661) );
  ANDN U13613 ( .A(n11669), .B(n6085), .Z(n11668) );
  XOR U13614 ( .A(n11670), .B(n11671), .Z(n6085) );
  IV U13615 ( .A(n11667), .Z(n11670) );
  XNOR U13616 ( .A(n6086), .B(n11667), .Z(n11669) );
  NAND U13617 ( .A(n11672), .B(nreg[105]), .Z(n6086) );
  NAND U13618 ( .A(n6107), .B(nreg[105]), .Z(n11672) );
  XOR U13619 ( .A(n11673), .B(n11674), .Z(n11667) );
  ANDN U13620 ( .A(n11675), .B(n6087), .Z(n11674) );
  XOR U13621 ( .A(n11676), .B(n11677), .Z(n6087) );
  IV U13622 ( .A(n11673), .Z(n11676) );
  XNOR U13623 ( .A(n6088), .B(n11673), .Z(n11675) );
  NAND U13624 ( .A(n11678), .B(nreg[104]), .Z(n6088) );
  NAND U13625 ( .A(n6107), .B(nreg[104]), .Z(n11678) );
  XOR U13626 ( .A(n11679), .B(n11680), .Z(n11673) );
  ANDN U13627 ( .A(n11681), .B(n6089), .Z(n11680) );
  XOR U13628 ( .A(n11682), .B(n11683), .Z(n6089) );
  IV U13629 ( .A(n11679), .Z(n11682) );
  XNOR U13630 ( .A(n6090), .B(n11679), .Z(n11681) );
  NAND U13631 ( .A(n11684), .B(nreg[103]), .Z(n6090) );
  NAND U13632 ( .A(n6107), .B(nreg[103]), .Z(n11684) );
  XOR U13633 ( .A(n11685), .B(n11686), .Z(n11679) );
  ANDN U13634 ( .A(n11687), .B(n6091), .Z(n11686) );
  XOR U13635 ( .A(n11688), .B(n11689), .Z(n6091) );
  IV U13636 ( .A(n11685), .Z(n11688) );
  XNOR U13637 ( .A(n6092), .B(n11685), .Z(n11687) );
  NAND U13638 ( .A(n11690), .B(nreg[102]), .Z(n6092) );
  NAND U13639 ( .A(n6107), .B(nreg[102]), .Z(n11690) );
  XOR U13640 ( .A(n11691), .B(n11692), .Z(n11685) );
  ANDN U13641 ( .A(n11693), .B(n6093), .Z(n11692) );
  XOR U13642 ( .A(n11694), .B(n11695), .Z(n6093) );
  IV U13643 ( .A(n11691), .Z(n11694) );
  XNOR U13644 ( .A(n6094), .B(n11691), .Z(n11693) );
  NAND U13645 ( .A(n11696), .B(nreg[101]), .Z(n6094) );
  NAND U13646 ( .A(n6107), .B(nreg[101]), .Z(n11696) );
  XOR U13647 ( .A(n11697), .B(n11698), .Z(n11691) );
  ANDN U13648 ( .A(n11699), .B(n6095), .Z(n11698) );
  XOR U13649 ( .A(n11700), .B(n11701), .Z(n6095) );
  IV U13650 ( .A(n11697), .Z(n11700) );
  XNOR U13651 ( .A(n6096), .B(n11697), .Z(n11699) );
  NAND U13652 ( .A(n11702), .B(nreg[100]), .Z(n6096) );
  NAND U13653 ( .A(n6107), .B(nreg[100]), .Z(n11702) );
  XOR U13654 ( .A(n11703), .B(n11704), .Z(n11697) );
  ANDN U13655 ( .A(n11705), .B(n6162), .Z(n11704) );
  XOR U13656 ( .A(n11706), .B(n11707), .Z(n6162) );
  IV U13657 ( .A(n11703), .Z(n11706) );
  XNOR U13658 ( .A(n6163), .B(n11703), .Z(n11705) );
  NAND U13659 ( .A(n11708), .B(nreg[99]), .Z(n6163) );
  NAND U13660 ( .A(n6107), .B(nreg[99]), .Z(n11708) );
  XOR U13661 ( .A(n11709), .B(n11710), .Z(n11703) );
  ANDN U13662 ( .A(n11711), .B(n6244), .Z(n11710) );
  XOR U13663 ( .A(n11712), .B(n11713), .Z(n6244) );
  IV U13664 ( .A(n11709), .Z(n11712) );
  XNOR U13665 ( .A(n6245), .B(n11709), .Z(n11711) );
  NAND U13666 ( .A(n11714), .B(nreg[98]), .Z(n6245) );
  NAND U13667 ( .A(n6107), .B(nreg[98]), .Z(n11714) );
  XOR U13668 ( .A(n11715), .B(n11716), .Z(n11709) );
  ANDN U13669 ( .A(n11717), .B(n11718), .Z(n11716) );
  XNOR U13670 ( .A(n11719), .B(n11715), .Z(n11717) );
  ANDN U13671 ( .A(n4110), .B(n1104), .Z(\modmult_1/N100 ) );
  XOR U13672 ( .A(n11718), .B(n11719), .Z(n1104) );
  NAND U13673 ( .A(n11720), .B(nreg[97]), .Z(n11719) );
  NAND U13674 ( .A(n6107), .B(nreg[97]), .Z(n11720) );
  XOR U13675 ( .A(n11721), .B(n11722), .Z(n11718) );
  IV U13676 ( .A(n11715), .Z(n11721) );
  XOR U13677 ( .A(n11723), .B(n11724), .Z(n11715) );
  ANDN U13678 ( .A(n11725), .B(n4131), .Z(n11724) );
  XOR U13679 ( .A(n11726), .B(n11727), .Z(n4131) );
  IV U13680 ( .A(n11723), .Z(n11726) );
  XNOR U13681 ( .A(n4132), .B(n11723), .Z(n11725) );
  NAND U13682 ( .A(n11728), .B(nreg[96]), .Z(n4132) );
  NAND U13683 ( .A(n6107), .B(nreg[96]), .Z(n11728) );
  XOR U13684 ( .A(n11729), .B(n11730), .Z(n11723) );
  ANDN U13685 ( .A(n11731), .B(n4153), .Z(n11730) );
  XOR U13686 ( .A(n11732), .B(n11733), .Z(n4153) );
  IV U13687 ( .A(n11729), .Z(n11732) );
  XNOR U13688 ( .A(n4154), .B(n11729), .Z(n11731) );
  NAND U13689 ( .A(n11734), .B(nreg[95]), .Z(n4154) );
  NAND U13690 ( .A(n6107), .B(nreg[95]), .Z(n11734) );
  XOR U13691 ( .A(n11735), .B(n11736), .Z(n11729) );
  ANDN U13692 ( .A(n11737), .B(n4175), .Z(n11736) );
  XOR U13693 ( .A(n11738), .B(n11739), .Z(n4175) );
  IV U13694 ( .A(n11735), .Z(n11738) );
  XNOR U13695 ( .A(n4176), .B(n11735), .Z(n11737) );
  NAND U13696 ( .A(n11740), .B(nreg[94]), .Z(n4176) );
  NAND U13697 ( .A(n6107), .B(nreg[94]), .Z(n11740) );
  XOR U13698 ( .A(n11741), .B(n11742), .Z(n11735) );
  ANDN U13699 ( .A(n11743), .B(n4197), .Z(n11742) );
  XOR U13700 ( .A(n11744), .B(n11745), .Z(n4197) );
  IV U13701 ( .A(n11741), .Z(n11744) );
  XNOR U13702 ( .A(n4198), .B(n11741), .Z(n11743) );
  NAND U13703 ( .A(n11746), .B(nreg[93]), .Z(n4198) );
  NAND U13704 ( .A(n6107), .B(nreg[93]), .Z(n11746) );
  XOR U13705 ( .A(n11747), .B(n11748), .Z(n11741) );
  ANDN U13706 ( .A(n11749), .B(n4219), .Z(n11748) );
  XOR U13707 ( .A(n11750), .B(n11751), .Z(n4219) );
  IV U13708 ( .A(n11747), .Z(n11750) );
  XNOR U13709 ( .A(n4220), .B(n11747), .Z(n11749) );
  NAND U13710 ( .A(n11752), .B(nreg[92]), .Z(n4220) );
  NAND U13711 ( .A(n6107), .B(nreg[92]), .Z(n11752) );
  XOR U13712 ( .A(n11753), .B(n11754), .Z(n11747) );
  ANDN U13713 ( .A(n11755), .B(n4241), .Z(n11754) );
  XOR U13714 ( .A(n11756), .B(n11757), .Z(n4241) );
  IV U13715 ( .A(n11753), .Z(n11756) );
  XNOR U13716 ( .A(n4242), .B(n11753), .Z(n11755) );
  NAND U13717 ( .A(n11758), .B(nreg[91]), .Z(n4242) );
  NAND U13718 ( .A(n6107), .B(nreg[91]), .Z(n11758) );
  XOR U13719 ( .A(n11759), .B(n11760), .Z(n11753) );
  ANDN U13720 ( .A(n11761), .B(n4263), .Z(n11760) );
  XOR U13721 ( .A(n11762), .B(n11763), .Z(n4263) );
  IV U13722 ( .A(n11759), .Z(n11762) );
  XNOR U13723 ( .A(n4264), .B(n11759), .Z(n11761) );
  NAND U13724 ( .A(n11764), .B(nreg[90]), .Z(n4264) );
  NAND U13725 ( .A(n6107), .B(nreg[90]), .Z(n11764) );
  XOR U13726 ( .A(n11765), .B(n11766), .Z(n11759) );
  ANDN U13727 ( .A(n11767), .B(n4285), .Z(n11766) );
  XOR U13728 ( .A(n11768), .B(n11769), .Z(n4285) );
  IV U13729 ( .A(n11765), .Z(n11768) );
  XNOR U13730 ( .A(n4286), .B(n11765), .Z(n11767) );
  NAND U13731 ( .A(n11770), .B(nreg[89]), .Z(n4286) );
  NAND U13732 ( .A(n6107), .B(nreg[89]), .Z(n11770) );
  XOR U13733 ( .A(n11771), .B(n11772), .Z(n11765) );
  ANDN U13734 ( .A(n11773), .B(n4307), .Z(n11772) );
  XOR U13735 ( .A(n11774), .B(n11775), .Z(n4307) );
  IV U13736 ( .A(n11771), .Z(n11774) );
  XNOR U13737 ( .A(n4308), .B(n11771), .Z(n11773) );
  NAND U13738 ( .A(n11776), .B(nreg[88]), .Z(n4308) );
  NAND U13739 ( .A(n6107), .B(nreg[88]), .Z(n11776) );
  XOR U13740 ( .A(n11777), .B(n11778), .Z(n11771) );
  ANDN U13741 ( .A(n11779), .B(n4329), .Z(n11778) );
  XOR U13742 ( .A(n11780), .B(n11781), .Z(n4329) );
  IV U13743 ( .A(n11777), .Z(n11780) );
  XNOR U13744 ( .A(n4330), .B(n11777), .Z(n11779) );
  NAND U13745 ( .A(n11782), .B(nreg[87]), .Z(n4330) );
  NAND U13746 ( .A(n6107), .B(nreg[87]), .Z(n11782) );
  XOR U13747 ( .A(n11783), .B(n11784), .Z(n11777) );
  ANDN U13748 ( .A(n11785), .B(n4353), .Z(n11784) );
  XOR U13749 ( .A(n11786), .B(n11787), .Z(n4353) );
  IV U13750 ( .A(n11783), .Z(n11786) );
  XNOR U13751 ( .A(n4354), .B(n11783), .Z(n11785) );
  NAND U13752 ( .A(n11788), .B(nreg[86]), .Z(n4354) );
  NAND U13753 ( .A(n6107), .B(nreg[86]), .Z(n11788) );
  XOR U13754 ( .A(n11789), .B(n11790), .Z(n11783) );
  ANDN U13755 ( .A(n11791), .B(n4375), .Z(n11790) );
  XOR U13756 ( .A(n11792), .B(n11793), .Z(n4375) );
  IV U13757 ( .A(n11789), .Z(n11792) );
  XNOR U13758 ( .A(n4376), .B(n11789), .Z(n11791) );
  NAND U13759 ( .A(n11794), .B(nreg[85]), .Z(n4376) );
  NAND U13760 ( .A(n6107), .B(nreg[85]), .Z(n11794) );
  XOR U13761 ( .A(n11795), .B(n11796), .Z(n11789) );
  ANDN U13762 ( .A(n11797), .B(n4397), .Z(n11796) );
  XOR U13763 ( .A(n11798), .B(n11799), .Z(n4397) );
  IV U13764 ( .A(n11795), .Z(n11798) );
  XNOR U13765 ( .A(n4398), .B(n11795), .Z(n11797) );
  NAND U13766 ( .A(n11800), .B(nreg[84]), .Z(n4398) );
  NAND U13767 ( .A(n6107), .B(nreg[84]), .Z(n11800) );
  XOR U13768 ( .A(n11801), .B(n11802), .Z(n11795) );
  ANDN U13769 ( .A(n11803), .B(n4419), .Z(n11802) );
  XOR U13770 ( .A(n11804), .B(n11805), .Z(n4419) );
  IV U13771 ( .A(n11801), .Z(n11804) );
  XNOR U13772 ( .A(n4420), .B(n11801), .Z(n11803) );
  NAND U13773 ( .A(n11806), .B(nreg[83]), .Z(n4420) );
  NAND U13774 ( .A(n6107), .B(nreg[83]), .Z(n11806) );
  XOR U13775 ( .A(n11807), .B(n11808), .Z(n11801) );
  ANDN U13776 ( .A(n11809), .B(n4441), .Z(n11808) );
  XOR U13777 ( .A(n11810), .B(n11811), .Z(n4441) );
  IV U13778 ( .A(n11807), .Z(n11810) );
  XNOR U13779 ( .A(n4442), .B(n11807), .Z(n11809) );
  NAND U13780 ( .A(n11812), .B(nreg[82]), .Z(n4442) );
  NAND U13781 ( .A(n6107), .B(nreg[82]), .Z(n11812) );
  XOR U13782 ( .A(n11813), .B(n11814), .Z(n11807) );
  ANDN U13783 ( .A(n11815), .B(n4463), .Z(n11814) );
  XOR U13784 ( .A(n11816), .B(n11817), .Z(n4463) );
  IV U13785 ( .A(n11813), .Z(n11816) );
  XNOR U13786 ( .A(n4464), .B(n11813), .Z(n11815) );
  NAND U13787 ( .A(n11818), .B(nreg[81]), .Z(n4464) );
  NAND U13788 ( .A(n6107), .B(nreg[81]), .Z(n11818) );
  XOR U13789 ( .A(n11819), .B(n11820), .Z(n11813) );
  ANDN U13790 ( .A(n11821), .B(n4485), .Z(n11820) );
  XOR U13791 ( .A(n11822), .B(n11823), .Z(n4485) );
  IV U13792 ( .A(n11819), .Z(n11822) );
  XNOR U13793 ( .A(n4486), .B(n11819), .Z(n11821) );
  NAND U13794 ( .A(n11824), .B(nreg[80]), .Z(n4486) );
  NAND U13795 ( .A(n6107), .B(nreg[80]), .Z(n11824) );
  XOR U13796 ( .A(n11825), .B(n11826), .Z(n11819) );
  ANDN U13797 ( .A(n11827), .B(n4507), .Z(n11826) );
  XOR U13798 ( .A(n11828), .B(n11829), .Z(n4507) );
  IV U13799 ( .A(n11825), .Z(n11828) );
  XNOR U13800 ( .A(n4508), .B(n11825), .Z(n11827) );
  NAND U13801 ( .A(n11830), .B(nreg[79]), .Z(n4508) );
  NAND U13802 ( .A(n6107), .B(nreg[79]), .Z(n11830) );
  XOR U13803 ( .A(n11831), .B(n11832), .Z(n11825) );
  ANDN U13804 ( .A(n11833), .B(n4529), .Z(n11832) );
  XOR U13805 ( .A(n11834), .B(n11835), .Z(n4529) );
  IV U13806 ( .A(n11831), .Z(n11834) );
  XNOR U13807 ( .A(n4530), .B(n11831), .Z(n11833) );
  NAND U13808 ( .A(n11836), .B(nreg[78]), .Z(n4530) );
  NAND U13809 ( .A(n6107), .B(nreg[78]), .Z(n11836) );
  XOR U13810 ( .A(n11837), .B(n11838), .Z(n11831) );
  ANDN U13811 ( .A(n11839), .B(n4551), .Z(n11838) );
  XOR U13812 ( .A(n11840), .B(n11841), .Z(n4551) );
  IV U13813 ( .A(n11837), .Z(n11840) );
  XNOR U13814 ( .A(n4552), .B(n11837), .Z(n11839) );
  NAND U13815 ( .A(n11842), .B(nreg[77]), .Z(n4552) );
  NAND U13816 ( .A(n6107), .B(nreg[77]), .Z(n11842) );
  XOR U13817 ( .A(n11843), .B(n11844), .Z(n11837) );
  ANDN U13818 ( .A(n11845), .B(n4575), .Z(n11844) );
  XOR U13819 ( .A(n11846), .B(n11847), .Z(n4575) );
  IV U13820 ( .A(n11843), .Z(n11846) );
  XNOR U13821 ( .A(n4576), .B(n11843), .Z(n11845) );
  NAND U13822 ( .A(n11848), .B(nreg[76]), .Z(n4576) );
  NAND U13823 ( .A(n6107), .B(nreg[76]), .Z(n11848) );
  XOR U13824 ( .A(n11849), .B(n11850), .Z(n11843) );
  ANDN U13825 ( .A(n11851), .B(n4597), .Z(n11850) );
  XOR U13826 ( .A(n11852), .B(n11853), .Z(n4597) );
  IV U13827 ( .A(n11849), .Z(n11852) );
  XNOR U13828 ( .A(n4598), .B(n11849), .Z(n11851) );
  NAND U13829 ( .A(n11854), .B(nreg[75]), .Z(n4598) );
  NAND U13830 ( .A(n6107), .B(nreg[75]), .Z(n11854) );
  XOR U13831 ( .A(n11855), .B(n11856), .Z(n11849) );
  ANDN U13832 ( .A(n11857), .B(n4619), .Z(n11856) );
  XOR U13833 ( .A(n11858), .B(n11859), .Z(n4619) );
  IV U13834 ( .A(n11855), .Z(n11858) );
  XNOR U13835 ( .A(n4620), .B(n11855), .Z(n11857) );
  NAND U13836 ( .A(n11860), .B(nreg[74]), .Z(n4620) );
  NAND U13837 ( .A(n6107), .B(nreg[74]), .Z(n11860) );
  XOR U13838 ( .A(n11861), .B(n11862), .Z(n11855) );
  ANDN U13839 ( .A(n11863), .B(n4641), .Z(n11862) );
  XOR U13840 ( .A(n11864), .B(n11865), .Z(n4641) );
  IV U13841 ( .A(n11861), .Z(n11864) );
  XNOR U13842 ( .A(n4642), .B(n11861), .Z(n11863) );
  NAND U13843 ( .A(n11866), .B(nreg[73]), .Z(n4642) );
  NAND U13844 ( .A(n6107), .B(nreg[73]), .Z(n11866) );
  XOR U13845 ( .A(n11867), .B(n11868), .Z(n11861) );
  ANDN U13846 ( .A(n11869), .B(n4663), .Z(n11868) );
  XOR U13847 ( .A(n11870), .B(n11871), .Z(n4663) );
  IV U13848 ( .A(n11867), .Z(n11870) );
  XNOR U13849 ( .A(n4664), .B(n11867), .Z(n11869) );
  NAND U13850 ( .A(n11872), .B(nreg[72]), .Z(n4664) );
  NAND U13851 ( .A(n6107), .B(nreg[72]), .Z(n11872) );
  XOR U13852 ( .A(n11873), .B(n11874), .Z(n11867) );
  ANDN U13853 ( .A(n11875), .B(n4685), .Z(n11874) );
  XOR U13854 ( .A(n11876), .B(n11877), .Z(n4685) );
  IV U13855 ( .A(n11873), .Z(n11876) );
  XNOR U13856 ( .A(n4686), .B(n11873), .Z(n11875) );
  NAND U13857 ( .A(n11878), .B(nreg[71]), .Z(n4686) );
  NAND U13858 ( .A(n6107), .B(nreg[71]), .Z(n11878) );
  XOR U13859 ( .A(n11879), .B(n11880), .Z(n11873) );
  ANDN U13860 ( .A(n11881), .B(n4707), .Z(n11880) );
  XOR U13861 ( .A(n11882), .B(n11883), .Z(n4707) );
  IV U13862 ( .A(n11879), .Z(n11882) );
  XNOR U13863 ( .A(n4708), .B(n11879), .Z(n11881) );
  NAND U13864 ( .A(n11884), .B(nreg[70]), .Z(n4708) );
  NAND U13865 ( .A(n6107), .B(nreg[70]), .Z(n11884) );
  XOR U13866 ( .A(n11885), .B(n11886), .Z(n11879) );
  ANDN U13867 ( .A(n11887), .B(n4729), .Z(n11886) );
  XOR U13868 ( .A(n11888), .B(n11889), .Z(n4729) );
  IV U13869 ( .A(n11885), .Z(n11888) );
  XNOR U13870 ( .A(n4730), .B(n11885), .Z(n11887) );
  NAND U13871 ( .A(n11890), .B(nreg[69]), .Z(n4730) );
  NAND U13872 ( .A(n6107), .B(nreg[69]), .Z(n11890) );
  XOR U13873 ( .A(n11891), .B(n11892), .Z(n11885) );
  ANDN U13874 ( .A(n11893), .B(n4751), .Z(n11892) );
  XOR U13875 ( .A(n11894), .B(n11895), .Z(n4751) );
  IV U13876 ( .A(n11891), .Z(n11894) );
  XNOR U13877 ( .A(n4752), .B(n11891), .Z(n11893) );
  NAND U13878 ( .A(n11896), .B(nreg[68]), .Z(n4752) );
  NAND U13879 ( .A(n6107), .B(nreg[68]), .Z(n11896) );
  XOR U13880 ( .A(n11897), .B(n11898), .Z(n11891) );
  ANDN U13881 ( .A(n11899), .B(n4773), .Z(n11898) );
  XOR U13882 ( .A(n11900), .B(n11901), .Z(n4773) );
  IV U13883 ( .A(n11897), .Z(n11900) );
  XNOR U13884 ( .A(n4774), .B(n11897), .Z(n11899) );
  NAND U13885 ( .A(n11902), .B(nreg[67]), .Z(n4774) );
  NAND U13886 ( .A(n6107), .B(nreg[67]), .Z(n11902) );
  XOR U13887 ( .A(n11903), .B(n11904), .Z(n11897) );
  ANDN U13888 ( .A(n11905), .B(n4797), .Z(n11904) );
  XOR U13889 ( .A(n11906), .B(n11907), .Z(n4797) );
  IV U13890 ( .A(n11903), .Z(n11906) );
  XNOR U13891 ( .A(n4798), .B(n11903), .Z(n11905) );
  NAND U13892 ( .A(n11908), .B(nreg[66]), .Z(n4798) );
  NAND U13893 ( .A(n6107), .B(nreg[66]), .Z(n11908) );
  XOR U13894 ( .A(n11909), .B(n11910), .Z(n11903) );
  ANDN U13895 ( .A(n11911), .B(n4819), .Z(n11910) );
  XOR U13896 ( .A(n11912), .B(n11913), .Z(n4819) );
  IV U13897 ( .A(n11909), .Z(n11912) );
  XNOR U13898 ( .A(n4820), .B(n11909), .Z(n11911) );
  NAND U13899 ( .A(n11914), .B(nreg[65]), .Z(n4820) );
  NAND U13900 ( .A(n6107), .B(nreg[65]), .Z(n11914) );
  XOR U13901 ( .A(n11915), .B(n11916), .Z(n11909) );
  ANDN U13902 ( .A(n11917), .B(n4841), .Z(n11916) );
  XOR U13903 ( .A(n11918), .B(n11919), .Z(n4841) );
  IV U13904 ( .A(n11915), .Z(n11918) );
  XNOR U13905 ( .A(n4842), .B(n11915), .Z(n11917) );
  NAND U13906 ( .A(n11920), .B(nreg[64]), .Z(n4842) );
  NAND U13907 ( .A(n6107), .B(nreg[64]), .Z(n11920) );
  XOR U13908 ( .A(n11921), .B(n11922), .Z(n11915) );
  ANDN U13909 ( .A(n11923), .B(n4863), .Z(n11922) );
  XOR U13910 ( .A(n11924), .B(n11925), .Z(n4863) );
  IV U13911 ( .A(n11921), .Z(n11924) );
  XNOR U13912 ( .A(n4864), .B(n11921), .Z(n11923) );
  NAND U13913 ( .A(n11926), .B(nreg[63]), .Z(n4864) );
  NAND U13914 ( .A(n6107), .B(nreg[63]), .Z(n11926) );
  XOR U13915 ( .A(n11927), .B(n11928), .Z(n11921) );
  ANDN U13916 ( .A(n11929), .B(n4885), .Z(n11928) );
  XOR U13917 ( .A(n11930), .B(n11931), .Z(n4885) );
  IV U13918 ( .A(n11927), .Z(n11930) );
  XNOR U13919 ( .A(n4886), .B(n11927), .Z(n11929) );
  NAND U13920 ( .A(n11932), .B(nreg[62]), .Z(n4886) );
  NAND U13921 ( .A(n6107), .B(nreg[62]), .Z(n11932) );
  XOR U13922 ( .A(n11933), .B(n11934), .Z(n11927) );
  ANDN U13923 ( .A(n11935), .B(n4907), .Z(n11934) );
  XOR U13924 ( .A(n11936), .B(n11937), .Z(n4907) );
  IV U13925 ( .A(n11933), .Z(n11936) );
  XNOR U13926 ( .A(n4908), .B(n11933), .Z(n11935) );
  NAND U13927 ( .A(n11938), .B(nreg[61]), .Z(n4908) );
  NAND U13928 ( .A(n6107), .B(nreg[61]), .Z(n11938) );
  XOR U13929 ( .A(n11939), .B(n11940), .Z(n11933) );
  ANDN U13930 ( .A(n11941), .B(n4929), .Z(n11940) );
  XOR U13931 ( .A(n11942), .B(n11943), .Z(n4929) );
  IV U13932 ( .A(n11939), .Z(n11942) );
  XNOR U13933 ( .A(n4930), .B(n11939), .Z(n11941) );
  NAND U13934 ( .A(n11944), .B(nreg[60]), .Z(n4930) );
  NAND U13935 ( .A(n6107), .B(nreg[60]), .Z(n11944) );
  XOR U13936 ( .A(n11945), .B(n11946), .Z(n11939) );
  ANDN U13937 ( .A(n11947), .B(n4951), .Z(n11946) );
  XOR U13938 ( .A(n11948), .B(n11949), .Z(n4951) );
  IV U13939 ( .A(n11945), .Z(n11948) );
  XNOR U13940 ( .A(n4952), .B(n11945), .Z(n11947) );
  NAND U13941 ( .A(n11950), .B(nreg[59]), .Z(n4952) );
  NAND U13942 ( .A(n6107), .B(nreg[59]), .Z(n11950) );
  XOR U13943 ( .A(n11951), .B(n11952), .Z(n11945) );
  ANDN U13944 ( .A(n11953), .B(n4973), .Z(n11952) );
  XOR U13945 ( .A(n11954), .B(n11955), .Z(n4973) );
  IV U13946 ( .A(n11951), .Z(n11954) );
  XNOR U13947 ( .A(n4974), .B(n11951), .Z(n11953) );
  NAND U13948 ( .A(n11956), .B(nreg[58]), .Z(n4974) );
  NAND U13949 ( .A(n6107), .B(nreg[58]), .Z(n11956) );
  XOR U13950 ( .A(n11957), .B(n11958), .Z(n11951) );
  ANDN U13951 ( .A(n11959), .B(n4995), .Z(n11958) );
  XOR U13952 ( .A(n11960), .B(n11961), .Z(n4995) );
  IV U13953 ( .A(n11957), .Z(n11960) );
  XNOR U13954 ( .A(n4996), .B(n11957), .Z(n11959) );
  NAND U13955 ( .A(n11962), .B(nreg[57]), .Z(n4996) );
  NAND U13956 ( .A(n6107), .B(nreg[57]), .Z(n11962) );
  XOR U13957 ( .A(n11963), .B(n11964), .Z(n11957) );
  ANDN U13958 ( .A(n11965), .B(n5019), .Z(n11964) );
  XOR U13959 ( .A(n11966), .B(n11967), .Z(n5019) );
  IV U13960 ( .A(n11963), .Z(n11966) );
  XNOR U13961 ( .A(n5020), .B(n11963), .Z(n11965) );
  NAND U13962 ( .A(n11968), .B(nreg[56]), .Z(n5020) );
  NAND U13963 ( .A(n6107), .B(nreg[56]), .Z(n11968) );
  XOR U13964 ( .A(n11969), .B(n11970), .Z(n11963) );
  ANDN U13965 ( .A(n11971), .B(n5041), .Z(n11970) );
  XOR U13966 ( .A(n11972), .B(n11973), .Z(n5041) );
  IV U13967 ( .A(n11969), .Z(n11972) );
  XNOR U13968 ( .A(n5042), .B(n11969), .Z(n11971) );
  NAND U13969 ( .A(n11974), .B(nreg[55]), .Z(n5042) );
  NAND U13970 ( .A(n6107), .B(nreg[55]), .Z(n11974) );
  XOR U13971 ( .A(n11975), .B(n11976), .Z(n11969) );
  ANDN U13972 ( .A(n11977), .B(n5063), .Z(n11976) );
  XOR U13973 ( .A(n11978), .B(n11979), .Z(n5063) );
  IV U13974 ( .A(n11975), .Z(n11978) );
  XNOR U13975 ( .A(n5064), .B(n11975), .Z(n11977) );
  NAND U13976 ( .A(n11980), .B(nreg[54]), .Z(n5064) );
  NAND U13977 ( .A(n6107), .B(nreg[54]), .Z(n11980) );
  XOR U13978 ( .A(n11981), .B(n11982), .Z(n11975) );
  ANDN U13979 ( .A(n11983), .B(n5085), .Z(n11982) );
  XOR U13980 ( .A(n11984), .B(n11985), .Z(n5085) );
  IV U13981 ( .A(n11981), .Z(n11984) );
  XNOR U13982 ( .A(n5086), .B(n11981), .Z(n11983) );
  NAND U13983 ( .A(n11986), .B(nreg[53]), .Z(n5086) );
  NAND U13984 ( .A(n6107), .B(nreg[53]), .Z(n11986) );
  XOR U13985 ( .A(n11987), .B(n11988), .Z(n11981) );
  ANDN U13986 ( .A(n11989), .B(n5107), .Z(n11988) );
  XOR U13987 ( .A(n11990), .B(n11991), .Z(n5107) );
  IV U13988 ( .A(n11987), .Z(n11990) );
  XNOR U13989 ( .A(n5108), .B(n11987), .Z(n11989) );
  NAND U13990 ( .A(n11992), .B(nreg[52]), .Z(n5108) );
  NAND U13991 ( .A(n6107), .B(nreg[52]), .Z(n11992) );
  XOR U13992 ( .A(n11993), .B(n11994), .Z(n11987) );
  ANDN U13993 ( .A(n11995), .B(n5129), .Z(n11994) );
  XOR U13994 ( .A(n11996), .B(n11997), .Z(n5129) );
  IV U13995 ( .A(n11993), .Z(n11996) );
  XNOR U13996 ( .A(n5130), .B(n11993), .Z(n11995) );
  NAND U13997 ( .A(n11998), .B(nreg[51]), .Z(n5130) );
  NAND U13998 ( .A(n6107), .B(nreg[51]), .Z(n11998) );
  XOR U13999 ( .A(n11999), .B(n12000), .Z(n11993) );
  ANDN U14000 ( .A(n12001), .B(n5151), .Z(n12000) );
  XOR U14001 ( .A(n12002), .B(n12003), .Z(n5151) );
  IV U14002 ( .A(n11999), .Z(n12002) );
  XNOR U14003 ( .A(n5152), .B(n11999), .Z(n12001) );
  NAND U14004 ( .A(n12004), .B(nreg[50]), .Z(n5152) );
  NAND U14005 ( .A(n6107), .B(nreg[50]), .Z(n12004) );
  XOR U14006 ( .A(n12005), .B(n12006), .Z(n11999) );
  ANDN U14007 ( .A(n12007), .B(n5173), .Z(n12006) );
  XOR U14008 ( .A(n12008), .B(n12009), .Z(n5173) );
  IV U14009 ( .A(n12005), .Z(n12008) );
  XNOR U14010 ( .A(n5174), .B(n12005), .Z(n12007) );
  NAND U14011 ( .A(n12010), .B(nreg[49]), .Z(n5174) );
  NAND U14012 ( .A(n6107), .B(nreg[49]), .Z(n12010) );
  XOR U14013 ( .A(n12011), .B(n12012), .Z(n12005) );
  ANDN U14014 ( .A(n12013), .B(n5195), .Z(n12012) );
  XOR U14015 ( .A(n12014), .B(n12015), .Z(n5195) );
  IV U14016 ( .A(n12011), .Z(n12014) );
  XNOR U14017 ( .A(n5196), .B(n12011), .Z(n12013) );
  NAND U14018 ( .A(n12016), .B(nreg[48]), .Z(n5196) );
  NAND U14019 ( .A(n6107), .B(nreg[48]), .Z(n12016) );
  XOR U14020 ( .A(n12017), .B(n12018), .Z(n12011) );
  ANDN U14021 ( .A(n12019), .B(n5217), .Z(n12018) );
  XOR U14022 ( .A(n12020), .B(n12021), .Z(n5217) );
  IV U14023 ( .A(n12017), .Z(n12020) );
  XNOR U14024 ( .A(n5218), .B(n12017), .Z(n12019) );
  NAND U14025 ( .A(n12022), .B(nreg[47]), .Z(n5218) );
  NAND U14026 ( .A(n6107), .B(nreg[47]), .Z(n12022) );
  XOR U14027 ( .A(n12023), .B(n12024), .Z(n12017) );
  ANDN U14028 ( .A(n12025), .B(n5241), .Z(n12024) );
  XOR U14029 ( .A(n12026), .B(n12027), .Z(n5241) );
  IV U14030 ( .A(n12023), .Z(n12026) );
  XNOR U14031 ( .A(n5242), .B(n12023), .Z(n12025) );
  NAND U14032 ( .A(n12028), .B(nreg[46]), .Z(n5242) );
  NAND U14033 ( .A(n6107), .B(nreg[46]), .Z(n12028) );
  XOR U14034 ( .A(n12029), .B(n12030), .Z(n12023) );
  ANDN U14035 ( .A(n12031), .B(n5263), .Z(n12030) );
  XOR U14036 ( .A(n12032), .B(n12033), .Z(n5263) );
  IV U14037 ( .A(n12029), .Z(n12032) );
  XNOR U14038 ( .A(n5264), .B(n12029), .Z(n12031) );
  NAND U14039 ( .A(n12034), .B(nreg[45]), .Z(n5264) );
  NAND U14040 ( .A(n6107), .B(nreg[45]), .Z(n12034) );
  XOR U14041 ( .A(n12035), .B(n12036), .Z(n12029) );
  ANDN U14042 ( .A(n12037), .B(n5285), .Z(n12036) );
  XOR U14043 ( .A(n12038), .B(n12039), .Z(n5285) );
  IV U14044 ( .A(n12035), .Z(n12038) );
  XNOR U14045 ( .A(n5286), .B(n12035), .Z(n12037) );
  NAND U14046 ( .A(n12040), .B(nreg[44]), .Z(n5286) );
  NAND U14047 ( .A(n6107), .B(nreg[44]), .Z(n12040) );
  XOR U14048 ( .A(n12041), .B(n12042), .Z(n12035) );
  ANDN U14049 ( .A(n12043), .B(n5307), .Z(n12042) );
  XOR U14050 ( .A(n12044), .B(n12045), .Z(n5307) );
  IV U14051 ( .A(n12041), .Z(n12044) );
  XNOR U14052 ( .A(n5308), .B(n12041), .Z(n12043) );
  NAND U14053 ( .A(n12046), .B(nreg[43]), .Z(n5308) );
  NAND U14054 ( .A(n6107), .B(nreg[43]), .Z(n12046) );
  XOR U14055 ( .A(n12047), .B(n12048), .Z(n12041) );
  ANDN U14056 ( .A(n12049), .B(n5329), .Z(n12048) );
  XOR U14057 ( .A(n12050), .B(n12051), .Z(n5329) );
  IV U14058 ( .A(n12047), .Z(n12050) );
  XNOR U14059 ( .A(n5330), .B(n12047), .Z(n12049) );
  NAND U14060 ( .A(n12052), .B(nreg[42]), .Z(n5330) );
  NAND U14061 ( .A(n6107), .B(nreg[42]), .Z(n12052) );
  XOR U14062 ( .A(n12053), .B(n12054), .Z(n12047) );
  ANDN U14063 ( .A(n12055), .B(n5351), .Z(n12054) );
  XOR U14064 ( .A(n12056), .B(n12057), .Z(n5351) );
  IV U14065 ( .A(n12053), .Z(n12056) );
  XNOR U14066 ( .A(n5352), .B(n12053), .Z(n12055) );
  NAND U14067 ( .A(n12058), .B(nreg[41]), .Z(n5352) );
  NAND U14068 ( .A(n6107), .B(nreg[41]), .Z(n12058) );
  XOR U14069 ( .A(n12059), .B(n12060), .Z(n12053) );
  ANDN U14070 ( .A(n12061), .B(n5373), .Z(n12060) );
  XOR U14071 ( .A(n12062), .B(n12063), .Z(n5373) );
  IV U14072 ( .A(n12059), .Z(n12062) );
  XNOR U14073 ( .A(n5374), .B(n12059), .Z(n12061) );
  NAND U14074 ( .A(n12064), .B(nreg[40]), .Z(n5374) );
  NAND U14075 ( .A(n6107), .B(nreg[40]), .Z(n12064) );
  XOR U14076 ( .A(n12065), .B(n12066), .Z(n12059) );
  ANDN U14077 ( .A(n12067), .B(n5395), .Z(n12066) );
  XOR U14078 ( .A(n12068), .B(n12069), .Z(n5395) );
  IV U14079 ( .A(n12065), .Z(n12068) );
  XNOR U14080 ( .A(n5396), .B(n12065), .Z(n12067) );
  NAND U14081 ( .A(n12070), .B(nreg[39]), .Z(n5396) );
  NAND U14082 ( .A(n6107), .B(nreg[39]), .Z(n12070) );
  XOR U14083 ( .A(n12071), .B(n12072), .Z(n12065) );
  ANDN U14084 ( .A(n12073), .B(n5417), .Z(n12072) );
  XOR U14085 ( .A(n12074), .B(n12075), .Z(n5417) );
  IV U14086 ( .A(n12071), .Z(n12074) );
  XNOR U14087 ( .A(n5418), .B(n12071), .Z(n12073) );
  NAND U14088 ( .A(n12076), .B(nreg[38]), .Z(n5418) );
  NAND U14089 ( .A(n6107), .B(nreg[38]), .Z(n12076) );
  XOR U14090 ( .A(n12077), .B(n12078), .Z(n12071) );
  ANDN U14091 ( .A(n12079), .B(n5439), .Z(n12078) );
  XOR U14092 ( .A(n12080), .B(n12081), .Z(n5439) );
  IV U14093 ( .A(n12077), .Z(n12080) );
  XNOR U14094 ( .A(n5440), .B(n12077), .Z(n12079) );
  NAND U14095 ( .A(n12082), .B(nreg[37]), .Z(n5440) );
  NAND U14096 ( .A(n6107), .B(nreg[37]), .Z(n12082) );
  XOR U14097 ( .A(n12083), .B(n12084), .Z(n12077) );
  ANDN U14098 ( .A(n12085), .B(n5463), .Z(n12084) );
  XOR U14099 ( .A(n12086), .B(n12087), .Z(n5463) );
  IV U14100 ( .A(n12083), .Z(n12086) );
  XNOR U14101 ( .A(n5464), .B(n12083), .Z(n12085) );
  NAND U14102 ( .A(n12088), .B(nreg[36]), .Z(n5464) );
  NAND U14103 ( .A(n6107), .B(nreg[36]), .Z(n12088) );
  XOR U14104 ( .A(n12089), .B(n12090), .Z(n12083) );
  ANDN U14105 ( .A(n12091), .B(n5485), .Z(n12090) );
  XOR U14106 ( .A(n12092), .B(n12093), .Z(n5485) );
  IV U14107 ( .A(n12089), .Z(n12092) );
  XNOR U14108 ( .A(n5486), .B(n12089), .Z(n12091) );
  NAND U14109 ( .A(n12094), .B(nreg[35]), .Z(n5486) );
  NAND U14110 ( .A(n6107), .B(nreg[35]), .Z(n12094) );
  XOR U14111 ( .A(n12095), .B(n12096), .Z(n12089) );
  ANDN U14112 ( .A(n12097), .B(n5507), .Z(n12096) );
  XOR U14113 ( .A(n12098), .B(n12099), .Z(n5507) );
  IV U14114 ( .A(n12095), .Z(n12098) );
  XNOR U14115 ( .A(n5508), .B(n12095), .Z(n12097) );
  NAND U14116 ( .A(n12100), .B(nreg[34]), .Z(n5508) );
  NAND U14117 ( .A(n6107), .B(nreg[34]), .Z(n12100) );
  XOR U14118 ( .A(n12101), .B(n12102), .Z(n12095) );
  ANDN U14119 ( .A(n12103), .B(n5529), .Z(n12102) );
  XOR U14120 ( .A(n12104), .B(n12105), .Z(n5529) );
  IV U14121 ( .A(n12101), .Z(n12104) );
  XNOR U14122 ( .A(n5530), .B(n12101), .Z(n12103) );
  NAND U14123 ( .A(n12106), .B(nreg[33]), .Z(n5530) );
  NAND U14124 ( .A(n6107), .B(nreg[33]), .Z(n12106) );
  XOR U14125 ( .A(n12107), .B(n12108), .Z(n12101) );
  ANDN U14126 ( .A(n12109), .B(n5551), .Z(n12108) );
  XOR U14127 ( .A(n12110), .B(n12111), .Z(n5551) );
  IV U14128 ( .A(n12107), .Z(n12110) );
  XNOR U14129 ( .A(n5552), .B(n12107), .Z(n12109) );
  NAND U14130 ( .A(n12112), .B(nreg[32]), .Z(n5552) );
  NAND U14131 ( .A(n6107), .B(nreg[32]), .Z(n12112) );
  XOR U14132 ( .A(n12113), .B(n12114), .Z(n12107) );
  ANDN U14133 ( .A(n12115), .B(n5573), .Z(n12114) );
  XOR U14134 ( .A(n12116), .B(n12117), .Z(n5573) );
  IV U14135 ( .A(n12113), .Z(n12116) );
  XNOR U14136 ( .A(n5574), .B(n12113), .Z(n12115) );
  NAND U14137 ( .A(n12118), .B(nreg[31]), .Z(n5574) );
  NAND U14138 ( .A(n6107), .B(nreg[31]), .Z(n12118) );
  XOR U14139 ( .A(n12119), .B(n12120), .Z(n12113) );
  ANDN U14140 ( .A(n12121), .B(n5595), .Z(n12120) );
  XOR U14141 ( .A(n12122), .B(n12123), .Z(n5595) );
  IV U14142 ( .A(n12119), .Z(n12122) );
  XNOR U14143 ( .A(n5596), .B(n12119), .Z(n12121) );
  NAND U14144 ( .A(n12124), .B(nreg[30]), .Z(n5596) );
  NAND U14145 ( .A(n6107), .B(nreg[30]), .Z(n12124) );
  XOR U14146 ( .A(n12125), .B(n12126), .Z(n12119) );
  ANDN U14147 ( .A(n12127), .B(n5617), .Z(n12126) );
  XOR U14148 ( .A(n12128), .B(n12129), .Z(n5617) );
  IV U14149 ( .A(n12125), .Z(n12128) );
  XNOR U14150 ( .A(n5618), .B(n12125), .Z(n12127) );
  NAND U14151 ( .A(n12130), .B(nreg[29]), .Z(n5618) );
  NAND U14152 ( .A(n6107), .B(nreg[29]), .Z(n12130) );
  XOR U14153 ( .A(n12131), .B(n12132), .Z(n12125) );
  ANDN U14154 ( .A(n12133), .B(n5639), .Z(n12132) );
  XOR U14155 ( .A(n12134), .B(n12135), .Z(n5639) );
  IV U14156 ( .A(n12131), .Z(n12134) );
  XNOR U14157 ( .A(n5640), .B(n12131), .Z(n12133) );
  NAND U14158 ( .A(n12136), .B(nreg[28]), .Z(n5640) );
  NAND U14159 ( .A(n6107), .B(nreg[28]), .Z(n12136) );
  XOR U14160 ( .A(n12137), .B(n12138), .Z(n12131) );
  ANDN U14161 ( .A(n12139), .B(n5661), .Z(n12138) );
  XOR U14162 ( .A(n12140), .B(n12141), .Z(n5661) );
  IV U14163 ( .A(n12137), .Z(n12140) );
  XNOR U14164 ( .A(n5662), .B(n12137), .Z(n12139) );
  NAND U14165 ( .A(n12142), .B(nreg[27]), .Z(n5662) );
  NAND U14166 ( .A(n6107), .B(nreg[27]), .Z(n12142) );
  XOR U14167 ( .A(n12143), .B(n12144), .Z(n12137) );
  ANDN U14168 ( .A(n12145), .B(n5685), .Z(n12144) );
  XOR U14169 ( .A(n12146), .B(n12147), .Z(n5685) );
  IV U14170 ( .A(n12143), .Z(n12146) );
  XNOR U14171 ( .A(n5686), .B(n12143), .Z(n12145) );
  NAND U14172 ( .A(n12148), .B(nreg[26]), .Z(n5686) );
  NAND U14173 ( .A(n6107), .B(nreg[26]), .Z(n12148) );
  XOR U14174 ( .A(n12149), .B(n12150), .Z(n12143) );
  ANDN U14175 ( .A(n12151), .B(n5707), .Z(n12150) );
  XOR U14176 ( .A(n12152), .B(n12153), .Z(n5707) );
  IV U14177 ( .A(n12149), .Z(n12152) );
  XNOR U14178 ( .A(n5708), .B(n12149), .Z(n12151) );
  NAND U14179 ( .A(n12154), .B(nreg[25]), .Z(n5708) );
  NAND U14180 ( .A(n6107), .B(nreg[25]), .Z(n12154) );
  XOR U14181 ( .A(n12155), .B(n12156), .Z(n12149) );
  ANDN U14182 ( .A(n12157), .B(n5729), .Z(n12156) );
  XOR U14183 ( .A(n12158), .B(n12159), .Z(n5729) );
  IV U14184 ( .A(n12155), .Z(n12158) );
  XNOR U14185 ( .A(n5730), .B(n12155), .Z(n12157) );
  NAND U14186 ( .A(n12160), .B(nreg[24]), .Z(n5730) );
  NAND U14187 ( .A(n6107), .B(nreg[24]), .Z(n12160) );
  XOR U14188 ( .A(n12161), .B(n12162), .Z(n12155) );
  ANDN U14189 ( .A(n12163), .B(n5751), .Z(n12162) );
  XOR U14190 ( .A(n12164), .B(n12165), .Z(n5751) );
  IV U14191 ( .A(n12161), .Z(n12164) );
  XNOR U14192 ( .A(n5752), .B(n12161), .Z(n12163) );
  NAND U14193 ( .A(n12166), .B(nreg[23]), .Z(n5752) );
  NAND U14194 ( .A(n6107), .B(nreg[23]), .Z(n12166) );
  XOR U14195 ( .A(n12167), .B(n12168), .Z(n12161) );
  ANDN U14196 ( .A(n12169), .B(n5773), .Z(n12168) );
  XOR U14197 ( .A(n12170), .B(n12171), .Z(n5773) );
  IV U14198 ( .A(n12167), .Z(n12170) );
  XNOR U14199 ( .A(n5774), .B(n12167), .Z(n12169) );
  NAND U14200 ( .A(n12172), .B(nreg[22]), .Z(n5774) );
  NAND U14201 ( .A(n6107), .B(nreg[22]), .Z(n12172) );
  XOR U14202 ( .A(n12173), .B(n12174), .Z(n12167) );
  ANDN U14203 ( .A(n12175), .B(n5795), .Z(n12174) );
  XOR U14204 ( .A(n12176), .B(n12177), .Z(n5795) );
  IV U14205 ( .A(n12173), .Z(n12176) );
  XNOR U14206 ( .A(n5796), .B(n12173), .Z(n12175) );
  NAND U14207 ( .A(n12178), .B(nreg[21]), .Z(n5796) );
  NAND U14208 ( .A(n6107), .B(nreg[21]), .Z(n12178) );
  XOR U14209 ( .A(n12179), .B(n12180), .Z(n12173) );
  ANDN U14210 ( .A(n12181), .B(n5817), .Z(n12180) );
  XOR U14211 ( .A(n12182), .B(n12183), .Z(n5817) );
  IV U14212 ( .A(n12179), .Z(n12182) );
  XNOR U14213 ( .A(n5818), .B(n12179), .Z(n12181) );
  NAND U14214 ( .A(n12184), .B(nreg[20]), .Z(n5818) );
  NAND U14215 ( .A(n6107), .B(nreg[20]), .Z(n12184) );
  XOR U14216 ( .A(n12185), .B(n12186), .Z(n12179) );
  ANDN U14217 ( .A(n12187), .B(n5839), .Z(n12186) );
  XOR U14218 ( .A(n12188), .B(n12189), .Z(n5839) );
  IV U14219 ( .A(n12185), .Z(n12188) );
  XNOR U14220 ( .A(n5840), .B(n12185), .Z(n12187) );
  NAND U14221 ( .A(n12190), .B(nreg[19]), .Z(n5840) );
  NAND U14222 ( .A(n6107), .B(nreg[19]), .Z(n12190) );
  XOR U14223 ( .A(n12191), .B(n12192), .Z(n12185) );
  ANDN U14224 ( .A(n12193), .B(n5861), .Z(n12192) );
  XOR U14225 ( .A(n12194), .B(n12195), .Z(n5861) );
  IV U14226 ( .A(n12191), .Z(n12194) );
  XNOR U14227 ( .A(n5862), .B(n12191), .Z(n12193) );
  NAND U14228 ( .A(n12196), .B(nreg[18]), .Z(n5862) );
  NAND U14229 ( .A(n6107), .B(nreg[18]), .Z(n12196) );
  XOR U14230 ( .A(n12197), .B(n12198), .Z(n12191) );
  ANDN U14231 ( .A(n12199), .B(n5883), .Z(n12198) );
  XOR U14232 ( .A(n12200), .B(n12201), .Z(n5883) );
  IV U14233 ( .A(n12197), .Z(n12200) );
  XNOR U14234 ( .A(n5884), .B(n12197), .Z(n12199) );
  NAND U14235 ( .A(n12202), .B(nreg[17]), .Z(n5884) );
  NAND U14236 ( .A(n6107), .B(nreg[17]), .Z(n12202) );
  XOR U14237 ( .A(n12203), .B(n12204), .Z(n12197) );
  ANDN U14238 ( .A(n12205), .B(n5905), .Z(n12204) );
  XOR U14239 ( .A(n12206), .B(n12207), .Z(n5905) );
  IV U14240 ( .A(n12203), .Z(n12206) );
  XNOR U14241 ( .A(n5906), .B(n12203), .Z(n12205) );
  NAND U14242 ( .A(n12208), .B(nreg[16]), .Z(n5906) );
  NAND U14243 ( .A(n6107), .B(nreg[16]), .Z(n12208) );
  XOR U14244 ( .A(n12209), .B(n12210), .Z(n12203) );
  ANDN U14245 ( .A(n12211), .B(n5927), .Z(n12210) );
  XOR U14246 ( .A(n12212), .B(n12213), .Z(n5927) );
  IV U14247 ( .A(n12209), .Z(n12212) );
  XNOR U14248 ( .A(n5928), .B(n12209), .Z(n12211) );
  NAND U14249 ( .A(n12214), .B(nreg[15]), .Z(n5928) );
  NAND U14250 ( .A(n6107), .B(nreg[15]), .Z(n12214) );
  XOR U14251 ( .A(n12215), .B(n12216), .Z(n12209) );
  ANDN U14252 ( .A(n12217), .B(n5949), .Z(n12216) );
  XOR U14253 ( .A(n12218), .B(n12219), .Z(n5949) );
  IV U14254 ( .A(n12215), .Z(n12218) );
  XNOR U14255 ( .A(n5950), .B(n12215), .Z(n12217) );
  NAND U14256 ( .A(n12220), .B(nreg[14]), .Z(n5950) );
  NAND U14257 ( .A(n6107), .B(nreg[14]), .Z(n12220) );
  XOR U14258 ( .A(n12221), .B(n12222), .Z(n12215) );
  ANDN U14259 ( .A(n12223), .B(n5971), .Z(n12222) );
  XOR U14260 ( .A(n12224), .B(n12225), .Z(n5971) );
  IV U14261 ( .A(n12221), .Z(n12224) );
  XNOR U14262 ( .A(n5972), .B(n12221), .Z(n12223) );
  NAND U14263 ( .A(n12226), .B(nreg[13]), .Z(n5972) );
  NAND U14264 ( .A(n6107), .B(nreg[13]), .Z(n12226) );
  XOR U14265 ( .A(n12227), .B(n12228), .Z(n12221) );
  ANDN U14266 ( .A(n12229), .B(n5993), .Z(n12228) );
  XOR U14267 ( .A(n12230), .B(n12231), .Z(n5993) );
  IV U14268 ( .A(n12227), .Z(n12230) );
  XNOR U14269 ( .A(n5994), .B(n12227), .Z(n12229) );
  NAND U14270 ( .A(n12232), .B(nreg[12]), .Z(n5994) );
  NAND U14271 ( .A(n6107), .B(nreg[12]), .Z(n12232) );
  XOR U14272 ( .A(n12233), .B(n12234), .Z(n12227) );
  ANDN U14273 ( .A(n12235), .B(n6015), .Z(n12234) );
  XOR U14274 ( .A(n12236), .B(n12237), .Z(n6015) );
  IV U14275 ( .A(n12233), .Z(n12236) );
  XNOR U14276 ( .A(n6016), .B(n12233), .Z(n12235) );
  NAND U14277 ( .A(n12238), .B(nreg[11]), .Z(n6016) );
  NAND U14278 ( .A(n6107), .B(nreg[11]), .Z(n12238) );
  XOR U14279 ( .A(n12239), .B(n12240), .Z(n12233) );
  ANDN U14280 ( .A(n12241), .B(n6037), .Z(n12240) );
  XOR U14281 ( .A(n12242), .B(n12243), .Z(n6037) );
  IV U14282 ( .A(n12239), .Z(n12242) );
  XNOR U14283 ( .A(n6038), .B(n12239), .Z(n12241) );
  NAND U14284 ( .A(n12244), .B(nreg[10]), .Z(n6038) );
  NAND U14285 ( .A(n6107), .B(nreg[10]), .Z(n12244) );
  XOR U14286 ( .A(n12245), .B(n12246), .Z(n12239) );
  ANDN U14287 ( .A(n12247), .B(n6059), .Z(n12246) );
  XOR U14288 ( .A(n12248), .B(n12249), .Z(n6059) );
  IV U14289 ( .A(n12245), .Z(n12248) );
  XNOR U14290 ( .A(n6060), .B(n12245), .Z(n12247) );
  NAND U14291 ( .A(n12250), .B(nreg[9]), .Z(n6060) );
  NAND U14292 ( .A(n6107), .B(nreg[9]), .Z(n12250) );
  XOR U14293 ( .A(n12251), .B(n12252), .Z(n12245) );
  ANDN U14294 ( .A(n12253), .B(n6081), .Z(n12252) );
  XOR U14295 ( .A(n12254), .B(n12255), .Z(n6081) );
  IV U14296 ( .A(n12251), .Z(n12254) );
  XNOR U14297 ( .A(n6082), .B(n12251), .Z(n12253) );
  NAND U14298 ( .A(n12256), .B(nreg[8]), .Z(n6082) );
  NAND U14299 ( .A(n6107), .B(nreg[8]), .Z(n12256) );
  XOR U14300 ( .A(n12257), .B(n12258), .Z(n12251) );
  ANDN U14301 ( .A(n12259), .B(n12260), .Z(n12258) );
  XNOR U14302 ( .A(n12261), .B(n12257), .Z(n12259) );
  ANDN U14303 ( .A(n4110), .B(n1701), .Z(\modmult_1/N10 ) );
  XOR U14304 ( .A(n12260), .B(n12261), .Z(n1701) );
  NAND U14305 ( .A(n12262), .B(nreg[7]), .Z(n12261) );
  NAND U14306 ( .A(n6107), .B(nreg[7]), .Z(n12262) );
  XOR U14307 ( .A(n12263), .B(n12264), .Z(n12260) );
  IV U14308 ( .A(n12257), .Z(n12263) );
  XOR U14309 ( .A(n12265), .B(n12266), .Z(n12257) );
  ANDN U14310 ( .A(n12267), .B(n4331), .Z(n12266) );
  XOR U14311 ( .A(n12268), .B(n12269), .Z(n4331) );
  IV U14312 ( .A(n12265), .Z(n12268) );
  XNOR U14313 ( .A(n4332), .B(n12265), .Z(n12267) );
  NAND U14314 ( .A(n12270), .B(nreg[6]), .Z(n4332) );
  NAND U14315 ( .A(n6107), .B(nreg[6]), .Z(n12270) );
  XOR U14316 ( .A(n12271), .B(n12272), .Z(n12265) );
  ANDN U14317 ( .A(n12273), .B(n4553), .Z(n12272) );
  XOR U14318 ( .A(n12274), .B(n12275), .Z(n4553) );
  IV U14319 ( .A(n12271), .Z(n12274) );
  XNOR U14320 ( .A(n4554), .B(n12271), .Z(n12273) );
  NAND U14321 ( .A(n12276), .B(nreg[5]), .Z(n4554) );
  NAND U14322 ( .A(n6107), .B(nreg[5]), .Z(n12276) );
  XOR U14323 ( .A(n12277), .B(n12278), .Z(n12271) );
  ANDN U14324 ( .A(n12279), .B(n4775), .Z(n12278) );
  XOR U14325 ( .A(n12280), .B(n12281), .Z(n4775) );
  IV U14326 ( .A(n12277), .Z(n12280) );
  XNOR U14327 ( .A(n4776), .B(n12277), .Z(n12279) );
  NAND U14328 ( .A(n12282), .B(nreg[4]), .Z(n4776) );
  NAND U14329 ( .A(n6107), .B(nreg[4]), .Z(n12282) );
  XOR U14330 ( .A(n12283), .B(n12284), .Z(n12277) );
  ANDN U14331 ( .A(n12285), .B(n4997), .Z(n12284) );
  XOR U14332 ( .A(n12286), .B(n12287), .Z(n4997) );
  IV U14333 ( .A(n12283), .Z(n12286) );
  XNOR U14334 ( .A(n4998), .B(n12283), .Z(n12285) );
  NAND U14335 ( .A(n12288), .B(nreg[3]), .Z(n4998) );
  NAND U14336 ( .A(n6107), .B(nreg[3]), .Z(n12288) );
  XNOR U14337 ( .A(n12289), .B(n12290), .Z(n12283) );
  ANDN U14338 ( .A(n12291), .B(n5219), .Z(n12290) );
  XOR U14339 ( .A(n12289), .B(n12292), .Z(n5219) );
  XOR U14340 ( .A(n5220), .B(n12289), .Z(n12291) );
  NAND U14341 ( .A(n12293), .B(nreg[2]), .Z(n5220) );
  NAND U14342 ( .A(n6107), .B(nreg[2]), .Z(n12293) );
  XOR U14343 ( .A(n12294), .B(n12295), .Z(n12289) );
  NANDN U14344 ( .B(n5441), .A(n12296), .Z(n12294) );
  XOR U14345 ( .A(n12297), .B(n5442), .Z(n12296) );
  NAND U14346 ( .A(n12298), .B(nreg[1]), .Z(n5442) );
  NAND U14347 ( .A(n6107), .B(nreg[1]), .Z(n12298) );
  XNOR U14348 ( .A(n12299), .B(n12297), .Z(n5441) );
  IV U14349 ( .A(n12295), .Z(n12297) );
  ANDN U14350 ( .A(n5663), .B(n5664), .Z(n12295) );
  NAND U14351 ( .A(n12300), .B(nreg[0]), .Z(n5664) );
  NAND U14352 ( .A(n6107), .B(nreg[0]), .Z(n12300) );
  XOR U14353 ( .A(n12301), .B(n12302), .Z(n6107) );
  AND U14354 ( .A(n12303), .B(n12304), .Z(n12302) );
  IV U14355 ( .A(n12301), .Z(n12304) );
  XOR U14356 ( .A(n12305), .B(n12306), .Z(n12303) );
  XOR U14357 ( .A(n12307), .B(n12301), .Z(n12306) );
  XNOR U14358 ( .A(n12308), .B(n12309), .Z(n12305) );
  NOR U14359 ( .A(n12310), .B(n6101), .Z(n12308) );
  XOR U14360 ( .A(n12311), .B(n12312), .Z(n12301) );
  AND U14361 ( .A(n12313), .B(n12314), .Z(n12312) );
  IV U14362 ( .A(n12311), .Z(n12314) );
  XOR U14363 ( .A(n12311), .B(n6101), .Z(n12313) );
  XNOR U14364 ( .A(n12310), .B(n12315), .Z(n6101) );
  IV U14365 ( .A(n12307), .Z(n12310) );
  XOR U14366 ( .A(n12316), .B(n12317), .Z(n12307) );
  AND U14367 ( .A(n12318), .B(n12319), .Z(n12317) );
  XNOR U14368 ( .A(n12320), .B(n12316), .Z(n12319) );
  XOR U14369 ( .A(n12321), .B(n12322), .Z(n12311) );
  AND U14370 ( .A(n12323), .B(n12324), .Z(n12322) );
  XNOR U14371 ( .A(n12321), .B(n6108), .Z(n12324) );
  XNOR U14372 ( .A(n12318), .B(n12320), .Z(n6108) );
  NAND U14373 ( .A(n12325), .B(nreg[1023]), .Z(n12320) );
  NAND U14374 ( .A(n12326), .B(nreg[1023]), .Z(n12325) );
  XNOR U14375 ( .A(n12316), .B(n12327), .Z(n12318) );
  XOR U14376 ( .A(n12328), .B(n12329), .Z(n12316) );
  AND U14377 ( .A(n12330), .B(n12331), .Z(n12329) );
  XNOR U14378 ( .A(n12332), .B(n12328), .Z(n12331) );
  XOR U14379 ( .A(n12333), .B(nreg[1023]), .Z(n12323) );
  IV U14380 ( .A(n12321), .Z(n12333) );
  XOR U14381 ( .A(n12334), .B(n12335), .Z(n12321) );
  AND U14382 ( .A(n12336), .B(n12337), .Z(n12335) );
  XNOR U14383 ( .A(n12334), .B(n6116), .Z(n12337) );
  XNOR U14384 ( .A(n12330), .B(n12332), .Z(n6116) );
  NAND U14385 ( .A(n12338), .B(nreg[1022]), .Z(n12332) );
  NAND U14386 ( .A(n12326), .B(nreg[1022]), .Z(n12338) );
  XNOR U14387 ( .A(n12328), .B(n12339), .Z(n12330) );
  XOR U14388 ( .A(n12340), .B(n12341), .Z(n12328) );
  AND U14389 ( .A(n12342), .B(n12343), .Z(n12341) );
  XNOR U14390 ( .A(n12344), .B(n12340), .Z(n12343) );
  XOR U14391 ( .A(n12345), .B(nreg[1022]), .Z(n12336) );
  IV U14392 ( .A(n12334), .Z(n12345) );
  XOR U14393 ( .A(n12346), .B(n12347), .Z(n12334) );
  AND U14394 ( .A(n12348), .B(n12349), .Z(n12347) );
  XNOR U14395 ( .A(n12346), .B(n6124), .Z(n12349) );
  XNOR U14396 ( .A(n12342), .B(n12344), .Z(n6124) );
  NAND U14397 ( .A(n12350), .B(nreg[1021]), .Z(n12344) );
  NAND U14398 ( .A(n12326), .B(nreg[1021]), .Z(n12350) );
  XNOR U14399 ( .A(n12340), .B(n12351), .Z(n12342) );
  XOR U14400 ( .A(n12352), .B(n12353), .Z(n12340) );
  AND U14401 ( .A(n12354), .B(n12355), .Z(n12353) );
  XNOR U14402 ( .A(n12356), .B(n12352), .Z(n12355) );
  XOR U14403 ( .A(n12357), .B(nreg[1021]), .Z(n12348) );
  IV U14404 ( .A(n12346), .Z(n12357) );
  XOR U14405 ( .A(n12358), .B(n12359), .Z(n12346) );
  AND U14406 ( .A(n12360), .B(n12361), .Z(n12359) );
  XNOR U14407 ( .A(n12358), .B(n6132), .Z(n12361) );
  XNOR U14408 ( .A(n12354), .B(n12356), .Z(n6132) );
  NAND U14409 ( .A(n12362), .B(nreg[1020]), .Z(n12356) );
  NAND U14410 ( .A(n12326), .B(nreg[1020]), .Z(n12362) );
  XNOR U14411 ( .A(n12352), .B(n12363), .Z(n12354) );
  XOR U14412 ( .A(n12364), .B(n12365), .Z(n12352) );
  AND U14413 ( .A(n12366), .B(n12367), .Z(n12365) );
  XNOR U14414 ( .A(n12368), .B(n12364), .Z(n12367) );
  XOR U14415 ( .A(n12369), .B(nreg[1020]), .Z(n12360) );
  IV U14416 ( .A(n12358), .Z(n12369) );
  XOR U14417 ( .A(n12370), .B(n12371), .Z(n12358) );
  AND U14418 ( .A(n12372), .B(n12373), .Z(n12371) );
  XNOR U14419 ( .A(n12370), .B(n6140), .Z(n12373) );
  XNOR U14420 ( .A(n12366), .B(n12368), .Z(n6140) );
  NAND U14421 ( .A(n12374), .B(nreg[1019]), .Z(n12368) );
  NAND U14422 ( .A(n12326), .B(nreg[1019]), .Z(n12374) );
  XNOR U14423 ( .A(n12364), .B(n12375), .Z(n12366) );
  XOR U14424 ( .A(n12376), .B(n12377), .Z(n12364) );
  AND U14425 ( .A(n12378), .B(n12379), .Z(n12377) );
  XNOR U14426 ( .A(n12380), .B(n12376), .Z(n12379) );
  XOR U14427 ( .A(n12381), .B(nreg[1019]), .Z(n12372) );
  IV U14428 ( .A(n12370), .Z(n12381) );
  XOR U14429 ( .A(n12382), .B(n12383), .Z(n12370) );
  AND U14430 ( .A(n12384), .B(n12385), .Z(n12383) );
  XNOR U14431 ( .A(n12382), .B(n6148), .Z(n12385) );
  XNOR U14432 ( .A(n12378), .B(n12380), .Z(n6148) );
  NAND U14433 ( .A(n12386), .B(nreg[1018]), .Z(n12380) );
  NAND U14434 ( .A(n12326), .B(nreg[1018]), .Z(n12386) );
  XNOR U14435 ( .A(n12376), .B(n12387), .Z(n12378) );
  XOR U14436 ( .A(n12388), .B(n12389), .Z(n12376) );
  AND U14437 ( .A(n12390), .B(n12391), .Z(n12389) );
  XNOR U14438 ( .A(n12392), .B(n12388), .Z(n12391) );
  XOR U14439 ( .A(n12393), .B(nreg[1018]), .Z(n12384) );
  IV U14440 ( .A(n12382), .Z(n12393) );
  XOR U14441 ( .A(n12394), .B(n12395), .Z(n12382) );
  AND U14442 ( .A(n12396), .B(n12397), .Z(n12395) );
  XNOR U14443 ( .A(n12394), .B(n6156), .Z(n12397) );
  XNOR U14444 ( .A(n12390), .B(n12392), .Z(n6156) );
  NAND U14445 ( .A(n12398), .B(nreg[1017]), .Z(n12392) );
  NAND U14446 ( .A(n12326), .B(nreg[1017]), .Z(n12398) );
  XNOR U14447 ( .A(n12388), .B(n12399), .Z(n12390) );
  XOR U14448 ( .A(n12400), .B(n12401), .Z(n12388) );
  AND U14449 ( .A(n12402), .B(n12403), .Z(n12401) );
  XNOR U14450 ( .A(n12404), .B(n12400), .Z(n12403) );
  XOR U14451 ( .A(n12405), .B(nreg[1017]), .Z(n12396) );
  IV U14452 ( .A(n12394), .Z(n12405) );
  XOR U14453 ( .A(n12406), .B(n12407), .Z(n12394) );
  AND U14454 ( .A(n12408), .B(n12409), .Z(n12407) );
  XNOR U14455 ( .A(n12406), .B(n6166), .Z(n12409) );
  XNOR U14456 ( .A(n12402), .B(n12404), .Z(n6166) );
  NAND U14457 ( .A(n12410), .B(nreg[1016]), .Z(n12404) );
  NAND U14458 ( .A(n12326), .B(nreg[1016]), .Z(n12410) );
  XNOR U14459 ( .A(n12400), .B(n12411), .Z(n12402) );
  XOR U14460 ( .A(n12412), .B(n12413), .Z(n12400) );
  AND U14461 ( .A(n12414), .B(n12415), .Z(n12413) );
  XNOR U14462 ( .A(n12416), .B(n12412), .Z(n12415) );
  XOR U14463 ( .A(n12417), .B(nreg[1016]), .Z(n12408) );
  IV U14464 ( .A(n12406), .Z(n12417) );
  XOR U14465 ( .A(n12418), .B(n12419), .Z(n12406) );
  AND U14466 ( .A(n12420), .B(n12421), .Z(n12419) );
  XNOR U14467 ( .A(n12418), .B(n6174), .Z(n12421) );
  XNOR U14468 ( .A(n12414), .B(n12416), .Z(n6174) );
  NAND U14469 ( .A(n12422), .B(nreg[1015]), .Z(n12416) );
  NAND U14470 ( .A(n12326), .B(nreg[1015]), .Z(n12422) );
  XNOR U14471 ( .A(n12412), .B(n12423), .Z(n12414) );
  XOR U14472 ( .A(n12424), .B(n12425), .Z(n12412) );
  AND U14473 ( .A(n12426), .B(n12427), .Z(n12425) );
  XNOR U14474 ( .A(n12428), .B(n12424), .Z(n12427) );
  XOR U14475 ( .A(n12429), .B(nreg[1015]), .Z(n12420) );
  IV U14476 ( .A(n12418), .Z(n12429) );
  XOR U14477 ( .A(n12430), .B(n12431), .Z(n12418) );
  AND U14478 ( .A(n12432), .B(n12433), .Z(n12431) );
  XNOR U14479 ( .A(n12430), .B(n6182), .Z(n12433) );
  XNOR U14480 ( .A(n12426), .B(n12428), .Z(n6182) );
  NAND U14481 ( .A(n12434), .B(nreg[1014]), .Z(n12428) );
  NAND U14482 ( .A(n12326), .B(nreg[1014]), .Z(n12434) );
  XNOR U14483 ( .A(n12424), .B(n12435), .Z(n12426) );
  XOR U14484 ( .A(n12436), .B(n12437), .Z(n12424) );
  AND U14485 ( .A(n12438), .B(n12439), .Z(n12437) );
  XNOR U14486 ( .A(n12440), .B(n12436), .Z(n12439) );
  XOR U14487 ( .A(n12441), .B(nreg[1014]), .Z(n12432) );
  IV U14488 ( .A(n12430), .Z(n12441) );
  XOR U14489 ( .A(n12442), .B(n12443), .Z(n12430) );
  AND U14490 ( .A(n12444), .B(n12445), .Z(n12443) );
  XNOR U14491 ( .A(n12442), .B(n6190), .Z(n12445) );
  XNOR U14492 ( .A(n12438), .B(n12440), .Z(n6190) );
  NAND U14493 ( .A(n12446), .B(nreg[1013]), .Z(n12440) );
  NAND U14494 ( .A(n12326), .B(nreg[1013]), .Z(n12446) );
  XNOR U14495 ( .A(n12436), .B(n12447), .Z(n12438) );
  XOR U14496 ( .A(n12448), .B(n12449), .Z(n12436) );
  AND U14497 ( .A(n12450), .B(n12451), .Z(n12449) );
  XNOR U14498 ( .A(n12452), .B(n12448), .Z(n12451) );
  XOR U14499 ( .A(n12453), .B(nreg[1013]), .Z(n12444) );
  IV U14500 ( .A(n12442), .Z(n12453) );
  XOR U14501 ( .A(n12454), .B(n12455), .Z(n12442) );
  AND U14502 ( .A(n12456), .B(n12457), .Z(n12455) );
  XNOR U14503 ( .A(n12454), .B(n6198), .Z(n12457) );
  XNOR U14504 ( .A(n12450), .B(n12452), .Z(n6198) );
  NAND U14505 ( .A(n12458), .B(nreg[1012]), .Z(n12452) );
  NAND U14506 ( .A(n12326), .B(nreg[1012]), .Z(n12458) );
  XNOR U14507 ( .A(n12448), .B(n12459), .Z(n12450) );
  XOR U14508 ( .A(n12460), .B(n12461), .Z(n12448) );
  AND U14509 ( .A(n12462), .B(n12463), .Z(n12461) );
  XNOR U14510 ( .A(n12464), .B(n12460), .Z(n12463) );
  XOR U14511 ( .A(n12465), .B(nreg[1012]), .Z(n12456) );
  IV U14512 ( .A(n12454), .Z(n12465) );
  XOR U14513 ( .A(n12466), .B(n12467), .Z(n12454) );
  AND U14514 ( .A(n12468), .B(n12469), .Z(n12467) );
  XNOR U14515 ( .A(n12466), .B(n6206), .Z(n12469) );
  XNOR U14516 ( .A(n12462), .B(n12464), .Z(n6206) );
  NAND U14517 ( .A(n12470), .B(nreg[1011]), .Z(n12464) );
  NAND U14518 ( .A(n12326), .B(nreg[1011]), .Z(n12470) );
  XNOR U14519 ( .A(n12460), .B(n12471), .Z(n12462) );
  XOR U14520 ( .A(n12472), .B(n12473), .Z(n12460) );
  AND U14521 ( .A(n12474), .B(n12475), .Z(n12473) );
  XNOR U14522 ( .A(n12476), .B(n12472), .Z(n12475) );
  XOR U14523 ( .A(n12477), .B(nreg[1011]), .Z(n12468) );
  IV U14524 ( .A(n12466), .Z(n12477) );
  XOR U14525 ( .A(n12478), .B(n12479), .Z(n12466) );
  AND U14526 ( .A(n12480), .B(n12481), .Z(n12479) );
  XNOR U14527 ( .A(n12478), .B(n6214), .Z(n12481) );
  XNOR U14528 ( .A(n12474), .B(n12476), .Z(n6214) );
  NAND U14529 ( .A(n12482), .B(nreg[1010]), .Z(n12476) );
  NAND U14530 ( .A(n12326), .B(nreg[1010]), .Z(n12482) );
  XNOR U14531 ( .A(n12472), .B(n12483), .Z(n12474) );
  XOR U14532 ( .A(n12484), .B(n12485), .Z(n12472) );
  AND U14533 ( .A(n12486), .B(n12487), .Z(n12485) );
  XNOR U14534 ( .A(n12488), .B(n12484), .Z(n12487) );
  XOR U14535 ( .A(n12489), .B(nreg[1010]), .Z(n12480) );
  IV U14536 ( .A(n12478), .Z(n12489) );
  XOR U14537 ( .A(n12490), .B(n12491), .Z(n12478) );
  AND U14538 ( .A(n12492), .B(n12493), .Z(n12491) );
  XNOR U14539 ( .A(n12490), .B(n6222), .Z(n12493) );
  XNOR U14540 ( .A(n12486), .B(n12488), .Z(n6222) );
  NAND U14541 ( .A(n12494), .B(nreg[1009]), .Z(n12488) );
  NAND U14542 ( .A(n12326), .B(nreg[1009]), .Z(n12494) );
  XNOR U14543 ( .A(n12484), .B(n12495), .Z(n12486) );
  XOR U14544 ( .A(n12496), .B(n12497), .Z(n12484) );
  AND U14545 ( .A(n12498), .B(n12499), .Z(n12497) );
  XNOR U14546 ( .A(n12500), .B(n12496), .Z(n12499) );
  XOR U14547 ( .A(n12501), .B(nreg[1009]), .Z(n12492) );
  IV U14548 ( .A(n12490), .Z(n12501) );
  XOR U14549 ( .A(n12502), .B(n12503), .Z(n12490) );
  AND U14550 ( .A(n12504), .B(n12505), .Z(n12503) );
  XNOR U14551 ( .A(n12502), .B(n6230), .Z(n12505) );
  XNOR U14552 ( .A(n12498), .B(n12500), .Z(n6230) );
  NAND U14553 ( .A(n12506), .B(nreg[1008]), .Z(n12500) );
  NAND U14554 ( .A(n12326), .B(nreg[1008]), .Z(n12506) );
  XNOR U14555 ( .A(n12496), .B(n12507), .Z(n12498) );
  XOR U14556 ( .A(n12508), .B(n12509), .Z(n12496) );
  AND U14557 ( .A(n12510), .B(n12511), .Z(n12509) );
  XNOR U14558 ( .A(n12512), .B(n12508), .Z(n12511) );
  XOR U14559 ( .A(n12513), .B(nreg[1008]), .Z(n12504) );
  IV U14560 ( .A(n12502), .Z(n12513) );
  XOR U14561 ( .A(n12514), .B(n12515), .Z(n12502) );
  AND U14562 ( .A(n12516), .B(n12517), .Z(n12515) );
  XNOR U14563 ( .A(n12514), .B(n6238), .Z(n12517) );
  XNOR U14564 ( .A(n12510), .B(n12512), .Z(n6238) );
  NAND U14565 ( .A(n12518), .B(nreg[1007]), .Z(n12512) );
  NAND U14566 ( .A(n12326), .B(nreg[1007]), .Z(n12518) );
  XNOR U14567 ( .A(n12508), .B(n12519), .Z(n12510) );
  XOR U14568 ( .A(n12520), .B(n12521), .Z(n12508) );
  AND U14569 ( .A(n12522), .B(n12523), .Z(n12521) );
  XNOR U14570 ( .A(n12524), .B(n12520), .Z(n12523) );
  XOR U14571 ( .A(n12525), .B(nreg[1007]), .Z(n12516) );
  IV U14572 ( .A(n12514), .Z(n12525) );
  XOR U14573 ( .A(n12526), .B(n12527), .Z(n12514) );
  AND U14574 ( .A(n12528), .B(n12529), .Z(n12527) );
  XNOR U14575 ( .A(n12526), .B(n6248), .Z(n12529) );
  XNOR U14576 ( .A(n12522), .B(n12524), .Z(n6248) );
  NAND U14577 ( .A(n12530), .B(nreg[1006]), .Z(n12524) );
  NAND U14578 ( .A(n12326), .B(nreg[1006]), .Z(n12530) );
  XNOR U14579 ( .A(n12520), .B(n12531), .Z(n12522) );
  XOR U14580 ( .A(n12532), .B(n12533), .Z(n12520) );
  AND U14581 ( .A(n12534), .B(n12535), .Z(n12533) );
  XNOR U14582 ( .A(n12536), .B(n12532), .Z(n12535) );
  XOR U14583 ( .A(n12537), .B(nreg[1006]), .Z(n12528) );
  IV U14584 ( .A(n12526), .Z(n12537) );
  XOR U14585 ( .A(n12538), .B(n12539), .Z(n12526) );
  AND U14586 ( .A(n12540), .B(n12541), .Z(n12539) );
  XNOR U14587 ( .A(n12538), .B(n6256), .Z(n12541) );
  XNOR U14588 ( .A(n12534), .B(n12536), .Z(n6256) );
  NAND U14589 ( .A(n12542), .B(nreg[1005]), .Z(n12536) );
  NAND U14590 ( .A(n12326), .B(nreg[1005]), .Z(n12542) );
  XNOR U14591 ( .A(n12532), .B(n12543), .Z(n12534) );
  XOR U14592 ( .A(n12544), .B(n12545), .Z(n12532) );
  AND U14593 ( .A(n12546), .B(n12547), .Z(n12545) );
  XNOR U14594 ( .A(n12548), .B(n12544), .Z(n12547) );
  XOR U14595 ( .A(n12549), .B(nreg[1005]), .Z(n12540) );
  IV U14596 ( .A(n12538), .Z(n12549) );
  XOR U14597 ( .A(n12550), .B(n12551), .Z(n12538) );
  AND U14598 ( .A(n12552), .B(n12553), .Z(n12551) );
  XNOR U14599 ( .A(n12550), .B(n6264), .Z(n12553) );
  XNOR U14600 ( .A(n12546), .B(n12548), .Z(n6264) );
  NAND U14601 ( .A(n12554), .B(nreg[1004]), .Z(n12548) );
  NAND U14602 ( .A(n12326), .B(nreg[1004]), .Z(n12554) );
  XNOR U14603 ( .A(n12544), .B(n12555), .Z(n12546) );
  XOR U14604 ( .A(n12556), .B(n12557), .Z(n12544) );
  AND U14605 ( .A(n12558), .B(n12559), .Z(n12557) );
  XNOR U14606 ( .A(n12560), .B(n12556), .Z(n12559) );
  XOR U14607 ( .A(n12561), .B(nreg[1004]), .Z(n12552) );
  IV U14608 ( .A(n12550), .Z(n12561) );
  XOR U14609 ( .A(n12562), .B(n12563), .Z(n12550) );
  AND U14610 ( .A(n12564), .B(n12565), .Z(n12563) );
  XNOR U14611 ( .A(n12562), .B(n6272), .Z(n12565) );
  XNOR U14612 ( .A(n12558), .B(n12560), .Z(n6272) );
  NAND U14613 ( .A(n12566), .B(nreg[1003]), .Z(n12560) );
  NAND U14614 ( .A(n12326), .B(nreg[1003]), .Z(n12566) );
  XNOR U14615 ( .A(n12556), .B(n12567), .Z(n12558) );
  XOR U14616 ( .A(n12568), .B(n12569), .Z(n12556) );
  AND U14617 ( .A(n12570), .B(n12571), .Z(n12569) );
  XNOR U14618 ( .A(n12572), .B(n12568), .Z(n12571) );
  XOR U14619 ( .A(n12573), .B(nreg[1003]), .Z(n12564) );
  IV U14620 ( .A(n12562), .Z(n12573) );
  XOR U14621 ( .A(n12574), .B(n12575), .Z(n12562) );
  AND U14622 ( .A(n12576), .B(n12577), .Z(n12575) );
  XNOR U14623 ( .A(n12574), .B(n6280), .Z(n12577) );
  XNOR U14624 ( .A(n12570), .B(n12572), .Z(n6280) );
  NAND U14625 ( .A(n12578), .B(nreg[1002]), .Z(n12572) );
  NAND U14626 ( .A(n12326), .B(nreg[1002]), .Z(n12578) );
  XNOR U14627 ( .A(n12568), .B(n12579), .Z(n12570) );
  XOR U14628 ( .A(n12580), .B(n12581), .Z(n12568) );
  AND U14629 ( .A(n12582), .B(n12583), .Z(n12581) );
  XNOR U14630 ( .A(n12584), .B(n12580), .Z(n12583) );
  XOR U14631 ( .A(n12585), .B(nreg[1002]), .Z(n12576) );
  IV U14632 ( .A(n12574), .Z(n12585) );
  XOR U14633 ( .A(n12586), .B(n12587), .Z(n12574) );
  AND U14634 ( .A(n12588), .B(n12589), .Z(n12587) );
  XNOR U14635 ( .A(n12586), .B(n6288), .Z(n12589) );
  XNOR U14636 ( .A(n12582), .B(n12584), .Z(n6288) );
  NAND U14637 ( .A(n12590), .B(nreg[1001]), .Z(n12584) );
  NAND U14638 ( .A(n12326), .B(nreg[1001]), .Z(n12590) );
  XNOR U14639 ( .A(n12580), .B(n12591), .Z(n12582) );
  XOR U14640 ( .A(n12592), .B(n12593), .Z(n12580) );
  AND U14641 ( .A(n12594), .B(n12595), .Z(n12593) );
  XNOR U14642 ( .A(n12596), .B(n12592), .Z(n12595) );
  XOR U14643 ( .A(n12597), .B(nreg[1001]), .Z(n12588) );
  IV U14644 ( .A(n12586), .Z(n12597) );
  XOR U14645 ( .A(n12598), .B(n12599), .Z(n12586) );
  AND U14646 ( .A(n12600), .B(n12601), .Z(n12599) );
  XNOR U14647 ( .A(n12598), .B(n6296), .Z(n12601) );
  XNOR U14648 ( .A(n12594), .B(n12596), .Z(n6296) );
  NAND U14649 ( .A(n12602), .B(nreg[1000]), .Z(n12596) );
  NAND U14650 ( .A(n12326), .B(nreg[1000]), .Z(n12602) );
  XNOR U14651 ( .A(n12592), .B(n12603), .Z(n12594) );
  XOR U14652 ( .A(n12604), .B(n12605), .Z(n12592) );
  AND U14653 ( .A(n12606), .B(n12607), .Z(n12605) );
  XNOR U14654 ( .A(n12608), .B(n12604), .Z(n12607) );
  XOR U14655 ( .A(n12609), .B(nreg[1000]), .Z(n12600) );
  IV U14656 ( .A(n12598), .Z(n12609) );
  XOR U14657 ( .A(n12610), .B(n12611), .Z(n12598) );
  AND U14658 ( .A(n12612), .B(n12613), .Z(n12611) );
  XNOR U14659 ( .A(n12610), .B(n6304), .Z(n12613) );
  XNOR U14660 ( .A(n12606), .B(n12608), .Z(n6304) );
  NAND U14661 ( .A(n12614), .B(nreg[999]), .Z(n12608) );
  NAND U14662 ( .A(n12326), .B(nreg[999]), .Z(n12614) );
  XNOR U14663 ( .A(n12604), .B(n12615), .Z(n12606) );
  XOR U14664 ( .A(n12616), .B(n12617), .Z(n12604) );
  AND U14665 ( .A(n12618), .B(n12619), .Z(n12617) );
  XNOR U14666 ( .A(n12620), .B(n12616), .Z(n12619) );
  XOR U14667 ( .A(n12621), .B(nreg[999]), .Z(n12612) );
  IV U14668 ( .A(n12610), .Z(n12621) );
  XOR U14669 ( .A(n12622), .B(n12623), .Z(n12610) );
  AND U14670 ( .A(n12624), .B(n12625), .Z(n12623) );
  XNOR U14671 ( .A(n12622), .B(n6312), .Z(n12625) );
  XNOR U14672 ( .A(n12618), .B(n12620), .Z(n6312) );
  NAND U14673 ( .A(n12626), .B(nreg[998]), .Z(n12620) );
  NAND U14674 ( .A(n12326), .B(nreg[998]), .Z(n12626) );
  XNOR U14675 ( .A(n12616), .B(n12627), .Z(n12618) );
  XOR U14676 ( .A(n12628), .B(n12629), .Z(n12616) );
  AND U14677 ( .A(n12630), .B(n12631), .Z(n12629) );
  XNOR U14678 ( .A(n12632), .B(n12628), .Z(n12631) );
  XOR U14679 ( .A(n12633), .B(nreg[998]), .Z(n12624) );
  IV U14680 ( .A(n12622), .Z(n12633) );
  XOR U14681 ( .A(n12634), .B(n12635), .Z(n12622) );
  AND U14682 ( .A(n12636), .B(n12637), .Z(n12635) );
  XNOR U14683 ( .A(n12634), .B(n6320), .Z(n12637) );
  XNOR U14684 ( .A(n12630), .B(n12632), .Z(n6320) );
  NAND U14685 ( .A(n12638), .B(nreg[997]), .Z(n12632) );
  NAND U14686 ( .A(n12326), .B(nreg[997]), .Z(n12638) );
  XNOR U14687 ( .A(n12628), .B(n12639), .Z(n12630) );
  XOR U14688 ( .A(n12640), .B(n12641), .Z(n12628) );
  AND U14689 ( .A(n12642), .B(n12643), .Z(n12641) );
  XNOR U14690 ( .A(n12644), .B(n12640), .Z(n12643) );
  XOR U14691 ( .A(n12645), .B(nreg[997]), .Z(n12636) );
  IV U14692 ( .A(n12634), .Z(n12645) );
  XOR U14693 ( .A(n12646), .B(n12647), .Z(n12634) );
  AND U14694 ( .A(n12648), .B(n12649), .Z(n12647) );
  XNOR U14695 ( .A(n12646), .B(n6325), .Z(n12649) );
  XNOR U14696 ( .A(n12642), .B(n12644), .Z(n6325) );
  NAND U14697 ( .A(n12650), .B(nreg[996]), .Z(n12644) );
  NAND U14698 ( .A(n12326), .B(nreg[996]), .Z(n12650) );
  XNOR U14699 ( .A(n12640), .B(n12651), .Z(n12642) );
  XOR U14700 ( .A(n12652), .B(n12653), .Z(n12640) );
  AND U14701 ( .A(n12654), .B(n12655), .Z(n12653) );
  XNOR U14702 ( .A(n12656), .B(n12652), .Z(n12655) );
  XOR U14703 ( .A(n12657), .B(nreg[996]), .Z(n12648) );
  IV U14704 ( .A(n12646), .Z(n12657) );
  XOR U14705 ( .A(n12658), .B(n12659), .Z(n12646) );
  AND U14706 ( .A(n12660), .B(n12661), .Z(n12659) );
  XNOR U14707 ( .A(n12658), .B(n6331), .Z(n12661) );
  XNOR U14708 ( .A(n12654), .B(n12656), .Z(n6331) );
  NAND U14709 ( .A(n12662), .B(nreg[995]), .Z(n12656) );
  NAND U14710 ( .A(n12326), .B(nreg[995]), .Z(n12662) );
  XNOR U14711 ( .A(n12652), .B(n12663), .Z(n12654) );
  XOR U14712 ( .A(n12664), .B(n12665), .Z(n12652) );
  AND U14713 ( .A(n12666), .B(n12667), .Z(n12665) );
  XNOR U14714 ( .A(n12668), .B(n12664), .Z(n12667) );
  XOR U14715 ( .A(n12669), .B(nreg[995]), .Z(n12660) );
  IV U14716 ( .A(n12658), .Z(n12669) );
  XOR U14717 ( .A(n12670), .B(n12671), .Z(n12658) );
  AND U14718 ( .A(n12672), .B(n12673), .Z(n12671) );
  XNOR U14719 ( .A(n12670), .B(n6337), .Z(n12673) );
  XNOR U14720 ( .A(n12666), .B(n12668), .Z(n6337) );
  NAND U14721 ( .A(n12674), .B(nreg[994]), .Z(n12668) );
  NAND U14722 ( .A(n12326), .B(nreg[994]), .Z(n12674) );
  XNOR U14723 ( .A(n12664), .B(n12675), .Z(n12666) );
  XOR U14724 ( .A(n12676), .B(n12677), .Z(n12664) );
  AND U14725 ( .A(n12678), .B(n12679), .Z(n12677) );
  XNOR U14726 ( .A(n12680), .B(n12676), .Z(n12679) );
  XOR U14727 ( .A(n12681), .B(nreg[994]), .Z(n12672) );
  IV U14728 ( .A(n12670), .Z(n12681) );
  XOR U14729 ( .A(n12682), .B(n12683), .Z(n12670) );
  AND U14730 ( .A(n12684), .B(n12685), .Z(n12683) );
  XNOR U14731 ( .A(n12682), .B(n6343), .Z(n12685) );
  XNOR U14732 ( .A(n12678), .B(n12680), .Z(n6343) );
  NAND U14733 ( .A(n12686), .B(nreg[993]), .Z(n12680) );
  NAND U14734 ( .A(n12326), .B(nreg[993]), .Z(n12686) );
  XNOR U14735 ( .A(n12676), .B(n12687), .Z(n12678) );
  XOR U14736 ( .A(n12688), .B(n12689), .Z(n12676) );
  AND U14737 ( .A(n12690), .B(n12691), .Z(n12689) );
  XNOR U14738 ( .A(n12692), .B(n12688), .Z(n12691) );
  XOR U14739 ( .A(n12693), .B(nreg[993]), .Z(n12684) );
  IV U14740 ( .A(n12682), .Z(n12693) );
  XOR U14741 ( .A(n12694), .B(n12695), .Z(n12682) );
  AND U14742 ( .A(n12696), .B(n12697), .Z(n12695) );
  XNOR U14743 ( .A(n12694), .B(n6349), .Z(n12697) );
  XNOR U14744 ( .A(n12690), .B(n12692), .Z(n6349) );
  NAND U14745 ( .A(n12698), .B(nreg[992]), .Z(n12692) );
  NAND U14746 ( .A(n12326), .B(nreg[992]), .Z(n12698) );
  XNOR U14747 ( .A(n12688), .B(n12699), .Z(n12690) );
  XOR U14748 ( .A(n12700), .B(n12701), .Z(n12688) );
  AND U14749 ( .A(n12702), .B(n12703), .Z(n12701) );
  XNOR U14750 ( .A(n12704), .B(n12700), .Z(n12703) );
  XOR U14751 ( .A(n12705), .B(nreg[992]), .Z(n12696) );
  IV U14752 ( .A(n12694), .Z(n12705) );
  XOR U14753 ( .A(n12706), .B(n12707), .Z(n12694) );
  AND U14754 ( .A(n12708), .B(n12709), .Z(n12707) );
  XNOR U14755 ( .A(n12706), .B(n6355), .Z(n12709) );
  XNOR U14756 ( .A(n12702), .B(n12704), .Z(n6355) );
  NAND U14757 ( .A(n12710), .B(nreg[991]), .Z(n12704) );
  NAND U14758 ( .A(n12326), .B(nreg[991]), .Z(n12710) );
  XNOR U14759 ( .A(n12700), .B(n12711), .Z(n12702) );
  XOR U14760 ( .A(n12712), .B(n12713), .Z(n12700) );
  AND U14761 ( .A(n12714), .B(n12715), .Z(n12713) );
  XNOR U14762 ( .A(n12716), .B(n12712), .Z(n12715) );
  XOR U14763 ( .A(n12717), .B(nreg[991]), .Z(n12708) );
  IV U14764 ( .A(n12706), .Z(n12717) );
  XOR U14765 ( .A(n12718), .B(n12719), .Z(n12706) );
  AND U14766 ( .A(n12720), .B(n12721), .Z(n12719) );
  XNOR U14767 ( .A(n12718), .B(n6361), .Z(n12721) );
  XNOR U14768 ( .A(n12714), .B(n12716), .Z(n6361) );
  NAND U14769 ( .A(n12722), .B(nreg[990]), .Z(n12716) );
  NAND U14770 ( .A(n12326), .B(nreg[990]), .Z(n12722) );
  XNOR U14771 ( .A(n12712), .B(n12723), .Z(n12714) );
  XOR U14772 ( .A(n12724), .B(n12725), .Z(n12712) );
  AND U14773 ( .A(n12726), .B(n12727), .Z(n12725) );
  XNOR U14774 ( .A(n12728), .B(n12724), .Z(n12727) );
  XOR U14775 ( .A(n12729), .B(nreg[990]), .Z(n12720) );
  IV U14776 ( .A(n12718), .Z(n12729) );
  XOR U14777 ( .A(n12730), .B(n12731), .Z(n12718) );
  AND U14778 ( .A(n12732), .B(n12733), .Z(n12731) );
  XNOR U14779 ( .A(n12730), .B(n6367), .Z(n12733) );
  XNOR U14780 ( .A(n12726), .B(n12728), .Z(n6367) );
  NAND U14781 ( .A(n12734), .B(nreg[989]), .Z(n12728) );
  NAND U14782 ( .A(n12326), .B(nreg[989]), .Z(n12734) );
  XNOR U14783 ( .A(n12724), .B(n12735), .Z(n12726) );
  XOR U14784 ( .A(n12736), .B(n12737), .Z(n12724) );
  AND U14785 ( .A(n12738), .B(n12739), .Z(n12737) );
  XNOR U14786 ( .A(n12740), .B(n12736), .Z(n12739) );
  XOR U14787 ( .A(n12741), .B(nreg[989]), .Z(n12732) );
  IV U14788 ( .A(n12730), .Z(n12741) );
  XOR U14789 ( .A(n12742), .B(n12743), .Z(n12730) );
  AND U14790 ( .A(n12744), .B(n12745), .Z(n12743) );
  XNOR U14791 ( .A(n12742), .B(n6373), .Z(n12745) );
  XNOR U14792 ( .A(n12738), .B(n12740), .Z(n6373) );
  NAND U14793 ( .A(n12746), .B(nreg[988]), .Z(n12740) );
  NAND U14794 ( .A(n12326), .B(nreg[988]), .Z(n12746) );
  XNOR U14795 ( .A(n12736), .B(n12747), .Z(n12738) );
  XOR U14796 ( .A(n12748), .B(n12749), .Z(n12736) );
  AND U14797 ( .A(n12750), .B(n12751), .Z(n12749) );
  XNOR U14798 ( .A(n12752), .B(n12748), .Z(n12751) );
  XOR U14799 ( .A(n12753), .B(nreg[988]), .Z(n12744) );
  IV U14800 ( .A(n12742), .Z(n12753) );
  XOR U14801 ( .A(n12754), .B(n12755), .Z(n12742) );
  AND U14802 ( .A(n12756), .B(n12757), .Z(n12755) );
  XNOR U14803 ( .A(n12754), .B(n6379), .Z(n12757) );
  XNOR U14804 ( .A(n12750), .B(n12752), .Z(n6379) );
  NAND U14805 ( .A(n12758), .B(nreg[987]), .Z(n12752) );
  NAND U14806 ( .A(n12326), .B(nreg[987]), .Z(n12758) );
  XNOR U14807 ( .A(n12748), .B(n12759), .Z(n12750) );
  XOR U14808 ( .A(n12760), .B(n12761), .Z(n12748) );
  AND U14809 ( .A(n12762), .B(n12763), .Z(n12761) );
  XNOR U14810 ( .A(n12764), .B(n12760), .Z(n12763) );
  XOR U14811 ( .A(n12765), .B(nreg[987]), .Z(n12756) );
  IV U14812 ( .A(n12754), .Z(n12765) );
  XOR U14813 ( .A(n12766), .B(n12767), .Z(n12754) );
  AND U14814 ( .A(n12768), .B(n12769), .Z(n12767) );
  XNOR U14815 ( .A(n12766), .B(n6385), .Z(n12769) );
  XNOR U14816 ( .A(n12762), .B(n12764), .Z(n6385) );
  NAND U14817 ( .A(n12770), .B(nreg[986]), .Z(n12764) );
  NAND U14818 ( .A(n12326), .B(nreg[986]), .Z(n12770) );
  XNOR U14819 ( .A(n12760), .B(n12771), .Z(n12762) );
  XOR U14820 ( .A(n12772), .B(n12773), .Z(n12760) );
  AND U14821 ( .A(n12774), .B(n12775), .Z(n12773) );
  XNOR U14822 ( .A(n12776), .B(n12772), .Z(n12775) );
  XOR U14823 ( .A(n12777), .B(nreg[986]), .Z(n12768) );
  IV U14824 ( .A(n12766), .Z(n12777) );
  XOR U14825 ( .A(n12778), .B(n12779), .Z(n12766) );
  AND U14826 ( .A(n12780), .B(n12781), .Z(n12779) );
  XNOR U14827 ( .A(n12778), .B(n6391), .Z(n12781) );
  XNOR U14828 ( .A(n12774), .B(n12776), .Z(n6391) );
  NAND U14829 ( .A(n12782), .B(nreg[985]), .Z(n12776) );
  NAND U14830 ( .A(n12326), .B(nreg[985]), .Z(n12782) );
  XNOR U14831 ( .A(n12772), .B(n12783), .Z(n12774) );
  XOR U14832 ( .A(n12784), .B(n12785), .Z(n12772) );
  AND U14833 ( .A(n12786), .B(n12787), .Z(n12785) );
  XNOR U14834 ( .A(n12788), .B(n12784), .Z(n12787) );
  XOR U14835 ( .A(n12789), .B(nreg[985]), .Z(n12780) );
  IV U14836 ( .A(n12778), .Z(n12789) );
  XOR U14837 ( .A(n12790), .B(n12791), .Z(n12778) );
  AND U14838 ( .A(n12792), .B(n12793), .Z(n12791) );
  XNOR U14839 ( .A(n12790), .B(n6397), .Z(n12793) );
  XNOR U14840 ( .A(n12786), .B(n12788), .Z(n6397) );
  NAND U14841 ( .A(n12794), .B(nreg[984]), .Z(n12788) );
  NAND U14842 ( .A(n12326), .B(nreg[984]), .Z(n12794) );
  XNOR U14843 ( .A(n12784), .B(n12795), .Z(n12786) );
  XOR U14844 ( .A(n12796), .B(n12797), .Z(n12784) );
  AND U14845 ( .A(n12798), .B(n12799), .Z(n12797) );
  XNOR U14846 ( .A(n12800), .B(n12796), .Z(n12799) );
  XOR U14847 ( .A(n12801), .B(nreg[984]), .Z(n12792) );
  IV U14848 ( .A(n12790), .Z(n12801) );
  XOR U14849 ( .A(n12802), .B(n12803), .Z(n12790) );
  AND U14850 ( .A(n12804), .B(n12805), .Z(n12803) );
  XNOR U14851 ( .A(n12802), .B(n6403), .Z(n12805) );
  XNOR U14852 ( .A(n12798), .B(n12800), .Z(n6403) );
  NAND U14853 ( .A(n12806), .B(nreg[983]), .Z(n12800) );
  NAND U14854 ( .A(n12326), .B(nreg[983]), .Z(n12806) );
  XNOR U14855 ( .A(n12796), .B(n12807), .Z(n12798) );
  XOR U14856 ( .A(n12808), .B(n12809), .Z(n12796) );
  AND U14857 ( .A(n12810), .B(n12811), .Z(n12809) );
  XNOR U14858 ( .A(n12812), .B(n12808), .Z(n12811) );
  XOR U14859 ( .A(n12813), .B(nreg[983]), .Z(n12804) );
  IV U14860 ( .A(n12802), .Z(n12813) );
  XOR U14861 ( .A(n12814), .B(n12815), .Z(n12802) );
  AND U14862 ( .A(n12816), .B(n12817), .Z(n12815) );
  XNOR U14863 ( .A(n12814), .B(n6409), .Z(n12817) );
  XNOR U14864 ( .A(n12810), .B(n12812), .Z(n6409) );
  NAND U14865 ( .A(n12818), .B(nreg[982]), .Z(n12812) );
  NAND U14866 ( .A(n12326), .B(nreg[982]), .Z(n12818) );
  XNOR U14867 ( .A(n12808), .B(n12819), .Z(n12810) );
  XOR U14868 ( .A(n12820), .B(n12821), .Z(n12808) );
  AND U14869 ( .A(n12822), .B(n12823), .Z(n12821) );
  XNOR U14870 ( .A(n12824), .B(n12820), .Z(n12823) );
  XOR U14871 ( .A(n12825), .B(nreg[982]), .Z(n12816) );
  IV U14872 ( .A(n12814), .Z(n12825) );
  XOR U14873 ( .A(n12826), .B(n12827), .Z(n12814) );
  AND U14874 ( .A(n12828), .B(n12829), .Z(n12827) );
  XNOR U14875 ( .A(n12826), .B(n6415), .Z(n12829) );
  XNOR U14876 ( .A(n12822), .B(n12824), .Z(n6415) );
  NAND U14877 ( .A(n12830), .B(nreg[981]), .Z(n12824) );
  NAND U14878 ( .A(n12326), .B(nreg[981]), .Z(n12830) );
  XNOR U14879 ( .A(n12820), .B(n12831), .Z(n12822) );
  XOR U14880 ( .A(n12832), .B(n12833), .Z(n12820) );
  AND U14881 ( .A(n12834), .B(n12835), .Z(n12833) );
  XNOR U14882 ( .A(n12836), .B(n12832), .Z(n12835) );
  XOR U14883 ( .A(n12837), .B(nreg[981]), .Z(n12828) );
  IV U14884 ( .A(n12826), .Z(n12837) );
  XOR U14885 ( .A(n12838), .B(n12839), .Z(n12826) );
  AND U14886 ( .A(n12840), .B(n12841), .Z(n12839) );
  XNOR U14887 ( .A(n12838), .B(n6421), .Z(n12841) );
  XNOR U14888 ( .A(n12834), .B(n12836), .Z(n6421) );
  NAND U14889 ( .A(n12842), .B(nreg[980]), .Z(n12836) );
  NAND U14890 ( .A(n12326), .B(nreg[980]), .Z(n12842) );
  XNOR U14891 ( .A(n12832), .B(n12843), .Z(n12834) );
  XOR U14892 ( .A(n12844), .B(n12845), .Z(n12832) );
  AND U14893 ( .A(n12846), .B(n12847), .Z(n12845) );
  XNOR U14894 ( .A(n12848), .B(n12844), .Z(n12847) );
  XOR U14895 ( .A(n12849), .B(nreg[980]), .Z(n12840) );
  IV U14896 ( .A(n12838), .Z(n12849) );
  XOR U14897 ( .A(n12850), .B(n12851), .Z(n12838) );
  AND U14898 ( .A(n12852), .B(n12853), .Z(n12851) );
  XNOR U14899 ( .A(n12850), .B(n6427), .Z(n12853) );
  XNOR U14900 ( .A(n12846), .B(n12848), .Z(n6427) );
  NAND U14901 ( .A(n12854), .B(nreg[979]), .Z(n12848) );
  NAND U14902 ( .A(n12326), .B(nreg[979]), .Z(n12854) );
  XNOR U14903 ( .A(n12844), .B(n12855), .Z(n12846) );
  XOR U14904 ( .A(n12856), .B(n12857), .Z(n12844) );
  AND U14905 ( .A(n12858), .B(n12859), .Z(n12857) );
  XNOR U14906 ( .A(n12860), .B(n12856), .Z(n12859) );
  XOR U14907 ( .A(n12861), .B(nreg[979]), .Z(n12852) );
  IV U14908 ( .A(n12850), .Z(n12861) );
  XOR U14909 ( .A(n12862), .B(n12863), .Z(n12850) );
  AND U14910 ( .A(n12864), .B(n12865), .Z(n12863) );
  XNOR U14911 ( .A(n12862), .B(n6433), .Z(n12865) );
  XNOR U14912 ( .A(n12858), .B(n12860), .Z(n6433) );
  NAND U14913 ( .A(n12866), .B(nreg[978]), .Z(n12860) );
  NAND U14914 ( .A(n12326), .B(nreg[978]), .Z(n12866) );
  XNOR U14915 ( .A(n12856), .B(n12867), .Z(n12858) );
  XOR U14916 ( .A(n12868), .B(n12869), .Z(n12856) );
  AND U14917 ( .A(n12870), .B(n12871), .Z(n12869) );
  XNOR U14918 ( .A(n12872), .B(n12868), .Z(n12871) );
  XOR U14919 ( .A(n12873), .B(nreg[978]), .Z(n12864) );
  IV U14920 ( .A(n12862), .Z(n12873) );
  XOR U14921 ( .A(n12874), .B(n12875), .Z(n12862) );
  AND U14922 ( .A(n12876), .B(n12877), .Z(n12875) );
  XNOR U14923 ( .A(n12874), .B(n6439), .Z(n12877) );
  XNOR U14924 ( .A(n12870), .B(n12872), .Z(n6439) );
  NAND U14925 ( .A(n12878), .B(nreg[977]), .Z(n12872) );
  NAND U14926 ( .A(n12326), .B(nreg[977]), .Z(n12878) );
  XNOR U14927 ( .A(n12868), .B(n12879), .Z(n12870) );
  XOR U14928 ( .A(n12880), .B(n12881), .Z(n12868) );
  AND U14929 ( .A(n12882), .B(n12883), .Z(n12881) );
  XNOR U14930 ( .A(n12884), .B(n12880), .Z(n12883) );
  XOR U14931 ( .A(n12885), .B(nreg[977]), .Z(n12876) );
  IV U14932 ( .A(n12874), .Z(n12885) );
  XOR U14933 ( .A(n12886), .B(n12887), .Z(n12874) );
  AND U14934 ( .A(n12888), .B(n12889), .Z(n12887) );
  XNOR U14935 ( .A(n12886), .B(n6445), .Z(n12889) );
  XNOR U14936 ( .A(n12882), .B(n12884), .Z(n6445) );
  NAND U14937 ( .A(n12890), .B(nreg[976]), .Z(n12884) );
  NAND U14938 ( .A(n12326), .B(nreg[976]), .Z(n12890) );
  XNOR U14939 ( .A(n12880), .B(n12891), .Z(n12882) );
  XOR U14940 ( .A(n12892), .B(n12893), .Z(n12880) );
  AND U14941 ( .A(n12894), .B(n12895), .Z(n12893) );
  XNOR U14942 ( .A(n12896), .B(n12892), .Z(n12895) );
  XOR U14943 ( .A(n12897), .B(nreg[976]), .Z(n12888) );
  IV U14944 ( .A(n12886), .Z(n12897) );
  XOR U14945 ( .A(n12898), .B(n12899), .Z(n12886) );
  AND U14946 ( .A(n12900), .B(n12901), .Z(n12899) );
  XNOR U14947 ( .A(n12898), .B(n6451), .Z(n12901) );
  XNOR U14948 ( .A(n12894), .B(n12896), .Z(n6451) );
  NAND U14949 ( .A(n12902), .B(nreg[975]), .Z(n12896) );
  NAND U14950 ( .A(n12326), .B(nreg[975]), .Z(n12902) );
  XNOR U14951 ( .A(n12892), .B(n12903), .Z(n12894) );
  XOR U14952 ( .A(n12904), .B(n12905), .Z(n12892) );
  AND U14953 ( .A(n12906), .B(n12907), .Z(n12905) );
  XNOR U14954 ( .A(n12908), .B(n12904), .Z(n12907) );
  XOR U14955 ( .A(n12909), .B(nreg[975]), .Z(n12900) );
  IV U14956 ( .A(n12898), .Z(n12909) );
  XOR U14957 ( .A(n12910), .B(n12911), .Z(n12898) );
  AND U14958 ( .A(n12912), .B(n12913), .Z(n12911) );
  XNOR U14959 ( .A(n12910), .B(n6457), .Z(n12913) );
  XNOR U14960 ( .A(n12906), .B(n12908), .Z(n6457) );
  NAND U14961 ( .A(n12914), .B(nreg[974]), .Z(n12908) );
  NAND U14962 ( .A(n12326), .B(nreg[974]), .Z(n12914) );
  XNOR U14963 ( .A(n12904), .B(n12915), .Z(n12906) );
  XOR U14964 ( .A(n12916), .B(n12917), .Z(n12904) );
  AND U14965 ( .A(n12918), .B(n12919), .Z(n12917) );
  XNOR U14966 ( .A(n12920), .B(n12916), .Z(n12919) );
  XOR U14967 ( .A(n12921), .B(nreg[974]), .Z(n12912) );
  IV U14968 ( .A(n12910), .Z(n12921) );
  XOR U14969 ( .A(n12922), .B(n12923), .Z(n12910) );
  AND U14970 ( .A(n12924), .B(n12925), .Z(n12923) );
  XNOR U14971 ( .A(n12922), .B(n6463), .Z(n12925) );
  XNOR U14972 ( .A(n12918), .B(n12920), .Z(n6463) );
  NAND U14973 ( .A(n12926), .B(nreg[973]), .Z(n12920) );
  NAND U14974 ( .A(n12326), .B(nreg[973]), .Z(n12926) );
  XNOR U14975 ( .A(n12916), .B(n12927), .Z(n12918) );
  XOR U14976 ( .A(n12928), .B(n12929), .Z(n12916) );
  AND U14977 ( .A(n12930), .B(n12931), .Z(n12929) );
  XNOR U14978 ( .A(n12932), .B(n12928), .Z(n12931) );
  XOR U14979 ( .A(n12933), .B(nreg[973]), .Z(n12924) );
  IV U14980 ( .A(n12922), .Z(n12933) );
  XOR U14981 ( .A(n12934), .B(n12935), .Z(n12922) );
  AND U14982 ( .A(n12936), .B(n12937), .Z(n12935) );
  XNOR U14983 ( .A(n12934), .B(n6469), .Z(n12937) );
  XNOR U14984 ( .A(n12930), .B(n12932), .Z(n6469) );
  NAND U14985 ( .A(n12938), .B(nreg[972]), .Z(n12932) );
  NAND U14986 ( .A(n12326), .B(nreg[972]), .Z(n12938) );
  XNOR U14987 ( .A(n12928), .B(n12939), .Z(n12930) );
  XOR U14988 ( .A(n12940), .B(n12941), .Z(n12928) );
  AND U14989 ( .A(n12942), .B(n12943), .Z(n12941) );
  XNOR U14990 ( .A(n12944), .B(n12940), .Z(n12943) );
  XOR U14991 ( .A(n12945), .B(nreg[972]), .Z(n12936) );
  IV U14992 ( .A(n12934), .Z(n12945) );
  XOR U14993 ( .A(n12946), .B(n12947), .Z(n12934) );
  AND U14994 ( .A(n12948), .B(n12949), .Z(n12947) );
  XNOR U14995 ( .A(n12946), .B(n6475), .Z(n12949) );
  XNOR U14996 ( .A(n12942), .B(n12944), .Z(n6475) );
  NAND U14997 ( .A(n12950), .B(nreg[971]), .Z(n12944) );
  NAND U14998 ( .A(n12326), .B(nreg[971]), .Z(n12950) );
  XNOR U14999 ( .A(n12940), .B(n12951), .Z(n12942) );
  XOR U15000 ( .A(n12952), .B(n12953), .Z(n12940) );
  AND U15001 ( .A(n12954), .B(n12955), .Z(n12953) );
  XNOR U15002 ( .A(n12956), .B(n12952), .Z(n12955) );
  XOR U15003 ( .A(n12957), .B(nreg[971]), .Z(n12948) );
  IV U15004 ( .A(n12946), .Z(n12957) );
  XOR U15005 ( .A(n12958), .B(n12959), .Z(n12946) );
  AND U15006 ( .A(n12960), .B(n12961), .Z(n12959) );
  XNOR U15007 ( .A(n12958), .B(n6481), .Z(n12961) );
  XNOR U15008 ( .A(n12954), .B(n12956), .Z(n6481) );
  NAND U15009 ( .A(n12962), .B(nreg[970]), .Z(n12956) );
  NAND U15010 ( .A(n12326), .B(nreg[970]), .Z(n12962) );
  XNOR U15011 ( .A(n12952), .B(n12963), .Z(n12954) );
  XOR U15012 ( .A(n12964), .B(n12965), .Z(n12952) );
  AND U15013 ( .A(n12966), .B(n12967), .Z(n12965) );
  XNOR U15014 ( .A(n12968), .B(n12964), .Z(n12967) );
  XOR U15015 ( .A(n12969), .B(nreg[970]), .Z(n12960) );
  IV U15016 ( .A(n12958), .Z(n12969) );
  XOR U15017 ( .A(n12970), .B(n12971), .Z(n12958) );
  AND U15018 ( .A(n12972), .B(n12973), .Z(n12971) );
  XNOR U15019 ( .A(n12970), .B(n6487), .Z(n12973) );
  XNOR U15020 ( .A(n12966), .B(n12968), .Z(n6487) );
  NAND U15021 ( .A(n12974), .B(nreg[969]), .Z(n12968) );
  NAND U15022 ( .A(n12326), .B(nreg[969]), .Z(n12974) );
  XNOR U15023 ( .A(n12964), .B(n12975), .Z(n12966) );
  XOR U15024 ( .A(n12976), .B(n12977), .Z(n12964) );
  AND U15025 ( .A(n12978), .B(n12979), .Z(n12977) );
  XNOR U15026 ( .A(n12980), .B(n12976), .Z(n12979) );
  XOR U15027 ( .A(n12981), .B(nreg[969]), .Z(n12972) );
  IV U15028 ( .A(n12970), .Z(n12981) );
  XOR U15029 ( .A(n12982), .B(n12983), .Z(n12970) );
  AND U15030 ( .A(n12984), .B(n12985), .Z(n12983) );
  XNOR U15031 ( .A(n12982), .B(n6493), .Z(n12985) );
  XNOR U15032 ( .A(n12978), .B(n12980), .Z(n6493) );
  NAND U15033 ( .A(n12986), .B(nreg[968]), .Z(n12980) );
  NAND U15034 ( .A(n12326), .B(nreg[968]), .Z(n12986) );
  XNOR U15035 ( .A(n12976), .B(n12987), .Z(n12978) );
  XOR U15036 ( .A(n12988), .B(n12989), .Z(n12976) );
  AND U15037 ( .A(n12990), .B(n12991), .Z(n12989) );
  XNOR U15038 ( .A(n12992), .B(n12988), .Z(n12991) );
  XOR U15039 ( .A(n12993), .B(nreg[968]), .Z(n12984) );
  IV U15040 ( .A(n12982), .Z(n12993) );
  XOR U15041 ( .A(n12994), .B(n12995), .Z(n12982) );
  AND U15042 ( .A(n12996), .B(n12997), .Z(n12995) );
  XNOR U15043 ( .A(n12994), .B(n6499), .Z(n12997) );
  XNOR U15044 ( .A(n12990), .B(n12992), .Z(n6499) );
  NAND U15045 ( .A(n12998), .B(nreg[967]), .Z(n12992) );
  NAND U15046 ( .A(n12326), .B(nreg[967]), .Z(n12998) );
  XNOR U15047 ( .A(n12988), .B(n12999), .Z(n12990) );
  XOR U15048 ( .A(n13000), .B(n13001), .Z(n12988) );
  AND U15049 ( .A(n13002), .B(n13003), .Z(n13001) );
  XNOR U15050 ( .A(n13004), .B(n13000), .Z(n13003) );
  XOR U15051 ( .A(n13005), .B(nreg[967]), .Z(n12996) );
  IV U15052 ( .A(n12994), .Z(n13005) );
  XOR U15053 ( .A(n13006), .B(n13007), .Z(n12994) );
  AND U15054 ( .A(n13008), .B(n13009), .Z(n13007) );
  XNOR U15055 ( .A(n13006), .B(n6505), .Z(n13009) );
  XNOR U15056 ( .A(n13002), .B(n13004), .Z(n6505) );
  NAND U15057 ( .A(n13010), .B(nreg[966]), .Z(n13004) );
  NAND U15058 ( .A(n12326), .B(nreg[966]), .Z(n13010) );
  XNOR U15059 ( .A(n13000), .B(n13011), .Z(n13002) );
  XOR U15060 ( .A(n13012), .B(n13013), .Z(n13000) );
  AND U15061 ( .A(n13014), .B(n13015), .Z(n13013) );
  XNOR U15062 ( .A(n13016), .B(n13012), .Z(n13015) );
  XOR U15063 ( .A(n13017), .B(nreg[966]), .Z(n13008) );
  IV U15064 ( .A(n13006), .Z(n13017) );
  XOR U15065 ( .A(n13018), .B(n13019), .Z(n13006) );
  AND U15066 ( .A(n13020), .B(n13021), .Z(n13019) );
  XNOR U15067 ( .A(n13018), .B(n6511), .Z(n13021) );
  XNOR U15068 ( .A(n13014), .B(n13016), .Z(n6511) );
  NAND U15069 ( .A(n13022), .B(nreg[965]), .Z(n13016) );
  NAND U15070 ( .A(n12326), .B(nreg[965]), .Z(n13022) );
  XNOR U15071 ( .A(n13012), .B(n13023), .Z(n13014) );
  XOR U15072 ( .A(n13024), .B(n13025), .Z(n13012) );
  AND U15073 ( .A(n13026), .B(n13027), .Z(n13025) );
  XNOR U15074 ( .A(n13028), .B(n13024), .Z(n13027) );
  XOR U15075 ( .A(n13029), .B(nreg[965]), .Z(n13020) );
  IV U15076 ( .A(n13018), .Z(n13029) );
  XOR U15077 ( .A(n13030), .B(n13031), .Z(n13018) );
  AND U15078 ( .A(n13032), .B(n13033), .Z(n13031) );
  XNOR U15079 ( .A(n13030), .B(n6517), .Z(n13033) );
  XNOR U15080 ( .A(n13026), .B(n13028), .Z(n6517) );
  NAND U15081 ( .A(n13034), .B(nreg[964]), .Z(n13028) );
  NAND U15082 ( .A(n12326), .B(nreg[964]), .Z(n13034) );
  XNOR U15083 ( .A(n13024), .B(n13035), .Z(n13026) );
  XOR U15084 ( .A(n13036), .B(n13037), .Z(n13024) );
  AND U15085 ( .A(n13038), .B(n13039), .Z(n13037) );
  XNOR U15086 ( .A(n13040), .B(n13036), .Z(n13039) );
  XOR U15087 ( .A(n13041), .B(nreg[964]), .Z(n13032) );
  IV U15088 ( .A(n13030), .Z(n13041) );
  XOR U15089 ( .A(n13042), .B(n13043), .Z(n13030) );
  AND U15090 ( .A(n13044), .B(n13045), .Z(n13043) );
  XNOR U15091 ( .A(n13042), .B(n6523), .Z(n13045) );
  XNOR U15092 ( .A(n13038), .B(n13040), .Z(n6523) );
  NAND U15093 ( .A(n13046), .B(nreg[963]), .Z(n13040) );
  NAND U15094 ( .A(n12326), .B(nreg[963]), .Z(n13046) );
  XNOR U15095 ( .A(n13036), .B(n13047), .Z(n13038) );
  XOR U15096 ( .A(n13048), .B(n13049), .Z(n13036) );
  AND U15097 ( .A(n13050), .B(n13051), .Z(n13049) );
  XNOR U15098 ( .A(n13052), .B(n13048), .Z(n13051) );
  XOR U15099 ( .A(n13053), .B(nreg[963]), .Z(n13044) );
  IV U15100 ( .A(n13042), .Z(n13053) );
  XOR U15101 ( .A(n13054), .B(n13055), .Z(n13042) );
  AND U15102 ( .A(n13056), .B(n13057), .Z(n13055) );
  XNOR U15103 ( .A(n13054), .B(n6529), .Z(n13057) );
  XNOR U15104 ( .A(n13050), .B(n13052), .Z(n6529) );
  NAND U15105 ( .A(n13058), .B(nreg[962]), .Z(n13052) );
  NAND U15106 ( .A(n12326), .B(nreg[962]), .Z(n13058) );
  XNOR U15107 ( .A(n13048), .B(n13059), .Z(n13050) );
  XOR U15108 ( .A(n13060), .B(n13061), .Z(n13048) );
  AND U15109 ( .A(n13062), .B(n13063), .Z(n13061) );
  XNOR U15110 ( .A(n13064), .B(n13060), .Z(n13063) );
  XOR U15111 ( .A(n13065), .B(nreg[962]), .Z(n13056) );
  IV U15112 ( .A(n13054), .Z(n13065) );
  XOR U15113 ( .A(n13066), .B(n13067), .Z(n13054) );
  AND U15114 ( .A(n13068), .B(n13069), .Z(n13067) );
  XNOR U15115 ( .A(n13066), .B(n6535), .Z(n13069) );
  XNOR U15116 ( .A(n13062), .B(n13064), .Z(n6535) );
  NAND U15117 ( .A(n13070), .B(nreg[961]), .Z(n13064) );
  NAND U15118 ( .A(n12326), .B(nreg[961]), .Z(n13070) );
  XNOR U15119 ( .A(n13060), .B(n13071), .Z(n13062) );
  XOR U15120 ( .A(n13072), .B(n13073), .Z(n13060) );
  AND U15121 ( .A(n13074), .B(n13075), .Z(n13073) );
  XNOR U15122 ( .A(n13076), .B(n13072), .Z(n13075) );
  XOR U15123 ( .A(n13077), .B(nreg[961]), .Z(n13068) );
  IV U15124 ( .A(n13066), .Z(n13077) );
  XOR U15125 ( .A(n13078), .B(n13079), .Z(n13066) );
  AND U15126 ( .A(n13080), .B(n13081), .Z(n13079) );
  XNOR U15127 ( .A(n13078), .B(n6541), .Z(n13081) );
  XNOR U15128 ( .A(n13074), .B(n13076), .Z(n6541) );
  NAND U15129 ( .A(n13082), .B(nreg[960]), .Z(n13076) );
  NAND U15130 ( .A(n12326), .B(nreg[960]), .Z(n13082) );
  XNOR U15131 ( .A(n13072), .B(n13083), .Z(n13074) );
  XOR U15132 ( .A(n13084), .B(n13085), .Z(n13072) );
  AND U15133 ( .A(n13086), .B(n13087), .Z(n13085) );
  XNOR U15134 ( .A(n13088), .B(n13084), .Z(n13087) );
  XOR U15135 ( .A(n13089), .B(nreg[960]), .Z(n13080) );
  IV U15136 ( .A(n13078), .Z(n13089) );
  XOR U15137 ( .A(n13090), .B(n13091), .Z(n13078) );
  AND U15138 ( .A(n13092), .B(n13093), .Z(n13091) );
  XNOR U15139 ( .A(n13090), .B(n6547), .Z(n13093) );
  XNOR U15140 ( .A(n13086), .B(n13088), .Z(n6547) );
  NAND U15141 ( .A(n13094), .B(nreg[959]), .Z(n13088) );
  NAND U15142 ( .A(n12326), .B(nreg[959]), .Z(n13094) );
  XNOR U15143 ( .A(n13084), .B(n13095), .Z(n13086) );
  XOR U15144 ( .A(n13096), .B(n13097), .Z(n13084) );
  AND U15145 ( .A(n13098), .B(n13099), .Z(n13097) );
  XNOR U15146 ( .A(n13100), .B(n13096), .Z(n13099) );
  XOR U15147 ( .A(n13101), .B(nreg[959]), .Z(n13092) );
  IV U15148 ( .A(n13090), .Z(n13101) );
  XOR U15149 ( .A(n13102), .B(n13103), .Z(n13090) );
  AND U15150 ( .A(n13104), .B(n13105), .Z(n13103) );
  XNOR U15151 ( .A(n13102), .B(n6553), .Z(n13105) );
  XNOR U15152 ( .A(n13098), .B(n13100), .Z(n6553) );
  NAND U15153 ( .A(n13106), .B(nreg[958]), .Z(n13100) );
  NAND U15154 ( .A(n12326), .B(nreg[958]), .Z(n13106) );
  XNOR U15155 ( .A(n13096), .B(n13107), .Z(n13098) );
  XOR U15156 ( .A(n13108), .B(n13109), .Z(n13096) );
  AND U15157 ( .A(n13110), .B(n13111), .Z(n13109) );
  XNOR U15158 ( .A(n13112), .B(n13108), .Z(n13111) );
  XOR U15159 ( .A(n13113), .B(nreg[958]), .Z(n13104) );
  IV U15160 ( .A(n13102), .Z(n13113) );
  XOR U15161 ( .A(n13114), .B(n13115), .Z(n13102) );
  AND U15162 ( .A(n13116), .B(n13117), .Z(n13115) );
  XNOR U15163 ( .A(n13114), .B(n6559), .Z(n13117) );
  XNOR U15164 ( .A(n13110), .B(n13112), .Z(n6559) );
  NAND U15165 ( .A(n13118), .B(nreg[957]), .Z(n13112) );
  NAND U15166 ( .A(n12326), .B(nreg[957]), .Z(n13118) );
  XNOR U15167 ( .A(n13108), .B(n13119), .Z(n13110) );
  XOR U15168 ( .A(n13120), .B(n13121), .Z(n13108) );
  AND U15169 ( .A(n13122), .B(n13123), .Z(n13121) );
  XNOR U15170 ( .A(n13124), .B(n13120), .Z(n13123) );
  XOR U15171 ( .A(n13125), .B(nreg[957]), .Z(n13116) );
  IV U15172 ( .A(n13114), .Z(n13125) );
  XOR U15173 ( .A(n13126), .B(n13127), .Z(n13114) );
  AND U15174 ( .A(n13128), .B(n13129), .Z(n13127) );
  XNOR U15175 ( .A(n13126), .B(n6565), .Z(n13129) );
  XNOR U15176 ( .A(n13122), .B(n13124), .Z(n6565) );
  NAND U15177 ( .A(n13130), .B(nreg[956]), .Z(n13124) );
  NAND U15178 ( .A(n12326), .B(nreg[956]), .Z(n13130) );
  XNOR U15179 ( .A(n13120), .B(n13131), .Z(n13122) );
  XOR U15180 ( .A(n13132), .B(n13133), .Z(n13120) );
  AND U15181 ( .A(n13134), .B(n13135), .Z(n13133) );
  XNOR U15182 ( .A(n13136), .B(n13132), .Z(n13135) );
  XOR U15183 ( .A(n13137), .B(nreg[956]), .Z(n13128) );
  IV U15184 ( .A(n13126), .Z(n13137) );
  XOR U15185 ( .A(n13138), .B(n13139), .Z(n13126) );
  AND U15186 ( .A(n13140), .B(n13141), .Z(n13139) );
  XNOR U15187 ( .A(n13138), .B(n6571), .Z(n13141) );
  XNOR U15188 ( .A(n13134), .B(n13136), .Z(n6571) );
  NAND U15189 ( .A(n13142), .B(nreg[955]), .Z(n13136) );
  NAND U15190 ( .A(n12326), .B(nreg[955]), .Z(n13142) );
  XNOR U15191 ( .A(n13132), .B(n13143), .Z(n13134) );
  XOR U15192 ( .A(n13144), .B(n13145), .Z(n13132) );
  AND U15193 ( .A(n13146), .B(n13147), .Z(n13145) );
  XNOR U15194 ( .A(n13148), .B(n13144), .Z(n13147) );
  XOR U15195 ( .A(n13149), .B(nreg[955]), .Z(n13140) );
  IV U15196 ( .A(n13138), .Z(n13149) );
  XOR U15197 ( .A(n13150), .B(n13151), .Z(n13138) );
  AND U15198 ( .A(n13152), .B(n13153), .Z(n13151) );
  XNOR U15199 ( .A(n13150), .B(n6577), .Z(n13153) );
  XNOR U15200 ( .A(n13146), .B(n13148), .Z(n6577) );
  NAND U15201 ( .A(n13154), .B(nreg[954]), .Z(n13148) );
  NAND U15202 ( .A(n12326), .B(nreg[954]), .Z(n13154) );
  XNOR U15203 ( .A(n13144), .B(n13155), .Z(n13146) );
  XOR U15204 ( .A(n13156), .B(n13157), .Z(n13144) );
  AND U15205 ( .A(n13158), .B(n13159), .Z(n13157) );
  XNOR U15206 ( .A(n13160), .B(n13156), .Z(n13159) );
  XOR U15207 ( .A(n13161), .B(nreg[954]), .Z(n13152) );
  IV U15208 ( .A(n13150), .Z(n13161) );
  XOR U15209 ( .A(n13162), .B(n13163), .Z(n13150) );
  AND U15210 ( .A(n13164), .B(n13165), .Z(n13163) );
  XNOR U15211 ( .A(n13162), .B(n6583), .Z(n13165) );
  XNOR U15212 ( .A(n13158), .B(n13160), .Z(n6583) );
  NAND U15213 ( .A(n13166), .B(nreg[953]), .Z(n13160) );
  NAND U15214 ( .A(n12326), .B(nreg[953]), .Z(n13166) );
  XNOR U15215 ( .A(n13156), .B(n13167), .Z(n13158) );
  XOR U15216 ( .A(n13168), .B(n13169), .Z(n13156) );
  AND U15217 ( .A(n13170), .B(n13171), .Z(n13169) );
  XNOR U15218 ( .A(n13172), .B(n13168), .Z(n13171) );
  XOR U15219 ( .A(n13173), .B(nreg[953]), .Z(n13164) );
  IV U15220 ( .A(n13162), .Z(n13173) );
  XOR U15221 ( .A(n13174), .B(n13175), .Z(n13162) );
  AND U15222 ( .A(n13176), .B(n13177), .Z(n13175) );
  XNOR U15223 ( .A(n13174), .B(n6589), .Z(n13177) );
  XNOR U15224 ( .A(n13170), .B(n13172), .Z(n6589) );
  NAND U15225 ( .A(n13178), .B(nreg[952]), .Z(n13172) );
  NAND U15226 ( .A(n12326), .B(nreg[952]), .Z(n13178) );
  XNOR U15227 ( .A(n13168), .B(n13179), .Z(n13170) );
  XOR U15228 ( .A(n13180), .B(n13181), .Z(n13168) );
  AND U15229 ( .A(n13182), .B(n13183), .Z(n13181) );
  XNOR U15230 ( .A(n13184), .B(n13180), .Z(n13183) );
  XOR U15231 ( .A(n13185), .B(nreg[952]), .Z(n13176) );
  IV U15232 ( .A(n13174), .Z(n13185) );
  XOR U15233 ( .A(n13186), .B(n13187), .Z(n13174) );
  AND U15234 ( .A(n13188), .B(n13189), .Z(n13187) );
  XNOR U15235 ( .A(n13186), .B(n6595), .Z(n13189) );
  XNOR U15236 ( .A(n13182), .B(n13184), .Z(n6595) );
  NAND U15237 ( .A(n13190), .B(nreg[951]), .Z(n13184) );
  NAND U15238 ( .A(n12326), .B(nreg[951]), .Z(n13190) );
  XNOR U15239 ( .A(n13180), .B(n13191), .Z(n13182) );
  XOR U15240 ( .A(n13192), .B(n13193), .Z(n13180) );
  AND U15241 ( .A(n13194), .B(n13195), .Z(n13193) );
  XNOR U15242 ( .A(n13196), .B(n13192), .Z(n13195) );
  XOR U15243 ( .A(n13197), .B(nreg[951]), .Z(n13188) );
  IV U15244 ( .A(n13186), .Z(n13197) );
  XOR U15245 ( .A(n13198), .B(n13199), .Z(n13186) );
  AND U15246 ( .A(n13200), .B(n13201), .Z(n13199) );
  XNOR U15247 ( .A(n13198), .B(n6601), .Z(n13201) );
  XNOR U15248 ( .A(n13194), .B(n13196), .Z(n6601) );
  NAND U15249 ( .A(n13202), .B(nreg[950]), .Z(n13196) );
  NAND U15250 ( .A(n12326), .B(nreg[950]), .Z(n13202) );
  XNOR U15251 ( .A(n13192), .B(n13203), .Z(n13194) );
  XOR U15252 ( .A(n13204), .B(n13205), .Z(n13192) );
  AND U15253 ( .A(n13206), .B(n13207), .Z(n13205) );
  XNOR U15254 ( .A(n13208), .B(n13204), .Z(n13207) );
  XOR U15255 ( .A(n13209), .B(nreg[950]), .Z(n13200) );
  IV U15256 ( .A(n13198), .Z(n13209) );
  XOR U15257 ( .A(n13210), .B(n13211), .Z(n13198) );
  AND U15258 ( .A(n13212), .B(n13213), .Z(n13211) );
  XNOR U15259 ( .A(n13210), .B(n6607), .Z(n13213) );
  XNOR U15260 ( .A(n13206), .B(n13208), .Z(n6607) );
  NAND U15261 ( .A(n13214), .B(nreg[949]), .Z(n13208) );
  NAND U15262 ( .A(n12326), .B(nreg[949]), .Z(n13214) );
  XNOR U15263 ( .A(n13204), .B(n13215), .Z(n13206) );
  XOR U15264 ( .A(n13216), .B(n13217), .Z(n13204) );
  AND U15265 ( .A(n13218), .B(n13219), .Z(n13217) );
  XNOR U15266 ( .A(n13220), .B(n13216), .Z(n13219) );
  XOR U15267 ( .A(n13221), .B(nreg[949]), .Z(n13212) );
  IV U15268 ( .A(n13210), .Z(n13221) );
  XOR U15269 ( .A(n13222), .B(n13223), .Z(n13210) );
  AND U15270 ( .A(n13224), .B(n13225), .Z(n13223) );
  XNOR U15271 ( .A(n13222), .B(n6613), .Z(n13225) );
  XNOR U15272 ( .A(n13218), .B(n13220), .Z(n6613) );
  NAND U15273 ( .A(n13226), .B(nreg[948]), .Z(n13220) );
  NAND U15274 ( .A(n12326), .B(nreg[948]), .Z(n13226) );
  XNOR U15275 ( .A(n13216), .B(n13227), .Z(n13218) );
  XOR U15276 ( .A(n13228), .B(n13229), .Z(n13216) );
  AND U15277 ( .A(n13230), .B(n13231), .Z(n13229) );
  XNOR U15278 ( .A(n13232), .B(n13228), .Z(n13231) );
  XOR U15279 ( .A(n13233), .B(nreg[948]), .Z(n13224) );
  IV U15280 ( .A(n13222), .Z(n13233) );
  XOR U15281 ( .A(n13234), .B(n13235), .Z(n13222) );
  AND U15282 ( .A(n13236), .B(n13237), .Z(n13235) );
  XNOR U15283 ( .A(n13234), .B(n6619), .Z(n13237) );
  XNOR U15284 ( .A(n13230), .B(n13232), .Z(n6619) );
  NAND U15285 ( .A(n13238), .B(nreg[947]), .Z(n13232) );
  NAND U15286 ( .A(n12326), .B(nreg[947]), .Z(n13238) );
  XNOR U15287 ( .A(n13228), .B(n13239), .Z(n13230) );
  XOR U15288 ( .A(n13240), .B(n13241), .Z(n13228) );
  AND U15289 ( .A(n13242), .B(n13243), .Z(n13241) );
  XNOR U15290 ( .A(n13244), .B(n13240), .Z(n13243) );
  XOR U15291 ( .A(n13245), .B(nreg[947]), .Z(n13236) );
  IV U15292 ( .A(n13234), .Z(n13245) );
  XOR U15293 ( .A(n13246), .B(n13247), .Z(n13234) );
  AND U15294 ( .A(n13248), .B(n13249), .Z(n13247) );
  XNOR U15295 ( .A(n13246), .B(n6625), .Z(n13249) );
  XNOR U15296 ( .A(n13242), .B(n13244), .Z(n6625) );
  NAND U15297 ( .A(n13250), .B(nreg[946]), .Z(n13244) );
  NAND U15298 ( .A(n12326), .B(nreg[946]), .Z(n13250) );
  XNOR U15299 ( .A(n13240), .B(n13251), .Z(n13242) );
  XOR U15300 ( .A(n13252), .B(n13253), .Z(n13240) );
  AND U15301 ( .A(n13254), .B(n13255), .Z(n13253) );
  XNOR U15302 ( .A(n13256), .B(n13252), .Z(n13255) );
  XOR U15303 ( .A(n13257), .B(nreg[946]), .Z(n13248) );
  IV U15304 ( .A(n13246), .Z(n13257) );
  XOR U15305 ( .A(n13258), .B(n13259), .Z(n13246) );
  AND U15306 ( .A(n13260), .B(n13261), .Z(n13259) );
  XNOR U15307 ( .A(n13258), .B(n6631), .Z(n13261) );
  XNOR U15308 ( .A(n13254), .B(n13256), .Z(n6631) );
  NAND U15309 ( .A(n13262), .B(nreg[945]), .Z(n13256) );
  NAND U15310 ( .A(n12326), .B(nreg[945]), .Z(n13262) );
  XNOR U15311 ( .A(n13252), .B(n13263), .Z(n13254) );
  XOR U15312 ( .A(n13264), .B(n13265), .Z(n13252) );
  AND U15313 ( .A(n13266), .B(n13267), .Z(n13265) );
  XNOR U15314 ( .A(n13268), .B(n13264), .Z(n13267) );
  XOR U15315 ( .A(n13269), .B(nreg[945]), .Z(n13260) );
  IV U15316 ( .A(n13258), .Z(n13269) );
  XOR U15317 ( .A(n13270), .B(n13271), .Z(n13258) );
  AND U15318 ( .A(n13272), .B(n13273), .Z(n13271) );
  XNOR U15319 ( .A(n13270), .B(n6637), .Z(n13273) );
  XNOR U15320 ( .A(n13266), .B(n13268), .Z(n6637) );
  NAND U15321 ( .A(n13274), .B(nreg[944]), .Z(n13268) );
  NAND U15322 ( .A(n12326), .B(nreg[944]), .Z(n13274) );
  XNOR U15323 ( .A(n13264), .B(n13275), .Z(n13266) );
  XOR U15324 ( .A(n13276), .B(n13277), .Z(n13264) );
  AND U15325 ( .A(n13278), .B(n13279), .Z(n13277) );
  XNOR U15326 ( .A(n13280), .B(n13276), .Z(n13279) );
  XOR U15327 ( .A(n13281), .B(nreg[944]), .Z(n13272) );
  IV U15328 ( .A(n13270), .Z(n13281) );
  XOR U15329 ( .A(n13282), .B(n13283), .Z(n13270) );
  AND U15330 ( .A(n13284), .B(n13285), .Z(n13283) );
  XNOR U15331 ( .A(n13282), .B(n6643), .Z(n13285) );
  XNOR U15332 ( .A(n13278), .B(n13280), .Z(n6643) );
  NAND U15333 ( .A(n13286), .B(nreg[943]), .Z(n13280) );
  NAND U15334 ( .A(n12326), .B(nreg[943]), .Z(n13286) );
  XNOR U15335 ( .A(n13276), .B(n13287), .Z(n13278) );
  XOR U15336 ( .A(n13288), .B(n13289), .Z(n13276) );
  AND U15337 ( .A(n13290), .B(n13291), .Z(n13289) );
  XNOR U15338 ( .A(n13292), .B(n13288), .Z(n13291) );
  XOR U15339 ( .A(n13293), .B(nreg[943]), .Z(n13284) );
  IV U15340 ( .A(n13282), .Z(n13293) );
  XOR U15341 ( .A(n13294), .B(n13295), .Z(n13282) );
  AND U15342 ( .A(n13296), .B(n13297), .Z(n13295) );
  XNOR U15343 ( .A(n13294), .B(n6649), .Z(n13297) );
  XNOR U15344 ( .A(n13290), .B(n13292), .Z(n6649) );
  NAND U15345 ( .A(n13298), .B(nreg[942]), .Z(n13292) );
  NAND U15346 ( .A(n12326), .B(nreg[942]), .Z(n13298) );
  XNOR U15347 ( .A(n13288), .B(n13299), .Z(n13290) );
  XOR U15348 ( .A(n13300), .B(n13301), .Z(n13288) );
  AND U15349 ( .A(n13302), .B(n13303), .Z(n13301) );
  XNOR U15350 ( .A(n13304), .B(n13300), .Z(n13303) );
  XOR U15351 ( .A(n13305), .B(nreg[942]), .Z(n13296) );
  IV U15352 ( .A(n13294), .Z(n13305) );
  XOR U15353 ( .A(n13306), .B(n13307), .Z(n13294) );
  AND U15354 ( .A(n13308), .B(n13309), .Z(n13307) );
  XNOR U15355 ( .A(n13306), .B(n6655), .Z(n13309) );
  XNOR U15356 ( .A(n13302), .B(n13304), .Z(n6655) );
  NAND U15357 ( .A(n13310), .B(nreg[941]), .Z(n13304) );
  NAND U15358 ( .A(n12326), .B(nreg[941]), .Z(n13310) );
  XNOR U15359 ( .A(n13300), .B(n13311), .Z(n13302) );
  XOR U15360 ( .A(n13312), .B(n13313), .Z(n13300) );
  AND U15361 ( .A(n13314), .B(n13315), .Z(n13313) );
  XNOR U15362 ( .A(n13316), .B(n13312), .Z(n13315) );
  XOR U15363 ( .A(n13317), .B(nreg[941]), .Z(n13308) );
  IV U15364 ( .A(n13306), .Z(n13317) );
  XOR U15365 ( .A(n13318), .B(n13319), .Z(n13306) );
  AND U15366 ( .A(n13320), .B(n13321), .Z(n13319) );
  XNOR U15367 ( .A(n13318), .B(n6661), .Z(n13321) );
  XNOR U15368 ( .A(n13314), .B(n13316), .Z(n6661) );
  NAND U15369 ( .A(n13322), .B(nreg[940]), .Z(n13316) );
  NAND U15370 ( .A(n12326), .B(nreg[940]), .Z(n13322) );
  XNOR U15371 ( .A(n13312), .B(n13323), .Z(n13314) );
  XOR U15372 ( .A(n13324), .B(n13325), .Z(n13312) );
  AND U15373 ( .A(n13326), .B(n13327), .Z(n13325) );
  XNOR U15374 ( .A(n13328), .B(n13324), .Z(n13327) );
  XOR U15375 ( .A(n13329), .B(nreg[940]), .Z(n13320) );
  IV U15376 ( .A(n13318), .Z(n13329) );
  XOR U15377 ( .A(n13330), .B(n13331), .Z(n13318) );
  AND U15378 ( .A(n13332), .B(n13333), .Z(n13331) );
  XNOR U15379 ( .A(n13330), .B(n6667), .Z(n13333) );
  XNOR U15380 ( .A(n13326), .B(n13328), .Z(n6667) );
  NAND U15381 ( .A(n13334), .B(nreg[939]), .Z(n13328) );
  NAND U15382 ( .A(n12326), .B(nreg[939]), .Z(n13334) );
  XNOR U15383 ( .A(n13324), .B(n13335), .Z(n13326) );
  XOR U15384 ( .A(n13336), .B(n13337), .Z(n13324) );
  AND U15385 ( .A(n13338), .B(n13339), .Z(n13337) );
  XNOR U15386 ( .A(n13340), .B(n13336), .Z(n13339) );
  XOR U15387 ( .A(n13341), .B(nreg[939]), .Z(n13332) );
  IV U15388 ( .A(n13330), .Z(n13341) );
  XOR U15389 ( .A(n13342), .B(n13343), .Z(n13330) );
  AND U15390 ( .A(n13344), .B(n13345), .Z(n13343) );
  XNOR U15391 ( .A(n13342), .B(n6673), .Z(n13345) );
  XNOR U15392 ( .A(n13338), .B(n13340), .Z(n6673) );
  NAND U15393 ( .A(n13346), .B(nreg[938]), .Z(n13340) );
  NAND U15394 ( .A(n12326), .B(nreg[938]), .Z(n13346) );
  XNOR U15395 ( .A(n13336), .B(n13347), .Z(n13338) );
  XOR U15396 ( .A(n13348), .B(n13349), .Z(n13336) );
  AND U15397 ( .A(n13350), .B(n13351), .Z(n13349) );
  XNOR U15398 ( .A(n13352), .B(n13348), .Z(n13351) );
  XOR U15399 ( .A(n13353), .B(nreg[938]), .Z(n13344) );
  IV U15400 ( .A(n13342), .Z(n13353) );
  XOR U15401 ( .A(n13354), .B(n13355), .Z(n13342) );
  AND U15402 ( .A(n13356), .B(n13357), .Z(n13355) );
  XNOR U15403 ( .A(n13354), .B(n6679), .Z(n13357) );
  XNOR U15404 ( .A(n13350), .B(n13352), .Z(n6679) );
  NAND U15405 ( .A(n13358), .B(nreg[937]), .Z(n13352) );
  NAND U15406 ( .A(n12326), .B(nreg[937]), .Z(n13358) );
  XNOR U15407 ( .A(n13348), .B(n13359), .Z(n13350) );
  XOR U15408 ( .A(n13360), .B(n13361), .Z(n13348) );
  AND U15409 ( .A(n13362), .B(n13363), .Z(n13361) );
  XNOR U15410 ( .A(n13364), .B(n13360), .Z(n13363) );
  XOR U15411 ( .A(n13365), .B(nreg[937]), .Z(n13356) );
  IV U15412 ( .A(n13354), .Z(n13365) );
  XOR U15413 ( .A(n13366), .B(n13367), .Z(n13354) );
  AND U15414 ( .A(n13368), .B(n13369), .Z(n13367) );
  XNOR U15415 ( .A(n13366), .B(n6685), .Z(n13369) );
  XNOR U15416 ( .A(n13362), .B(n13364), .Z(n6685) );
  NAND U15417 ( .A(n13370), .B(nreg[936]), .Z(n13364) );
  NAND U15418 ( .A(n12326), .B(nreg[936]), .Z(n13370) );
  XNOR U15419 ( .A(n13360), .B(n13371), .Z(n13362) );
  XOR U15420 ( .A(n13372), .B(n13373), .Z(n13360) );
  AND U15421 ( .A(n13374), .B(n13375), .Z(n13373) );
  XNOR U15422 ( .A(n13376), .B(n13372), .Z(n13375) );
  XOR U15423 ( .A(n13377), .B(nreg[936]), .Z(n13368) );
  IV U15424 ( .A(n13366), .Z(n13377) );
  XOR U15425 ( .A(n13378), .B(n13379), .Z(n13366) );
  AND U15426 ( .A(n13380), .B(n13381), .Z(n13379) );
  XNOR U15427 ( .A(n13378), .B(n6691), .Z(n13381) );
  XNOR U15428 ( .A(n13374), .B(n13376), .Z(n6691) );
  NAND U15429 ( .A(n13382), .B(nreg[935]), .Z(n13376) );
  NAND U15430 ( .A(n12326), .B(nreg[935]), .Z(n13382) );
  XNOR U15431 ( .A(n13372), .B(n13383), .Z(n13374) );
  XOR U15432 ( .A(n13384), .B(n13385), .Z(n13372) );
  AND U15433 ( .A(n13386), .B(n13387), .Z(n13385) );
  XNOR U15434 ( .A(n13388), .B(n13384), .Z(n13387) );
  XOR U15435 ( .A(n13389), .B(nreg[935]), .Z(n13380) );
  IV U15436 ( .A(n13378), .Z(n13389) );
  XOR U15437 ( .A(n13390), .B(n13391), .Z(n13378) );
  AND U15438 ( .A(n13392), .B(n13393), .Z(n13391) );
  XNOR U15439 ( .A(n13390), .B(n6697), .Z(n13393) );
  XNOR U15440 ( .A(n13386), .B(n13388), .Z(n6697) );
  NAND U15441 ( .A(n13394), .B(nreg[934]), .Z(n13388) );
  NAND U15442 ( .A(n12326), .B(nreg[934]), .Z(n13394) );
  XNOR U15443 ( .A(n13384), .B(n13395), .Z(n13386) );
  XOR U15444 ( .A(n13396), .B(n13397), .Z(n13384) );
  AND U15445 ( .A(n13398), .B(n13399), .Z(n13397) );
  XNOR U15446 ( .A(n13400), .B(n13396), .Z(n13399) );
  XOR U15447 ( .A(n13401), .B(nreg[934]), .Z(n13392) );
  IV U15448 ( .A(n13390), .Z(n13401) );
  XOR U15449 ( .A(n13402), .B(n13403), .Z(n13390) );
  AND U15450 ( .A(n13404), .B(n13405), .Z(n13403) );
  XNOR U15451 ( .A(n13402), .B(n6703), .Z(n13405) );
  XNOR U15452 ( .A(n13398), .B(n13400), .Z(n6703) );
  NAND U15453 ( .A(n13406), .B(nreg[933]), .Z(n13400) );
  NAND U15454 ( .A(n12326), .B(nreg[933]), .Z(n13406) );
  XNOR U15455 ( .A(n13396), .B(n13407), .Z(n13398) );
  XOR U15456 ( .A(n13408), .B(n13409), .Z(n13396) );
  AND U15457 ( .A(n13410), .B(n13411), .Z(n13409) );
  XNOR U15458 ( .A(n13412), .B(n13408), .Z(n13411) );
  XOR U15459 ( .A(n13413), .B(nreg[933]), .Z(n13404) );
  IV U15460 ( .A(n13402), .Z(n13413) );
  XOR U15461 ( .A(n13414), .B(n13415), .Z(n13402) );
  AND U15462 ( .A(n13416), .B(n13417), .Z(n13415) );
  XNOR U15463 ( .A(n13414), .B(n6709), .Z(n13417) );
  XNOR U15464 ( .A(n13410), .B(n13412), .Z(n6709) );
  NAND U15465 ( .A(n13418), .B(nreg[932]), .Z(n13412) );
  NAND U15466 ( .A(n12326), .B(nreg[932]), .Z(n13418) );
  XNOR U15467 ( .A(n13408), .B(n13419), .Z(n13410) );
  XOR U15468 ( .A(n13420), .B(n13421), .Z(n13408) );
  AND U15469 ( .A(n13422), .B(n13423), .Z(n13421) );
  XNOR U15470 ( .A(n13424), .B(n13420), .Z(n13423) );
  XOR U15471 ( .A(n13425), .B(nreg[932]), .Z(n13416) );
  IV U15472 ( .A(n13414), .Z(n13425) );
  XOR U15473 ( .A(n13426), .B(n13427), .Z(n13414) );
  AND U15474 ( .A(n13428), .B(n13429), .Z(n13427) );
  XNOR U15475 ( .A(n13426), .B(n6715), .Z(n13429) );
  XNOR U15476 ( .A(n13422), .B(n13424), .Z(n6715) );
  NAND U15477 ( .A(n13430), .B(nreg[931]), .Z(n13424) );
  NAND U15478 ( .A(n12326), .B(nreg[931]), .Z(n13430) );
  XNOR U15479 ( .A(n13420), .B(n13431), .Z(n13422) );
  XOR U15480 ( .A(n13432), .B(n13433), .Z(n13420) );
  AND U15481 ( .A(n13434), .B(n13435), .Z(n13433) );
  XNOR U15482 ( .A(n13436), .B(n13432), .Z(n13435) );
  XOR U15483 ( .A(n13437), .B(nreg[931]), .Z(n13428) );
  IV U15484 ( .A(n13426), .Z(n13437) );
  XOR U15485 ( .A(n13438), .B(n13439), .Z(n13426) );
  AND U15486 ( .A(n13440), .B(n13441), .Z(n13439) );
  XNOR U15487 ( .A(n13438), .B(n6721), .Z(n13441) );
  XNOR U15488 ( .A(n13434), .B(n13436), .Z(n6721) );
  NAND U15489 ( .A(n13442), .B(nreg[930]), .Z(n13436) );
  NAND U15490 ( .A(n12326), .B(nreg[930]), .Z(n13442) );
  XNOR U15491 ( .A(n13432), .B(n13443), .Z(n13434) );
  XOR U15492 ( .A(n13444), .B(n13445), .Z(n13432) );
  AND U15493 ( .A(n13446), .B(n13447), .Z(n13445) );
  XNOR U15494 ( .A(n13448), .B(n13444), .Z(n13447) );
  XOR U15495 ( .A(n13449), .B(nreg[930]), .Z(n13440) );
  IV U15496 ( .A(n13438), .Z(n13449) );
  XOR U15497 ( .A(n13450), .B(n13451), .Z(n13438) );
  AND U15498 ( .A(n13452), .B(n13453), .Z(n13451) );
  XNOR U15499 ( .A(n13450), .B(n6727), .Z(n13453) );
  XNOR U15500 ( .A(n13446), .B(n13448), .Z(n6727) );
  NAND U15501 ( .A(n13454), .B(nreg[929]), .Z(n13448) );
  NAND U15502 ( .A(n12326), .B(nreg[929]), .Z(n13454) );
  XNOR U15503 ( .A(n13444), .B(n13455), .Z(n13446) );
  XOR U15504 ( .A(n13456), .B(n13457), .Z(n13444) );
  AND U15505 ( .A(n13458), .B(n13459), .Z(n13457) );
  XNOR U15506 ( .A(n13460), .B(n13456), .Z(n13459) );
  XOR U15507 ( .A(n13461), .B(nreg[929]), .Z(n13452) );
  IV U15508 ( .A(n13450), .Z(n13461) );
  XOR U15509 ( .A(n13462), .B(n13463), .Z(n13450) );
  AND U15510 ( .A(n13464), .B(n13465), .Z(n13463) );
  XNOR U15511 ( .A(n13462), .B(n6733), .Z(n13465) );
  XNOR U15512 ( .A(n13458), .B(n13460), .Z(n6733) );
  NAND U15513 ( .A(n13466), .B(nreg[928]), .Z(n13460) );
  NAND U15514 ( .A(n12326), .B(nreg[928]), .Z(n13466) );
  XNOR U15515 ( .A(n13456), .B(n13467), .Z(n13458) );
  XOR U15516 ( .A(n13468), .B(n13469), .Z(n13456) );
  AND U15517 ( .A(n13470), .B(n13471), .Z(n13469) );
  XNOR U15518 ( .A(n13472), .B(n13468), .Z(n13471) );
  XOR U15519 ( .A(n13473), .B(nreg[928]), .Z(n13464) );
  IV U15520 ( .A(n13462), .Z(n13473) );
  XOR U15521 ( .A(n13474), .B(n13475), .Z(n13462) );
  AND U15522 ( .A(n13476), .B(n13477), .Z(n13475) );
  XNOR U15523 ( .A(n13474), .B(n6739), .Z(n13477) );
  XNOR U15524 ( .A(n13470), .B(n13472), .Z(n6739) );
  NAND U15525 ( .A(n13478), .B(nreg[927]), .Z(n13472) );
  NAND U15526 ( .A(n12326), .B(nreg[927]), .Z(n13478) );
  XNOR U15527 ( .A(n13468), .B(n13479), .Z(n13470) );
  XOR U15528 ( .A(n13480), .B(n13481), .Z(n13468) );
  AND U15529 ( .A(n13482), .B(n13483), .Z(n13481) );
  XNOR U15530 ( .A(n13484), .B(n13480), .Z(n13483) );
  XOR U15531 ( .A(n13485), .B(nreg[927]), .Z(n13476) );
  IV U15532 ( .A(n13474), .Z(n13485) );
  XOR U15533 ( .A(n13486), .B(n13487), .Z(n13474) );
  AND U15534 ( .A(n13488), .B(n13489), .Z(n13487) );
  XNOR U15535 ( .A(n13486), .B(n6745), .Z(n13489) );
  XNOR U15536 ( .A(n13482), .B(n13484), .Z(n6745) );
  NAND U15537 ( .A(n13490), .B(nreg[926]), .Z(n13484) );
  NAND U15538 ( .A(n12326), .B(nreg[926]), .Z(n13490) );
  XNOR U15539 ( .A(n13480), .B(n13491), .Z(n13482) );
  XOR U15540 ( .A(n13492), .B(n13493), .Z(n13480) );
  AND U15541 ( .A(n13494), .B(n13495), .Z(n13493) );
  XNOR U15542 ( .A(n13496), .B(n13492), .Z(n13495) );
  XOR U15543 ( .A(n13497), .B(nreg[926]), .Z(n13488) );
  IV U15544 ( .A(n13486), .Z(n13497) );
  XOR U15545 ( .A(n13498), .B(n13499), .Z(n13486) );
  AND U15546 ( .A(n13500), .B(n13501), .Z(n13499) );
  XNOR U15547 ( .A(n13498), .B(n6751), .Z(n13501) );
  XNOR U15548 ( .A(n13494), .B(n13496), .Z(n6751) );
  NAND U15549 ( .A(n13502), .B(nreg[925]), .Z(n13496) );
  NAND U15550 ( .A(n12326), .B(nreg[925]), .Z(n13502) );
  XNOR U15551 ( .A(n13492), .B(n13503), .Z(n13494) );
  XOR U15552 ( .A(n13504), .B(n13505), .Z(n13492) );
  AND U15553 ( .A(n13506), .B(n13507), .Z(n13505) );
  XNOR U15554 ( .A(n13508), .B(n13504), .Z(n13507) );
  XOR U15555 ( .A(n13509), .B(nreg[925]), .Z(n13500) );
  IV U15556 ( .A(n13498), .Z(n13509) );
  XOR U15557 ( .A(n13510), .B(n13511), .Z(n13498) );
  AND U15558 ( .A(n13512), .B(n13513), .Z(n13511) );
  XNOR U15559 ( .A(n13510), .B(n6757), .Z(n13513) );
  XNOR U15560 ( .A(n13506), .B(n13508), .Z(n6757) );
  NAND U15561 ( .A(n13514), .B(nreg[924]), .Z(n13508) );
  NAND U15562 ( .A(n12326), .B(nreg[924]), .Z(n13514) );
  XNOR U15563 ( .A(n13504), .B(n13515), .Z(n13506) );
  XOR U15564 ( .A(n13516), .B(n13517), .Z(n13504) );
  AND U15565 ( .A(n13518), .B(n13519), .Z(n13517) );
  XNOR U15566 ( .A(n13520), .B(n13516), .Z(n13519) );
  XOR U15567 ( .A(n13521), .B(nreg[924]), .Z(n13512) );
  IV U15568 ( .A(n13510), .Z(n13521) );
  XOR U15569 ( .A(n13522), .B(n13523), .Z(n13510) );
  AND U15570 ( .A(n13524), .B(n13525), .Z(n13523) );
  XNOR U15571 ( .A(n13522), .B(n6763), .Z(n13525) );
  XNOR U15572 ( .A(n13518), .B(n13520), .Z(n6763) );
  NAND U15573 ( .A(n13526), .B(nreg[923]), .Z(n13520) );
  NAND U15574 ( .A(n12326), .B(nreg[923]), .Z(n13526) );
  XNOR U15575 ( .A(n13516), .B(n13527), .Z(n13518) );
  XOR U15576 ( .A(n13528), .B(n13529), .Z(n13516) );
  AND U15577 ( .A(n13530), .B(n13531), .Z(n13529) );
  XNOR U15578 ( .A(n13532), .B(n13528), .Z(n13531) );
  XOR U15579 ( .A(n13533), .B(nreg[923]), .Z(n13524) );
  IV U15580 ( .A(n13522), .Z(n13533) );
  XOR U15581 ( .A(n13534), .B(n13535), .Z(n13522) );
  AND U15582 ( .A(n13536), .B(n13537), .Z(n13535) );
  XNOR U15583 ( .A(n13534), .B(n6769), .Z(n13537) );
  XNOR U15584 ( .A(n13530), .B(n13532), .Z(n6769) );
  NAND U15585 ( .A(n13538), .B(nreg[922]), .Z(n13532) );
  NAND U15586 ( .A(n12326), .B(nreg[922]), .Z(n13538) );
  XNOR U15587 ( .A(n13528), .B(n13539), .Z(n13530) );
  XOR U15588 ( .A(n13540), .B(n13541), .Z(n13528) );
  AND U15589 ( .A(n13542), .B(n13543), .Z(n13541) );
  XNOR U15590 ( .A(n13544), .B(n13540), .Z(n13543) );
  XOR U15591 ( .A(n13545), .B(nreg[922]), .Z(n13536) );
  IV U15592 ( .A(n13534), .Z(n13545) );
  XOR U15593 ( .A(n13546), .B(n13547), .Z(n13534) );
  AND U15594 ( .A(n13548), .B(n13549), .Z(n13547) );
  XNOR U15595 ( .A(n13546), .B(n6775), .Z(n13549) );
  XNOR U15596 ( .A(n13542), .B(n13544), .Z(n6775) );
  NAND U15597 ( .A(n13550), .B(nreg[921]), .Z(n13544) );
  NAND U15598 ( .A(n12326), .B(nreg[921]), .Z(n13550) );
  XNOR U15599 ( .A(n13540), .B(n13551), .Z(n13542) );
  XOR U15600 ( .A(n13552), .B(n13553), .Z(n13540) );
  AND U15601 ( .A(n13554), .B(n13555), .Z(n13553) );
  XNOR U15602 ( .A(n13556), .B(n13552), .Z(n13555) );
  XOR U15603 ( .A(n13557), .B(nreg[921]), .Z(n13548) );
  IV U15604 ( .A(n13546), .Z(n13557) );
  XOR U15605 ( .A(n13558), .B(n13559), .Z(n13546) );
  AND U15606 ( .A(n13560), .B(n13561), .Z(n13559) );
  XNOR U15607 ( .A(n13558), .B(n6781), .Z(n13561) );
  XNOR U15608 ( .A(n13554), .B(n13556), .Z(n6781) );
  NAND U15609 ( .A(n13562), .B(nreg[920]), .Z(n13556) );
  NAND U15610 ( .A(n12326), .B(nreg[920]), .Z(n13562) );
  XNOR U15611 ( .A(n13552), .B(n13563), .Z(n13554) );
  XOR U15612 ( .A(n13564), .B(n13565), .Z(n13552) );
  AND U15613 ( .A(n13566), .B(n13567), .Z(n13565) );
  XNOR U15614 ( .A(n13568), .B(n13564), .Z(n13567) );
  XOR U15615 ( .A(n13569), .B(nreg[920]), .Z(n13560) );
  IV U15616 ( .A(n13558), .Z(n13569) );
  XOR U15617 ( .A(n13570), .B(n13571), .Z(n13558) );
  AND U15618 ( .A(n13572), .B(n13573), .Z(n13571) );
  XNOR U15619 ( .A(n13570), .B(n6787), .Z(n13573) );
  XNOR U15620 ( .A(n13566), .B(n13568), .Z(n6787) );
  NAND U15621 ( .A(n13574), .B(nreg[919]), .Z(n13568) );
  NAND U15622 ( .A(n12326), .B(nreg[919]), .Z(n13574) );
  XNOR U15623 ( .A(n13564), .B(n13575), .Z(n13566) );
  XOR U15624 ( .A(n13576), .B(n13577), .Z(n13564) );
  AND U15625 ( .A(n13578), .B(n13579), .Z(n13577) );
  XNOR U15626 ( .A(n13580), .B(n13576), .Z(n13579) );
  XOR U15627 ( .A(n13581), .B(nreg[919]), .Z(n13572) );
  IV U15628 ( .A(n13570), .Z(n13581) );
  XOR U15629 ( .A(n13582), .B(n13583), .Z(n13570) );
  AND U15630 ( .A(n13584), .B(n13585), .Z(n13583) );
  XNOR U15631 ( .A(n13582), .B(n6793), .Z(n13585) );
  XNOR U15632 ( .A(n13578), .B(n13580), .Z(n6793) );
  NAND U15633 ( .A(n13586), .B(nreg[918]), .Z(n13580) );
  NAND U15634 ( .A(n12326), .B(nreg[918]), .Z(n13586) );
  XNOR U15635 ( .A(n13576), .B(n13587), .Z(n13578) );
  XOR U15636 ( .A(n13588), .B(n13589), .Z(n13576) );
  AND U15637 ( .A(n13590), .B(n13591), .Z(n13589) );
  XNOR U15638 ( .A(n13592), .B(n13588), .Z(n13591) );
  XOR U15639 ( .A(n13593), .B(nreg[918]), .Z(n13584) );
  IV U15640 ( .A(n13582), .Z(n13593) );
  XOR U15641 ( .A(n13594), .B(n13595), .Z(n13582) );
  AND U15642 ( .A(n13596), .B(n13597), .Z(n13595) );
  XNOR U15643 ( .A(n13594), .B(n6799), .Z(n13597) );
  XNOR U15644 ( .A(n13590), .B(n13592), .Z(n6799) );
  NAND U15645 ( .A(n13598), .B(nreg[917]), .Z(n13592) );
  NAND U15646 ( .A(n12326), .B(nreg[917]), .Z(n13598) );
  XNOR U15647 ( .A(n13588), .B(n13599), .Z(n13590) );
  XOR U15648 ( .A(n13600), .B(n13601), .Z(n13588) );
  AND U15649 ( .A(n13602), .B(n13603), .Z(n13601) );
  XNOR U15650 ( .A(n13604), .B(n13600), .Z(n13603) );
  XOR U15651 ( .A(n13605), .B(nreg[917]), .Z(n13596) );
  IV U15652 ( .A(n13594), .Z(n13605) );
  XOR U15653 ( .A(n13606), .B(n13607), .Z(n13594) );
  AND U15654 ( .A(n13608), .B(n13609), .Z(n13607) );
  XNOR U15655 ( .A(n13606), .B(n6805), .Z(n13609) );
  XNOR U15656 ( .A(n13602), .B(n13604), .Z(n6805) );
  NAND U15657 ( .A(n13610), .B(nreg[916]), .Z(n13604) );
  NAND U15658 ( .A(n12326), .B(nreg[916]), .Z(n13610) );
  XNOR U15659 ( .A(n13600), .B(n13611), .Z(n13602) );
  XOR U15660 ( .A(n13612), .B(n13613), .Z(n13600) );
  AND U15661 ( .A(n13614), .B(n13615), .Z(n13613) );
  XNOR U15662 ( .A(n13616), .B(n13612), .Z(n13615) );
  XOR U15663 ( .A(n13617), .B(nreg[916]), .Z(n13608) );
  IV U15664 ( .A(n13606), .Z(n13617) );
  XOR U15665 ( .A(n13618), .B(n13619), .Z(n13606) );
  AND U15666 ( .A(n13620), .B(n13621), .Z(n13619) );
  XNOR U15667 ( .A(n13618), .B(n6811), .Z(n13621) );
  XNOR U15668 ( .A(n13614), .B(n13616), .Z(n6811) );
  NAND U15669 ( .A(n13622), .B(nreg[915]), .Z(n13616) );
  NAND U15670 ( .A(n12326), .B(nreg[915]), .Z(n13622) );
  XNOR U15671 ( .A(n13612), .B(n13623), .Z(n13614) );
  XOR U15672 ( .A(n13624), .B(n13625), .Z(n13612) );
  AND U15673 ( .A(n13626), .B(n13627), .Z(n13625) );
  XNOR U15674 ( .A(n13628), .B(n13624), .Z(n13627) );
  XOR U15675 ( .A(n13629), .B(nreg[915]), .Z(n13620) );
  IV U15676 ( .A(n13618), .Z(n13629) );
  XOR U15677 ( .A(n13630), .B(n13631), .Z(n13618) );
  AND U15678 ( .A(n13632), .B(n13633), .Z(n13631) );
  XNOR U15679 ( .A(n13630), .B(n6817), .Z(n13633) );
  XNOR U15680 ( .A(n13626), .B(n13628), .Z(n6817) );
  NAND U15681 ( .A(n13634), .B(nreg[914]), .Z(n13628) );
  NAND U15682 ( .A(n12326), .B(nreg[914]), .Z(n13634) );
  XNOR U15683 ( .A(n13624), .B(n13635), .Z(n13626) );
  XOR U15684 ( .A(n13636), .B(n13637), .Z(n13624) );
  AND U15685 ( .A(n13638), .B(n13639), .Z(n13637) );
  XNOR U15686 ( .A(n13640), .B(n13636), .Z(n13639) );
  XOR U15687 ( .A(n13641), .B(nreg[914]), .Z(n13632) );
  IV U15688 ( .A(n13630), .Z(n13641) );
  XOR U15689 ( .A(n13642), .B(n13643), .Z(n13630) );
  AND U15690 ( .A(n13644), .B(n13645), .Z(n13643) );
  XNOR U15691 ( .A(n13642), .B(n6823), .Z(n13645) );
  XNOR U15692 ( .A(n13638), .B(n13640), .Z(n6823) );
  NAND U15693 ( .A(n13646), .B(nreg[913]), .Z(n13640) );
  NAND U15694 ( .A(n12326), .B(nreg[913]), .Z(n13646) );
  XNOR U15695 ( .A(n13636), .B(n13647), .Z(n13638) );
  XOR U15696 ( .A(n13648), .B(n13649), .Z(n13636) );
  AND U15697 ( .A(n13650), .B(n13651), .Z(n13649) );
  XNOR U15698 ( .A(n13652), .B(n13648), .Z(n13651) );
  XOR U15699 ( .A(n13653), .B(nreg[913]), .Z(n13644) );
  IV U15700 ( .A(n13642), .Z(n13653) );
  XOR U15701 ( .A(n13654), .B(n13655), .Z(n13642) );
  AND U15702 ( .A(n13656), .B(n13657), .Z(n13655) );
  XNOR U15703 ( .A(n13654), .B(n6829), .Z(n13657) );
  XNOR U15704 ( .A(n13650), .B(n13652), .Z(n6829) );
  NAND U15705 ( .A(n13658), .B(nreg[912]), .Z(n13652) );
  NAND U15706 ( .A(n12326), .B(nreg[912]), .Z(n13658) );
  XNOR U15707 ( .A(n13648), .B(n13659), .Z(n13650) );
  XOR U15708 ( .A(n13660), .B(n13661), .Z(n13648) );
  AND U15709 ( .A(n13662), .B(n13663), .Z(n13661) );
  XNOR U15710 ( .A(n13664), .B(n13660), .Z(n13663) );
  XOR U15711 ( .A(n13665), .B(nreg[912]), .Z(n13656) );
  IV U15712 ( .A(n13654), .Z(n13665) );
  XOR U15713 ( .A(n13666), .B(n13667), .Z(n13654) );
  AND U15714 ( .A(n13668), .B(n13669), .Z(n13667) );
  XNOR U15715 ( .A(n13666), .B(n6835), .Z(n13669) );
  XNOR U15716 ( .A(n13662), .B(n13664), .Z(n6835) );
  NAND U15717 ( .A(n13670), .B(nreg[911]), .Z(n13664) );
  NAND U15718 ( .A(n12326), .B(nreg[911]), .Z(n13670) );
  XNOR U15719 ( .A(n13660), .B(n13671), .Z(n13662) );
  XOR U15720 ( .A(n13672), .B(n13673), .Z(n13660) );
  AND U15721 ( .A(n13674), .B(n13675), .Z(n13673) );
  XNOR U15722 ( .A(n13676), .B(n13672), .Z(n13675) );
  XOR U15723 ( .A(n13677), .B(nreg[911]), .Z(n13668) );
  IV U15724 ( .A(n13666), .Z(n13677) );
  XOR U15725 ( .A(n13678), .B(n13679), .Z(n13666) );
  AND U15726 ( .A(n13680), .B(n13681), .Z(n13679) );
  XNOR U15727 ( .A(n13678), .B(n6841), .Z(n13681) );
  XNOR U15728 ( .A(n13674), .B(n13676), .Z(n6841) );
  NAND U15729 ( .A(n13682), .B(nreg[910]), .Z(n13676) );
  NAND U15730 ( .A(n12326), .B(nreg[910]), .Z(n13682) );
  XNOR U15731 ( .A(n13672), .B(n13683), .Z(n13674) );
  XOR U15732 ( .A(n13684), .B(n13685), .Z(n13672) );
  AND U15733 ( .A(n13686), .B(n13687), .Z(n13685) );
  XNOR U15734 ( .A(n13688), .B(n13684), .Z(n13687) );
  XOR U15735 ( .A(n13689), .B(nreg[910]), .Z(n13680) );
  IV U15736 ( .A(n13678), .Z(n13689) );
  XOR U15737 ( .A(n13690), .B(n13691), .Z(n13678) );
  AND U15738 ( .A(n13692), .B(n13693), .Z(n13691) );
  XNOR U15739 ( .A(n13690), .B(n6847), .Z(n13693) );
  XNOR U15740 ( .A(n13686), .B(n13688), .Z(n6847) );
  NAND U15741 ( .A(n13694), .B(nreg[909]), .Z(n13688) );
  NAND U15742 ( .A(n12326), .B(nreg[909]), .Z(n13694) );
  XNOR U15743 ( .A(n13684), .B(n13695), .Z(n13686) );
  XOR U15744 ( .A(n13696), .B(n13697), .Z(n13684) );
  AND U15745 ( .A(n13698), .B(n13699), .Z(n13697) );
  XNOR U15746 ( .A(n13700), .B(n13696), .Z(n13699) );
  XOR U15747 ( .A(n13701), .B(nreg[909]), .Z(n13692) );
  IV U15748 ( .A(n13690), .Z(n13701) );
  XOR U15749 ( .A(n13702), .B(n13703), .Z(n13690) );
  AND U15750 ( .A(n13704), .B(n13705), .Z(n13703) );
  XNOR U15751 ( .A(n13702), .B(n6853), .Z(n13705) );
  XNOR U15752 ( .A(n13698), .B(n13700), .Z(n6853) );
  NAND U15753 ( .A(n13706), .B(nreg[908]), .Z(n13700) );
  NAND U15754 ( .A(n12326), .B(nreg[908]), .Z(n13706) );
  XNOR U15755 ( .A(n13696), .B(n13707), .Z(n13698) );
  XOR U15756 ( .A(n13708), .B(n13709), .Z(n13696) );
  AND U15757 ( .A(n13710), .B(n13711), .Z(n13709) );
  XNOR U15758 ( .A(n13712), .B(n13708), .Z(n13711) );
  XOR U15759 ( .A(n13713), .B(nreg[908]), .Z(n13704) );
  IV U15760 ( .A(n13702), .Z(n13713) );
  XOR U15761 ( .A(n13714), .B(n13715), .Z(n13702) );
  AND U15762 ( .A(n13716), .B(n13717), .Z(n13715) );
  XNOR U15763 ( .A(n13714), .B(n6859), .Z(n13717) );
  XNOR U15764 ( .A(n13710), .B(n13712), .Z(n6859) );
  NAND U15765 ( .A(n13718), .B(nreg[907]), .Z(n13712) );
  NAND U15766 ( .A(n12326), .B(nreg[907]), .Z(n13718) );
  XNOR U15767 ( .A(n13708), .B(n13719), .Z(n13710) );
  XOR U15768 ( .A(n13720), .B(n13721), .Z(n13708) );
  AND U15769 ( .A(n13722), .B(n13723), .Z(n13721) );
  XNOR U15770 ( .A(n13724), .B(n13720), .Z(n13723) );
  XOR U15771 ( .A(n13725), .B(nreg[907]), .Z(n13716) );
  IV U15772 ( .A(n13714), .Z(n13725) );
  XOR U15773 ( .A(n13726), .B(n13727), .Z(n13714) );
  AND U15774 ( .A(n13728), .B(n13729), .Z(n13727) );
  XNOR U15775 ( .A(n13726), .B(n6865), .Z(n13729) );
  XNOR U15776 ( .A(n13722), .B(n13724), .Z(n6865) );
  NAND U15777 ( .A(n13730), .B(nreg[906]), .Z(n13724) );
  NAND U15778 ( .A(n12326), .B(nreg[906]), .Z(n13730) );
  XNOR U15779 ( .A(n13720), .B(n13731), .Z(n13722) );
  XOR U15780 ( .A(n13732), .B(n13733), .Z(n13720) );
  AND U15781 ( .A(n13734), .B(n13735), .Z(n13733) );
  XNOR U15782 ( .A(n13736), .B(n13732), .Z(n13735) );
  XOR U15783 ( .A(n13737), .B(nreg[906]), .Z(n13728) );
  IV U15784 ( .A(n13726), .Z(n13737) );
  XOR U15785 ( .A(n13738), .B(n13739), .Z(n13726) );
  AND U15786 ( .A(n13740), .B(n13741), .Z(n13739) );
  XNOR U15787 ( .A(n13738), .B(n6871), .Z(n13741) );
  XNOR U15788 ( .A(n13734), .B(n13736), .Z(n6871) );
  NAND U15789 ( .A(n13742), .B(nreg[905]), .Z(n13736) );
  NAND U15790 ( .A(n12326), .B(nreg[905]), .Z(n13742) );
  XNOR U15791 ( .A(n13732), .B(n13743), .Z(n13734) );
  XOR U15792 ( .A(n13744), .B(n13745), .Z(n13732) );
  AND U15793 ( .A(n13746), .B(n13747), .Z(n13745) );
  XNOR U15794 ( .A(n13748), .B(n13744), .Z(n13747) );
  XOR U15795 ( .A(n13749), .B(nreg[905]), .Z(n13740) );
  IV U15796 ( .A(n13738), .Z(n13749) );
  XOR U15797 ( .A(n13750), .B(n13751), .Z(n13738) );
  AND U15798 ( .A(n13752), .B(n13753), .Z(n13751) );
  XNOR U15799 ( .A(n13750), .B(n6877), .Z(n13753) );
  XNOR U15800 ( .A(n13746), .B(n13748), .Z(n6877) );
  NAND U15801 ( .A(n13754), .B(nreg[904]), .Z(n13748) );
  NAND U15802 ( .A(n12326), .B(nreg[904]), .Z(n13754) );
  XNOR U15803 ( .A(n13744), .B(n13755), .Z(n13746) );
  XOR U15804 ( .A(n13756), .B(n13757), .Z(n13744) );
  AND U15805 ( .A(n13758), .B(n13759), .Z(n13757) );
  XNOR U15806 ( .A(n13760), .B(n13756), .Z(n13759) );
  XOR U15807 ( .A(n13761), .B(nreg[904]), .Z(n13752) );
  IV U15808 ( .A(n13750), .Z(n13761) );
  XOR U15809 ( .A(n13762), .B(n13763), .Z(n13750) );
  AND U15810 ( .A(n13764), .B(n13765), .Z(n13763) );
  XNOR U15811 ( .A(n13762), .B(n6883), .Z(n13765) );
  XNOR U15812 ( .A(n13758), .B(n13760), .Z(n6883) );
  NAND U15813 ( .A(n13766), .B(nreg[903]), .Z(n13760) );
  NAND U15814 ( .A(n12326), .B(nreg[903]), .Z(n13766) );
  XNOR U15815 ( .A(n13756), .B(n13767), .Z(n13758) );
  XOR U15816 ( .A(n13768), .B(n13769), .Z(n13756) );
  AND U15817 ( .A(n13770), .B(n13771), .Z(n13769) );
  XNOR U15818 ( .A(n13772), .B(n13768), .Z(n13771) );
  XOR U15819 ( .A(n13773), .B(nreg[903]), .Z(n13764) );
  IV U15820 ( .A(n13762), .Z(n13773) );
  XOR U15821 ( .A(n13774), .B(n13775), .Z(n13762) );
  AND U15822 ( .A(n13776), .B(n13777), .Z(n13775) );
  XNOR U15823 ( .A(n13774), .B(n6889), .Z(n13777) );
  XNOR U15824 ( .A(n13770), .B(n13772), .Z(n6889) );
  NAND U15825 ( .A(n13778), .B(nreg[902]), .Z(n13772) );
  NAND U15826 ( .A(n12326), .B(nreg[902]), .Z(n13778) );
  XNOR U15827 ( .A(n13768), .B(n13779), .Z(n13770) );
  XOR U15828 ( .A(n13780), .B(n13781), .Z(n13768) );
  AND U15829 ( .A(n13782), .B(n13783), .Z(n13781) );
  XNOR U15830 ( .A(n13784), .B(n13780), .Z(n13783) );
  XOR U15831 ( .A(n13785), .B(nreg[902]), .Z(n13776) );
  IV U15832 ( .A(n13774), .Z(n13785) );
  XOR U15833 ( .A(n13786), .B(n13787), .Z(n13774) );
  AND U15834 ( .A(n13788), .B(n13789), .Z(n13787) );
  XNOR U15835 ( .A(n13786), .B(n6895), .Z(n13789) );
  XNOR U15836 ( .A(n13782), .B(n13784), .Z(n6895) );
  NAND U15837 ( .A(n13790), .B(nreg[901]), .Z(n13784) );
  NAND U15838 ( .A(n12326), .B(nreg[901]), .Z(n13790) );
  XNOR U15839 ( .A(n13780), .B(n13791), .Z(n13782) );
  XOR U15840 ( .A(n13792), .B(n13793), .Z(n13780) );
  AND U15841 ( .A(n13794), .B(n13795), .Z(n13793) );
  XNOR U15842 ( .A(n13796), .B(n13792), .Z(n13795) );
  XOR U15843 ( .A(n13797), .B(nreg[901]), .Z(n13788) );
  IV U15844 ( .A(n13786), .Z(n13797) );
  XOR U15845 ( .A(n13798), .B(n13799), .Z(n13786) );
  AND U15846 ( .A(n13800), .B(n13801), .Z(n13799) );
  XNOR U15847 ( .A(n13798), .B(n6901), .Z(n13801) );
  XNOR U15848 ( .A(n13794), .B(n13796), .Z(n6901) );
  NAND U15849 ( .A(n13802), .B(nreg[900]), .Z(n13796) );
  NAND U15850 ( .A(n12326), .B(nreg[900]), .Z(n13802) );
  XNOR U15851 ( .A(n13792), .B(n13803), .Z(n13794) );
  XOR U15852 ( .A(n13804), .B(n13805), .Z(n13792) );
  AND U15853 ( .A(n13806), .B(n13807), .Z(n13805) );
  XNOR U15854 ( .A(n13808), .B(n13804), .Z(n13807) );
  XOR U15855 ( .A(n13809), .B(nreg[900]), .Z(n13800) );
  IV U15856 ( .A(n13798), .Z(n13809) );
  XOR U15857 ( .A(n13810), .B(n13811), .Z(n13798) );
  AND U15858 ( .A(n13812), .B(n13813), .Z(n13811) );
  XNOR U15859 ( .A(n13810), .B(n6907), .Z(n13813) );
  XNOR U15860 ( .A(n13806), .B(n13808), .Z(n6907) );
  NAND U15861 ( .A(n13814), .B(nreg[899]), .Z(n13808) );
  NAND U15862 ( .A(n12326), .B(nreg[899]), .Z(n13814) );
  XNOR U15863 ( .A(n13804), .B(n13815), .Z(n13806) );
  XOR U15864 ( .A(n13816), .B(n13817), .Z(n13804) );
  AND U15865 ( .A(n13818), .B(n13819), .Z(n13817) );
  XNOR U15866 ( .A(n13820), .B(n13816), .Z(n13819) );
  XOR U15867 ( .A(n13821), .B(nreg[899]), .Z(n13812) );
  IV U15868 ( .A(n13810), .Z(n13821) );
  XOR U15869 ( .A(n13822), .B(n13823), .Z(n13810) );
  AND U15870 ( .A(n13824), .B(n13825), .Z(n13823) );
  XNOR U15871 ( .A(n13822), .B(n6913), .Z(n13825) );
  XNOR U15872 ( .A(n13818), .B(n13820), .Z(n6913) );
  NAND U15873 ( .A(n13826), .B(nreg[898]), .Z(n13820) );
  NAND U15874 ( .A(n12326), .B(nreg[898]), .Z(n13826) );
  XNOR U15875 ( .A(n13816), .B(n13827), .Z(n13818) );
  XOR U15876 ( .A(n13828), .B(n13829), .Z(n13816) );
  AND U15877 ( .A(n13830), .B(n13831), .Z(n13829) );
  XNOR U15878 ( .A(n13832), .B(n13828), .Z(n13831) );
  XOR U15879 ( .A(n13833), .B(nreg[898]), .Z(n13824) );
  IV U15880 ( .A(n13822), .Z(n13833) );
  XOR U15881 ( .A(n13834), .B(n13835), .Z(n13822) );
  AND U15882 ( .A(n13836), .B(n13837), .Z(n13835) );
  XNOR U15883 ( .A(n13834), .B(n6919), .Z(n13837) );
  XNOR U15884 ( .A(n13830), .B(n13832), .Z(n6919) );
  NAND U15885 ( .A(n13838), .B(nreg[897]), .Z(n13832) );
  NAND U15886 ( .A(n12326), .B(nreg[897]), .Z(n13838) );
  XNOR U15887 ( .A(n13828), .B(n13839), .Z(n13830) );
  XOR U15888 ( .A(n13840), .B(n13841), .Z(n13828) );
  AND U15889 ( .A(n13842), .B(n13843), .Z(n13841) );
  XNOR U15890 ( .A(n13844), .B(n13840), .Z(n13843) );
  XOR U15891 ( .A(n13845), .B(nreg[897]), .Z(n13836) );
  IV U15892 ( .A(n13834), .Z(n13845) );
  XOR U15893 ( .A(n13846), .B(n13847), .Z(n13834) );
  AND U15894 ( .A(n13848), .B(n13849), .Z(n13847) );
  XNOR U15895 ( .A(n13846), .B(n6925), .Z(n13849) );
  XNOR U15896 ( .A(n13842), .B(n13844), .Z(n6925) );
  NAND U15897 ( .A(n13850), .B(nreg[896]), .Z(n13844) );
  NAND U15898 ( .A(n12326), .B(nreg[896]), .Z(n13850) );
  XNOR U15899 ( .A(n13840), .B(n13851), .Z(n13842) );
  XOR U15900 ( .A(n13852), .B(n13853), .Z(n13840) );
  AND U15901 ( .A(n13854), .B(n13855), .Z(n13853) );
  XNOR U15902 ( .A(n13856), .B(n13852), .Z(n13855) );
  XOR U15903 ( .A(n13857), .B(nreg[896]), .Z(n13848) );
  IV U15904 ( .A(n13846), .Z(n13857) );
  XOR U15905 ( .A(n13858), .B(n13859), .Z(n13846) );
  AND U15906 ( .A(n13860), .B(n13861), .Z(n13859) );
  XNOR U15907 ( .A(n13858), .B(n6931), .Z(n13861) );
  XNOR U15908 ( .A(n13854), .B(n13856), .Z(n6931) );
  NAND U15909 ( .A(n13862), .B(nreg[895]), .Z(n13856) );
  NAND U15910 ( .A(n12326), .B(nreg[895]), .Z(n13862) );
  XNOR U15911 ( .A(n13852), .B(n13863), .Z(n13854) );
  XOR U15912 ( .A(n13864), .B(n13865), .Z(n13852) );
  AND U15913 ( .A(n13866), .B(n13867), .Z(n13865) );
  XNOR U15914 ( .A(n13868), .B(n13864), .Z(n13867) );
  XOR U15915 ( .A(n13869), .B(nreg[895]), .Z(n13860) );
  IV U15916 ( .A(n13858), .Z(n13869) );
  XOR U15917 ( .A(n13870), .B(n13871), .Z(n13858) );
  AND U15918 ( .A(n13872), .B(n13873), .Z(n13871) );
  XNOR U15919 ( .A(n13870), .B(n6937), .Z(n13873) );
  XNOR U15920 ( .A(n13866), .B(n13868), .Z(n6937) );
  NAND U15921 ( .A(n13874), .B(nreg[894]), .Z(n13868) );
  NAND U15922 ( .A(n12326), .B(nreg[894]), .Z(n13874) );
  XNOR U15923 ( .A(n13864), .B(n13875), .Z(n13866) );
  XOR U15924 ( .A(n13876), .B(n13877), .Z(n13864) );
  AND U15925 ( .A(n13878), .B(n13879), .Z(n13877) );
  XNOR U15926 ( .A(n13880), .B(n13876), .Z(n13879) );
  XOR U15927 ( .A(n13881), .B(nreg[894]), .Z(n13872) );
  IV U15928 ( .A(n13870), .Z(n13881) );
  XOR U15929 ( .A(n13882), .B(n13883), .Z(n13870) );
  AND U15930 ( .A(n13884), .B(n13885), .Z(n13883) );
  XNOR U15931 ( .A(n13882), .B(n6943), .Z(n13885) );
  XNOR U15932 ( .A(n13878), .B(n13880), .Z(n6943) );
  NAND U15933 ( .A(n13886), .B(nreg[893]), .Z(n13880) );
  NAND U15934 ( .A(n12326), .B(nreg[893]), .Z(n13886) );
  XNOR U15935 ( .A(n13876), .B(n13887), .Z(n13878) );
  XOR U15936 ( .A(n13888), .B(n13889), .Z(n13876) );
  AND U15937 ( .A(n13890), .B(n13891), .Z(n13889) );
  XNOR U15938 ( .A(n13892), .B(n13888), .Z(n13891) );
  XOR U15939 ( .A(n13893), .B(nreg[893]), .Z(n13884) );
  IV U15940 ( .A(n13882), .Z(n13893) );
  XOR U15941 ( .A(n13894), .B(n13895), .Z(n13882) );
  AND U15942 ( .A(n13896), .B(n13897), .Z(n13895) );
  XNOR U15943 ( .A(n13894), .B(n6949), .Z(n13897) );
  XNOR U15944 ( .A(n13890), .B(n13892), .Z(n6949) );
  NAND U15945 ( .A(n13898), .B(nreg[892]), .Z(n13892) );
  NAND U15946 ( .A(n12326), .B(nreg[892]), .Z(n13898) );
  XNOR U15947 ( .A(n13888), .B(n13899), .Z(n13890) );
  XOR U15948 ( .A(n13900), .B(n13901), .Z(n13888) );
  AND U15949 ( .A(n13902), .B(n13903), .Z(n13901) );
  XNOR U15950 ( .A(n13904), .B(n13900), .Z(n13903) );
  XOR U15951 ( .A(n13905), .B(nreg[892]), .Z(n13896) );
  IV U15952 ( .A(n13894), .Z(n13905) );
  XOR U15953 ( .A(n13906), .B(n13907), .Z(n13894) );
  AND U15954 ( .A(n13908), .B(n13909), .Z(n13907) );
  XNOR U15955 ( .A(n13906), .B(n6955), .Z(n13909) );
  XNOR U15956 ( .A(n13902), .B(n13904), .Z(n6955) );
  NAND U15957 ( .A(n13910), .B(nreg[891]), .Z(n13904) );
  NAND U15958 ( .A(n12326), .B(nreg[891]), .Z(n13910) );
  XNOR U15959 ( .A(n13900), .B(n13911), .Z(n13902) );
  XOR U15960 ( .A(n13912), .B(n13913), .Z(n13900) );
  AND U15961 ( .A(n13914), .B(n13915), .Z(n13913) );
  XNOR U15962 ( .A(n13916), .B(n13912), .Z(n13915) );
  XOR U15963 ( .A(n13917), .B(nreg[891]), .Z(n13908) );
  IV U15964 ( .A(n13906), .Z(n13917) );
  XOR U15965 ( .A(n13918), .B(n13919), .Z(n13906) );
  AND U15966 ( .A(n13920), .B(n13921), .Z(n13919) );
  XNOR U15967 ( .A(n13918), .B(n6961), .Z(n13921) );
  XNOR U15968 ( .A(n13914), .B(n13916), .Z(n6961) );
  NAND U15969 ( .A(n13922), .B(nreg[890]), .Z(n13916) );
  NAND U15970 ( .A(n12326), .B(nreg[890]), .Z(n13922) );
  XNOR U15971 ( .A(n13912), .B(n13923), .Z(n13914) );
  XOR U15972 ( .A(n13924), .B(n13925), .Z(n13912) );
  AND U15973 ( .A(n13926), .B(n13927), .Z(n13925) );
  XNOR U15974 ( .A(n13928), .B(n13924), .Z(n13927) );
  XOR U15975 ( .A(n13929), .B(nreg[890]), .Z(n13920) );
  IV U15976 ( .A(n13918), .Z(n13929) );
  XOR U15977 ( .A(n13930), .B(n13931), .Z(n13918) );
  AND U15978 ( .A(n13932), .B(n13933), .Z(n13931) );
  XNOR U15979 ( .A(n13930), .B(n6967), .Z(n13933) );
  XNOR U15980 ( .A(n13926), .B(n13928), .Z(n6967) );
  NAND U15981 ( .A(n13934), .B(nreg[889]), .Z(n13928) );
  NAND U15982 ( .A(n12326), .B(nreg[889]), .Z(n13934) );
  XNOR U15983 ( .A(n13924), .B(n13935), .Z(n13926) );
  XOR U15984 ( .A(n13936), .B(n13937), .Z(n13924) );
  AND U15985 ( .A(n13938), .B(n13939), .Z(n13937) );
  XNOR U15986 ( .A(n13940), .B(n13936), .Z(n13939) );
  XOR U15987 ( .A(n13941), .B(nreg[889]), .Z(n13932) );
  IV U15988 ( .A(n13930), .Z(n13941) );
  XOR U15989 ( .A(n13942), .B(n13943), .Z(n13930) );
  AND U15990 ( .A(n13944), .B(n13945), .Z(n13943) );
  XNOR U15991 ( .A(n13942), .B(n6973), .Z(n13945) );
  XNOR U15992 ( .A(n13938), .B(n13940), .Z(n6973) );
  NAND U15993 ( .A(n13946), .B(nreg[888]), .Z(n13940) );
  NAND U15994 ( .A(n12326), .B(nreg[888]), .Z(n13946) );
  XNOR U15995 ( .A(n13936), .B(n13947), .Z(n13938) );
  XOR U15996 ( .A(n13948), .B(n13949), .Z(n13936) );
  AND U15997 ( .A(n13950), .B(n13951), .Z(n13949) );
  XNOR U15998 ( .A(n13952), .B(n13948), .Z(n13951) );
  XOR U15999 ( .A(n13953), .B(nreg[888]), .Z(n13944) );
  IV U16000 ( .A(n13942), .Z(n13953) );
  XOR U16001 ( .A(n13954), .B(n13955), .Z(n13942) );
  AND U16002 ( .A(n13956), .B(n13957), .Z(n13955) );
  XNOR U16003 ( .A(n13954), .B(n6979), .Z(n13957) );
  XNOR U16004 ( .A(n13950), .B(n13952), .Z(n6979) );
  NAND U16005 ( .A(n13958), .B(nreg[887]), .Z(n13952) );
  NAND U16006 ( .A(n12326), .B(nreg[887]), .Z(n13958) );
  XNOR U16007 ( .A(n13948), .B(n13959), .Z(n13950) );
  XOR U16008 ( .A(n13960), .B(n13961), .Z(n13948) );
  AND U16009 ( .A(n13962), .B(n13963), .Z(n13961) );
  XNOR U16010 ( .A(n13964), .B(n13960), .Z(n13963) );
  XOR U16011 ( .A(n13965), .B(nreg[887]), .Z(n13956) );
  IV U16012 ( .A(n13954), .Z(n13965) );
  XOR U16013 ( .A(n13966), .B(n13967), .Z(n13954) );
  AND U16014 ( .A(n13968), .B(n13969), .Z(n13967) );
  XNOR U16015 ( .A(n13966), .B(n6985), .Z(n13969) );
  XNOR U16016 ( .A(n13962), .B(n13964), .Z(n6985) );
  NAND U16017 ( .A(n13970), .B(nreg[886]), .Z(n13964) );
  NAND U16018 ( .A(n12326), .B(nreg[886]), .Z(n13970) );
  XNOR U16019 ( .A(n13960), .B(n13971), .Z(n13962) );
  XOR U16020 ( .A(n13972), .B(n13973), .Z(n13960) );
  AND U16021 ( .A(n13974), .B(n13975), .Z(n13973) );
  XNOR U16022 ( .A(n13976), .B(n13972), .Z(n13975) );
  XOR U16023 ( .A(n13977), .B(nreg[886]), .Z(n13968) );
  IV U16024 ( .A(n13966), .Z(n13977) );
  XOR U16025 ( .A(n13978), .B(n13979), .Z(n13966) );
  AND U16026 ( .A(n13980), .B(n13981), .Z(n13979) );
  XNOR U16027 ( .A(n13978), .B(n6991), .Z(n13981) );
  XNOR U16028 ( .A(n13974), .B(n13976), .Z(n6991) );
  NAND U16029 ( .A(n13982), .B(nreg[885]), .Z(n13976) );
  NAND U16030 ( .A(n12326), .B(nreg[885]), .Z(n13982) );
  XNOR U16031 ( .A(n13972), .B(n13983), .Z(n13974) );
  XOR U16032 ( .A(n13984), .B(n13985), .Z(n13972) );
  AND U16033 ( .A(n13986), .B(n13987), .Z(n13985) );
  XNOR U16034 ( .A(n13988), .B(n13984), .Z(n13987) );
  XOR U16035 ( .A(n13989), .B(nreg[885]), .Z(n13980) );
  IV U16036 ( .A(n13978), .Z(n13989) );
  XOR U16037 ( .A(n13990), .B(n13991), .Z(n13978) );
  AND U16038 ( .A(n13992), .B(n13993), .Z(n13991) );
  XNOR U16039 ( .A(n13990), .B(n6997), .Z(n13993) );
  XNOR U16040 ( .A(n13986), .B(n13988), .Z(n6997) );
  NAND U16041 ( .A(n13994), .B(nreg[884]), .Z(n13988) );
  NAND U16042 ( .A(n12326), .B(nreg[884]), .Z(n13994) );
  XNOR U16043 ( .A(n13984), .B(n13995), .Z(n13986) );
  XOR U16044 ( .A(n13996), .B(n13997), .Z(n13984) );
  AND U16045 ( .A(n13998), .B(n13999), .Z(n13997) );
  XNOR U16046 ( .A(n14000), .B(n13996), .Z(n13999) );
  XOR U16047 ( .A(n14001), .B(nreg[884]), .Z(n13992) );
  IV U16048 ( .A(n13990), .Z(n14001) );
  XOR U16049 ( .A(n14002), .B(n14003), .Z(n13990) );
  AND U16050 ( .A(n14004), .B(n14005), .Z(n14003) );
  XNOR U16051 ( .A(n14002), .B(n7003), .Z(n14005) );
  XNOR U16052 ( .A(n13998), .B(n14000), .Z(n7003) );
  NAND U16053 ( .A(n14006), .B(nreg[883]), .Z(n14000) );
  NAND U16054 ( .A(n12326), .B(nreg[883]), .Z(n14006) );
  XNOR U16055 ( .A(n13996), .B(n14007), .Z(n13998) );
  XOR U16056 ( .A(n14008), .B(n14009), .Z(n13996) );
  AND U16057 ( .A(n14010), .B(n14011), .Z(n14009) );
  XNOR U16058 ( .A(n14012), .B(n14008), .Z(n14011) );
  XOR U16059 ( .A(n14013), .B(nreg[883]), .Z(n14004) );
  IV U16060 ( .A(n14002), .Z(n14013) );
  XOR U16061 ( .A(n14014), .B(n14015), .Z(n14002) );
  AND U16062 ( .A(n14016), .B(n14017), .Z(n14015) );
  XNOR U16063 ( .A(n14014), .B(n7009), .Z(n14017) );
  XNOR U16064 ( .A(n14010), .B(n14012), .Z(n7009) );
  NAND U16065 ( .A(n14018), .B(nreg[882]), .Z(n14012) );
  NAND U16066 ( .A(n12326), .B(nreg[882]), .Z(n14018) );
  XNOR U16067 ( .A(n14008), .B(n14019), .Z(n14010) );
  XOR U16068 ( .A(n14020), .B(n14021), .Z(n14008) );
  AND U16069 ( .A(n14022), .B(n14023), .Z(n14021) );
  XNOR U16070 ( .A(n14024), .B(n14020), .Z(n14023) );
  XOR U16071 ( .A(n14025), .B(nreg[882]), .Z(n14016) );
  IV U16072 ( .A(n14014), .Z(n14025) );
  XOR U16073 ( .A(n14026), .B(n14027), .Z(n14014) );
  AND U16074 ( .A(n14028), .B(n14029), .Z(n14027) );
  XNOR U16075 ( .A(n14026), .B(n7015), .Z(n14029) );
  XNOR U16076 ( .A(n14022), .B(n14024), .Z(n7015) );
  NAND U16077 ( .A(n14030), .B(nreg[881]), .Z(n14024) );
  NAND U16078 ( .A(n12326), .B(nreg[881]), .Z(n14030) );
  XNOR U16079 ( .A(n14020), .B(n14031), .Z(n14022) );
  XOR U16080 ( .A(n14032), .B(n14033), .Z(n14020) );
  AND U16081 ( .A(n14034), .B(n14035), .Z(n14033) );
  XNOR U16082 ( .A(n14036), .B(n14032), .Z(n14035) );
  XOR U16083 ( .A(n14037), .B(nreg[881]), .Z(n14028) );
  IV U16084 ( .A(n14026), .Z(n14037) );
  XOR U16085 ( .A(n14038), .B(n14039), .Z(n14026) );
  AND U16086 ( .A(n14040), .B(n14041), .Z(n14039) );
  XNOR U16087 ( .A(n14038), .B(n7021), .Z(n14041) );
  XNOR U16088 ( .A(n14034), .B(n14036), .Z(n7021) );
  NAND U16089 ( .A(n14042), .B(nreg[880]), .Z(n14036) );
  NAND U16090 ( .A(n12326), .B(nreg[880]), .Z(n14042) );
  XNOR U16091 ( .A(n14032), .B(n14043), .Z(n14034) );
  XOR U16092 ( .A(n14044), .B(n14045), .Z(n14032) );
  AND U16093 ( .A(n14046), .B(n14047), .Z(n14045) );
  XNOR U16094 ( .A(n14048), .B(n14044), .Z(n14047) );
  XOR U16095 ( .A(n14049), .B(nreg[880]), .Z(n14040) );
  IV U16096 ( .A(n14038), .Z(n14049) );
  XOR U16097 ( .A(n14050), .B(n14051), .Z(n14038) );
  AND U16098 ( .A(n14052), .B(n14053), .Z(n14051) );
  XNOR U16099 ( .A(n14050), .B(n7027), .Z(n14053) );
  XNOR U16100 ( .A(n14046), .B(n14048), .Z(n7027) );
  NAND U16101 ( .A(n14054), .B(nreg[879]), .Z(n14048) );
  NAND U16102 ( .A(n12326), .B(nreg[879]), .Z(n14054) );
  XNOR U16103 ( .A(n14044), .B(n14055), .Z(n14046) );
  XOR U16104 ( .A(n14056), .B(n14057), .Z(n14044) );
  AND U16105 ( .A(n14058), .B(n14059), .Z(n14057) );
  XNOR U16106 ( .A(n14060), .B(n14056), .Z(n14059) );
  XOR U16107 ( .A(n14061), .B(nreg[879]), .Z(n14052) );
  IV U16108 ( .A(n14050), .Z(n14061) );
  XOR U16109 ( .A(n14062), .B(n14063), .Z(n14050) );
  AND U16110 ( .A(n14064), .B(n14065), .Z(n14063) );
  XNOR U16111 ( .A(n14062), .B(n7033), .Z(n14065) );
  XNOR U16112 ( .A(n14058), .B(n14060), .Z(n7033) );
  NAND U16113 ( .A(n14066), .B(nreg[878]), .Z(n14060) );
  NAND U16114 ( .A(n12326), .B(nreg[878]), .Z(n14066) );
  XNOR U16115 ( .A(n14056), .B(n14067), .Z(n14058) );
  XOR U16116 ( .A(n14068), .B(n14069), .Z(n14056) );
  AND U16117 ( .A(n14070), .B(n14071), .Z(n14069) );
  XNOR U16118 ( .A(n14072), .B(n14068), .Z(n14071) );
  XOR U16119 ( .A(n14073), .B(nreg[878]), .Z(n14064) );
  IV U16120 ( .A(n14062), .Z(n14073) );
  XOR U16121 ( .A(n14074), .B(n14075), .Z(n14062) );
  AND U16122 ( .A(n14076), .B(n14077), .Z(n14075) );
  XNOR U16123 ( .A(n14074), .B(n7039), .Z(n14077) );
  XNOR U16124 ( .A(n14070), .B(n14072), .Z(n7039) );
  NAND U16125 ( .A(n14078), .B(nreg[877]), .Z(n14072) );
  NAND U16126 ( .A(n12326), .B(nreg[877]), .Z(n14078) );
  XNOR U16127 ( .A(n14068), .B(n14079), .Z(n14070) );
  XOR U16128 ( .A(n14080), .B(n14081), .Z(n14068) );
  AND U16129 ( .A(n14082), .B(n14083), .Z(n14081) );
  XNOR U16130 ( .A(n14084), .B(n14080), .Z(n14083) );
  XOR U16131 ( .A(n14085), .B(nreg[877]), .Z(n14076) );
  IV U16132 ( .A(n14074), .Z(n14085) );
  XOR U16133 ( .A(n14086), .B(n14087), .Z(n14074) );
  AND U16134 ( .A(n14088), .B(n14089), .Z(n14087) );
  XNOR U16135 ( .A(n14086), .B(n7045), .Z(n14089) );
  XNOR U16136 ( .A(n14082), .B(n14084), .Z(n7045) );
  NAND U16137 ( .A(n14090), .B(nreg[876]), .Z(n14084) );
  NAND U16138 ( .A(n12326), .B(nreg[876]), .Z(n14090) );
  XNOR U16139 ( .A(n14080), .B(n14091), .Z(n14082) );
  XOR U16140 ( .A(n14092), .B(n14093), .Z(n14080) );
  AND U16141 ( .A(n14094), .B(n14095), .Z(n14093) );
  XNOR U16142 ( .A(n14096), .B(n14092), .Z(n14095) );
  XOR U16143 ( .A(n14097), .B(nreg[876]), .Z(n14088) );
  IV U16144 ( .A(n14086), .Z(n14097) );
  XOR U16145 ( .A(n14098), .B(n14099), .Z(n14086) );
  AND U16146 ( .A(n14100), .B(n14101), .Z(n14099) );
  XNOR U16147 ( .A(n14098), .B(n7051), .Z(n14101) );
  XNOR U16148 ( .A(n14094), .B(n14096), .Z(n7051) );
  NAND U16149 ( .A(n14102), .B(nreg[875]), .Z(n14096) );
  NAND U16150 ( .A(n12326), .B(nreg[875]), .Z(n14102) );
  XNOR U16151 ( .A(n14092), .B(n14103), .Z(n14094) );
  XOR U16152 ( .A(n14104), .B(n14105), .Z(n14092) );
  AND U16153 ( .A(n14106), .B(n14107), .Z(n14105) );
  XNOR U16154 ( .A(n14108), .B(n14104), .Z(n14107) );
  XOR U16155 ( .A(n14109), .B(nreg[875]), .Z(n14100) );
  IV U16156 ( .A(n14098), .Z(n14109) );
  XOR U16157 ( .A(n14110), .B(n14111), .Z(n14098) );
  AND U16158 ( .A(n14112), .B(n14113), .Z(n14111) );
  XNOR U16159 ( .A(n14110), .B(n7057), .Z(n14113) );
  XNOR U16160 ( .A(n14106), .B(n14108), .Z(n7057) );
  NAND U16161 ( .A(n14114), .B(nreg[874]), .Z(n14108) );
  NAND U16162 ( .A(n12326), .B(nreg[874]), .Z(n14114) );
  XNOR U16163 ( .A(n14104), .B(n14115), .Z(n14106) );
  XOR U16164 ( .A(n14116), .B(n14117), .Z(n14104) );
  AND U16165 ( .A(n14118), .B(n14119), .Z(n14117) );
  XNOR U16166 ( .A(n14120), .B(n14116), .Z(n14119) );
  XOR U16167 ( .A(n14121), .B(nreg[874]), .Z(n14112) );
  IV U16168 ( .A(n14110), .Z(n14121) );
  XOR U16169 ( .A(n14122), .B(n14123), .Z(n14110) );
  AND U16170 ( .A(n14124), .B(n14125), .Z(n14123) );
  XNOR U16171 ( .A(n14122), .B(n7063), .Z(n14125) );
  XNOR U16172 ( .A(n14118), .B(n14120), .Z(n7063) );
  NAND U16173 ( .A(n14126), .B(nreg[873]), .Z(n14120) );
  NAND U16174 ( .A(n12326), .B(nreg[873]), .Z(n14126) );
  XNOR U16175 ( .A(n14116), .B(n14127), .Z(n14118) );
  XOR U16176 ( .A(n14128), .B(n14129), .Z(n14116) );
  AND U16177 ( .A(n14130), .B(n14131), .Z(n14129) );
  XNOR U16178 ( .A(n14132), .B(n14128), .Z(n14131) );
  XOR U16179 ( .A(n14133), .B(nreg[873]), .Z(n14124) );
  IV U16180 ( .A(n14122), .Z(n14133) );
  XOR U16181 ( .A(n14134), .B(n14135), .Z(n14122) );
  AND U16182 ( .A(n14136), .B(n14137), .Z(n14135) );
  XNOR U16183 ( .A(n14134), .B(n7069), .Z(n14137) );
  XNOR U16184 ( .A(n14130), .B(n14132), .Z(n7069) );
  NAND U16185 ( .A(n14138), .B(nreg[872]), .Z(n14132) );
  NAND U16186 ( .A(n12326), .B(nreg[872]), .Z(n14138) );
  XNOR U16187 ( .A(n14128), .B(n14139), .Z(n14130) );
  XOR U16188 ( .A(n14140), .B(n14141), .Z(n14128) );
  AND U16189 ( .A(n14142), .B(n14143), .Z(n14141) );
  XNOR U16190 ( .A(n14144), .B(n14140), .Z(n14143) );
  XOR U16191 ( .A(n14145), .B(nreg[872]), .Z(n14136) );
  IV U16192 ( .A(n14134), .Z(n14145) );
  XOR U16193 ( .A(n14146), .B(n14147), .Z(n14134) );
  AND U16194 ( .A(n14148), .B(n14149), .Z(n14147) );
  XNOR U16195 ( .A(n14146), .B(n7075), .Z(n14149) );
  XNOR U16196 ( .A(n14142), .B(n14144), .Z(n7075) );
  NAND U16197 ( .A(n14150), .B(nreg[871]), .Z(n14144) );
  NAND U16198 ( .A(n12326), .B(nreg[871]), .Z(n14150) );
  XNOR U16199 ( .A(n14140), .B(n14151), .Z(n14142) );
  XOR U16200 ( .A(n14152), .B(n14153), .Z(n14140) );
  AND U16201 ( .A(n14154), .B(n14155), .Z(n14153) );
  XNOR U16202 ( .A(n14156), .B(n14152), .Z(n14155) );
  XOR U16203 ( .A(n14157), .B(nreg[871]), .Z(n14148) );
  IV U16204 ( .A(n14146), .Z(n14157) );
  XOR U16205 ( .A(n14158), .B(n14159), .Z(n14146) );
  AND U16206 ( .A(n14160), .B(n14161), .Z(n14159) );
  XNOR U16207 ( .A(n14158), .B(n7081), .Z(n14161) );
  XNOR U16208 ( .A(n14154), .B(n14156), .Z(n7081) );
  NAND U16209 ( .A(n14162), .B(nreg[870]), .Z(n14156) );
  NAND U16210 ( .A(n12326), .B(nreg[870]), .Z(n14162) );
  XNOR U16211 ( .A(n14152), .B(n14163), .Z(n14154) );
  XOR U16212 ( .A(n14164), .B(n14165), .Z(n14152) );
  AND U16213 ( .A(n14166), .B(n14167), .Z(n14165) );
  XNOR U16214 ( .A(n14168), .B(n14164), .Z(n14167) );
  XOR U16215 ( .A(n14169), .B(nreg[870]), .Z(n14160) );
  IV U16216 ( .A(n14158), .Z(n14169) );
  XOR U16217 ( .A(n14170), .B(n14171), .Z(n14158) );
  AND U16218 ( .A(n14172), .B(n14173), .Z(n14171) );
  XNOR U16219 ( .A(n14170), .B(n7087), .Z(n14173) );
  XNOR U16220 ( .A(n14166), .B(n14168), .Z(n7087) );
  NAND U16221 ( .A(n14174), .B(nreg[869]), .Z(n14168) );
  NAND U16222 ( .A(n12326), .B(nreg[869]), .Z(n14174) );
  XNOR U16223 ( .A(n14164), .B(n14175), .Z(n14166) );
  XOR U16224 ( .A(n14176), .B(n14177), .Z(n14164) );
  AND U16225 ( .A(n14178), .B(n14179), .Z(n14177) );
  XNOR U16226 ( .A(n14180), .B(n14176), .Z(n14179) );
  XOR U16227 ( .A(n14181), .B(nreg[869]), .Z(n14172) );
  IV U16228 ( .A(n14170), .Z(n14181) );
  XOR U16229 ( .A(n14182), .B(n14183), .Z(n14170) );
  AND U16230 ( .A(n14184), .B(n14185), .Z(n14183) );
  XNOR U16231 ( .A(n14182), .B(n7093), .Z(n14185) );
  XNOR U16232 ( .A(n14178), .B(n14180), .Z(n7093) );
  NAND U16233 ( .A(n14186), .B(nreg[868]), .Z(n14180) );
  NAND U16234 ( .A(n12326), .B(nreg[868]), .Z(n14186) );
  XNOR U16235 ( .A(n14176), .B(n14187), .Z(n14178) );
  XOR U16236 ( .A(n14188), .B(n14189), .Z(n14176) );
  AND U16237 ( .A(n14190), .B(n14191), .Z(n14189) );
  XNOR U16238 ( .A(n14192), .B(n14188), .Z(n14191) );
  XOR U16239 ( .A(n14193), .B(nreg[868]), .Z(n14184) );
  IV U16240 ( .A(n14182), .Z(n14193) );
  XOR U16241 ( .A(n14194), .B(n14195), .Z(n14182) );
  AND U16242 ( .A(n14196), .B(n14197), .Z(n14195) );
  XNOR U16243 ( .A(n14194), .B(n7099), .Z(n14197) );
  XNOR U16244 ( .A(n14190), .B(n14192), .Z(n7099) );
  NAND U16245 ( .A(n14198), .B(nreg[867]), .Z(n14192) );
  NAND U16246 ( .A(n12326), .B(nreg[867]), .Z(n14198) );
  XNOR U16247 ( .A(n14188), .B(n14199), .Z(n14190) );
  XOR U16248 ( .A(n14200), .B(n14201), .Z(n14188) );
  AND U16249 ( .A(n14202), .B(n14203), .Z(n14201) );
  XNOR U16250 ( .A(n14204), .B(n14200), .Z(n14203) );
  XOR U16251 ( .A(n14205), .B(nreg[867]), .Z(n14196) );
  IV U16252 ( .A(n14194), .Z(n14205) );
  XOR U16253 ( .A(n14206), .B(n14207), .Z(n14194) );
  AND U16254 ( .A(n14208), .B(n14209), .Z(n14207) );
  XNOR U16255 ( .A(n14206), .B(n7105), .Z(n14209) );
  XNOR U16256 ( .A(n14202), .B(n14204), .Z(n7105) );
  NAND U16257 ( .A(n14210), .B(nreg[866]), .Z(n14204) );
  NAND U16258 ( .A(n12326), .B(nreg[866]), .Z(n14210) );
  XNOR U16259 ( .A(n14200), .B(n14211), .Z(n14202) );
  XOR U16260 ( .A(n14212), .B(n14213), .Z(n14200) );
  AND U16261 ( .A(n14214), .B(n14215), .Z(n14213) );
  XNOR U16262 ( .A(n14216), .B(n14212), .Z(n14215) );
  XOR U16263 ( .A(n14217), .B(nreg[866]), .Z(n14208) );
  IV U16264 ( .A(n14206), .Z(n14217) );
  XOR U16265 ( .A(n14218), .B(n14219), .Z(n14206) );
  AND U16266 ( .A(n14220), .B(n14221), .Z(n14219) );
  XNOR U16267 ( .A(n14218), .B(n7111), .Z(n14221) );
  XNOR U16268 ( .A(n14214), .B(n14216), .Z(n7111) );
  NAND U16269 ( .A(n14222), .B(nreg[865]), .Z(n14216) );
  NAND U16270 ( .A(n12326), .B(nreg[865]), .Z(n14222) );
  XNOR U16271 ( .A(n14212), .B(n14223), .Z(n14214) );
  XOR U16272 ( .A(n14224), .B(n14225), .Z(n14212) );
  AND U16273 ( .A(n14226), .B(n14227), .Z(n14225) );
  XNOR U16274 ( .A(n14228), .B(n14224), .Z(n14227) );
  XOR U16275 ( .A(n14229), .B(nreg[865]), .Z(n14220) );
  IV U16276 ( .A(n14218), .Z(n14229) );
  XOR U16277 ( .A(n14230), .B(n14231), .Z(n14218) );
  AND U16278 ( .A(n14232), .B(n14233), .Z(n14231) );
  XNOR U16279 ( .A(n14230), .B(n7117), .Z(n14233) );
  XNOR U16280 ( .A(n14226), .B(n14228), .Z(n7117) );
  NAND U16281 ( .A(n14234), .B(nreg[864]), .Z(n14228) );
  NAND U16282 ( .A(n12326), .B(nreg[864]), .Z(n14234) );
  XNOR U16283 ( .A(n14224), .B(n14235), .Z(n14226) );
  XOR U16284 ( .A(n14236), .B(n14237), .Z(n14224) );
  AND U16285 ( .A(n14238), .B(n14239), .Z(n14237) );
  XNOR U16286 ( .A(n14240), .B(n14236), .Z(n14239) );
  XOR U16287 ( .A(n14241), .B(nreg[864]), .Z(n14232) );
  IV U16288 ( .A(n14230), .Z(n14241) );
  XOR U16289 ( .A(n14242), .B(n14243), .Z(n14230) );
  AND U16290 ( .A(n14244), .B(n14245), .Z(n14243) );
  XNOR U16291 ( .A(n14242), .B(n7123), .Z(n14245) );
  XNOR U16292 ( .A(n14238), .B(n14240), .Z(n7123) );
  NAND U16293 ( .A(n14246), .B(nreg[863]), .Z(n14240) );
  NAND U16294 ( .A(n12326), .B(nreg[863]), .Z(n14246) );
  XNOR U16295 ( .A(n14236), .B(n14247), .Z(n14238) );
  XOR U16296 ( .A(n14248), .B(n14249), .Z(n14236) );
  AND U16297 ( .A(n14250), .B(n14251), .Z(n14249) );
  XNOR U16298 ( .A(n14252), .B(n14248), .Z(n14251) );
  XOR U16299 ( .A(n14253), .B(nreg[863]), .Z(n14244) );
  IV U16300 ( .A(n14242), .Z(n14253) );
  XOR U16301 ( .A(n14254), .B(n14255), .Z(n14242) );
  AND U16302 ( .A(n14256), .B(n14257), .Z(n14255) );
  XNOR U16303 ( .A(n14254), .B(n7129), .Z(n14257) );
  XNOR U16304 ( .A(n14250), .B(n14252), .Z(n7129) );
  NAND U16305 ( .A(n14258), .B(nreg[862]), .Z(n14252) );
  NAND U16306 ( .A(n12326), .B(nreg[862]), .Z(n14258) );
  XNOR U16307 ( .A(n14248), .B(n14259), .Z(n14250) );
  XOR U16308 ( .A(n14260), .B(n14261), .Z(n14248) );
  AND U16309 ( .A(n14262), .B(n14263), .Z(n14261) );
  XNOR U16310 ( .A(n14264), .B(n14260), .Z(n14263) );
  XOR U16311 ( .A(n14265), .B(nreg[862]), .Z(n14256) );
  IV U16312 ( .A(n14254), .Z(n14265) );
  XOR U16313 ( .A(n14266), .B(n14267), .Z(n14254) );
  AND U16314 ( .A(n14268), .B(n14269), .Z(n14267) );
  XNOR U16315 ( .A(n14266), .B(n7135), .Z(n14269) );
  XNOR U16316 ( .A(n14262), .B(n14264), .Z(n7135) );
  NAND U16317 ( .A(n14270), .B(nreg[861]), .Z(n14264) );
  NAND U16318 ( .A(n12326), .B(nreg[861]), .Z(n14270) );
  XNOR U16319 ( .A(n14260), .B(n14271), .Z(n14262) );
  XOR U16320 ( .A(n14272), .B(n14273), .Z(n14260) );
  AND U16321 ( .A(n14274), .B(n14275), .Z(n14273) );
  XNOR U16322 ( .A(n14276), .B(n14272), .Z(n14275) );
  XOR U16323 ( .A(n14277), .B(nreg[861]), .Z(n14268) );
  IV U16324 ( .A(n14266), .Z(n14277) );
  XOR U16325 ( .A(n14278), .B(n14279), .Z(n14266) );
  AND U16326 ( .A(n14280), .B(n14281), .Z(n14279) );
  XNOR U16327 ( .A(n14278), .B(n7141), .Z(n14281) );
  XNOR U16328 ( .A(n14274), .B(n14276), .Z(n7141) );
  NAND U16329 ( .A(n14282), .B(nreg[860]), .Z(n14276) );
  NAND U16330 ( .A(n12326), .B(nreg[860]), .Z(n14282) );
  XNOR U16331 ( .A(n14272), .B(n14283), .Z(n14274) );
  XOR U16332 ( .A(n14284), .B(n14285), .Z(n14272) );
  AND U16333 ( .A(n14286), .B(n14287), .Z(n14285) );
  XNOR U16334 ( .A(n14288), .B(n14284), .Z(n14287) );
  XOR U16335 ( .A(n14289), .B(nreg[860]), .Z(n14280) );
  IV U16336 ( .A(n14278), .Z(n14289) );
  XOR U16337 ( .A(n14290), .B(n14291), .Z(n14278) );
  AND U16338 ( .A(n14292), .B(n14293), .Z(n14291) );
  XNOR U16339 ( .A(n14290), .B(n7147), .Z(n14293) );
  XNOR U16340 ( .A(n14286), .B(n14288), .Z(n7147) );
  NAND U16341 ( .A(n14294), .B(nreg[859]), .Z(n14288) );
  NAND U16342 ( .A(n12326), .B(nreg[859]), .Z(n14294) );
  XNOR U16343 ( .A(n14284), .B(n14295), .Z(n14286) );
  XOR U16344 ( .A(n14296), .B(n14297), .Z(n14284) );
  AND U16345 ( .A(n14298), .B(n14299), .Z(n14297) );
  XNOR U16346 ( .A(n14300), .B(n14296), .Z(n14299) );
  XOR U16347 ( .A(n14301), .B(nreg[859]), .Z(n14292) );
  IV U16348 ( .A(n14290), .Z(n14301) );
  XOR U16349 ( .A(n14302), .B(n14303), .Z(n14290) );
  AND U16350 ( .A(n14304), .B(n14305), .Z(n14303) );
  XNOR U16351 ( .A(n14302), .B(n7153), .Z(n14305) );
  XNOR U16352 ( .A(n14298), .B(n14300), .Z(n7153) );
  NAND U16353 ( .A(n14306), .B(nreg[858]), .Z(n14300) );
  NAND U16354 ( .A(n12326), .B(nreg[858]), .Z(n14306) );
  XNOR U16355 ( .A(n14296), .B(n14307), .Z(n14298) );
  XOR U16356 ( .A(n14308), .B(n14309), .Z(n14296) );
  AND U16357 ( .A(n14310), .B(n14311), .Z(n14309) );
  XNOR U16358 ( .A(n14312), .B(n14308), .Z(n14311) );
  XOR U16359 ( .A(n14313), .B(nreg[858]), .Z(n14304) );
  IV U16360 ( .A(n14302), .Z(n14313) );
  XOR U16361 ( .A(n14314), .B(n14315), .Z(n14302) );
  AND U16362 ( .A(n14316), .B(n14317), .Z(n14315) );
  XNOR U16363 ( .A(n14314), .B(n7159), .Z(n14317) );
  XNOR U16364 ( .A(n14310), .B(n14312), .Z(n7159) );
  NAND U16365 ( .A(n14318), .B(nreg[857]), .Z(n14312) );
  NAND U16366 ( .A(n12326), .B(nreg[857]), .Z(n14318) );
  XNOR U16367 ( .A(n14308), .B(n14319), .Z(n14310) );
  XOR U16368 ( .A(n14320), .B(n14321), .Z(n14308) );
  AND U16369 ( .A(n14322), .B(n14323), .Z(n14321) );
  XNOR U16370 ( .A(n14324), .B(n14320), .Z(n14323) );
  XOR U16371 ( .A(n14325), .B(nreg[857]), .Z(n14316) );
  IV U16372 ( .A(n14314), .Z(n14325) );
  XOR U16373 ( .A(n14326), .B(n14327), .Z(n14314) );
  AND U16374 ( .A(n14328), .B(n14329), .Z(n14327) );
  XNOR U16375 ( .A(n14326), .B(n7165), .Z(n14329) );
  XNOR U16376 ( .A(n14322), .B(n14324), .Z(n7165) );
  NAND U16377 ( .A(n14330), .B(nreg[856]), .Z(n14324) );
  NAND U16378 ( .A(n12326), .B(nreg[856]), .Z(n14330) );
  XNOR U16379 ( .A(n14320), .B(n14331), .Z(n14322) );
  XOR U16380 ( .A(n14332), .B(n14333), .Z(n14320) );
  AND U16381 ( .A(n14334), .B(n14335), .Z(n14333) );
  XNOR U16382 ( .A(n14336), .B(n14332), .Z(n14335) );
  XOR U16383 ( .A(n14337), .B(nreg[856]), .Z(n14328) );
  IV U16384 ( .A(n14326), .Z(n14337) );
  XOR U16385 ( .A(n14338), .B(n14339), .Z(n14326) );
  AND U16386 ( .A(n14340), .B(n14341), .Z(n14339) );
  XNOR U16387 ( .A(n14338), .B(n7171), .Z(n14341) );
  XNOR U16388 ( .A(n14334), .B(n14336), .Z(n7171) );
  NAND U16389 ( .A(n14342), .B(nreg[855]), .Z(n14336) );
  NAND U16390 ( .A(n12326), .B(nreg[855]), .Z(n14342) );
  XNOR U16391 ( .A(n14332), .B(n14343), .Z(n14334) );
  XOR U16392 ( .A(n14344), .B(n14345), .Z(n14332) );
  AND U16393 ( .A(n14346), .B(n14347), .Z(n14345) );
  XNOR U16394 ( .A(n14348), .B(n14344), .Z(n14347) );
  XOR U16395 ( .A(n14349), .B(nreg[855]), .Z(n14340) );
  IV U16396 ( .A(n14338), .Z(n14349) );
  XOR U16397 ( .A(n14350), .B(n14351), .Z(n14338) );
  AND U16398 ( .A(n14352), .B(n14353), .Z(n14351) );
  XNOR U16399 ( .A(n14350), .B(n7177), .Z(n14353) );
  XNOR U16400 ( .A(n14346), .B(n14348), .Z(n7177) );
  NAND U16401 ( .A(n14354), .B(nreg[854]), .Z(n14348) );
  NAND U16402 ( .A(n12326), .B(nreg[854]), .Z(n14354) );
  XNOR U16403 ( .A(n14344), .B(n14355), .Z(n14346) );
  XOR U16404 ( .A(n14356), .B(n14357), .Z(n14344) );
  AND U16405 ( .A(n14358), .B(n14359), .Z(n14357) );
  XNOR U16406 ( .A(n14360), .B(n14356), .Z(n14359) );
  XOR U16407 ( .A(n14361), .B(nreg[854]), .Z(n14352) );
  IV U16408 ( .A(n14350), .Z(n14361) );
  XOR U16409 ( .A(n14362), .B(n14363), .Z(n14350) );
  AND U16410 ( .A(n14364), .B(n14365), .Z(n14363) );
  XNOR U16411 ( .A(n14362), .B(n7183), .Z(n14365) );
  XNOR U16412 ( .A(n14358), .B(n14360), .Z(n7183) );
  NAND U16413 ( .A(n14366), .B(nreg[853]), .Z(n14360) );
  NAND U16414 ( .A(n12326), .B(nreg[853]), .Z(n14366) );
  XNOR U16415 ( .A(n14356), .B(n14367), .Z(n14358) );
  XOR U16416 ( .A(n14368), .B(n14369), .Z(n14356) );
  AND U16417 ( .A(n14370), .B(n14371), .Z(n14369) );
  XNOR U16418 ( .A(n14372), .B(n14368), .Z(n14371) );
  XOR U16419 ( .A(n14373), .B(nreg[853]), .Z(n14364) );
  IV U16420 ( .A(n14362), .Z(n14373) );
  XOR U16421 ( .A(n14374), .B(n14375), .Z(n14362) );
  AND U16422 ( .A(n14376), .B(n14377), .Z(n14375) );
  XNOR U16423 ( .A(n14374), .B(n7189), .Z(n14377) );
  XNOR U16424 ( .A(n14370), .B(n14372), .Z(n7189) );
  NAND U16425 ( .A(n14378), .B(nreg[852]), .Z(n14372) );
  NAND U16426 ( .A(n12326), .B(nreg[852]), .Z(n14378) );
  XNOR U16427 ( .A(n14368), .B(n14379), .Z(n14370) );
  XOR U16428 ( .A(n14380), .B(n14381), .Z(n14368) );
  AND U16429 ( .A(n14382), .B(n14383), .Z(n14381) );
  XNOR U16430 ( .A(n14384), .B(n14380), .Z(n14383) );
  XOR U16431 ( .A(n14385), .B(nreg[852]), .Z(n14376) );
  IV U16432 ( .A(n14374), .Z(n14385) );
  XOR U16433 ( .A(n14386), .B(n14387), .Z(n14374) );
  AND U16434 ( .A(n14388), .B(n14389), .Z(n14387) );
  XNOR U16435 ( .A(n14386), .B(n7195), .Z(n14389) );
  XNOR U16436 ( .A(n14382), .B(n14384), .Z(n7195) );
  NAND U16437 ( .A(n14390), .B(nreg[851]), .Z(n14384) );
  NAND U16438 ( .A(n12326), .B(nreg[851]), .Z(n14390) );
  XNOR U16439 ( .A(n14380), .B(n14391), .Z(n14382) );
  XOR U16440 ( .A(n14392), .B(n14393), .Z(n14380) );
  AND U16441 ( .A(n14394), .B(n14395), .Z(n14393) );
  XNOR U16442 ( .A(n14396), .B(n14392), .Z(n14395) );
  XOR U16443 ( .A(n14397), .B(nreg[851]), .Z(n14388) );
  IV U16444 ( .A(n14386), .Z(n14397) );
  XOR U16445 ( .A(n14398), .B(n14399), .Z(n14386) );
  AND U16446 ( .A(n14400), .B(n14401), .Z(n14399) );
  XNOR U16447 ( .A(n14398), .B(n7201), .Z(n14401) );
  XNOR U16448 ( .A(n14394), .B(n14396), .Z(n7201) );
  NAND U16449 ( .A(n14402), .B(nreg[850]), .Z(n14396) );
  NAND U16450 ( .A(n12326), .B(nreg[850]), .Z(n14402) );
  XNOR U16451 ( .A(n14392), .B(n14403), .Z(n14394) );
  XOR U16452 ( .A(n14404), .B(n14405), .Z(n14392) );
  AND U16453 ( .A(n14406), .B(n14407), .Z(n14405) );
  XNOR U16454 ( .A(n14408), .B(n14404), .Z(n14407) );
  XOR U16455 ( .A(n14409), .B(nreg[850]), .Z(n14400) );
  IV U16456 ( .A(n14398), .Z(n14409) );
  XOR U16457 ( .A(n14410), .B(n14411), .Z(n14398) );
  AND U16458 ( .A(n14412), .B(n14413), .Z(n14411) );
  XNOR U16459 ( .A(n14410), .B(n7207), .Z(n14413) );
  XNOR U16460 ( .A(n14406), .B(n14408), .Z(n7207) );
  NAND U16461 ( .A(n14414), .B(nreg[849]), .Z(n14408) );
  NAND U16462 ( .A(n12326), .B(nreg[849]), .Z(n14414) );
  XNOR U16463 ( .A(n14404), .B(n14415), .Z(n14406) );
  XOR U16464 ( .A(n14416), .B(n14417), .Z(n14404) );
  AND U16465 ( .A(n14418), .B(n14419), .Z(n14417) );
  XNOR U16466 ( .A(n14420), .B(n14416), .Z(n14419) );
  XOR U16467 ( .A(n14421), .B(nreg[849]), .Z(n14412) );
  IV U16468 ( .A(n14410), .Z(n14421) );
  XOR U16469 ( .A(n14422), .B(n14423), .Z(n14410) );
  AND U16470 ( .A(n14424), .B(n14425), .Z(n14423) );
  XNOR U16471 ( .A(n14422), .B(n7213), .Z(n14425) );
  XNOR U16472 ( .A(n14418), .B(n14420), .Z(n7213) );
  NAND U16473 ( .A(n14426), .B(nreg[848]), .Z(n14420) );
  NAND U16474 ( .A(n12326), .B(nreg[848]), .Z(n14426) );
  XNOR U16475 ( .A(n14416), .B(n14427), .Z(n14418) );
  XOR U16476 ( .A(n14428), .B(n14429), .Z(n14416) );
  AND U16477 ( .A(n14430), .B(n14431), .Z(n14429) );
  XNOR U16478 ( .A(n14432), .B(n14428), .Z(n14431) );
  XOR U16479 ( .A(n14433), .B(nreg[848]), .Z(n14424) );
  IV U16480 ( .A(n14422), .Z(n14433) );
  XOR U16481 ( .A(n14434), .B(n14435), .Z(n14422) );
  AND U16482 ( .A(n14436), .B(n14437), .Z(n14435) );
  XNOR U16483 ( .A(n14434), .B(n7219), .Z(n14437) );
  XNOR U16484 ( .A(n14430), .B(n14432), .Z(n7219) );
  NAND U16485 ( .A(n14438), .B(nreg[847]), .Z(n14432) );
  NAND U16486 ( .A(n12326), .B(nreg[847]), .Z(n14438) );
  XNOR U16487 ( .A(n14428), .B(n14439), .Z(n14430) );
  XOR U16488 ( .A(n14440), .B(n14441), .Z(n14428) );
  AND U16489 ( .A(n14442), .B(n14443), .Z(n14441) );
  XNOR U16490 ( .A(n14444), .B(n14440), .Z(n14443) );
  XOR U16491 ( .A(n14445), .B(nreg[847]), .Z(n14436) );
  IV U16492 ( .A(n14434), .Z(n14445) );
  XOR U16493 ( .A(n14446), .B(n14447), .Z(n14434) );
  AND U16494 ( .A(n14448), .B(n14449), .Z(n14447) );
  XNOR U16495 ( .A(n14446), .B(n7225), .Z(n14449) );
  XNOR U16496 ( .A(n14442), .B(n14444), .Z(n7225) );
  NAND U16497 ( .A(n14450), .B(nreg[846]), .Z(n14444) );
  NAND U16498 ( .A(n12326), .B(nreg[846]), .Z(n14450) );
  XNOR U16499 ( .A(n14440), .B(n14451), .Z(n14442) );
  XOR U16500 ( .A(n14452), .B(n14453), .Z(n14440) );
  AND U16501 ( .A(n14454), .B(n14455), .Z(n14453) );
  XNOR U16502 ( .A(n14456), .B(n14452), .Z(n14455) );
  XOR U16503 ( .A(n14457), .B(nreg[846]), .Z(n14448) );
  IV U16504 ( .A(n14446), .Z(n14457) );
  XOR U16505 ( .A(n14458), .B(n14459), .Z(n14446) );
  AND U16506 ( .A(n14460), .B(n14461), .Z(n14459) );
  XNOR U16507 ( .A(n14458), .B(n7231), .Z(n14461) );
  XNOR U16508 ( .A(n14454), .B(n14456), .Z(n7231) );
  NAND U16509 ( .A(n14462), .B(nreg[845]), .Z(n14456) );
  NAND U16510 ( .A(n12326), .B(nreg[845]), .Z(n14462) );
  XNOR U16511 ( .A(n14452), .B(n14463), .Z(n14454) );
  XOR U16512 ( .A(n14464), .B(n14465), .Z(n14452) );
  AND U16513 ( .A(n14466), .B(n14467), .Z(n14465) );
  XNOR U16514 ( .A(n14468), .B(n14464), .Z(n14467) );
  XOR U16515 ( .A(n14469), .B(nreg[845]), .Z(n14460) );
  IV U16516 ( .A(n14458), .Z(n14469) );
  XOR U16517 ( .A(n14470), .B(n14471), .Z(n14458) );
  AND U16518 ( .A(n14472), .B(n14473), .Z(n14471) );
  XNOR U16519 ( .A(n14470), .B(n7237), .Z(n14473) );
  XNOR U16520 ( .A(n14466), .B(n14468), .Z(n7237) );
  NAND U16521 ( .A(n14474), .B(nreg[844]), .Z(n14468) );
  NAND U16522 ( .A(n12326), .B(nreg[844]), .Z(n14474) );
  XNOR U16523 ( .A(n14464), .B(n14475), .Z(n14466) );
  XOR U16524 ( .A(n14476), .B(n14477), .Z(n14464) );
  AND U16525 ( .A(n14478), .B(n14479), .Z(n14477) );
  XNOR U16526 ( .A(n14480), .B(n14476), .Z(n14479) );
  XOR U16527 ( .A(n14481), .B(nreg[844]), .Z(n14472) );
  IV U16528 ( .A(n14470), .Z(n14481) );
  XOR U16529 ( .A(n14482), .B(n14483), .Z(n14470) );
  AND U16530 ( .A(n14484), .B(n14485), .Z(n14483) );
  XNOR U16531 ( .A(n14482), .B(n7243), .Z(n14485) );
  XNOR U16532 ( .A(n14478), .B(n14480), .Z(n7243) );
  NAND U16533 ( .A(n14486), .B(nreg[843]), .Z(n14480) );
  NAND U16534 ( .A(n12326), .B(nreg[843]), .Z(n14486) );
  XNOR U16535 ( .A(n14476), .B(n14487), .Z(n14478) );
  XOR U16536 ( .A(n14488), .B(n14489), .Z(n14476) );
  AND U16537 ( .A(n14490), .B(n14491), .Z(n14489) );
  XNOR U16538 ( .A(n14492), .B(n14488), .Z(n14491) );
  XOR U16539 ( .A(n14493), .B(nreg[843]), .Z(n14484) );
  IV U16540 ( .A(n14482), .Z(n14493) );
  XOR U16541 ( .A(n14494), .B(n14495), .Z(n14482) );
  AND U16542 ( .A(n14496), .B(n14497), .Z(n14495) );
  XNOR U16543 ( .A(n14494), .B(n7249), .Z(n14497) );
  XNOR U16544 ( .A(n14490), .B(n14492), .Z(n7249) );
  NAND U16545 ( .A(n14498), .B(nreg[842]), .Z(n14492) );
  NAND U16546 ( .A(n12326), .B(nreg[842]), .Z(n14498) );
  XNOR U16547 ( .A(n14488), .B(n14499), .Z(n14490) );
  XOR U16548 ( .A(n14500), .B(n14501), .Z(n14488) );
  AND U16549 ( .A(n14502), .B(n14503), .Z(n14501) );
  XNOR U16550 ( .A(n14504), .B(n14500), .Z(n14503) );
  XOR U16551 ( .A(n14505), .B(nreg[842]), .Z(n14496) );
  IV U16552 ( .A(n14494), .Z(n14505) );
  XOR U16553 ( .A(n14506), .B(n14507), .Z(n14494) );
  AND U16554 ( .A(n14508), .B(n14509), .Z(n14507) );
  XNOR U16555 ( .A(n14506), .B(n7255), .Z(n14509) );
  XNOR U16556 ( .A(n14502), .B(n14504), .Z(n7255) );
  NAND U16557 ( .A(n14510), .B(nreg[841]), .Z(n14504) );
  NAND U16558 ( .A(n12326), .B(nreg[841]), .Z(n14510) );
  XNOR U16559 ( .A(n14500), .B(n14511), .Z(n14502) );
  XOR U16560 ( .A(n14512), .B(n14513), .Z(n14500) );
  AND U16561 ( .A(n14514), .B(n14515), .Z(n14513) );
  XNOR U16562 ( .A(n14516), .B(n14512), .Z(n14515) );
  XOR U16563 ( .A(n14517), .B(nreg[841]), .Z(n14508) );
  IV U16564 ( .A(n14506), .Z(n14517) );
  XOR U16565 ( .A(n14518), .B(n14519), .Z(n14506) );
  AND U16566 ( .A(n14520), .B(n14521), .Z(n14519) );
  XNOR U16567 ( .A(n14518), .B(n7261), .Z(n14521) );
  XNOR U16568 ( .A(n14514), .B(n14516), .Z(n7261) );
  NAND U16569 ( .A(n14522), .B(nreg[840]), .Z(n14516) );
  NAND U16570 ( .A(n12326), .B(nreg[840]), .Z(n14522) );
  XNOR U16571 ( .A(n14512), .B(n14523), .Z(n14514) );
  XOR U16572 ( .A(n14524), .B(n14525), .Z(n14512) );
  AND U16573 ( .A(n14526), .B(n14527), .Z(n14525) );
  XNOR U16574 ( .A(n14528), .B(n14524), .Z(n14527) );
  XOR U16575 ( .A(n14529), .B(nreg[840]), .Z(n14520) );
  IV U16576 ( .A(n14518), .Z(n14529) );
  XOR U16577 ( .A(n14530), .B(n14531), .Z(n14518) );
  AND U16578 ( .A(n14532), .B(n14533), .Z(n14531) );
  XNOR U16579 ( .A(n14530), .B(n7267), .Z(n14533) );
  XNOR U16580 ( .A(n14526), .B(n14528), .Z(n7267) );
  NAND U16581 ( .A(n14534), .B(nreg[839]), .Z(n14528) );
  NAND U16582 ( .A(n12326), .B(nreg[839]), .Z(n14534) );
  XNOR U16583 ( .A(n14524), .B(n14535), .Z(n14526) );
  XOR U16584 ( .A(n14536), .B(n14537), .Z(n14524) );
  AND U16585 ( .A(n14538), .B(n14539), .Z(n14537) );
  XNOR U16586 ( .A(n14540), .B(n14536), .Z(n14539) );
  XOR U16587 ( .A(n14541), .B(nreg[839]), .Z(n14532) );
  IV U16588 ( .A(n14530), .Z(n14541) );
  XOR U16589 ( .A(n14542), .B(n14543), .Z(n14530) );
  AND U16590 ( .A(n14544), .B(n14545), .Z(n14543) );
  XNOR U16591 ( .A(n14542), .B(n7273), .Z(n14545) );
  XNOR U16592 ( .A(n14538), .B(n14540), .Z(n7273) );
  NAND U16593 ( .A(n14546), .B(nreg[838]), .Z(n14540) );
  NAND U16594 ( .A(n12326), .B(nreg[838]), .Z(n14546) );
  XNOR U16595 ( .A(n14536), .B(n14547), .Z(n14538) );
  XOR U16596 ( .A(n14548), .B(n14549), .Z(n14536) );
  AND U16597 ( .A(n14550), .B(n14551), .Z(n14549) );
  XNOR U16598 ( .A(n14552), .B(n14548), .Z(n14551) );
  XOR U16599 ( .A(n14553), .B(nreg[838]), .Z(n14544) );
  IV U16600 ( .A(n14542), .Z(n14553) );
  XOR U16601 ( .A(n14554), .B(n14555), .Z(n14542) );
  AND U16602 ( .A(n14556), .B(n14557), .Z(n14555) );
  XNOR U16603 ( .A(n14554), .B(n7279), .Z(n14557) );
  XNOR U16604 ( .A(n14550), .B(n14552), .Z(n7279) );
  NAND U16605 ( .A(n14558), .B(nreg[837]), .Z(n14552) );
  NAND U16606 ( .A(n12326), .B(nreg[837]), .Z(n14558) );
  XNOR U16607 ( .A(n14548), .B(n14559), .Z(n14550) );
  XOR U16608 ( .A(n14560), .B(n14561), .Z(n14548) );
  AND U16609 ( .A(n14562), .B(n14563), .Z(n14561) );
  XNOR U16610 ( .A(n14564), .B(n14560), .Z(n14563) );
  XOR U16611 ( .A(n14565), .B(nreg[837]), .Z(n14556) );
  IV U16612 ( .A(n14554), .Z(n14565) );
  XOR U16613 ( .A(n14566), .B(n14567), .Z(n14554) );
  AND U16614 ( .A(n14568), .B(n14569), .Z(n14567) );
  XNOR U16615 ( .A(n14566), .B(n7285), .Z(n14569) );
  XNOR U16616 ( .A(n14562), .B(n14564), .Z(n7285) );
  NAND U16617 ( .A(n14570), .B(nreg[836]), .Z(n14564) );
  NAND U16618 ( .A(n12326), .B(nreg[836]), .Z(n14570) );
  XNOR U16619 ( .A(n14560), .B(n14571), .Z(n14562) );
  XOR U16620 ( .A(n14572), .B(n14573), .Z(n14560) );
  AND U16621 ( .A(n14574), .B(n14575), .Z(n14573) );
  XNOR U16622 ( .A(n14576), .B(n14572), .Z(n14575) );
  XOR U16623 ( .A(n14577), .B(nreg[836]), .Z(n14568) );
  IV U16624 ( .A(n14566), .Z(n14577) );
  XOR U16625 ( .A(n14578), .B(n14579), .Z(n14566) );
  AND U16626 ( .A(n14580), .B(n14581), .Z(n14579) );
  XNOR U16627 ( .A(n14578), .B(n7291), .Z(n14581) );
  XNOR U16628 ( .A(n14574), .B(n14576), .Z(n7291) );
  NAND U16629 ( .A(n14582), .B(nreg[835]), .Z(n14576) );
  NAND U16630 ( .A(n12326), .B(nreg[835]), .Z(n14582) );
  XNOR U16631 ( .A(n14572), .B(n14583), .Z(n14574) );
  XOR U16632 ( .A(n14584), .B(n14585), .Z(n14572) );
  AND U16633 ( .A(n14586), .B(n14587), .Z(n14585) );
  XNOR U16634 ( .A(n14588), .B(n14584), .Z(n14587) );
  XOR U16635 ( .A(n14589), .B(nreg[835]), .Z(n14580) );
  IV U16636 ( .A(n14578), .Z(n14589) );
  XOR U16637 ( .A(n14590), .B(n14591), .Z(n14578) );
  AND U16638 ( .A(n14592), .B(n14593), .Z(n14591) );
  XNOR U16639 ( .A(n14590), .B(n7297), .Z(n14593) );
  XNOR U16640 ( .A(n14586), .B(n14588), .Z(n7297) );
  NAND U16641 ( .A(n14594), .B(nreg[834]), .Z(n14588) );
  NAND U16642 ( .A(n12326), .B(nreg[834]), .Z(n14594) );
  XNOR U16643 ( .A(n14584), .B(n14595), .Z(n14586) );
  XOR U16644 ( .A(n14596), .B(n14597), .Z(n14584) );
  AND U16645 ( .A(n14598), .B(n14599), .Z(n14597) );
  XNOR U16646 ( .A(n14600), .B(n14596), .Z(n14599) );
  XOR U16647 ( .A(n14601), .B(nreg[834]), .Z(n14592) );
  IV U16648 ( .A(n14590), .Z(n14601) );
  XOR U16649 ( .A(n14602), .B(n14603), .Z(n14590) );
  AND U16650 ( .A(n14604), .B(n14605), .Z(n14603) );
  XNOR U16651 ( .A(n14602), .B(n7303), .Z(n14605) );
  XNOR U16652 ( .A(n14598), .B(n14600), .Z(n7303) );
  NAND U16653 ( .A(n14606), .B(nreg[833]), .Z(n14600) );
  NAND U16654 ( .A(n12326), .B(nreg[833]), .Z(n14606) );
  XNOR U16655 ( .A(n14596), .B(n14607), .Z(n14598) );
  XOR U16656 ( .A(n14608), .B(n14609), .Z(n14596) );
  AND U16657 ( .A(n14610), .B(n14611), .Z(n14609) );
  XNOR U16658 ( .A(n14612), .B(n14608), .Z(n14611) );
  XOR U16659 ( .A(n14613), .B(nreg[833]), .Z(n14604) );
  IV U16660 ( .A(n14602), .Z(n14613) );
  XOR U16661 ( .A(n14614), .B(n14615), .Z(n14602) );
  AND U16662 ( .A(n14616), .B(n14617), .Z(n14615) );
  XNOR U16663 ( .A(n14614), .B(n7309), .Z(n14617) );
  XNOR U16664 ( .A(n14610), .B(n14612), .Z(n7309) );
  NAND U16665 ( .A(n14618), .B(nreg[832]), .Z(n14612) );
  NAND U16666 ( .A(n12326), .B(nreg[832]), .Z(n14618) );
  XNOR U16667 ( .A(n14608), .B(n14619), .Z(n14610) );
  XOR U16668 ( .A(n14620), .B(n14621), .Z(n14608) );
  AND U16669 ( .A(n14622), .B(n14623), .Z(n14621) );
  XNOR U16670 ( .A(n14624), .B(n14620), .Z(n14623) );
  XOR U16671 ( .A(n14625), .B(nreg[832]), .Z(n14616) );
  IV U16672 ( .A(n14614), .Z(n14625) );
  XOR U16673 ( .A(n14626), .B(n14627), .Z(n14614) );
  AND U16674 ( .A(n14628), .B(n14629), .Z(n14627) );
  XNOR U16675 ( .A(n14626), .B(n7315), .Z(n14629) );
  XNOR U16676 ( .A(n14622), .B(n14624), .Z(n7315) );
  NAND U16677 ( .A(n14630), .B(nreg[831]), .Z(n14624) );
  NAND U16678 ( .A(n12326), .B(nreg[831]), .Z(n14630) );
  XNOR U16679 ( .A(n14620), .B(n14631), .Z(n14622) );
  XOR U16680 ( .A(n14632), .B(n14633), .Z(n14620) );
  AND U16681 ( .A(n14634), .B(n14635), .Z(n14633) );
  XNOR U16682 ( .A(n14636), .B(n14632), .Z(n14635) );
  XOR U16683 ( .A(n14637), .B(nreg[831]), .Z(n14628) );
  IV U16684 ( .A(n14626), .Z(n14637) );
  XOR U16685 ( .A(n14638), .B(n14639), .Z(n14626) );
  AND U16686 ( .A(n14640), .B(n14641), .Z(n14639) );
  XNOR U16687 ( .A(n14638), .B(n7321), .Z(n14641) );
  XNOR U16688 ( .A(n14634), .B(n14636), .Z(n7321) );
  NAND U16689 ( .A(n14642), .B(nreg[830]), .Z(n14636) );
  NAND U16690 ( .A(n12326), .B(nreg[830]), .Z(n14642) );
  XNOR U16691 ( .A(n14632), .B(n14643), .Z(n14634) );
  XOR U16692 ( .A(n14644), .B(n14645), .Z(n14632) );
  AND U16693 ( .A(n14646), .B(n14647), .Z(n14645) );
  XNOR U16694 ( .A(n14648), .B(n14644), .Z(n14647) );
  XOR U16695 ( .A(n14649), .B(nreg[830]), .Z(n14640) );
  IV U16696 ( .A(n14638), .Z(n14649) );
  XOR U16697 ( .A(n14650), .B(n14651), .Z(n14638) );
  AND U16698 ( .A(n14652), .B(n14653), .Z(n14651) );
  XNOR U16699 ( .A(n14650), .B(n7327), .Z(n14653) );
  XNOR U16700 ( .A(n14646), .B(n14648), .Z(n7327) );
  NAND U16701 ( .A(n14654), .B(nreg[829]), .Z(n14648) );
  NAND U16702 ( .A(n12326), .B(nreg[829]), .Z(n14654) );
  XNOR U16703 ( .A(n14644), .B(n14655), .Z(n14646) );
  XOR U16704 ( .A(n14656), .B(n14657), .Z(n14644) );
  AND U16705 ( .A(n14658), .B(n14659), .Z(n14657) );
  XNOR U16706 ( .A(n14660), .B(n14656), .Z(n14659) );
  XOR U16707 ( .A(n14661), .B(nreg[829]), .Z(n14652) );
  IV U16708 ( .A(n14650), .Z(n14661) );
  XOR U16709 ( .A(n14662), .B(n14663), .Z(n14650) );
  AND U16710 ( .A(n14664), .B(n14665), .Z(n14663) );
  XNOR U16711 ( .A(n14662), .B(n7333), .Z(n14665) );
  XNOR U16712 ( .A(n14658), .B(n14660), .Z(n7333) );
  NAND U16713 ( .A(n14666), .B(nreg[828]), .Z(n14660) );
  NAND U16714 ( .A(n12326), .B(nreg[828]), .Z(n14666) );
  XNOR U16715 ( .A(n14656), .B(n14667), .Z(n14658) );
  XOR U16716 ( .A(n14668), .B(n14669), .Z(n14656) );
  AND U16717 ( .A(n14670), .B(n14671), .Z(n14669) );
  XNOR U16718 ( .A(n14672), .B(n14668), .Z(n14671) );
  XOR U16719 ( .A(n14673), .B(nreg[828]), .Z(n14664) );
  IV U16720 ( .A(n14662), .Z(n14673) );
  XOR U16721 ( .A(n14674), .B(n14675), .Z(n14662) );
  AND U16722 ( .A(n14676), .B(n14677), .Z(n14675) );
  XNOR U16723 ( .A(n14674), .B(n7339), .Z(n14677) );
  XNOR U16724 ( .A(n14670), .B(n14672), .Z(n7339) );
  NAND U16725 ( .A(n14678), .B(nreg[827]), .Z(n14672) );
  NAND U16726 ( .A(n12326), .B(nreg[827]), .Z(n14678) );
  XNOR U16727 ( .A(n14668), .B(n14679), .Z(n14670) );
  XOR U16728 ( .A(n14680), .B(n14681), .Z(n14668) );
  AND U16729 ( .A(n14682), .B(n14683), .Z(n14681) );
  XNOR U16730 ( .A(n14684), .B(n14680), .Z(n14683) );
  XOR U16731 ( .A(n14685), .B(nreg[827]), .Z(n14676) );
  IV U16732 ( .A(n14674), .Z(n14685) );
  XOR U16733 ( .A(n14686), .B(n14687), .Z(n14674) );
  AND U16734 ( .A(n14688), .B(n14689), .Z(n14687) );
  XNOR U16735 ( .A(n14686), .B(n7345), .Z(n14689) );
  XNOR U16736 ( .A(n14682), .B(n14684), .Z(n7345) );
  NAND U16737 ( .A(n14690), .B(nreg[826]), .Z(n14684) );
  NAND U16738 ( .A(n12326), .B(nreg[826]), .Z(n14690) );
  XNOR U16739 ( .A(n14680), .B(n14691), .Z(n14682) );
  XOR U16740 ( .A(n14692), .B(n14693), .Z(n14680) );
  AND U16741 ( .A(n14694), .B(n14695), .Z(n14693) );
  XNOR U16742 ( .A(n14696), .B(n14692), .Z(n14695) );
  XOR U16743 ( .A(n14697), .B(nreg[826]), .Z(n14688) );
  IV U16744 ( .A(n14686), .Z(n14697) );
  XOR U16745 ( .A(n14698), .B(n14699), .Z(n14686) );
  AND U16746 ( .A(n14700), .B(n14701), .Z(n14699) );
  XNOR U16747 ( .A(n14698), .B(n7351), .Z(n14701) );
  XNOR U16748 ( .A(n14694), .B(n14696), .Z(n7351) );
  NAND U16749 ( .A(n14702), .B(nreg[825]), .Z(n14696) );
  NAND U16750 ( .A(n12326), .B(nreg[825]), .Z(n14702) );
  XNOR U16751 ( .A(n14692), .B(n14703), .Z(n14694) );
  XOR U16752 ( .A(n14704), .B(n14705), .Z(n14692) );
  AND U16753 ( .A(n14706), .B(n14707), .Z(n14705) );
  XNOR U16754 ( .A(n14708), .B(n14704), .Z(n14707) );
  XOR U16755 ( .A(n14709), .B(nreg[825]), .Z(n14700) );
  IV U16756 ( .A(n14698), .Z(n14709) );
  XOR U16757 ( .A(n14710), .B(n14711), .Z(n14698) );
  AND U16758 ( .A(n14712), .B(n14713), .Z(n14711) );
  XNOR U16759 ( .A(n14710), .B(n7357), .Z(n14713) );
  XNOR U16760 ( .A(n14706), .B(n14708), .Z(n7357) );
  NAND U16761 ( .A(n14714), .B(nreg[824]), .Z(n14708) );
  NAND U16762 ( .A(n12326), .B(nreg[824]), .Z(n14714) );
  XNOR U16763 ( .A(n14704), .B(n14715), .Z(n14706) );
  XOR U16764 ( .A(n14716), .B(n14717), .Z(n14704) );
  AND U16765 ( .A(n14718), .B(n14719), .Z(n14717) );
  XNOR U16766 ( .A(n14720), .B(n14716), .Z(n14719) );
  XOR U16767 ( .A(n14721), .B(nreg[824]), .Z(n14712) );
  IV U16768 ( .A(n14710), .Z(n14721) );
  XOR U16769 ( .A(n14722), .B(n14723), .Z(n14710) );
  AND U16770 ( .A(n14724), .B(n14725), .Z(n14723) );
  XNOR U16771 ( .A(n14722), .B(n7363), .Z(n14725) );
  XNOR U16772 ( .A(n14718), .B(n14720), .Z(n7363) );
  NAND U16773 ( .A(n14726), .B(nreg[823]), .Z(n14720) );
  NAND U16774 ( .A(n12326), .B(nreg[823]), .Z(n14726) );
  XNOR U16775 ( .A(n14716), .B(n14727), .Z(n14718) );
  XOR U16776 ( .A(n14728), .B(n14729), .Z(n14716) );
  AND U16777 ( .A(n14730), .B(n14731), .Z(n14729) );
  XNOR U16778 ( .A(n14732), .B(n14728), .Z(n14731) );
  XOR U16779 ( .A(n14733), .B(nreg[823]), .Z(n14724) );
  IV U16780 ( .A(n14722), .Z(n14733) );
  XOR U16781 ( .A(n14734), .B(n14735), .Z(n14722) );
  AND U16782 ( .A(n14736), .B(n14737), .Z(n14735) );
  XNOR U16783 ( .A(n14734), .B(n7369), .Z(n14737) );
  XNOR U16784 ( .A(n14730), .B(n14732), .Z(n7369) );
  NAND U16785 ( .A(n14738), .B(nreg[822]), .Z(n14732) );
  NAND U16786 ( .A(n12326), .B(nreg[822]), .Z(n14738) );
  XNOR U16787 ( .A(n14728), .B(n14739), .Z(n14730) );
  XOR U16788 ( .A(n14740), .B(n14741), .Z(n14728) );
  AND U16789 ( .A(n14742), .B(n14743), .Z(n14741) );
  XNOR U16790 ( .A(n14744), .B(n14740), .Z(n14743) );
  XOR U16791 ( .A(n14745), .B(nreg[822]), .Z(n14736) );
  IV U16792 ( .A(n14734), .Z(n14745) );
  XOR U16793 ( .A(n14746), .B(n14747), .Z(n14734) );
  AND U16794 ( .A(n14748), .B(n14749), .Z(n14747) );
  XNOR U16795 ( .A(n14746), .B(n7375), .Z(n14749) );
  XNOR U16796 ( .A(n14742), .B(n14744), .Z(n7375) );
  NAND U16797 ( .A(n14750), .B(nreg[821]), .Z(n14744) );
  NAND U16798 ( .A(n12326), .B(nreg[821]), .Z(n14750) );
  XNOR U16799 ( .A(n14740), .B(n14751), .Z(n14742) );
  XOR U16800 ( .A(n14752), .B(n14753), .Z(n14740) );
  AND U16801 ( .A(n14754), .B(n14755), .Z(n14753) );
  XNOR U16802 ( .A(n14756), .B(n14752), .Z(n14755) );
  XOR U16803 ( .A(n14757), .B(nreg[821]), .Z(n14748) );
  IV U16804 ( .A(n14746), .Z(n14757) );
  XOR U16805 ( .A(n14758), .B(n14759), .Z(n14746) );
  AND U16806 ( .A(n14760), .B(n14761), .Z(n14759) );
  XNOR U16807 ( .A(n14758), .B(n7381), .Z(n14761) );
  XNOR U16808 ( .A(n14754), .B(n14756), .Z(n7381) );
  NAND U16809 ( .A(n14762), .B(nreg[820]), .Z(n14756) );
  NAND U16810 ( .A(n12326), .B(nreg[820]), .Z(n14762) );
  XNOR U16811 ( .A(n14752), .B(n14763), .Z(n14754) );
  XOR U16812 ( .A(n14764), .B(n14765), .Z(n14752) );
  AND U16813 ( .A(n14766), .B(n14767), .Z(n14765) );
  XNOR U16814 ( .A(n14768), .B(n14764), .Z(n14767) );
  XOR U16815 ( .A(n14769), .B(nreg[820]), .Z(n14760) );
  IV U16816 ( .A(n14758), .Z(n14769) );
  XOR U16817 ( .A(n14770), .B(n14771), .Z(n14758) );
  AND U16818 ( .A(n14772), .B(n14773), .Z(n14771) );
  XNOR U16819 ( .A(n14770), .B(n7387), .Z(n14773) );
  XNOR U16820 ( .A(n14766), .B(n14768), .Z(n7387) );
  NAND U16821 ( .A(n14774), .B(nreg[819]), .Z(n14768) );
  NAND U16822 ( .A(n12326), .B(nreg[819]), .Z(n14774) );
  XNOR U16823 ( .A(n14764), .B(n14775), .Z(n14766) );
  XOR U16824 ( .A(n14776), .B(n14777), .Z(n14764) );
  AND U16825 ( .A(n14778), .B(n14779), .Z(n14777) );
  XNOR U16826 ( .A(n14780), .B(n14776), .Z(n14779) );
  XOR U16827 ( .A(n14781), .B(nreg[819]), .Z(n14772) );
  IV U16828 ( .A(n14770), .Z(n14781) );
  XOR U16829 ( .A(n14782), .B(n14783), .Z(n14770) );
  AND U16830 ( .A(n14784), .B(n14785), .Z(n14783) );
  XNOR U16831 ( .A(n14782), .B(n7393), .Z(n14785) );
  XNOR U16832 ( .A(n14778), .B(n14780), .Z(n7393) );
  NAND U16833 ( .A(n14786), .B(nreg[818]), .Z(n14780) );
  NAND U16834 ( .A(n12326), .B(nreg[818]), .Z(n14786) );
  XNOR U16835 ( .A(n14776), .B(n14787), .Z(n14778) );
  XOR U16836 ( .A(n14788), .B(n14789), .Z(n14776) );
  AND U16837 ( .A(n14790), .B(n14791), .Z(n14789) );
  XNOR U16838 ( .A(n14792), .B(n14788), .Z(n14791) );
  XOR U16839 ( .A(n14793), .B(nreg[818]), .Z(n14784) );
  IV U16840 ( .A(n14782), .Z(n14793) );
  XOR U16841 ( .A(n14794), .B(n14795), .Z(n14782) );
  AND U16842 ( .A(n14796), .B(n14797), .Z(n14795) );
  XNOR U16843 ( .A(n14794), .B(n7399), .Z(n14797) );
  XNOR U16844 ( .A(n14790), .B(n14792), .Z(n7399) );
  NAND U16845 ( .A(n14798), .B(nreg[817]), .Z(n14792) );
  NAND U16846 ( .A(n12326), .B(nreg[817]), .Z(n14798) );
  XNOR U16847 ( .A(n14788), .B(n14799), .Z(n14790) );
  XOR U16848 ( .A(n14800), .B(n14801), .Z(n14788) );
  AND U16849 ( .A(n14802), .B(n14803), .Z(n14801) );
  XNOR U16850 ( .A(n14804), .B(n14800), .Z(n14803) );
  XOR U16851 ( .A(n14805), .B(nreg[817]), .Z(n14796) );
  IV U16852 ( .A(n14794), .Z(n14805) );
  XOR U16853 ( .A(n14806), .B(n14807), .Z(n14794) );
  AND U16854 ( .A(n14808), .B(n14809), .Z(n14807) );
  XNOR U16855 ( .A(n14806), .B(n7405), .Z(n14809) );
  XNOR U16856 ( .A(n14802), .B(n14804), .Z(n7405) );
  NAND U16857 ( .A(n14810), .B(nreg[816]), .Z(n14804) );
  NAND U16858 ( .A(n12326), .B(nreg[816]), .Z(n14810) );
  XNOR U16859 ( .A(n14800), .B(n14811), .Z(n14802) );
  XOR U16860 ( .A(n14812), .B(n14813), .Z(n14800) );
  AND U16861 ( .A(n14814), .B(n14815), .Z(n14813) );
  XNOR U16862 ( .A(n14816), .B(n14812), .Z(n14815) );
  XOR U16863 ( .A(n14817), .B(nreg[816]), .Z(n14808) );
  IV U16864 ( .A(n14806), .Z(n14817) );
  XOR U16865 ( .A(n14818), .B(n14819), .Z(n14806) );
  AND U16866 ( .A(n14820), .B(n14821), .Z(n14819) );
  XNOR U16867 ( .A(n14818), .B(n7411), .Z(n14821) );
  XNOR U16868 ( .A(n14814), .B(n14816), .Z(n7411) );
  NAND U16869 ( .A(n14822), .B(nreg[815]), .Z(n14816) );
  NAND U16870 ( .A(n12326), .B(nreg[815]), .Z(n14822) );
  XNOR U16871 ( .A(n14812), .B(n14823), .Z(n14814) );
  XOR U16872 ( .A(n14824), .B(n14825), .Z(n14812) );
  AND U16873 ( .A(n14826), .B(n14827), .Z(n14825) );
  XNOR U16874 ( .A(n14828), .B(n14824), .Z(n14827) );
  XOR U16875 ( .A(n14829), .B(nreg[815]), .Z(n14820) );
  IV U16876 ( .A(n14818), .Z(n14829) );
  XOR U16877 ( .A(n14830), .B(n14831), .Z(n14818) );
  AND U16878 ( .A(n14832), .B(n14833), .Z(n14831) );
  XNOR U16879 ( .A(n14830), .B(n7417), .Z(n14833) );
  XNOR U16880 ( .A(n14826), .B(n14828), .Z(n7417) );
  NAND U16881 ( .A(n14834), .B(nreg[814]), .Z(n14828) );
  NAND U16882 ( .A(n12326), .B(nreg[814]), .Z(n14834) );
  XNOR U16883 ( .A(n14824), .B(n14835), .Z(n14826) );
  XOR U16884 ( .A(n14836), .B(n14837), .Z(n14824) );
  AND U16885 ( .A(n14838), .B(n14839), .Z(n14837) );
  XNOR U16886 ( .A(n14840), .B(n14836), .Z(n14839) );
  XOR U16887 ( .A(n14841), .B(nreg[814]), .Z(n14832) );
  IV U16888 ( .A(n14830), .Z(n14841) );
  XOR U16889 ( .A(n14842), .B(n14843), .Z(n14830) );
  AND U16890 ( .A(n14844), .B(n14845), .Z(n14843) );
  XNOR U16891 ( .A(n14842), .B(n7423), .Z(n14845) );
  XNOR U16892 ( .A(n14838), .B(n14840), .Z(n7423) );
  NAND U16893 ( .A(n14846), .B(nreg[813]), .Z(n14840) );
  NAND U16894 ( .A(n12326), .B(nreg[813]), .Z(n14846) );
  XNOR U16895 ( .A(n14836), .B(n14847), .Z(n14838) );
  XOR U16896 ( .A(n14848), .B(n14849), .Z(n14836) );
  AND U16897 ( .A(n14850), .B(n14851), .Z(n14849) );
  XNOR U16898 ( .A(n14852), .B(n14848), .Z(n14851) );
  XOR U16899 ( .A(n14853), .B(nreg[813]), .Z(n14844) );
  IV U16900 ( .A(n14842), .Z(n14853) );
  XOR U16901 ( .A(n14854), .B(n14855), .Z(n14842) );
  AND U16902 ( .A(n14856), .B(n14857), .Z(n14855) );
  XNOR U16903 ( .A(n14854), .B(n7429), .Z(n14857) );
  XNOR U16904 ( .A(n14850), .B(n14852), .Z(n7429) );
  NAND U16905 ( .A(n14858), .B(nreg[812]), .Z(n14852) );
  NAND U16906 ( .A(n12326), .B(nreg[812]), .Z(n14858) );
  XNOR U16907 ( .A(n14848), .B(n14859), .Z(n14850) );
  XOR U16908 ( .A(n14860), .B(n14861), .Z(n14848) );
  AND U16909 ( .A(n14862), .B(n14863), .Z(n14861) );
  XNOR U16910 ( .A(n14864), .B(n14860), .Z(n14863) );
  XOR U16911 ( .A(n14865), .B(nreg[812]), .Z(n14856) );
  IV U16912 ( .A(n14854), .Z(n14865) );
  XOR U16913 ( .A(n14866), .B(n14867), .Z(n14854) );
  AND U16914 ( .A(n14868), .B(n14869), .Z(n14867) );
  XNOR U16915 ( .A(n14866), .B(n7435), .Z(n14869) );
  XNOR U16916 ( .A(n14862), .B(n14864), .Z(n7435) );
  NAND U16917 ( .A(n14870), .B(nreg[811]), .Z(n14864) );
  NAND U16918 ( .A(n12326), .B(nreg[811]), .Z(n14870) );
  XNOR U16919 ( .A(n14860), .B(n14871), .Z(n14862) );
  XOR U16920 ( .A(n14872), .B(n14873), .Z(n14860) );
  AND U16921 ( .A(n14874), .B(n14875), .Z(n14873) );
  XNOR U16922 ( .A(n14876), .B(n14872), .Z(n14875) );
  XOR U16923 ( .A(n14877), .B(nreg[811]), .Z(n14868) );
  IV U16924 ( .A(n14866), .Z(n14877) );
  XOR U16925 ( .A(n14878), .B(n14879), .Z(n14866) );
  AND U16926 ( .A(n14880), .B(n14881), .Z(n14879) );
  XNOR U16927 ( .A(n14878), .B(n7441), .Z(n14881) );
  XNOR U16928 ( .A(n14874), .B(n14876), .Z(n7441) );
  NAND U16929 ( .A(n14882), .B(nreg[810]), .Z(n14876) );
  NAND U16930 ( .A(n12326), .B(nreg[810]), .Z(n14882) );
  XNOR U16931 ( .A(n14872), .B(n14883), .Z(n14874) );
  XOR U16932 ( .A(n14884), .B(n14885), .Z(n14872) );
  AND U16933 ( .A(n14886), .B(n14887), .Z(n14885) );
  XNOR U16934 ( .A(n14888), .B(n14884), .Z(n14887) );
  XOR U16935 ( .A(n14889), .B(nreg[810]), .Z(n14880) );
  IV U16936 ( .A(n14878), .Z(n14889) );
  XOR U16937 ( .A(n14890), .B(n14891), .Z(n14878) );
  AND U16938 ( .A(n14892), .B(n14893), .Z(n14891) );
  XNOR U16939 ( .A(n14890), .B(n7447), .Z(n14893) );
  XNOR U16940 ( .A(n14886), .B(n14888), .Z(n7447) );
  NAND U16941 ( .A(n14894), .B(nreg[809]), .Z(n14888) );
  NAND U16942 ( .A(n12326), .B(nreg[809]), .Z(n14894) );
  XNOR U16943 ( .A(n14884), .B(n14895), .Z(n14886) );
  XOR U16944 ( .A(n14896), .B(n14897), .Z(n14884) );
  AND U16945 ( .A(n14898), .B(n14899), .Z(n14897) );
  XNOR U16946 ( .A(n14900), .B(n14896), .Z(n14899) );
  XOR U16947 ( .A(n14901), .B(nreg[809]), .Z(n14892) );
  IV U16948 ( .A(n14890), .Z(n14901) );
  XOR U16949 ( .A(n14902), .B(n14903), .Z(n14890) );
  AND U16950 ( .A(n14904), .B(n14905), .Z(n14903) );
  XNOR U16951 ( .A(n14902), .B(n7453), .Z(n14905) );
  XNOR U16952 ( .A(n14898), .B(n14900), .Z(n7453) );
  NAND U16953 ( .A(n14906), .B(nreg[808]), .Z(n14900) );
  NAND U16954 ( .A(n12326), .B(nreg[808]), .Z(n14906) );
  XNOR U16955 ( .A(n14896), .B(n14907), .Z(n14898) );
  XOR U16956 ( .A(n14908), .B(n14909), .Z(n14896) );
  AND U16957 ( .A(n14910), .B(n14911), .Z(n14909) );
  XNOR U16958 ( .A(n14912), .B(n14908), .Z(n14911) );
  XOR U16959 ( .A(n14913), .B(nreg[808]), .Z(n14904) );
  IV U16960 ( .A(n14902), .Z(n14913) );
  XOR U16961 ( .A(n14914), .B(n14915), .Z(n14902) );
  AND U16962 ( .A(n14916), .B(n14917), .Z(n14915) );
  XNOR U16963 ( .A(n14914), .B(n7459), .Z(n14917) );
  XNOR U16964 ( .A(n14910), .B(n14912), .Z(n7459) );
  NAND U16965 ( .A(n14918), .B(nreg[807]), .Z(n14912) );
  NAND U16966 ( .A(n12326), .B(nreg[807]), .Z(n14918) );
  XNOR U16967 ( .A(n14908), .B(n14919), .Z(n14910) );
  XOR U16968 ( .A(n14920), .B(n14921), .Z(n14908) );
  AND U16969 ( .A(n14922), .B(n14923), .Z(n14921) );
  XNOR U16970 ( .A(n14924), .B(n14920), .Z(n14923) );
  XOR U16971 ( .A(n14925), .B(nreg[807]), .Z(n14916) );
  IV U16972 ( .A(n14914), .Z(n14925) );
  XOR U16973 ( .A(n14926), .B(n14927), .Z(n14914) );
  AND U16974 ( .A(n14928), .B(n14929), .Z(n14927) );
  XNOR U16975 ( .A(n14926), .B(n7465), .Z(n14929) );
  XNOR U16976 ( .A(n14922), .B(n14924), .Z(n7465) );
  NAND U16977 ( .A(n14930), .B(nreg[806]), .Z(n14924) );
  NAND U16978 ( .A(n12326), .B(nreg[806]), .Z(n14930) );
  XNOR U16979 ( .A(n14920), .B(n14931), .Z(n14922) );
  XOR U16980 ( .A(n14932), .B(n14933), .Z(n14920) );
  AND U16981 ( .A(n14934), .B(n14935), .Z(n14933) );
  XNOR U16982 ( .A(n14936), .B(n14932), .Z(n14935) );
  XOR U16983 ( .A(n14937), .B(nreg[806]), .Z(n14928) );
  IV U16984 ( .A(n14926), .Z(n14937) );
  XOR U16985 ( .A(n14938), .B(n14939), .Z(n14926) );
  AND U16986 ( .A(n14940), .B(n14941), .Z(n14939) );
  XNOR U16987 ( .A(n14938), .B(n7471), .Z(n14941) );
  XNOR U16988 ( .A(n14934), .B(n14936), .Z(n7471) );
  NAND U16989 ( .A(n14942), .B(nreg[805]), .Z(n14936) );
  NAND U16990 ( .A(n12326), .B(nreg[805]), .Z(n14942) );
  XNOR U16991 ( .A(n14932), .B(n14943), .Z(n14934) );
  XOR U16992 ( .A(n14944), .B(n14945), .Z(n14932) );
  AND U16993 ( .A(n14946), .B(n14947), .Z(n14945) );
  XNOR U16994 ( .A(n14948), .B(n14944), .Z(n14947) );
  XOR U16995 ( .A(n14949), .B(nreg[805]), .Z(n14940) );
  IV U16996 ( .A(n14938), .Z(n14949) );
  XOR U16997 ( .A(n14950), .B(n14951), .Z(n14938) );
  AND U16998 ( .A(n14952), .B(n14953), .Z(n14951) );
  XNOR U16999 ( .A(n14950), .B(n7477), .Z(n14953) );
  XNOR U17000 ( .A(n14946), .B(n14948), .Z(n7477) );
  NAND U17001 ( .A(n14954), .B(nreg[804]), .Z(n14948) );
  NAND U17002 ( .A(n12326), .B(nreg[804]), .Z(n14954) );
  XNOR U17003 ( .A(n14944), .B(n14955), .Z(n14946) );
  XOR U17004 ( .A(n14956), .B(n14957), .Z(n14944) );
  AND U17005 ( .A(n14958), .B(n14959), .Z(n14957) );
  XNOR U17006 ( .A(n14960), .B(n14956), .Z(n14959) );
  XOR U17007 ( .A(n14961), .B(nreg[804]), .Z(n14952) );
  IV U17008 ( .A(n14950), .Z(n14961) );
  XOR U17009 ( .A(n14962), .B(n14963), .Z(n14950) );
  AND U17010 ( .A(n14964), .B(n14965), .Z(n14963) );
  XNOR U17011 ( .A(n14962), .B(n7483), .Z(n14965) );
  XNOR U17012 ( .A(n14958), .B(n14960), .Z(n7483) );
  NAND U17013 ( .A(n14966), .B(nreg[803]), .Z(n14960) );
  NAND U17014 ( .A(n12326), .B(nreg[803]), .Z(n14966) );
  XNOR U17015 ( .A(n14956), .B(n14967), .Z(n14958) );
  XOR U17016 ( .A(n14968), .B(n14969), .Z(n14956) );
  AND U17017 ( .A(n14970), .B(n14971), .Z(n14969) );
  XNOR U17018 ( .A(n14972), .B(n14968), .Z(n14971) );
  XOR U17019 ( .A(n14973), .B(nreg[803]), .Z(n14964) );
  IV U17020 ( .A(n14962), .Z(n14973) );
  XOR U17021 ( .A(n14974), .B(n14975), .Z(n14962) );
  AND U17022 ( .A(n14976), .B(n14977), .Z(n14975) );
  XNOR U17023 ( .A(n14974), .B(n7489), .Z(n14977) );
  XNOR U17024 ( .A(n14970), .B(n14972), .Z(n7489) );
  NAND U17025 ( .A(n14978), .B(nreg[802]), .Z(n14972) );
  NAND U17026 ( .A(n12326), .B(nreg[802]), .Z(n14978) );
  XNOR U17027 ( .A(n14968), .B(n14979), .Z(n14970) );
  XOR U17028 ( .A(n14980), .B(n14981), .Z(n14968) );
  AND U17029 ( .A(n14982), .B(n14983), .Z(n14981) );
  XNOR U17030 ( .A(n14984), .B(n14980), .Z(n14983) );
  XOR U17031 ( .A(n14985), .B(nreg[802]), .Z(n14976) );
  IV U17032 ( .A(n14974), .Z(n14985) );
  XOR U17033 ( .A(n14986), .B(n14987), .Z(n14974) );
  AND U17034 ( .A(n14988), .B(n14989), .Z(n14987) );
  XNOR U17035 ( .A(n14986), .B(n7495), .Z(n14989) );
  XNOR U17036 ( .A(n14982), .B(n14984), .Z(n7495) );
  NAND U17037 ( .A(n14990), .B(nreg[801]), .Z(n14984) );
  NAND U17038 ( .A(n12326), .B(nreg[801]), .Z(n14990) );
  XNOR U17039 ( .A(n14980), .B(n14991), .Z(n14982) );
  XOR U17040 ( .A(n14992), .B(n14993), .Z(n14980) );
  AND U17041 ( .A(n14994), .B(n14995), .Z(n14993) );
  XNOR U17042 ( .A(n14996), .B(n14992), .Z(n14995) );
  XOR U17043 ( .A(n14997), .B(nreg[801]), .Z(n14988) );
  IV U17044 ( .A(n14986), .Z(n14997) );
  XOR U17045 ( .A(n14998), .B(n14999), .Z(n14986) );
  AND U17046 ( .A(n15000), .B(n15001), .Z(n14999) );
  XNOR U17047 ( .A(n14998), .B(n7501), .Z(n15001) );
  XNOR U17048 ( .A(n14994), .B(n14996), .Z(n7501) );
  NAND U17049 ( .A(n15002), .B(nreg[800]), .Z(n14996) );
  NAND U17050 ( .A(n12326), .B(nreg[800]), .Z(n15002) );
  XNOR U17051 ( .A(n14992), .B(n15003), .Z(n14994) );
  XOR U17052 ( .A(n15004), .B(n15005), .Z(n14992) );
  AND U17053 ( .A(n15006), .B(n15007), .Z(n15005) );
  XNOR U17054 ( .A(n15008), .B(n15004), .Z(n15007) );
  XOR U17055 ( .A(n15009), .B(nreg[800]), .Z(n15000) );
  IV U17056 ( .A(n14998), .Z(n15009) );
  XOR U17057 ( .A(n15010), .B(n15011), .Z(n14998) );
  AND U17058 ( .A(n15012), .B(n15013), .Z(n15011) );
  XNOR U17059 ( .A(n15010), .B(n7507), .Z(n15013) );
  XNOR U17060 ( .A(n15006), .B(n15008), .Z(n7507) );
  NAND U17061 ( .A(n15014), .B(nreg[799]), .Z(n15008) );
  NAND U17062 ( .A(n12326), .B(nreg[799]), .Z(n15014) );
  XNOR U17063 ( .A(n15004), .B(n15015), .Z(n15006) );
  XOR U17064 ( .A(n15016), .B(n15017), .Z(n15004) );
  AND U17065 ( .A(n15018), .B(n15019), .Z(n15017) );
  XNOR U17066 ( .A(n15020), .B(n15016), .Z(n15019) );
  XOR U17067 ( .A(n15021), .B(nreg[799]), .Z(n15012) );
  IV U17068 ( .A(n15010), .Z(n15021) );
  XOR U17069 ( .A(n15022), .B(n15023), .Z(n15010) );
  AND U17070 ( .A(n15024), .B(n15025), .Z(n15023) );
  XNOR U17071 ( .A(n15022), .B(n7513), .Z(n15025) );
  XNOR U17072 ( .A(n15018), .B(n15020), .Z(n7513) );
  NAND U17073 ( .A(n15026), .B(nreg[798]), .Z(n15020) );
  NAND U17074 ( .A(n12326), .B(nreg[798]), .Z(n15026) );
  XNOR U17075 ( .A(n15016), .B(n15027), .Z(n15018) );
  XOR U17076 ( .A(n15028), .B(n15029), .Z(n15016) );
  AND U17077 ( .A(n15030), .B(n15031), .Z(n15029) );
  XNOR U17078 ( .A(n15032), .B(n15028), .Z(n15031) );
  XOR U17079 ( .A(n15033), .B(nreg[798]), .Z(n15024) );
  IV U17080 ( .A(n15022), .Z(n15033) );
  XOR U17081 ( .A(n15034), .B(n15035), .Z(n15022) );
  AND U17082 ( .A(n15036), .B(n15037), .Z(n15035) );
  XNOR U17083 ( .A(n15034), .B(n7519), .Z(n15037) );
  XNOR U17084 ( .A(n15030), .B(n15032), .Z(n7519) );
  NAND U17085 ( .A(n15038), .B(nreg[797]), .Z(n15032) );
  NAND U17086 ( .A(n12326), .B(nreg[797]), .Z(n15038) );
  XNOR U17087 ( .A(n15028), .B(n15039), .Z(n15030) );
  XOR U17088 ( .A(n15040), .B(n15041), .Z(n15028) );
  AND U17089 ( .A(n15042), .B(n15043), .Z(n15041) );
  XNOR U17090 ( .A(n15044), .B(n15040), .Z(n15043) );
  XOR U17091 ( .A(n15045), .B(nreg[797]), .Z(n15036) );
  IV U17092 ( .A(n15034), .Z(n15045) );
  XOR U17093 ( .A(n15046), .B(n15047), .Z(n15034) );
  AND U17094 ( .A(n15048), .B(n15049), .Z(n15047) );
  XNOR U17095 ( .A(n15046), .B(n7525), .Z(n15049) );
  XNOR U17096 ( .A(n15042), .B(n15044), .Z(n7525) );
  NAND U17097 ( .A(n15050), .B(nreg[796]), .Z(n15044) );
  NAND U17098 ( .A(n12326), .B(nreg[796]), .Z(n15050) );
  XNOR U17099 ( .A(n15040), .B(n15051), .Z(n15042) );
  XOR U17100 ( .A(n15052), .B(n15053), .Z(n15040) );
  AND U17101 ( .A(n15054), .B(n15055), .Z(n15053) );
  XNOR U17102 ( .A(n15056), .B(n15052), .Z(n15055) );
  XOR U17103 ( .A(n15057), .B(nreg[796]), .Z(n15048) );
  IV U17104 ( .A(n15046), .Z(n15057) );
  XOR U17105 ( .A(n15058), .B(n15059), .Z(n15046) );
  AND U17106 ( .A(n15060), .B(n15061), .Z(n15059) );
  XNOR U17107 ( .A(n15058), .B(n7531), .Z(n15061) );
  XNOR U17108 ( .A(n15054), .B(n15056), .Z(n7531) );
  NAND U17109 ( .A(n15062), .B(nreg[795]), .Z(n15056) );
  NAND U17110 ( .A(n12326), .B(nreg[795]), .Z(n15062) );
  XNOR U17111 ( .A(n15052), .B(n15063), .Z(n15054) );
  XOR U17112 ( .A(n15064), .B(n15065), .Z(n15052) );
  AND U17113 ( .A(n15066), .B(n15067), .Z(n15065) );
  XNOR U17114 ( .A(n15068), .B(n15064), .Z(n15067) );
  XOR U17115 ( .A(n15069), .B(nreg[795]), .Z(n15060) );
  IV U17116 ( .A(n15058), .Z(n15069) );
  XOR U17117 ( .A(n15070), .B(n15071), .Z(n15058) );
  AND U17118 ( .A(n15072), .B(n15073), .Z(n15071) );
  XNOR U17119 ( .A(n15070), .B(n7537), .Z(n15073) );
  XNOR U17120 ( .A(n15066), .B(n15068), .Z(n7537) );
  NAND U17121 ( .A(n15074), .B(nreg[794]), .Z(n15068) );
  NAND U17122 ( .A(n12326), .B(nreg[794]), .Z(n15074) );
  XNOR U17123 ( .A(n15064), .B(n15075), .Z(n15066) );
  XOR U17124 ( .A(n15076), .B(n15077), .Z(n15064) );
  AND U17125 ( .A(n15078), .B(n15079), .Z(n15077) );
  XNOR U17126 ( .A(n15080), .B(n15076), .Z(n15079) );
  XOR U17127 ( .A(n15081), .B(nreg[794]), .Z(n15072) );
  IV U17128 ( .A(n15070), .Z(n15081) );
  XOR U17129 ( .A(n15082), .B(n15083), .Z(n15070) );
  AND U17130 ( .A(n15084), .B(n15085), .Z(n15083) );
  XNOR U17131 ( .A(n15082), .B(n7543), .Z(n15085) );
  XNOR U17132 ( .A(n15078), .B(n15080), .Z(n7543) );
  NAND U17133 ( .A(n15086), .B(nreg[793]), .Z(n15080) );
  NAND U17134 ( .A(n12326), .B(nreg[793]), .Z(n15086) );
  XNOR U17135 ( .A(n15076), .B(n15087), .Z(n15078) );
  XOR U17136 ( .A(n15088), .B(n15089), .Z(n15076) );
  AND U17137 ( .A(n15090), .B(n15091), .Z(n15089) );
  XNOR U17138 ( .A(n15092), .B(n15088), .Z(n15091) );
  XOR U17139 ( .A(n15093), .B(nreg[793]), .Z(n15084) );
  IV U17140 ( .A(n15082), .Z(n15093) );
  XOR U17141 ( .A(n15094), .B(n15095), .Z(n15082) );
  AND U17142 ( .A(n15096), .B(n15097), .Z(n15095) );
  XNOR U17143 ( .A(n15094), .B(n7549), .Z(n15097) );
  XNOR U17144 ( .A(n15090), .B(n15092), .Z(n7549) );
  NAND U17145 ( .A(n15098), .B(nreg[792]), .Z(n15092) );
  NAND U17146 ( .A(n12326), .B(nreg[792]), .Z(n15098) );
  XNOR U17147 ( .A(n15088), .B(n15099), .Z(n15090) );
  XOR U17148 ( .A(n15100), .B(n15101), .Z(n15088) );
  AND U17149 ( .A(n15102), .B(n15103), .Z(n15101) );
  XNOR U17150 ( .A(n15104), .B(n15100), .Z(n15103) );
  XOR U17151 ( .A(n15105), .B(nreg[792]), .Z(n15096) );
  IV U17152 ( .A(n15094), .Z(n15105) );
  XOR U17153 ( .A(n15106), .B(n15107), .Z(n15094) );
  AND U17154 ( .A(n15108), .B(n15109), .Z(n15107) );
  XNOR U17155 ( .A(n15106), .B(n7555), .Z(n15109) );
  XNOR U17156 ( .A(n15102), .B(n15104), .Z(n7555) );
  NAND U17157 ( .A(n15110), .B(nreg[791]), .Z(n15104) );
  NAND U17158 ( .A(n12326), .B(nreg[791]), .Z(n15110) );
  XNOR U17159 ( .A(n15100), .B(n15111), .Z(n15102) );
  XOR U17160 ( .A(n15112), .B(n15113), .Z(n15100) );
  AND U17161 ( .A(n15114), .B(n15115), .Z(n15113) );
  XNOR U17162 ( .A(n15116), .B(n15112), .Z(n15115) );
  XOR U17163 ( .A(n15117), .B(nreg[791]), .Z(n15108) );
  IV U17164 ( .A(n15106), .Z(n15117) );
  XOR U17165 ( .A(n15118), .B(n15119), .Z(n15106) );
  AND U17166 ( .A(n15120), .B(n15121), .Z(n15119) );
  XNOR U17167 ( .A(n15118), .B(n7561), .Z(n15121) );
  XNOR U17168 ( .A(n15114), .B(n15116), .Z(n7561) );
  NAND U17169 ( .A(n15122), .B(nreg[790]), .Z(n15116) );
  NAND U17170 ( .A(n12326), .B(nreg[790]), .Z(n15122) );
  XNOR U17171 ( .A(n15112), .B(n15123), .Z(n15114) );
  XOR U17172 ( .A(n15124), .B(n15125), .Z(n15112) );
  AND U17173 ( .A(n15126), .B(n15127), .Z(n15125) );
  XNOR U17174 ( .A(n15128), .B(n15124), .Z(n15127) );
  XOR U17175 ( .A(n15129), .B(nreg[790]), .Z(n15120) );
  IV U17176 ( .A(n15118), .Z(n15129) );
  XOR U17177 ( .A(n15130), .B(n15131), .Z(n15118) );
  AND U17178 ( .A(n15132), .B(n15133), .Z(n15131) );
  XNOR U17179 ( .A(n15130), .B(n7567), .Z(n15133) );
  XNOR U17180 ( .A(n15126), .B(n15128), .Z(n7567) );
  NAND U17181 ( .A(n15134), .B(nreg[789]), .Z(n15128) );
  NAND U17182 ( .A(n12326), .B(nreg[789]), .Z(n15134) );
  XNOR U17183 ( .A(n15124), .B(n15135), .Z(n15126) );
  XOR U17184 ( .A(n15136), .B(n15137), .Z(n15124) );
  AND U17185 ( .A(n15138), .B(n15139), .Z(n15137) );
  XNOR U17186 ( .A(n15140), .B(n15136), .Z(n15139) );
  XOR U17187 ( .A(n15141), .B(nreg[789]), .Z(n15132) );
  IV U17188 ( .A(n15130), .Z(n15141) );
  XOR U17189 ( .A(n15142), .B(n15143), .Z(n15130) );
  AND U17190 ( .A(n15144), .B(n15145), .Z(n15143) );
  XNOR U17191 ( .A(n15142), .B(n7573), .Z(n15145) );
  XNOR U17192 ( .A(n15138), .B(n15140), .Z(n7573) );
  NAND U17193 ( .A(n15146), .B(nreg[788]), .Z(n15140) );
  NAND U17194 ( .A(n12326), .B(nreg[788]), .Z(n15146) );
  XNOR U17195 ( .A(n15136), .B(n15147), .Z(n15138) );
  XOR U17196 ( .A(n15148), .B(n15149), .Z(n15136) );
  AND U17197 ( .A(n15150), .B(n15151), .Z(n15149) );
  XNOR U17198 ( .A(n15152), .B(n15148), .Z(n15151) );
  XOR U17199 ( .A(n15153), .B(nreg[788]), .Z(n15144) );
  IV U17200 ( .A(n15142), .Z(n15153) );
  XOR U17201 ( .A(n15154), .B(n15155), .Z(n15142) );
  AND U17202 ( .A(n15156), .B(n15157), .Z(n15155) );
  XNOR U17203 ( .A(n15154), .B(n7579), .Z(n15157) );
  XNOR U17204 ( .A(n15150), .B(n15152), .Z(n7579) );
  NAND U17205 ( .A(n15158), .B(nreg[787]), .Z(n15152) );
  NAND U17206 ( .A(n12326), .B(nreg[787]), .Z(n15158) );
  XNOR U17207 ( .A(n15148), .B(n15159), .Z(n15150) );
  XOR U17208 ( .A(n15160), .B(n15161), .Z(n15148) );
  AND U17209 ( .A(n15162), .B(n15163), .Z(n15161) );
  XNOR U17210 ( .A(n15164), .B(n15160), .Z(n15163) );
  XOR U17211 ( .A(n15165), .B(nreg[787]), .Z(n15156) );
  IV U17212 ( .A(n15154), .Z(n15165) );
  XOR U17213 ( .A(n15166), .B(n15167), .Z(n15154) );
  AND U17214 ( .A(n15168), .B(n15169), .Z(n15167) );
  XNOR U17215 ( .A(n15166), .B(n7585), .Z(n15169) );
  XNOR U17216 ( .A(n15162), .B(n15164), .Z(n7585) );
  NAND U17217 ( .A(n15170), .B(nreg[786]), .Z(n15164) );
  NAND U17218 ( .A(n12326), .B(nreg[786]), .Z(n15170) );
  XNOR U17219 ( .A(n15160), .B(n15171), .Z(n15162) );
  XOR U17220 ( .A(n15172), .B(n15173), .Z(n15160) );
  AND U17221 ( .A(n15174), .B(n15175), .Z(n15173) );
  XNOR U17222 ( .A(n15176), .B(n15172), .Z(n15175) );
  XOR U17223 ( .A(n15177), .B(nreg[786]), .Z(n15168) );
  IV U17224 ( .A(n15166), .Z(n15177) );
  XOR U17225 ( .A(n15178), .B(n15179), .Z(n15166) );
  AND U17226 ( .A(n15180), .B(n15181), .Z(n15179) );
  XNOR U17227 ( .A(n15178), .B(n7591), .Z(n15181) );
  XNOR U17228 ( .A(n15174), .B(n15176), .Z(n7591) );
  NAND U17229 ( .A(n15182), .B(nreg[785]), .Z(n15176) );
  NAND U17230 ( .A(n12326), .B(nreg[785]), .Z(n15182) );
  XNOR U17231 ( .A(n15172), .B(n15183), .Z(n15174) );
  XOR U17232 ( .A(n15184), .B(n15185), .Z(n15172) );
  AND U17233 ( .A(n15186), .B(n15187), .Z(n15185) );
  XNOR U17234 ( .A(n15188), .B(n15184), .Z(n15187) );
  XOR U17235 ( .A(n15189), .B(nreg[785]), .Z(n15180) );
  IV U17236 ( .A(n15178), .Z(n15189) );
  XOR U17237 ( .A(n15190), .B(n15191), .Z(n15178) );
  AND U17238 ( .A(n15192), .B(n15193), .Z(n15191) );
  XNOR U17239 ( .A(n15190), .B(n7597), .Z(n15193) );
  XNOR U17240 ( .A(n15186), .B(n15188), .Z(n7597) );
  NAND U17241 ( .A(n15194), .B(nreg[784]), .Z(n15188) );
  NAND U17242 ( .A(n12326), .B(nreg[784]), .Z(n15194) );
  XNOR U17243 ( .A(n15184), .B(n15195), .Z(n15186) );
  XOR U17244 ( .A(n15196), .B(n15197), .Z(n15184) );
  AND U17245 ( .A(n15198), .B(n15199), .Z(n15197) );
  XNOR U17246 ( .A(n15200), .B(n15196), .Z(n15199) );
  XOR U17247 ( .A(n15201), .B(nreg[784]), .Z(n15192) );
  IV U17248 ( .A(n15190), .Z(n15201) );
  XOR U17249 ( .A(n15202), .B(n15203), .Z(n15190) );
  AND U17250 ( .A(n15204), .B(n15205), .Z(n15203) );
  XNOR U17251 ( .A(n15202), .B(n7603), .Z(n15205) );
  XNOR U17252 ( .A(n15198), .B(n15200), .Z(n7603) );
  NAND U17253 ( .A(n15206), .B(nreg[783]), .Z(n15200) );
  NAND U17254 ( .A(n12326), .B(nreg[783]), .Z(n15206) );
  XNOR U17255 ( .A(n15196), .B(n15207), .Z(n15198) );
  XOR U17256 ( .A(n15208), .B(n15209), .Z(n15196) );
  AND U17257 ( .A(n15210), .B(n15211), .Z(n15209) );
  XNOR U17258 ( .A(n15212), .B(n15208), .Z(n15211) );
  XOR U17259 ( .A(n15213), .B(nreg[783]), .Z(n15204) );
  IV U17260 ( .A(n15202), .Z(n15213) );
  XOR U17261 ( .A(n15214), .B(n15215), .Z(n15202) );
  AND U17262 ( .A(n15216), .B(n15217), .Z(n15215) );
  XNOR U17263 ( .A(n15214), .B(n7609), .Z(n15217) );
  XNOR U17264 ( .A(n15210), .B(n15212), .Z(n7609) );
  NAND U17265 ( .A(n15218), .B(nreg[782]), .Z(n15212) );
  NAND U17266 ( .A(n12326), .B(nreg[782]), .Z(n15218) );
  XNOR U17267 ( .A(n15208), .B(n15219), .Z(n15210) );
  XOR U17268 ( .A(n15220), .B(n15221), .Z(n15208) );
  AND U17269 ( .A(n15222), .B(n15223), .Z(n15221) );
  XNOR U17270 ( .A(n15224), .B(n15220), .Z(n15223) );
  XOR U17271 ( .A(n15225), .B(nreg[782]), .Z(n15216) );
  IV U17272 ( .A(n15214), .Z(n15225) );
  XOR U17273 ( .A(n15226), .B(n15227), .Z(n15214) );
  AND U17274 ( .A(n15228), .B(n15229), .Z(n15227) );
  XNOR U17275 ( .A(n15226), .B(n7615), .Z(n15229) );
  XNOR U17276 ( .A(n15222), .B(n15224), .Z(n7615) );
  NAND U17277 ( .A(n15230), .B(nreg[781]), .Z(n15224) );
  NAND U17278 ( .A(n12326), .B(nreg[781]), .Z(n15230) );
  XNOR U17279 ( .A(n15220), .B(n15231), .Z(n15222) );
  XOR U17280 ( .A(n15232), .B(n15233), .Z(n15220) );
  AND U17281 ( .A(n15234), .B(n15235), .Z(n15233) );
  XNOR U17282 ( .A(n15236), .B(n15232), .Z(n15235) );
  XOR U17283 ( .A(n15237), .B(nreg[781]), .Z(n15228) );
  IV U17284 ( .A(n15226), .Z(n15237) );
  XOR U17285 ( .A(n15238), .B(n15239), .Z(n15226) );
  AND U17286 ( .A(n15240), .B(n15241), .Z(n15239) );
  XNOR U17287 ( .A(n15238), .B(n7621), .Z(n15241) );
  XNOR U17288 ( .A(n15234), .B(n15236), .Z(n7621) );
  NAND U17289 ( .A(n15242), .B(nreg[780]), .Z(n15236) );
  NAND U17290 ( .A(n12326), .B(nreg[780]), .Z(n15242) );
  XNOR U17291 ( .A(n15232), .B(n15243), .Z(n15234) );
  XOR U17292 ( .A(n15244), .B(n15245), .Z(n15232) );
  AND U17293 ( .A(n15246), .B(n15247), .Z(n15245) );
  XNOR U17294 ( .A(n15248), .B(n15244), .Z(n15247) );
  XOR U17295 ( .A(n15249), .B(nreg[780]), .Z(n15240) );
  IV U17296 ( .A(n15238), .Z(n15249) );
  XOR U17297 ( .A(n15250), .B(n15251), .Z(n15238) );
  AND U17298 ( .A(n15252), .B(n15253), .Z(n15251) );
  XNOR U17299 ( .A(n15250), .B(n7627), .Z(n15253) );
  XNOR U17300 ( .A(n15246), .B(n15248), .Z(n7627) );
  NAND U17301 ( .A(n15254), .B(nreg[779]), .Z(n15248) );
  NAND U17302 ( .A(n12326), .B(nreg[779]), .Z(n15254) );
  XNOR U17303 ( .A(n15244), .B(n15255), .Z(n15246) );
  XOR U17304 ( .A(n15256), .B(n15257), .Z(n15244) );
  AND U17305 ( .A(n15258), .B(n15259), .Z(n15257) );
  XNOR U17306 ( .A(n15260), .B(n15256), .Z(n15259) );
  XOR U17307 ( .A(n15261), .B(nreg[779]), .Z(n15252) );
  IV U17308 ( .A(n15250), .Z(n15261) );
  XOR U17309 ( .A(n15262), .B(n15263), .Z(n15250) );
  AND U17310 ( .A(n15264), .B(n15265), .Z(n15263) );
  XNOR U17311 ( .A(n15262), .B(n7633), .Z(n15265) );
  XNOR U17312 ( .A(n15258), .B(n15260), .Z(n7633) );
  NAND U17313 ( .A(n15266), .B(nreg[778]), .Z(n15260) );
  NAND U17314 ( .A(n12326), .B(nreg[778]), .Z(n15266) );
  XNOR U17315 ( .A(n15256), .B(n15267), .Z(n15258) );
  XOR U17316 ( .A(n15268), .B(n15269), .Z(n15256) );
  AND U17317 ( .A(n15270), .B(n15271), .Z(n15269) );
  XNOR U17318 ( .A(n15272), .B(n15268), .Z(n15271) );
  XOR U17319 ( .A(n15273), .B(nreg[778]), .Z(n15264) );
  IV U17320 ( .A(n15262), .Z(n15273) );
  XOR U17321 ( .A(n15274), .B(n15275), .Z(n15262) );
  AND U17322 ( .A(n15276), .B(n15277), .Z(n15275) );
  XNOR U17323 ( .A(n15274), .B(n7639), .Z(n15277) );
  XNOR U17324 ( .A(n15270), .B(n15272), .Z(n7639) );
  NAND U17325 ( .A(n15278), .B(nreg[777]), .Z(n15272) );
  NAND U17326 ( .A(n12326), .B(nreg[777]), .Z(n15278) );
  XNOR U17327 ( .A(n15268), .B(n15279), .Z(n15270) );
  XOR U17328 ( .A(n15280), .B(n15281), .Z(n15268) );
  AND U17329 ( .A(n15282), .B(n15283), .Z(n15281) );
  XNOR U17330 ( .A(n15284), .B(n15280), .Z(n15283) );
  XOR U17331 ( .A(n15285), .B(nreg[777]), .Z(n15276) );
  IV U17332 ( .A(n15274), .Z(n15285) );
  XOR U17333 ( .A(n15286), .B(n15287), .Z(n15274) );
  AND U17334 ( .A(n15288), .B(n15289), .Z(n15287) );
  XNOR U17335 ( .A(n15286), .B(n7645), .Z(n15289) );
  XNOR U17336 ( .A(n15282), .B(n15284), .Z(n7645) );
  NAND U17337 ( .A(n15290), .B(nreg[776]), .Z(n15284) );
  NAND U17338 ( .A(n12326), .B(nreg[776]), .Z(n15290) );
  XNOR U17339 ( .A(n15280), .B(n15291), .Z(n15282) );
  XOR U17340 ( .A(n15292), .B(n15293), .Z(n15280) );
  AND U17341 ( .A(n15294), .B(n15295), .Z(n15293) );
  XNOR U17342 ( .A(n15296), .B(n15292), .Z(n15295) );
  XOR U17343 ( .A(n15297), .B(nreg[776]), .Z(n15288) );
  IV U17344 ( .A(n15286), .Z(n15297) );
  XOR U17345 ( .A(n15298), .B(n15299), .Z(n15286) );
  AND U17346 ( .A(n15300), .B(n15301), .Z(n15299) );
  XNOR U17347 ( .A(n15298), .B(n7651), .Z(n15301) );
  XNOR U17348 ( .A(n15294), .B(n15296), .Z(n7651) );
  NAND U17349 ( .A(n15302), .B(nreg[775]), .Z(n15296) );
  NAND U17350 ( .A(n12326), .B(nreg[775]), .Z(n15302) );
  XNOR U17351 ( .A(n15292), .B(n15303), .Z(n15294) );
  XOR U17352 ( .A(n15304), .B(n15305), .Z(n15292) );
  AND U17353 ( .A(n15306), .B(n15307), .Z(n15305) );
  XNOR U17354 ( .A(n15308), .B(n15304), .Z(n15307) );
  XOR U17355 ( .A(n15309), .B(nreg[775]), .Z(n15300) );
  IV U17356 ( .A(n15298), .Z(n15309) );
  XOR U17357 ( .A(n15310), .B(n15311), .Z(n15298) );
  AND U17358 ( .A(n15312), .B(n15313), .Z(n15311) );
  XNOR U17359 ( .A(n15310), .B(n7657), .Z(n15313) );
  XNOR U17360 ( .A(n15306), .B(n15308), .Z(n7657) );
  NAND U17361 ( .A(n15314), .B(nreg[774]), .Z(n15308) );
  NAND U17362 ( .A(n12326), .B(nreg[774]), .Z(n15314) );
  XNOR U17363 ( .A(n15304), .B(n15315), .Z(n15306) );
  XOR U17364 ( .A(n15316), .B(n15317), .Z(n15304) );
  AND U17365 ( .A(n15318), .B(n15319), .Z(n15317) );
  XNOR U17366 ( .A(n15320), .B(n15316), .Z(n15319) );
  XOR U17367 ( .A(n15321), .B(nreg[774]), .Z(n15312) );
  IV U17368 ( .A(n15310), .Z(n15321) );
  XOR U17369 ( .A(n15322), .B(n15323), .Z(n15310) );
  AND U17370 ( .A(n15324), .B(n15325), .Z(n15323) );
  XNOR U17371 ( .A(n15322), .B(n7663), .Z(n15325) );
  XNOR U17372 ( .A(n15318), .B(n15320), .Z(n7663) );
  NAND U17373 ( .A(n15326), .B(nreg[773]), .Z(n15320) );
  NAND U17374 ( .A(n12326), .B(nreg[773]), .Z(n15326) );
  XNOR U17375 ( .A(n15316), .B(n15327), .Z(n15318) );
  XOR U17376 ( .A(n15328), .B(n15329), .Z(n15316) );
  AND U17377 ( .A(n15330), .B(n15331), .Z(n15329) );
  XNOR U17378 ( .A(n15332), .B(n15328), .Z(n15331) );
  XOR U17379 ( .A(n15333), .B(nreg[773]), .Z(n15324) );
  IV U17380 ( .A(n15322), .Z(n15333) );
  XOR U17381 ( .A(n15334), .B(n15335), .Z(n15322) );
  AND U17382 ( .A(n15336), .B(n15337), .Z(n15335) );
  XNOR U17383 ( .A(n15334), .B(n7669), .Z(n15337) );
  XNOR U17384 ( .A(n15330), .B(n15332), .Z(n7669) );
  NAND U17385 ( .A(n15338), .B(nreg[772]), .Z(n15332) );
  NAND U17386 ( .A(n12326), .B(nreg[772]), .Z(n15338) );
  XNOR U17387 ( .A(n15328), .B(n15339), .Z(n15330) );
  XOR U17388 ( .A(n15340), .B(n15341), .Z(n15328) );
  AND U17389 ( .A(n15342), .B(n15343), .Z(n15341) );
  XNOR U17390 ( .A(n15344), .B(n15340), .Z(n15343) );
  XOR U17391 ( .A(n15345), .B(nreg[772]), .Z(n15336) );
  IV U17392 ( .A(n15334), .Z(n15345) );
  XOR U17393 ( .A(n15346), .B(n15347), .Z(n15334) );
  AND U17394 ( .A(n15348), .B(n15349), .Z(n15347) );
  XNOR U17395 ( .A(n15346), .B(n7675), .Z(n15349) );
  XNOR U17396 ( .A(n15342), .B(n15344), .Z(n7675) );
  NAND U17397 ( .A(n15350), .B(nreg[771]), .Z(n15344) );
  NAND U17398 ( .A(n12326), .B(nreg[771]), .Z(n15350) );
  XNOR U17399 ( .A(n15340), .B(n15351), .Z(n15342) );
  XOR U17400 ( .A(n15352), .B(n15353), .Z(n15340) );
  AND U17401 ( .A(n15354), .B(n15355), .Z(n15353) );
  XNOR U17402 ( .A(n15356), .B(n15352), .Z(n15355) );
  XOR U17403 ( .A(n15357), .B(nreg[771]), .Z(n15348) );
  IV U17404 ( .A(n15346), .Z(n15357) );
  XOR U17405 ( .A(n15358), .B(n15359), .Z(n15346) );
  AND U17406 ( .A(n15360), .B(n15361), .Z(n15359) );
  XNOR U17407 ( .A(n15358), .B(n7681), .Z(n15361) );
  XNOR U17408 ( .A(n15354), .B(n15356), .Z(n7681) );
  NAND U17409 ( .A(n15362), .B(nreg[770]), .Z(n15356) );
  NAND U17410 ( .A(n12326), .B(nreg[770]), .Z(n15362) );
  XNOR U17411 ( .A(n15352), .B(n15363), .Z(n15354) );
  XOR U17412 ( .A(n15364), .B(n15365), .Z(n15352) );
  AND U17413 ( .A(n15366), .B(n15367), .Z(n15365) );
  XNOR U17414 ( .A(n15368), .B(n15364), .Z(n15367) );
  XOR U17415 ( .A(n15369), .B(nreg[770]), .Z(n15360) );
  IV U17416 ( .A(n15358), .Z(n15369) );
  XOR U17417 ( .A(n15370), .B(n15371), .Z(n15358) );
  AND U17418 ( .A(n15372), .B(n15373), .Z(n15371) );
  XNOR U17419 ( .A(n15370), .B(n7687), .Z(n15373) );
  XNOR U17420 ( .A(n15366), .B(n15368), .Z(n7687) );
  NAND U17421 ( .A(n15374), .B(nreg[769]), .Z(n15368) );
  NAND U17422 ( .A(n12326), .B(nreg[769]), .Z(n15374) );
  XNOR U17423 ( .A(n15364), .B(n15375), .Z(n15366) );
  XOR U17424 ( .A(n15376), .B(n15377), .Z(n15364) );
  AND U17425 ( .A(n15378), .B(n15379), .Z(n15377) );
  XNOR U17426 ( .A(n15380), .B(n15376), .Z(n15379) );
  XOR U17427 ( .A(n15381), .B(nreg[769]), .Z(n15372) );
  IV U17428 ( .A(n15370), .Z(n15381) );
  XOR U17429 ( .A(n15382), .B(n15383), .Z(n15370) );
  AND U17430 ( .A(n15384), .B(n15385), .Z(n15383) );
  XNOR U17431 ( .A(n15382), .B(n7693), .Z(n15385) );
  XNOR U17432 ( .A(n15378), .B(n15380), .Z(n7693) );
  NAND U17433 ( .A(n15386), .B(nreg[768]), .Z(n15380) );
  NAND U17434 ( .A(n12326), .B(nreg[768]), .Z(n15386) );
  XNOR U17435 ( .A(n15376), .B(n15387), .Z(n15378) );
  XOR U17436 ( .A(n15388), .B(n15389), .Z(n15376) );
  AND U17437 ( .A(n15390), .B(n15391), .Z(n15389) );
  XNOR U17438 ( .A(n15392), .B(n15388), .Z(n15391) );
  XOR U17439 ( .A(n15393), .B(nreg[768]), .Z(n15384) );
  IV U17440 ( .A(n15382), .Z(n15393) );
  XOR U17441 ( .A(n15394), .B(n15395), .Z(n15382) );
  AND U17442 ( .A(n15396), .B(n15397), .Z(n15395) );
  XNOR U17443 ( .A(n15394), .B(n7699), .Z(n15397) );
  XNOR U17444 ( .A(n15390), .B(n15392), .Z(n7699) );
  NAND U17445 ( .A(n15398), .B(nreg[767]), .Z(n15392) );
  NAND U17446 ( .A(n12326), .B(nreg[767]), .Z(n15398) );
  XNOR U17447 ( .A(n15388), .B(n15399), .Z(n15390) );
  XOR U17448 ( .A(n15400), .B(n15401), .Z(n15388) );
  AND U17449 ( .A(n15402), .B(n15403), .Z(n15401) );
  XNOR U17450 ( .A(n15404), .B(n15400), .Z(n15403) );
  XOR U17451 ( .A(n15405), .B(nreg[767]), .Z(n15396) );
  IV U17452 ( .A(n15394), .Z(n15405) );
  XOR U17453 ( .A(n15406), .B(n15407), .Z(n15394) );
  AND U17454 ( .A(n15408), .B(n15409), .Z(n15407) );
  XNOR U17455 ( .A(n15406), .B(n7705), .Z(n15409) );
  XNOR U17456 ( .A(n15402), .B(n15404), .Z(n7705) );
  NAND U17457 ( .A(n15410), .B(nreg[766]), .Z(n15404) );
  NAND U17458 ( .A(n12326), .B(nreg[766]), .Z(n15410) );
  XNOR U17459 ( .A(n15400), .B(n15411), .Z(n15402) );
  XOR U17460 ( .A(n15412), .B(n15413), .Z(n15400) );
  AND U17461 ( .A(n15414), .B(n15415), .Z(n15413) );
  XNOR U17462 ( .A(n15416), .B(n15412), .Z(n15415) );
  XOR U17463 ( .A(n15417), .B(nreg[766]), .Z(n15408) );
  IV U17464 ( .A(n15406), .Z(n15417) );
  XOR U17465 ( .A(n15418), .B(n15419), .Z(n15406) );
  AND U17466 ( .A(n15420), .B(n15421), .Z(n15419) );
  XNOR U17467 ( .A(n15418), .B(n7711), .Z(n15421) );
  XNOR U17468 ( .A(n15414), .B(n15416), .Z(n7711) );
  NAND U17469 ( .A(n15422), .B(nreg[765]), .Z(n15416) );
  NAND U17470 ( .A(n12326), .B(nreg[765]), .Z(n15422) );
  XNOR U17471 ( .A(n15412), .B(n15423), .Z(n15414) );
  XOR U17472 ( .A(n15424), .B(n15425), .Z(n15412) );
  AND U17473 ( .A(n15426), .B(n15427), .Z(n15425) );
  XNOR U17474 ( .A(n15428), .B(n15424), .Z(n15427) );
  XOR U17475 ( .A(n15429), .B(nreg[765]), .Z(n15420) );
  IV U17476 ( .A(n15418), .Z(n15429) );
  XOR U17477 ( .A(n15430), .B(n15431), .Z(n15418) );
  AND U17478 ( .A(n15432), .B(n15433), .Z(n15431) );
  XNOR U17479 ( .A(n15430), .B(n7717), .Z(n15433) );
  XNOR U17480 ( .A(n15426), .B(n15428), .Z(n7717) );
  NAND U17481 ( .A(n15434), .B(nreg[764]), .Z(n15428) );
  NAND U17482 ( .A(n12326), .B(nreg[764]), .Z(n15434) );
  XNOR U17483 ( .A(n15424), .B(n15435), .Z(n15426) );
  XOR U17484 ( .A(n15436), .B(n15437), .Z(n15424) );
  AND U17485 ( .A(n15438), .B(n15439), .Z(n15437) );
  XNOR U17486 ( .A(n15440), .B(n15436), .Z(n15439) );
  XOR U17487 ( .A(n15441), .B(nreg[764]), .Z(n15432) );
  IV U17488 ( .A(n15430), .Z(n15441) );
  XOR U17489 ( .A(n15442), .B(n15443), .Z(n15430) );
  AND U17490 ( .A(n15444), .B(n15445), .Z(n15443) );
  XNOR U17491 ( .A(n15442), .B(n7723), .Z(n15445) );
  XNOR U17492 ( .A(n15438), .B(n15440), .Z(n7723) );
  NAND U17493 ( .A(n15446), .B(nreg[763]), .Z(n15440) );
  NAND U17494 ( .A(n12326), .B(nreg[763]), .Z(n15446) );
  XNOR U17495 ( .A(n15436), .B(n15447), .Z(n15438) );
  XOR U17496 ( .A(n15448), .B(n15449), .Z(n15436) );
  AND U17497 ( .A(n15450), .B(n15451), .Z(n15449) );
  XNOR U17498 ( .A(n15452), .B(n15448), .Z(n15451) );
  XOR U17499 ( .A(n15453), .B(nreg[763]), .Z(n15444) );
  IV U17500 ( .A(n15442), .Z(n15453) );
  XOR U17501 ( .A(n15454), .B(n15455), .Z(n15442) );
  AND U17502 ( .A(n15456), .B(n15457), .Z(n15455) );
  XNOR U17503 ( .A(n15454), .B(n7729), .Z(n15457) );
  XNOR U17504 ( .A(n15450), .B(n15452), .Z(n7729) );
  NAND U17505 ( .A(n15458), .B(nreg[762]), .Z(n15452) );
  NAND U17506 ( .A(n12326), .B(nreg[762]), .Z(n15458) );
  XNOR U17507 ( .A(n15448), .B(n15459), .Z(n15450) );
  XOR U17508 ( .A(n15460), .B(n15461), .Z(n15448) );
  AND U17509 ( .A(n15462), .B(n15463), .Z(n15461) );
  XNOR U17510 ( .A(n15464), .B(n15460), .Z(n15463) );
  XOR U17511 ( .A(n15465), .B(nreg[762]), .Z(n15456) );
  IV U17512 ( .A(n15454), .Z(n15465) );
  XOR U17513 ( .A(n15466), .B(n15467), .Z(n15454) );
  AND U17514 ( .A(n15468), .B(n15469), .Z(n15467) );
  XNOR U17515 ( .A(n15466), .B(n7735), .Z(n15469) );
  XNOR U17516 ( .A(n15462), .B(n15464), .Z(n7735) );
  NAND U17517 ( .A(n15470), .B(nreg[761]), .Z(n15464) );
  NAND U17518 ( .A(n12326), .B(nreg[761]), .Z(n15470) );
  XNOR U17519 ( .A(n15460), .B(n15471), .Z(n15462) );
  XOR U17520 ( .A(n15472), .B(n15473), .Z(n15460) );
  AND U17521 ( .A(n15474), .B(n15475), .Z(n15473) );
  XNOR U17522 ( .A(n15476), .B(n15472), .Z(n15475) );
  XOR U17523 ( .A(n15477), .B(nreg[761]), .Z(n15468) );
  IV U17524 ( .A(n15466), .Z(n15477) );
  XOR U17525 ( .A(n15478), .B(n15479), .Z(n15466) );
  AND U17526 ( .A(n15480), .B(n15481), .Z(n15479) );
  XNOR U17527 ( .A(n15478), .B(n7741), .Z(n15481) );
  XNOR U17528 ( .A(n15474), .B(n15476), .Z(n7741) );
  NAND U17529 ( .A(n15482), .B(nreg[760]), .Z(n15476) );
  NAND U17530 ( .A(n12326), .B(nreg[760]), .Z(n15482) );
  XNOR U17531 ( .A(n15472), .B(n15483), .Z(n15474) );
  XOR U17532 ( .A(n15484), .B(n15485), .Z(n15472) );
  AND U17533 ( .A(n15486), .B(n15487), .Z(n15485) );
  XNOR U17534 ( .A(n15488), .B(n15484), .Z(n15487) );
  XOR U17535 ( .A(n15489), .B(nreg[760]), .Z(n15480) );
  IV U17536 ( .A(n15478), .Z(n15489) );
  XOR U17537 ( .A(n15490), .B(n15491), .Z(n15478) );
  AND U17538 ( .A(n15492), .B(n15493), .Z(n15491) );
  XNOR U17539 ( .A(n15490), .B(n7747), .Z(n15493) );
  XNOR U17540 ( .A(n15486), .B(n15488), .Z(n7747) );
  NAND U17541 ( .A(n15494), .B(nreg[759]), .Z(n15488) );
  NAND U17542 ( .A(n12326), .B(nreg[759]), .Z(n15494) );
  XNOR U17543 ( .A(n15484), .B(n15495), .Z(n15486) );
  XOR U17544 ( .A(n15496), .B(n15497), .Z(n15484) );
  AND U17545 ( .A(n15498), .B(n15499), .Z(n15497) );
  XNOR U17546 ( .A(n15500), .B(n15496), .Z(n15499) );
  XOR U17547 ( .A(n15501), .B(nreg[759]), .Z(n15492) );
  IV U17548 ( .A(n15490), .Z(n15501) );
  XOR U17549 ( .A(n15502), .B(n15503), .Z(n15490) );
  AND U17550 ( .A(n15504), .B(n15505), .Z(n15503) );
  XNOR U17551 ( .A(n15502), .B(n7753), .Z(n15505) );
  XNOR U17552 ( .A(n15498), .B(n15500), .Z(n7753) );
  NAND U17553 ( .A(n15506), .B(nreg[758]), .Z(n15500) );
  NAND U17554 ( .A(n12326), .B(nreg[758]), .Z(n15506) );
  XNOR U17555 ( .A(n15496), .B(n15507), .Z(n15498) );
  XOR U17556 ( .A(n15508), .B(n15509), .Z(n15496) );
  AND U17557 ( .A(n15510), .B(n15511), .Z(n15509) );
  XNOR U17558 ( .A(n15512), .B(n15508), .Z(n15511) );
  XOR U17559 ( .A(n15513), .B(nreg[758]), .Z(n15504) );
  IV U17560 ( .A(n15502), .Z(n15513) );
  XOR U17561 ( .A(n15514), .B(n15515), .Z(n15502) );
  AND U17562 ( .A(n15516), .B(n15517), .Z(n15515) );
  XNOR U17563 ( .A(n15514), .B(n7759), .Z(n15517) );
  XNOR U17564 ( .A(n15510), .B(n15512), .Z(n7759) );
  NAND U17565 ( .A(n15518), .B(nreg[757]), .Z(n15512) );
  NAND U17566 ( .A(n12326), .B(nreg[757]), .Z(n15518) );
  XNOR U17567 ( .A(n15508), .B(n15519), .Z(n15510) );
  XOR U17568 ( .A(n15520), .B(n15521), .Z(n15508) );
  AND U17569 ( .A(n15522), .B(n15523), .Z(n15521) );
  XNOR U17570 ( .A(n15524), .B(n15520), .Z(n15523) );
  XOR U17571 ( .A(n15525), .B(nreg[757]), .Z(n15516) );
  IV U17572 ( .A(n15514), .Z(n15525) );
  XOR U17573 ( .A(n15526), .B(n15527), .Z(n15514) );
  AND U17574 ( .A(n15528), .B(n15529), .Z(n15527) );
  XNOR U17575 ( .A(n15526), .B(n7765), .Z(n15529) );
  XNOR U17576 ( .A(n15522), .B(n15524), .Z(n7765) );
  NAND U17577 ( .A(n15530), .B(nreg[756]), .Z(n15524) );
  NAND U17578 ( .A(n12326), .B(nreg[756]), .Z(n15530) );
  XNOR U17579 ( .A(n15520), .B(n15531), .Z(n15522) );
  XOR U17580 ( .A(n15532), .B(n15533), .Z(n15520) );
  AND U17581 ( .A(n15534), .B(n15535), .Z(n15533) );
  XNOR U17582 ( .A(n15536), .B(n15532), .Z(n15535) );
  XOR U17583 ( .A(n15537), .B(nreg[756]), .Z(n15528) );
  IV U17584 ( .A(n15526), .Z(n15537) );
  XOR U17585 ( .A(n15538), .B(n15539), .Z(n15526) );
  AND U17586 ( .A(n15540), .B(n15541), .Z(n15539) );
  XNOR U17587 ( .A(n15538), .B(n7771), .Z(n15541) );
  XNOR U17588 ( .A(n15534), .B(n15536), .Z(n7771) );
  NAND U17589 ( .A(n15542), .B(nreg[755]), .Z(n15536) );
  NAND U17590 ( .A(n12326), .B(nreg[755]), .Z(n15542) );
  XNOR U17591 ( .A(n15532), .B(n15543), .Z(n15534) );
  XOR U17592 ( .A(n15544), .B(n15545), .Z(n15532) );
  AND U17593 ( .A(n15546), .B(n15547), .Z(n15545) );
  XNOR U17594 ( .A(n15548), .B(n15544), .Z(n15547) );
  XOR U17595 ( .A(n15549), .B(nreg[755]), .Z(n15540) );
  IV U17596 ( .A(n15538), .Z(n15549) );
  XOR U17597 ( .A(n15550), .B(n15551), .Z(n15538) );
  AND U17598 ( .A(n15552), .B(n15553), .Z(n15551) );
  XNOR U17599 ( .A(n15550), .B(n7777), .Z(n15553) );
  XNOR U17600 ( .A(n15546), .B(n15548), .Z(n7777) );
  NAND U17601 ( .A(n15554), .B(nreg[754]), .Z(n15548) );
  NAND U17602 ( .A(n12326), .B(nreg[754]), .Z(n15554) );
  XNOR U17603 ( .A(n15544), .B(n15555), .Z(n15546) );
  XOR U17604 ( .A(n15556), .B(n15557), .Z(n15544) );
  AND U17605 ( .A(n15558), .B(n15559), .Z(n15557) );
  XNOR U17606 ( .A(n15560), .B(n15556), .Z(n15559) );
  XOR U17607 ( .A(n15561), .B(nreg[754]), .Z(n15552) );
  IV U17608 ( .A(n15550), .Z(n15561) );
  XOR U17609 ( .A(n15562), .B(n15563), .Z(n15550) );
  AND U17610 ( .A(n15564), .B(n15565), .Z(n15563) );
  XNOR U17611 ( .A(n15562), .B(n7783), .Z(n15565) );
  XNOR U17612 ( .A(n15558), .B(n15560), .Z(n7783) );
  NAND U17613 ( .A(n15566), .B(nreg[753]), .Z(n15560) );
  NAND U17614 ( .A(n12326), .B(nreg[753]), .Z(n15566) );
  XNOR U17615 ( .A(n15556), .B(n15567), .Z(n15558) );
  XOR U17616 ( .A(n15568), .B(n15569), .Z(n15556) );
  AND U17617 ( .A(n15570), .B(n15571), .Z(n15569) );
  XNOR U17618 ( .A(n15572), .B(n15568), .Z(n15571) );
  XOR U17619 ( .A(n15573), .B(nreg[753]), .Z(n15564) );
  IV U17620 ( .A(n15562), .Z(n15573) );
  XOR U17621 ( .A(n15574), .B(n15575), .Z(n15562) );
  AND U17622 ( .A(n15576), .B(n15577), .Z(n15575) );
  XNOR U17623 ( .A(n15574), .B(n7789), .Z(n15577) );
  XNOR U17624 ( .A(n15570), .B(n15572), .Z(n7789) );
  NAND U17625 ( .A(n15578), .B(nreg[752]), .Z(n15572) );
  NAND U17626 ( .A(n12326), .B(nreg[752]), .Z(n15578) );
  XNOR U17627 ( .A(n15568), .B(n15579), .Z(n15570) );
  XOR U17628 ( .A(n15580), .B(n15581), .Z(n15568) );
  AND U17629 ( .A(n15582), .B(n15583), .Z(n15581) );
  XNOR U17630 ( .A(n15584), .B(n15580), .Z(n15583) );
  XOR U17631 ( .A(n15585), .B(nreg[752]), .Z(n15576) );
  IV U17632 ( .A(n15574), .Z(n15585) );
  XOR U17633 ( .A(n15586), .B(n15587), .Z(n15574) );
  AND U17634 ( .A(n15588), .B(n15589), .Z(n15587) );
  XNOR U17635 ( .A(n15586), .B(n7795), .Z(n15589) );
  XNOR U17636 ( .A(n15582), .B(n15584), .Z(n7795) );
  NAND U17637 ( .A(n15590), .B(nreg[751]), .Z(n15584) );
  NAND U17638 ( .A(n12326), .B(nreg[751]), .Z(n15590) );
  XNOR U17639 ( .A(n15580), .B(n15591), .Z(n15582) );
  XOR U17640 ( .A(n15592), .B(n15593), .Z(n15580) );
  AND U17641 ( .A(n15594), .B(n15595), .Z(n15593) );
  XNOR U17642 ( .A(n15596), .B(n15592), .Z(n15595) );
  XOR U17643 ( .A(n15597), .B(nreg[751]), .Z(n15588) );
  IV U17644 ( .A(n15586), .Z(n15597) );
  XOR U17645 ( .A(n15598), .B(n15599), .Z(n15586) );
  AND U17646 ( .A(n15600), .B(n15601), .Z(n15599) );
  XNOR U17647 ( .A(n15598), .B(n7801), .Z(n15601) );
  XNOR U17648 ( .A(n15594), .B(n15596), .Z(n7801) );
  NAND U17649 ( .A(n15602), .B(nreg[750]), .Z(n15596) );
  NAND U17650 ( .A(n12326), .B(nreg[750]), .Z(n15602) );
  XNOR U17651 ( .A(n15592), .B(n15603), .Z(n15594) );
  XOR U17652 ( .A(n15604), .B(n15605), .Z(n15592) );
  AND U17653 ( .A(n15606), .B(n15607), .Z(n15605) );
  XNOR U17654 ( .A(n15608), .B(n15604), .Z(n15607) );
  XOR U17655 ( .A(n15609), .B(nreg[750]), .Z(n15600) );
  IV U17656 ( .A(n15598), .Z(n15609) );
  XOR U17657 ( .A(n15610), .B(n15611), .Z(n15598) );
  AND U17658 ( .A(n15612), .B(n15613), .Z(n15611) );
  XNOR U17659 ( .A(n15610), .B(n7807), .Z(n15613) );
  XNOR U17660 ( .A(n15606), .B(n15608), .Z(n7807) );
  NAND U17661 ( .A(n15614), .B(nreg[749]), .Z(n15608) );
  NAND U17662 ( .A(n12326), .B(nreg[749]), .Z(n15614) );
  XNOR U17663 ( .A(n15604), .B(n15615), .Z(n15606) );
  XOR U17664 ( .A(n15616), .B(n15617), .Z(n15604) );
  AND U17665 ( .A(n15618), .B(n15619), .Z(n15617) );
  XNOR U17666 ( .A(n15620), .B(n15616), .Z(n15619) );
  XOR U17667 ( .A(n15621), .B(nreg[749]), .Z(n15612) );
  IV U17668 ( .A(n15610), .Z(n15621) );
  XOR U17669 ( .A(n15622), .B(n15623), .Z(n15610) );
  AND U17670 ( .A(n15624), .B(n15625), .Z(n15623) );
  XNOR U17671 ( .A(n15622), .B(n7813), .Z(n15625) );
  XNOR U17672 ( .A(n15618), .B(n15620), .Z(n7813) );
  NAND U17673 ( .A(n15626), .B(nreg[748]), .Z(n15620) );
  NAND U17674 ( .A(n12326), .B(nreg[748]), .Z(n15626) );
  XNOR U17675 ( .A(n15616), .B(n15627), .Z(n15618) );
  XOR U17676 ( .A(n15628), .B(n15629), .Z(n15616) );
  AND U17677 ( .A(n15630), .B(n15631), .Z(n15629) );
  XNOR U17678 ( .A(n15632), .B(n15628), .Z(n15631) );
  XOR U17679 ( .A(n15633), .B(nreg[748]), .Z(n15624) );
  IV U17680 ( .A(n15622), .Z(n15633) );
  XOR U17681 ( .A(n15634), .B(n15635), .Z(n15622) );
  AND U17682 ( .A(n15636), .B(n15637), .Z(n15635) );
  XNOR U17683 ( .A(n15634), .B(n7819), .Z(n15637) );
  XNOR U17684 ( .A(n15630), .B(n15632), .Z(n7819) );
  NAND U17685 ( .A(n15638), .B(nreg[747]), .Z(n15632) );
  NAND U17686 ( .A(n12326), .B(nreg[747]), .Z(n15638) );
  XNOR U17687 ( .A(n15628), .B(n15639), .Z(n15630) );
  XOR U17688 ( .A(n15640), .B(n15641), .Z(n15628) );
  AND U17689 ( .A(n15642), .B(n15643), .Z(n15641) );
  XNOR U17690 ( .A(n15644), .B(n15640), .Z(n15643) );
  XOR U17691 ( .A(n15645), .B(nreg[747]), .Z(n15636) );
  IV U17692 ( .A(n15634), .Z(n15645) );
  XOR U17693 ( .A(n15646), .B(n15647), .Z(n15634) );
  AND U17694 ( .A(n15648), .B(n15649), .Z(n15647) );
  XNOR U17695 ( .A(n15646), .B(n7825), .Z(n15649) );
  XNOR U17696 ( .A(n15642), .B(n15644), .Z(n7825) );
  NAND U17697 ( .A(n15650), .B(nreg[746]), .Z(n15644) );
  NAND U17698 ( .A(n12326), .B(nreg[746]), .Z(n15650) );
  XNOR U17699 ( .A(n15640), .B(n15651), .Z(n15642) );
  XOR U17700 ( .A(n15652), .B(n15653), .Z(n15640) );
  AND U17701 ( .A(n15654), .B(n15655), .Z(n15653) );
  XNOR U17702 ( .A(n15656), .B(n15652), .Z(n15655) );
  XOR U17703 ( .A(n15657), .B(nreg[746]), .Z(n15648) );
  IV U17704 ( .A(n15646), .Z(n15657) );
  XOR U17705 ( .A(n15658), .B(n15659), .Z(n15646) );
  AND U17706 ( .A(n15660), .B(n15661), .Z(n15659) );
  XNOR U17707 ( .A(n15658), .B(n7831), .Z(n15661) );
  XNOR U17708 ( .A(n15654), .B(n15656), .Z(n7831) );
  NAND U17709 ( .A(n15662), .B(nreg[745]), .Z(n15656) );
  NAND U17710 ( .A(n12326), .B(nreg[745]), .Z(n15662) );
  XNOR U17711 ( .A(n15652), .B(n15663), .Z(n15654) );
  XOR U17712 ( .A(n15664), .B(n15665), .Z(n15652) );
  AND U17713 ( .A(n15666), .B(n15667), .Z(n15665) );
  XNOR U17714 ( .A(n15668), .B(n15664), .Z(n15667) );
  XOR U17715 ( .A(n15669), .B(nreg[745]), .Z(n15660) );
  IV U17716 ( .A(n15658), .Z(n15669) );
  XOR U17717 ( .A(n15670), .B(n15671), .Z(n15658) );
  AND U17718 ( .A(n15672), .B(n15673), .Z(n15671) );
  XNOR U17719 ( .A(n15670), .B(n7837), .Z(n15673) );
  XNOR U17720 ( .A(n15666), .B(n15668), .Z(n7837) );
  NAND U17721 ( .A(n15674), .B(nreg[744]), .Z(n15668) );
  NAND U17722 ( .A(n12326), .B(nreg[744]), .Z(n15674) );
  XNOR U17723 ( .A(n15664), .B(n15675), .Z(n15666) );
  XOR U17724 ( .A(n15676), .B(n15677), .Z(n15664) );
  AND U17725 ( .A(n15678), .B(n15679), .Z(n15677) );
  XNOR U17726 ( .A(n15680), .B(n15676), .Z(n15679) );
  XOR U17727 ( .A(n15681), .B(nreg[744]), .Z(n15672) );
  IV U17728 ( .A(n15670), .Z(n15681) );
  XOR U17729 ( .A(n15682), .B(n15683), .Z(n15670) );
  AND U17730 ( .A(n15684), .B(n15685), .Z(n15683) );
  XNOR U17731 ( .A(n15682), .B(n7843), .Z(n15685) );
  XNOR U17732 ( .A(n15678), .B(n15680), .Z(n7843) );
  NAND U17733 ( .A(n15686), .B(nreg[743]), .Z(n15680) );
  NAND U17734 ( .A(n12326), .B(nreg[743]), .Z(n15686) );
  XNOR U17735 ( .A(n15676), .B(n15687), .Z(n15678) );
  XOR U17736 ( .A(n15688), .B(n15689), .Z(n15676) );
  AND U17737 ( .A(n15690), .B(n15691), .Z(n15689) );
  XNOR U17738 ( .A(n15692), .B(n15688), .Z(n15691) );
  XOR U17739 ( .A(n15693), .B(nreg[743]), .Z(n15684) );
  IV U17740 ( .A(n15682), .Z(n15693) );
  XOR U17741 ( .A(n15694), .B(n15695), .Z(n15682) );
  AND U17742 ( .A(n15696), .B(n15697), .Z(n15695) );
  XNOR U17743 ( .A(n15694), .B(n7849), .Z(n15697) );
  XNOR U17744 ( .A(n15690), .B(n15692), .Z(n7849) );
  NAND U17745 ( .A(n15698), .B(nreg[742]), .Z(n15692) );
  NAND U17746 ( .A(n12326), .B(nreg[742]), .Z(n15698) );
  XNOR U17747 ( .A(n15688), .B(n15699), .Z(n15690) );
  XOR U17748 ( .A(n15700), .B(n15701), .Z(n15688) );
  AND U17749 ( .A(n15702), .B(n15703), .Z(n15701) );
  XNOR U17750 ( .A(n15704), .B(n15700), .Z(n15703) );
  XOR U17751 ( .A(n15705), .B(nreg[742]), .Z(n15696) );
  IV U17752 ( .A(n15694), .Z(n15705) );
  XOR U17753 ( .A(n15706), .B(n15707), .Z(n15694) );
  AND U17754 ( .A(n15708), .B(n15709), .Z(n15707) );
  XNOR U17755 ( .A(n15706), .B(n7855), .Z(n15709) );
  XNOR U17756 ( .A(n15702), .B(n15704), .Z(n7855) );
  NAND U17757 ( .A(n15710), .B(nreg[741]), .Z(n15704) );
  NAND U17758 ( .A(n12326), .B(nreg[741]), .Z(n15710) );
  XNOR U17759 ( .A(n15700), .B(n15711), .Z(n15702) );
  XOR U17760 ( .A(n15712), .B(n15713), .Z(n15700) );
  AND U17761 ( .A(n15714), .B(n15715), .Z(n15713) );
  XNOR U17762 ( .A(n15716), .B(n15712), .Z(n15715) );
  XOR U17763 ( .A(n15717), .B(nreg[741]), .Z(n15708) );
  IV U17764 ( .A(n15706), .Z(n15717) );
  XOR U17765 ( .A(n15718), .B(n15719), .Z(n15706) );
  AND U17766 ( .A(n15720), .B(n15721), .Z(n15719) );
  XNOR U17767 ( .A(n15718), .B(n7861), .Z(n15721) );
  XNOR U17768 ( .A(n15714), .B(n15716), .Z(n7861) );
  NAND U17769 ( .A(n15722), .B(nreg[740]), .Z(n15716) );
  NAND U17770 ( .A(n12326), .B(nreg[740]), .Z(n15722) );
  XNOR U17771 ( .A(n15712), .B(n15723), .Z(n15714) );
  XOR U17772 ( .A(n15724), .B(n15725), .Z(n15712) );
  AND U17773 ( .A(n15726), .B(n15727), .Z(n15725) );
  XNOR U17774 ( .A(n15728), .B(n15724), .Z(n15727) );
  XOR U17775 ( .A(n15729), .B(nreg[740]), .Z(n15720) );
  IV U17776 ( .A(n15718), .Z(n15729) );
  XOR U17777 ( .A(n15730), .B(n15731), .Z(n15718) );
  AND U17778 ( .A(n15732), .B(n15733), .Z(n15731) );
  XNOR U17779 ( .A(n15730), .B(n7867), .Z(n15733) );
  XNOR U17780 ( .A(n15726), .B(n15728), .Z(n7867) );
  NAND U17781 ( .A(n15734), .B(nreg[739]), .Z(n15728) );
  NAND U17782 ( .A(n12326), .B(nreg[739]), .Z(n15734) );
  XNOR U17783 ( .A(n15724), .B(n15735), .Z(n15726) );
  XOR U17784 ( .A(n15736), .B(n15737), .Z(n15724) );
  AND U17785 ( .A(n15738), .B(n15739), .Z(n15737) );
  XNOR U17786 ( .A(n15740), .B(n15736), .Z(n15739) );
  XOR U17787 ( .A(n15741), .B(nreg[739]), .Z(n15732) );
  IV U17788 ( .A(n15730), .Z(n15741) );
  XOR U17789 ( .A(n15742), .B(n15743), .Z(n15730) );
  AND U17790 ( .A(n15744), .B(n15745), .Z(n15743) );
  XNOR U17791 ( .A(n15742), .B(n7873), .Z(n15745) );
  XNOR U17792 ( .A(n15738), .B(n15740), .Z(n7873) );
  NAND U17793 ( .A(n15746), .B(nreg[738]), .Z(n15740) );
  NAND U17794 ( .A(n12326), .B(nreg[738]), .Z(n15746) );
  XNOR U17795 ( .A(n15736), .B(n15747), .Z(n15738) );
  XOR U17796 ( .A(n15748), .B(n15749), .Z(n15736) );
  AND U17797 ( .A(n15750), .B(n15751), .Z(n15749) );
  XNOR U17798 ( .A(n15752), .B(n15748), .Z(n15751) );
  XOR U17799 ( .A(n15753), .B(nreg[738]), .Z(n15744) );
  IV U17800 ( .A(n15742), .Z(n15753) );
  XOR U17801 ( .A(n15754), .B(n15755), .Z(n15742) );
  AND U17802 ( .A(n15756), .B(n15757), .Z(n15755) );
  XNOR U17803 ( .A(n15754), .B(n7879), .Z(n15757) );
  XNOR U17804 ( .A(n15750), .B(n15752), .Z(n7879) );
  NAND U17805 ( .A(n15758), .B(nreg[737]), .Z(n15752) );
  NAND U17806 ( .A(n12326), .B(nreg[737]), .Z(n15758) );
  XNOR U17807 ( .A(n15748), .B(n15759), .Z(n15750) );
  XOR U17808 ( .A(n15760), .B(n15761), .Z(n15748) );
  AND U17809 ( .A(n15762), .B(n15763), .Z(n15761) );
  XNOR U17810 ( .A(n15764), .B(n15760), .Z(n15763) );
  XOR U17811 ( .A(n15765), .B(nreg[737]), .Z(n15756) );
  IV U17812 ( .A(n15754), .Z(n15765) );
  XOR U17813 ( .A(n15766), .B(n15767), .Z(n15754) );
  AND U17814 ( .A(n15768), .B(n15769), .Z(n15767) );
  XNOR U17815 ( .A(n15766), .B(n7885), .Z(n15769) );
  XNOR U17816 ( .A(n15762), .B(n15764), .Z(n7885) );
  NAND U17817 ( .A(n15770), .B(nreg[736]), .Z(n15764) );
  NAND U17818 ( .A(n12326), .B(nreg[736]), .Z(n15770) );
  XNOR U17819 ( .A(n15760), .B(n15771), .Z(n15762) );
  XOR U17820 ( .A(n15772), .B(n15773), .Z(n15760) );
  AND U17821 ( .A(n15774), .B(n15775), .Z(n15773) );
  XNOR U17822 ( .A(n15776), .B(n15772), .Z(n15775) );
  XOR U17823 ( .A(n15777), .B(nreg[736]), .Z(n15768) );
  IV U17824 ( .A(n15766), .Z(n15777) );
  XOR U17825 ( .A(n15778), .B(n15779), .Z(n15766) );
  AND U17826 ( .A(n15780), .B(n15781), .Z(n15779) );
  XNOR U17827 ( .A(n15778), .B(n7891), .Z(n15781) );
  XNOR U17828 ( .A(n15774), .B(n15776), .Z(n7891) );
  NAND U17829 ( .A(n15782), .B(nreg[735]), .Z(n15776) );
  NAND U17830 ( .A(n12326), .B(nreg[735]), .Z(n15782) );
  XNOR U17831 ( .A(n15772), .B(n15783), .Z(n15774) );
  XOR U17832 ( .A(n15784), .B(n15785), .Z(n15772) );
  AND U17833 ( .A(n15786), .B(n15787), .Z(n15785) );
  XNOR U17834 ( .A(n15788), .B(n15784), .Z(n15787) );
  XOR U17835 ( .A(n15789), .B(nreg[735]), .Z(n15780) );
  IV U17836 ( .A(n15778), .Z(n15789) );
  XOR U17837 ( .A(n15790), .B(n15791), .Z(n15778) );
  AND U17838 ( .A(n15792), .B(n15793), .Z(n15791) );
  XNOR U17839 ( .A(n15790), .B(n7897), .Z(n15793) );
  XNOR U17840 ( .A(n15786), .B(n15788), .Z(n7897) );
  NAND U17841 ( .A(n15794), .B(nreg[734]), .Z(n15788) );
  NAND U17842 ( .A(n12326), .B(nreg[734]), .Z(n15794) );
  XNOR U17843 ( .A(n15784), .B(n15795), .Z(n15786) );
  XOR U17844 ( .A(n15796), .B(n15797), .Z(n15784) );
  AND U17845 ( .A(n15798), .B(n15799), .Z(n15797) );
  XNOR U17846 ( .A(n15800), .B(n15796), .Z(n15799) );
  XOR U17847 ( .A(n15801), .B(nreg[734]), .Z(n15792) );
  IV U17848 ( .A(n15790), .Z(n15801) );
  XOR U17849 ( .A(n15802), .B(n15803), .Z(n15790) );
  AND U17850 ( .A(n15804), .B(n15805), .Z(n15803) );
  XNOR U17851 ( .A(n15802), .B(n7903), .Z(n15805) );
  XNOR U17852 ( .A(n15798), .B(n15800), .Z(n7903) );
  NAND U17853 ( .A(n15806), .B(nreg[733]), .Z(n15800) );
  NAND U17854 ( .A(n12326), .B(nreg[733]), .Z(n15806) );
  XNOR U17855 ( .A(n15796), .B(n15807), .Z(n15798) );
  XOR U17856 ( .A(n15808), .B(n15809), .Z(n15796) );
  AND U17857 ( .A(n15810), .B(n15811), .Z(n15809) );
  XNOR U17858 ( .A(n15812), .B(n15808), .Z(n15811) );
  XOR U17859 ( .A(n15813), .B(nreg[733]), .Z(n15804) );
  IV U17860 ( .A(n15802), .Z(n15813) );
  XOR U17861 ( .A(n15814), .B(n15815), .Z(n15802) );
  AND U17862 ( .A(n15816), .B(n15817), .Z(n15815) );
  XNOR U17863 ( .A(n15814), .B(n7909), .Z(n15817) );
  XNOR U17864 ( .A(n15810), .B(n15812), .Z(n7909) );
  NAND U17865 ( .A(n15818), .B(nreg[732]), .Z(n15812) );
  NAND U17866 ( .A(n12326), .B(nreg[732]), .Z(n15818) );
  XNOR U17867 ( .A(n15808), .B(n15819), .Z(n15810) );
  XOR U17868 ( .A(n15820), .B(n15821), .Z(n15808) );
  AND U17869 ( .A(n15822), .B(n15823), .Z(n15821) );
  XNOR U17870 ( .A(n15824), .B(n15820), .Z(n15823) );
  XOR U17871 ( .A(n15825), .B(nreg[732]), .Z(n15816) );
  IV U17872 ( .A(n15814), .Z(n15825) );
  XOR U17873 ( .A(n15826), .B(n15827), .Z(n15814) );
  AND U17874 ( .A(n15828), .B(n15829), .Z(n15827) );
  XNOR U17875 ( .A(n15826), .B(n7915), .Z(n15829) );
  XNOR U17876 ( .A(n15822), .B(n15824), .Z(n7915) );
  NAND U17877 ( .A(n15830), .B(nreg[731]), .Z(n15824) );
  NAND U17878 ( .A(n12326), .B(nreg[731]), .Z(n15830) );
  XNOR U17879 ( .A(n15820), .B(n15831), .Z(n15822) );
  XOR U17880 ( .A(n15832), .B(n15833), .Z(n15820) );
  AND U17881 ( .A(n15834), .B(n15835), .Z(n15833) );
  XNOR U17882 ( .A(n15836), .B(n15832), .Z(n15835) );
  XOR U17883 ( .A(n15837), .B(nreg[731]), .Z(n15828) );
  IV U17884 ( .A(n15826), .Z(n15837) );
  XOR U17885 ( .A(n15838), .B(n15839), .Z(n15826) );
  AND U17886 ( .A(n15840), .B(n15841), .Z(n15839) );
  XNOR U17887 ( .A(n15838), .B(n7921), .Z(n15841) );
  XNOR U17888 ( .A(n15834), .B(n15836), .Z(n7921) );
  NAND U17889 ( .A(n15842), .B(nreg[730]), .Z(n15836) );
  NAND U17890 ( .A(n12326), .B(nreg[730]), .Z(n15842) );
  XNOR U17891 ( .A(n15832), .B(n15843), .Z(n15834) );
  XOR U17892 ( .A(n15844), .B(n15845), .Z(n15832) );
  AND U17893 ( .A(n15846), .B(n15847), .Z(n15845) );
  XNOR U17894 ( .A(n15848), .B(n15844), .Z(n15847) );
  XOR U17895 ( .A(n15849), .B(nreg[730]), .Z(n15840) );
  IV U17896 ( .A(n15838), .Z(n15849) );
  XOR U17897 ( .A(n15850), .B(n15851), .Z(n15838) );
  AND U17898 ( .A(n15852), .B(n15853), .Z(n15851) );
  XNOR U17899 ( .A(n15850), .B(n7927), .Z(n15853) );
  XNOR U17900 ( .A(n15846), .B(n15848), .Z(n7927) );
  NAND U17901 ( .A(n15854), .B(nreg[729]), .Z(n15848) );
  NAND U17902 ( .A(n12326), .B(nreg[729]), .Z(n15854) );
  XNOR U17903 ( .A(n15844), .B(n15855), .Z(n15846) );
  XOR U17904 ( .A(n15856), .B(n15857), .Z(n15844) );
  AND U17905 ( .A(n15858), .B(n15859), .Z(n15857) );
  XNOR U17906 ( .A(n15860), .B(n15856), .Z(n15859) );
  XOR U17907 ( .A(n15861), .B(nreg[729]), .Z(n15852) );
  IV U17908 ( .A(n15850), .Z(n15861) );
  XOR U17909 ( .A(n15862), .B(n15863), .Z(n15850) );
  AND U17910 ( .A(n15864), .B(n15865), .Z(n15863) );
  XNOR U17911 ( .A(n15862), .B(n7933), .Z(n15865) );
  XNOR U17912 ( .A(n15858), .B(n15860), .Z(n7933) );
  NAND U17913 ( .A(n15866), .B(nreg[728]), .Z(n15860) );
  NAND U17914 ( .A(n12326), .B(nreg[728]), .Z(n15866) );
  XNOR U17915 ( .A(n15856), .B(n15867), .Z(n15858) );
  XOR U17916 ( .A(n15868), .B(n15869), .Z(n15856) );
  AND U17917 ( .A(n15870), .B(n15871), .Z(n15869) );
  XNOR U17918 ( .A(n15872), .B(n15868), .Z(n15871) );
  XOR U17919 ( .A(n15873), .B(nreg[728]), .Z(n15864) );
  IV U17920 ( .A(n15862), .Z(n15873) );
  XOR U17921 ( .A(n15874), .B(n15875), .Z(n15862) );
  AND U17922 ( .A(n15876), .B(n15877), .Z(n15875) );
  XNOR U17923 ( .A(n15874), .B(n7939), .Z(n15877) );
  XNOR U17924 ( .A(n15870), .B(n15872), .Z(n7939) );
  NAND U17925 ( .A(n15878), .B(nreg[727]), .Z(n15872) );
  NAND U17926 ( .A(n12326), .B(nreg[727]), .Z(n15878) );
  XNOR U17927 ( .A(n15868), .B(n15879), .Z(n15870) );
  XOR U17928 ( .A(n15880), .B(n15881), .Z(n15868) );
  AND U17929 ( .A(n15882), .B(n15883), .Z(n15881) );
  XNOR U17930 ( .A(n15884), .B(n15880), .Z(n15883) );
  XOR U17931 ( .A(n15885), .B(nreg[727]), .Z(n15876) );
  IV U17932 ( .A(n15874), .Z(n15885) );
  XOR U17933 ( .A(n15886), .B(n15887), .Z(n15874) );
  AND U17934 ( .A(n15888), .B(n15889), .Z(n15887) );
  XNOR U17935 ( .A(n15886), .B(n7945), .Z(n15889) );
  XNOR U17936 ( .A(n15882), .B(n15884), .Z(n7945) );
  NAND U17937 ( .A(n15890), .B(nreg[726]), .Z(n15884) );
  NAND U17938 ( .A(n12326), .B(nreg[726]), .Z(n15890) );
  XNOR U17939 ( .A(n15880), .B(n15891), .Z(n15882) );
  XOR U17940 ( .A(n15892), .B(n15893), .Z(n15880) );
  AND U17941 ( .A(n15894), .B(n15895), .Z(n15893) );
  XNOR U17942 ( .A(n15896), .B(n15892), .Z(n15895) );
  XOR U17943 ( .A(n15897), .B(nreg[726]), .Z(n15888) );
  IV U17944 ( .A(n15886), .Z(n15897) );
  XOR U17945 ( .A(n15898), .B(n15899), .Z(n15886) );
  AND U17946 ( .A(n15900), .B(n15901), .Z(n15899) );
  XNOR U17947 ( .A(n15898), .B(n7951), .Z(n15901) );
  XNOR U17948 ( .A(n15894), .B(n15896), .Z(n7951) );
  NAND U17949 ( .A(n15902), .B(nreg[725]), .Z(n15896) );
  NAND U17950 ( .A(n12326), .B(nreg[725]), .Z(n15902) );
  XNOR U17951 ( .A(n15892), .B(n15903), .Z(n15894) );
  XOR U17952 ( .A(n15904), .B(n15905), .Z(n15892) );
  AND U17953 ( .A(n15906), .B(n15907), .Z(n15905) );
  XNOR U17954 ( .A(n15908), .B(n15904), .Z(n15907) );
  XOR U17955 ( .A(n15909), .B(nreg[725]), .Z(n15900) );
  IV U17956 ( .A(n15898), .Z(n15909) );
  XOR U17957 ( .A(n15910), .B(n15911), .Z(n15898) );
  AND U17958 ( .A(n15912), .B(n15913), .Z(n15911) );
  XNOR U17959 ( .A(n15910), .B(n7957), .Z(n15913) );
  XNOR U17960 ( .A(n15906), .B(n15908), .Z(n7957) );
  NAND U17961 ( .A(n15914), .B(nreg[724]), .Z(n15908) );
  NAND U17962 ( .A(n12326), .B(nreg[724]), .Z(n15914) );
  XNOR U17963 ( .A(n15904), .B(n15915), .Z(n15906) );
  XOR U17964 ( .A(n15916), .B(n15917), .Z(n15904) );
  AND U17965 ( .A(n15918), .B(n15919), .Z(n15917) );
  XNOR U17966 ( .A(n15920), .B(n15916), .Z(n15919) );
  XOR U17967 ( .A(n15921), .B(nreg[724]), .Z(n15912) );
  IV U17968 ( .A(n15910), .Z(n15921) );
  XOR U17969 ( .A(n15922), .B(n15923), .Z(n15910) );
  AND U17970 ( .A(n15924), .B(n15925), .Z(n15923) );
  XNOR U17971 ( .A(n15922), .B(n7963), .Z(n15925) );
  XNOR U17972 ( .A(n15918), .B(n15920), .Z(n7963) );
  NAND U17973 ( .A(n15926), .B(nreg[723]), .Z(n15920) );
  NAND U17974 ( .A(n12326), .B(nreg[723]), .Z(n15926) );
  XNOR U17975 ( .A(n15916), .B(n15927), .Z(n15918) );
  XOR U17976 ( .A(n15928), .B(n15929), .Z(n15916) );
  AND U17977 ( .A(n15930), .B(n15931), .Z(n15929) );
  XNOR U17978 ( .A(n15932), .B(n15928), .Z(n15931) );
  XOR U17979 ( .A(n15933), .B(nreg[723]), .Z(n15924) );
  IV U17980 ( .A(n15922), .Z(n15933) );
  XOR U17981 ( .A(n15934), .B(n15935), .Z(n15922) );
  AND U17982 ( .A(n15936), .B(n15937), .Z(n15935) );
  XNOR U17983 ( .A(n15934), .B(n7969), .Z(n15937) );
  XNOR U17984 ( .A(n15930), .B(n15932), .Z(n7969) );
  NAND U17985 ( .A(n15938), .B(nreg[722]), .Z(n15932) );
  NAND U17986 ( .A(n12326), .B(nreg[722]), .Z(n15938) );
  XNOR U17987 ( .A(n15928), .B(n15939), .Z(n15930) );
  XOR U17988 ( .A(n15940), .B(n15941), .Z(n15928) );
  AND U17989 ( .A(n15942), .B(n15943), .Z(n15941) );
  XNOR U17990 ( .A(n15944), .B(n15940), .Z(n15943) );
  XOR U17991 ( .A(n15945), .B(nreg[722]), .Z(n15936) );
  IV U17992 ( .A(n15934), .Z(n15945) );
  XOR U17993 ( .A(n15946), .B(n15947), .Z(n15934) );
  AND U17994 ( .A(n15948), .B(n15949), .Z(n15947) );
  XNOR U17995 ( .A(n15946), .B(n7975), .Z(n15949) );
  XNOR U17996 ( .A(n15942), .B(n15944), .Z(n7975) );
  NAND U17997 ( .A(n15950), .B(nreg[721]), .Z(n15944) );
  NAND U17998 ( .A(n12326), .B(nreg[721]), .Z(n15950) );
  XNOR U17999 ( .A(n15940), .B(n15951), .Z(n15942) );
  XOR U18000 ( .A(n15952), .B(n15953), .Z(n15940) );
  AND U18001 ( .A(n15954), .B(n15955), .Z(n15953) );
  XNOR U18002 ( .A(n15956), .B(n15952), .Z(n15955) );
  XOR U18003 ( .A(n15957), .B(nreg[721]), .Z(n15948) );
  IV U18004 ( .A(n15946), .Z(n15957) );
  XOR U18005 ( .A(n15958), .B(n15959), .Z(n15946) );
  AND U18006 ( .A(n15960), .B(n15961), .Z(n15959) );
  XNOR U18007 ( .A(n15958), .B(n7981), .Z(n15961) );
  XNOR U18008 ( .A(n15954), .B(n15956), .Z(n7981) );
  NAND U18009 ( .A(n15962), .B(nreg[720]), .Z(n15956) );
  NAND U18010 ( .A(n12326), .B(nreg[720]), .Z(n15962) );
  XNOR U18011 ( .A(n15952), .B(n15963), .Z(n15954) );
  XOR U18012 ( .A(n15964), .B(n15965), .Z(n15952) );
  AND U18013 ( .A(n15966), .B(n15967), .Z(n15965) );
  XNOR U18014 ( .A(n15968), .B(n15964), .Z(n15967) );
  XOR U18015 ( .A(n15969), .B(nreg[720]), .Z(n15960) );
  IV U18016 ( .A(n15958), .Z(n15969) );
  XOR U18017 ( .A(n15970), .B(n15971), .Z(n15958) );
  AND U18018 ( .A(n15972), .B(n15973), .Z(n15971) );
  XNOR U18019 ( .A(n15970), .B(n7987), .Z(n15973) );
  XNOR U18020 ( .A(n15966), .B(n15968), .Z(n7987) );
  NAND U18021 ( .A(n15974), .B(nreg[719]), .Z(n15968) );
  NAND U18022 ( .A(n12326), .B(nreg[719]), .Z(n15974) );
  XNOR U18023 ( .A(n15964), .B(n15975), .Z(n15966) );
  XOR U18024 ( .A(n15976), .B(n15977), .Z(n15964) );
  AND U18025 ( .A(n15978), .B(n15979), .Z(n15977) );
  XNOR U18026 ( .A(n15980), .B(n15976), .Z(n15979) );
  XOR U18027 ( .A(n15981), .B(nreg[719]), .Z(n15972) );
  IV U18028 ( .A(n15970), .Z(n15981) );
  XOR U18029 ( .A(n15982), .B(n15983), .Z(n15970) );
  AND U18030 ( .A(n15984), .B(n15985), .Z(n15983) );
  XNOR U18031 ( .A(n15982), .B(n7993), .Z(n15985) );
  XNOR U18032 ( .A(n15978), .B(n15980), .Z(n7993) );
  NAND U18033 ( .A(n15986), .B(nreg[718]), .Z(n15980) );
  NAND U18034 ( .A(n12326), .B(nreg[718]), .Z(n15986) );
  XNOR U18035 ( .A(n15976), .B(n15987), .Z(n15978) );
  XOR U18036 ( .A(n15988), .B(n15989), .Z(n15976) );
  AND U18037 ( .A(n15990), .B(n15991), .Z(n15989) );
  XNOR U18038 ( .A(n15992), .B(n15988), .Z(n15991) );
  XOR U18039 ( .A(n15993), .B(nreg[718]), .Z(n15984) );
  IV U18040 ( .A(n15982), .Z(n15993) );
  XOR U18041 ( .A(n15994), .B(n15995), .Z(n15982) );
  AND U18042 ( .A(n15996), .B(n15997), .Z(n15995) );
  XNOR U18043 ( .A(n15994), .B(n7999), .Z(n15997) );
  XNOR U18044 ( .A(n15990), .B(n15992), .Z(n7999) );
  NAND U18045 ( .A(n15998), .B(nreg[717]), .Z(n15992) );
  NAND U18046 ( .A(n12326), .B(nreg[717]), .Z(n15998) );
  XNOR U18047 ( .A(n15988), .B(n15999), .Z(n15990) );
  XOR U18048 ( .A(n16000), .B(n16001), .Z(n15988) );
  AND U18049 ( .A(n16002), .B(n16003), .Z(n16001) );
  XNOR U18050 ( .A(n16004), .B(n16000), .Z(n16003) );
  XOR U18051 ( .A(n16005), .B(nreg[717]), .Z(n15996) );
  IV U18052 ( .A(n15994), .Z(n16005) );
  XOR U18053 ( .A(n16006), .B(n16007), .Z(n15994) );
  AND U18054 ( .A(n16008), .B(n16009), .Z(n16007) );
  XNOR U18055 ( .A(n16006), .B(n8005), .Z(n16009) );
  XNOR U18056 ( .A(n16002), .B(n16004), .Z(n8005) );
  NAND U18057 ( .A(n16010), .B(nreg[716]), .Z(n16004) );
  NAND U18058 ( .A(n12326), .B(nreg[716]), .Z(n16010) );
  XNOR U18059 ( .A(n16000), .B(n16011), .Z(n16002) );
  XOR U18060 ( .A(n16012), .B(n16013), .Z(n16000) );
  AND U18061 ( .A(n16014), .B(n16015), .Z(n16013) );
  XNOR U18062 ( .A(n16016), .B(n16012), .Z(n16015) );
  XOR U18063 ( .A(n16017), .B(nreg[716]), .Z(n16008) );
  IV U18064 ( .A(n16006), .Z(n16017) );
  XOR U18065 ( .A(n16018), .B(n16019), .Z(n16006) );
  AND U18066 ( .A(n16020), .B(n16021), .Z(n16019) );
  XNOR U18067 ( .A(n16018), .B(n8011), .Z(n16021) );
  XNOR U18068 ( .A(n16014), .B(n16016), .Z(n8011) );
  NAND U18069 ( .A(n16022), .B(nreg[715]), .Z(n16016) );
  NAND U18070 ( .A(n12326), .B(nreg[715]), .Z(n16022) );
  XNOR U18071 ( .A(n16012), .B(n16023), .Z(n16014) );
  XOR U18072 ( .A(n16024), .B(n16025), .Z(n16012) );
  AND U18073 ( .A(n16026), .B(n16027), .Z(n16025) );
  XNOR U18074 ( .A(n16028), .B(n16024), .Z(n16027) );
  XOR U18075 ( .A(n16029), .B(nreg[715]), .Z(n16020) );
  IV U18076 ( .A(n16018), .Z(n16029) );
  XOR U18077 ( .A(n16030), .B(n16031), .Z(n16018) );
  AND U18078 ( .A(n16032), .B(n16033), .Z(n16031) );
  XNOR U18079 ( .A(n16030), .B(n8017), .Z(n16033) );
  XNOR U18080 ( .A(n16026), .B(n16028), .Z(n8017) );
  NAND U18081 ( .A(n16034), .B(nreg[714]), .Z(n16028) );
  NAND U18082 ( .A(n12326), .B(nreg[714]), .Z(n16034) );
  XNOR U18083 ( .A(n16024), .B(n16035), .Z(n16026) );
  XOR U18084 ( .A(n16036), .B(n16037), .Z(n16024) );
  AND U18085 ( .A(n16038), .B(n16039), .Z(n16037) );
  XNOR U18086 ( .A(n16040), .B(n16036), .Z(n16039) );
  XOR U18087 ( .A(n16041), .B(nreg[714]), .Z(n16032) );
  IV U18088 ( .A(n16030), .Z(n16041) );
  XOR U18089 ( .A(n16042), .B(n16043), .Z(n16030) );
  AND U18090 ( .A(n16044), .B(n16045), .Z(n16043) );
  XNOR U18091 ( .A(n16042), .B(n8023), .Z(n16045) );
  XNOR U18092 ( .A(n16038), .B(n16040), .Z(n8023) );
  NAND U18093 ( .A(n16046), .B(nreg[713]), .Z(n16040) );
  NAND U18094 ( .A(n12326), .B(nreg[713]), .Z(n16046) );
  XNOR U18095 ( .A(n16036), .B(n16047), .Z(n16038) );
  XOR U18096 ( .A(n16048), .B(n16049), .Z(n16036) );
  AND U18097 ( .A(n16050), .B(n16051), .Z(n16049) );
  XNOR U18098 ( .A(n16052), .B(n16048), .Z(n16051) );
  XOR U18099 ( .A(n16053), .B(nreg[713]), .Z(n16044) );
  IV U18100 ( .A(n16042), .Z(n16053) );
  XOR U18101 ( .A(n16054), .B(n16055), .Z(n16042) );
  AND U18102 ( .A(n16056), .B(n16057), .Z(n16055) );
  XNOR U18103 ( .A(n16054), .B(n8029), .Z(n16057) );
  XNOR U18104 ( .A(n16050), .B(n16052), .Z(n8029) );
  NAND U18105 ( .A(n16058), .B(nreg[712]), .Z(n16052) );
  NAND U18106 ( .A(n12326), .B(nreg[712]), .Z(n16058) );
  XNOR U18107 ( .A(n16048), .B(n16059), .Z(n16050) );
  XOR U18108 ( .A(n16060), .B(n16061), .Z(n16048) );
  AND U18109 ( .A(n16062), .B(n16063), .Z(n16061) );
  XNOR U18110 ( .A(n16064), .B(n16060), .Z(n16063) );
  XOR U18111 ( .A(n16065), .B(nreg[712]), .Z(n16056) );
  IV U18112 ( .A(n16054), .Z(n16065) );
  XOR U18113 ( .A(n16066), .B(n16067), .Z(n16054) );
  AND U18114 ( .A(n16068), .B(n16069), .Z(n16067) );
  XNOR U18115 ( .A(n16066), .B(n8035), .Z(n16069) );
  XNOR U18116 ( .A(n16062), .B(n16064), .Z(n8035) );
  NAND U18117 ( .A(n16070), .B(nreg[711]), .Z(n16064) );
  NAND U18118 ( .A(n12326), .B(nreg[711]), .Z(n16070) );
  XNOR U18119 ( .A(n16060), .B(n16071), .Z(n16062) );
  XOR U18120 ( .A(n16072), .B(n16073), .Z(n16060) );
  AND U18121 ( .A(n16074), .B(n16075), .Z(n16073) );
  XNOR U18122 ( .A(n16076), .B(n16072), .Z(n16075) );
  XOR U18123 ( .A(n16077), .B(nreg[711]), .Z(n16068) );
  IV U18124 ( .A(n16066), .Z(n16077) );
  XOR U18125 ( .A(n16078), .B(n16079), .Z(n16066) );
  AND U18126 ( .A(n16080), .B(n16081), .Z(n16079) );
  XNOR U18127 ( .A(n16078), .B(n8041), .Z(n16081) );
  XNOR U18128 ( .A(n16074), .B(n16076), .Z(n8041) );
  NAND U18129 ( .A(n16082), .B(nreg[710]), .Z(n16076) );
  NAND U18130 ( .A(n12326), .B(nreg[710]), .Z(n16082) );
  XNOR U18131 ( .A(n16072), .B(n16083), .Z(n16074) );
  XOR U18132 ( .A(n16084), .B(n16085), .Z(n16072) );
  AND U18133 ( .A(n16086), .B(n16087), .Z(n16085) );
  XNOR U18134 ( .A(n16088), .B(n16084), .Z(n16087) );
  XOR U18135 ( .A(n16089), .B(nreg[710]), .Z(n16080) );
  IV U18136 ( .A(n16078), .Z(n16089) );
  XOR U18137 ( .A(n16090), .B(n16091), .Z(n16078) );
  AND U18138 ( .A(n16092), .B(n16093), .Z(n16091) );
  XNOR U18139 ( .A(n16090), .B(n8047), .Z(n16093) );
  XNOR U18140 ( .A(n16086), .B(n16088), .Z(n8047) );
  NAND U18141 ( .A(n16094), .B(nreg[709]), .Z(n16088) );
  NAND U18142 ( .A(n12326), .B(nreg[709]), .Z(n16094) );
  XNOR U18143 ( .A(n16084), .B(n16095), .Z(n16086) );
  XOR U18144 ( .A(n16096), .B(n16097), .Z(n16084) );
  AND U18145 ( .A(n16098), .B(n16099), .Z(n16097) );
  XNOR U18146 ( .A(n16100), .B(n16096), .Z(n16099) );
  XOR U18147 ( .A(n16101), .B(nreg[709]), .Z(n16092) );
  IV U18148 ( .A(n16090), .Z(n16101) );
  XOR U18149 ( .A(n16102), .B(n16103), .Z(n16090) );
  AND U18150 ( .A(n16104), .B(n16105), .Z(n16103) );
  XNOR U18151 ( .A(n16102), .B(n8053), .Z(n16105) );
  XNOR U18152 ( .A(n16098), .B(n16100), .Z(n8053) );
  NAND U18153 ( .A(n16106), .B(nreg[708]), .Z(n16100) );
  NAND U18154 ( .A(n12326), .B(nreg[708]), .Z(n16106) );
  XNOR U18155 ( .A(n16096), .B(n16107), .Z(n16098) );
  XOR U18156 ( .A(n16108), .B(n16109), .Z(n16096) );
  AND U18157 ( .A(n16110), .B(n16111), .Z(n16109) );
  XNOR U18158 ( .A(n16112), .B(n16108), .Z(n16111) );
  XOR U18159 ( .A(n16113), .B(nreg[708]), .Z(n16104) );
  IV U18160 ( .A(n16102), .Z(n16113) );
  XOR U18161 ( .A(n16114), .B(n16115), .Z(n16102) );
  AND U18162 ( .A(n16116), .B(n16117), .Z(n16115) );
  XNOR U18163 ( .A(n16114), .B(n8059), .Z(n16117) );
  XNOR U18164 ( .A(n16110), .B(n16112), .Z(n8059) );
  NAND U18165 ( .A(n16118), .B(nreg[707]), .Z(n16112) );
  NAND U18166 ( .A(n12326), .B(nreg[707]), .Z(n16118) );
  XNOR U18167 ( .A(n16108), .B(n16119), .Z(n16110) );
  XOR U18168 ( .A(n16120), .B(n16121), .Z(n16108) );
  AND U18169 ( .A(n16122), .B(n16123), .Z(n16121) );
  XNOR U18170 ( .A(n16124), .B(n16120), .Z(n16123) );
  XOR U18171 ( .A(n16125), .B(nreg[707]), .Z(n16116) );
  IV U18172 ( .A(n16114), .Z(n16125) );
  XOR U18173 ( .A(n16126), .B(n16127), .Z(n16114) );
  AND U18174 ( .A(n16128), .B(n16129), .Z(n16127) );
  XNOR U18175 ( .A(n16126), .B(n8065), .Z(n16129) );
  XNOR U18176 ( .A(n16122), .B(n16124), .Z(n8065) );
  NAND U18177 ( .A(n16130), .B(nreg[706]), .Z(n16124) );
  NAND U18178 ( .A(n12326), .B(nreg[706]), .Z(n16130) );
  XNOR U18179 ( .A(n16120), .B(n16131), .Z(n16122) );
  XOR U18180 ( .A(n16132), .B(n16133), .Z(n16120) );
  AND U18181 ( .A(n16134), .B(n16135), .Z(n16133) );
  XNOR U18182 ( .A(n16136), .B(n16132), .Z(n16135) );
  XOR U18183 ( .A(n16137), .B(nreg[706]), .Z(n16128) );
  IV U18184 ( .A(n16126), .Z(n16137) );
  XOR U18185 ( .A(n16138), .B(n16139), .Z(n16126) );
  AND U18186 ( .A(n16140), .B(n16141), .Z(n16139) );
  XNOR U18187 ( .A(n16138), .B(n8071), .Z(n16141) );
  XNOR U18188 ( .A(n16134), .B(n16136), .Z(n8071) );
  NAND U18189 ( .A(n16142), .B(nreg[705]), .Z(n16136) );
  NAND U18190 ( .A(n12326), .B(nreg[705]), .Z(n16142) );
  XNOR U18191 ( .A(n16132), .B(n16143), .Z(n16134) );
  XOR U18192 ( .A(n16144), .B(n16145), .Z(n16132) );
  AND U18193 ( .A(n16146), .B(n16147), .Z(n16145) );
  XNOR U18194 ( .A(n16148), .B(n16144), .Z(n16147) );
  XOR U18195 ( .A(n16149), .B(nreg[705]), .Z(n16140) );
  IV U18196 ( .A(n16138), .Z(n16149) );
  XOR U18197 ( .A(n16150), .B(n16151), .Z(n16138) );
  AND U18198 ( .A(n16152), .B(n16153), .Z(n16151) );
  XNOR U18199 ( .A(n16150), .B(n8077), .Z(n16153) );
  XNOR U18200 ( .A(n16146), .B(n16148), .Z(n8077) );
  NAND U18201 ( .A(n16154), .B(nreg[704]), .Z(n16148) );
  NAND U18202 ( .A(n12326), .B(nreg[704]), .Z(n16154) );
  XNOR U18203 ( .A(n16144), .B(n16155), .Z(n16146) );
  XOR U18204 ( .A(n16156), .B(n16157), .Z(n16144) );
  AND U18205 ( .A(n16158), .B(n16159), .Z(n16157) );
  XNOR U18206 ( .A(n16160), .B(n16156), .Z(n16159) );
  XOR U18207 ( .A(n16161), .B(nreg[704]), .Z(n16152) );
  IV U18208 ( .A(n16150), .Z(n16161) );
  XOR U18209 ( .A(n16162), .B(n16163), .Z(n16150) );
  AND U18210 ( .A(n16164), .B(n16165), .Z(n16163) );
  XNOR U18211 ( .A(n16162), .B(n8083), .Z(n16165) );
  XNOR U18212 ( .A(n16158), .B(n16160), .Z(n8083) );
  NAND U18213 ( .A(n16166), .B(nreg[703]), .Z(n16160) );
  NAND U18214 ( .A(n12326), .B(nreg[703]), .Z(n16166) );
  XNOR U18215 ( .A(n16156), .B(n16167), .Z(n16158) );
  XOR U18216 ( .A(n16168), .B(n16169), .Z(n16156) );
  AND U18217 ( .A(n16170), .B(n16171), .Z(n16169) );
  XNOR U18218 ( .A(n16172), .B(n16168), .Z(n16171) );
  XOR U18219 ( .A(n16173), .B(nreg[703]), .Z(n16164) );
  IV U18220 ( .A(n16162), .Z(n16173) );
  XOR U18221 ( .A(n16174), .B(n16175), .Z(n16162) );
  AND U18222 ( .A(n16176), .B(n16177), .Z(n16175) );
  XNOR U18223 ( .A(n16174), .B(n8089), .Z(n16177) );
  XNOR U18224 ( .A(n16170), .B(n16172), .Z(n8089) );
  NAND U18225 ( .A(n16178), .B(nreg[702]), .Z(n16172) );
  NAND U18226 ( .A(n12326), .B(nreg[702]), .Z(n16178) );
  XNOR U18227 ( .A(n16168), .B(n16179), .Z(n16170) );
  XOR U18228 ( .A(n16180), .B(n16181), .Z(n16168) );
  AND U18229 ( .A(n16182), .B(n16183), .Z(n16181) );
  XNOR U18230 ( .A(n16184), .B(n16180), .Z(n16183) );
  XOR U18231 ( .A(n16185), .B(nreg[702]), .Z(n16176) );
  IV U18232 ( .A(n16174), .Z(n16185) );
  XOR U18233 ( .A(n16186), .B(n16187), .Z(n16174) );
  AND U18234 ( .A(n16188), .B(n16189), .Z(n16187) );
  XNOR U18235 ( .A(n16186), .B(n8095), .Z(n16189) );
  XNOR U18236 ( .A(n16182), .B(n16184), .Z(n8095) );
  NAND U18237 ( .A(n16190), .B(nreg[701]), .Z(n16184) );
  NAND U18238 ( .A(n12326), .B(nreg[701]), .Z(n16190) );
  XNOR U18239 ( .A(n16180), .B(n16191), .Z(n16182) );
  XOR U18240 ( .A(n16192), .B(n16193), .Z(n16180) );
  AND U18241 ( .A(n16194), .B(n16195), .Z(n16193) );
  XNOR U18242 ( .A(n16196), .B(n16192), .Z(n16195) );
  XOR U18243 ( .A(n16197), .B(nreg[701]), .Z(n16188) );
  IV U18244 ( .A(n16186), .Z(n16197) );
  XOR U18245 ( .A(n16198), .B(n16199), .Z(n16186) );
  AND U18246 ( .A(n16200), .B(n16201), .Z(n16199) );
  XNOR U18247 ( .A(n16198), .B(n8101), .Z(n16201) );
  XNOR U18248 ( .A(n16194), .B(n16196), .Z(n8101) );
  NAND U18249 ( .A(n16202), .B(nreg[700]), .Z(n16196) );
  NAND U18250 ( .A(n12326), .B(nreg[700]), .Z(n16202) );
  XNOR U18251 ( .A(n16192), .B(n16203), .Z(n16194) );
  XOR U18252 ( .A(n16204), .B(n16205), .Z(n16192) );
  AND U18253 ( .A(n16206), .B(n16207), .Z(n16205) );
  XNOR U18254 ( .A(n16208), .B(n16204), .Z(n16207) );
  XOR U18255 ( .A(n16209), .B(nreg[700]), .Z(n16200) );
  IV U18256 ( .A(n16198), .Z(n16209) );
  XOR U18257 ( .A(n16210), .B(n16211), .Z(n16198) );
  AND U18258 ( .A(n16212), .B(n16213), .Z(n16211) );
  XNOR U18259 ( .A(n16210), .B(n8107), .Z(n16213) );
  XNOR U18260 ( .A(n16206), .B(n16208), .Z(n8107) );
  NAND U18261 ( .A(n16214), .B(nreg[699]), .Z(n16208) );
  NAND U18262 ( .A(n12326), .B(nreg[699]), .Z(n16214) );
  XNOR U18263 ( .A(n16204), .B(n16215), .Z(n16206) );
  XOR U18264 ( .A(n16216), .B(n16217), .Z(n16204) );
  AND U18265 ( .A(n16218), .B(n16219), .Z(n16217) );
  XNOR U18266 ( .A(n16220), .B(n16216), .Z(n16219) );
  XOR U18267 ( .A(n16221), .B(nreg[699]), .Z(n16212) );
  IV U18268 ( .A(n16210), .Z(n16221) );
  XOR U18269 ( .A(n16222), .B(n16223), .Z(n16210) );
  AND U18270 ( .A(n16224), .B(n16225), .Z(n16223) );
  XNOR U18271 ( .A(n16222), .B(n8113), .Z(n16225) );
  XNOR U18272 ( .A(n16218), .B(n16220), .Z(n8113) );
  NAND U18273 ( .A(n16226), .B(nreg[698]), .Z(n16220) );
  NAND U18274 ( .A(n12326), .B(nreg[698]), .Z(n16226) );
  XNOR U18275 ( .A(n16216), .B(n16227), .Z(n16218) );
  XOR U18276 ( .A(n16228), .B(n16229), .Z(n16216) );
  AND U18277 ( .A(n16230), .B(n16231), .Z(n16229) );
  XNOR U18278 ( .A(n16232), .B(n16228), .Z(n16231) );
  XOR U18279 ( .A(n16233), .B(nreg[698]), .Z(n16224) );
  IV U18280 ( .A(n16222), .Z(n16233) );
  XOR U18281 ( .A(n16234), .B(n16235), .Z(n16222) );
  AND U18282 ( .A(n16236), .B(n16237), .Z(n16235) );
  XNOR U18283 ( .A(n16234), .B(n8119), .Z(n16237) );
  XNOR U18284 ( .A(n16230), .B(n16232), .Z(n8119) );
  NAND U18285 ( .A(n16238), .B(nreg[697]), .Z(n16232) );
  NAND U18286 ( .A(n12326), .B(nreg[697]), .Z(n16238) );
  XNOR U18287 ( .A(n16228), .B(n16239), .Z(n16230) );
  XOR U18288 ( .A(n16240), .B(n16241), .Z(n16228) );
  AND U18289 ( .A(n16242), .B(n16243), .Z(n16241) );
  XNOR U18290 ( .A(n16244), .B(n16240), .Z(n16243) );
  XOR U18291 ( .A(n16245), .B(nreg[697]), .Z(n16236) );
  IV U18292 ( .A(n16234), .Z(n16245) );
  XOR U18293 ( .A(n16246), .B(n16247), .Z(n16234) );
  AND U18294 ( .A(n16248), .B(n16249), .Z(n16247) );
  XNOR U18295 ( .A(n16246), .B(n8125), .Z(n16249) );
  XNOR U18296 ( .A(n16242), .B(n16244), .Z(n8125) );
  NAND U18297 ( .A(n16250), .B(nreg[696]), .Z(n16244) );
  NAND U18298 ( .A(n12326), .B(nreg[696]), .Z(n16250) );
  XNOR U18299 ( .A(n16240), .B(n16251), .Z(n16242) );
  XOR U18300 ( .A(n16252), .B(n16253), .Z(n16240) );
  AND U18301 ( .A(n16254), .B(n16255), .Z(n16253) );
  XNOR U18302 ( .A(n16256), .B(n16252), .Z(n16255) );
  XOR U18303 ( .A(n16257), .B(nreg[696]), .Z(n16248) );
  IV U18304 ( .A(n16246), .Z(n16257) );
  XOR U18305 ( .A(n16258), .B(n16259), .Z(n16246) );
  AND U18306 ( .A(n16260), .B(n16261), .Z(n16259) );
  XNOR U18307 ( .A(n16258), .B(n8131), .Z(n16261) );
  XNOR U18308 ( .A(n16254), .B(n16256), .Z(n8131) );
  NAND U18309 ( .A(n16262), .B(nreg[695]), .Z(n16256) );
  NAND U18310 ( .A(n12326), .B(nreg[695]), .Z(n16262) );
  XNOR U18311 ( .A(n16252), .B(n16263), .Z(n16254) );
  XOR U18312 ( .A(n16264), .B(n16265), .Z(n16252) );
  AND U18313 ( .A(n16266), .B(n16267), .Z(n16265) );
  XNOR U18314 ( .A(n16268), .B(n16264), .Z(n16267) );
  XOR U18315 ( .A(n16269), .B(nreg[695]), .Z(n16260) );
  IV U18316 ( .A(n16258), .Z(n16269) );
  XOR U18317 ( .A(n16270), .B(n16271), .Z(n16258) );
  AND U18318 ( .A(n16272), .B(n16273), .Z(n16271) );
  XNOR U18319 ( .A(n16270), .B(n8137), .Z(n16273) );
  XNOR U18320 ( .A(n16266), .B(n16268), .Z(n8137) );
  NAND U18321 ( .A(n16274), .B(nreg[694]), .Z(n16268) );
  NAND U18322 ( .A(n12326), .B(nreg[694]), .Z(n16274) );
  XNOR U18323 ( .A(n16264), .B(n16275), .Z(n16266) );
  XOR U18324 ( .A(n16276), .B(n16277), .Z(n16264) );
  AND U18325 ( .A(n16278), .B(n16279), .Z(n16277) );
  XNOR U18326 ( .A(n16280), .B(n16276), .Z(n16279) );
  XOR U18327 ( .A(n16281), .B(nreg[694]), .Z(n16272) );
  IV U18328 ( .A(n16270), .Z(n16281) );
  XOR U18329 ( .A(n16282), .B(n16283), .Z(n16270) );
  AND U18330 ( .A(n16284), .B(n16285), .Z(n16283) );
  XNOR U18331 ( .A(n16282), .B(n8143), .Z(n16285) );
  XNOR U18332 ( .A(n16278), .B(n16280), .Z(n8143) );
  NAND U18333 ( .A(n16286), .B(nreg[693]), .Z(n16280) );
  NAND U18334 ( .A(n12326), .B(nreg[693]), .Z(n16286) );
  XNOR U18335 ( .A(n16276), .B(n16287), .Z(n16278) );
  XOR U18336 ( .A(n16288), .B(n16289), .Z(n16276) );
  AND U18337 ( .A(n16290), .B(n16291), .Z(n16289) );
  XNOR U18338 ( .A(n16292), .B(n16288), .Z(n16291) );
  XOR U18339 ( .A(n16293), .B(nreg[693]), .Z(n16284) );
  IV U18340 ( .A(n16282), .Z(n16293) );
  XOR U18341 ( .A(n16294), .B(n16295), .Z(n16282) );
  AND U18342 ( .A(n16296), .B(n16297), .Z(n16295) );
  XNOR U18343 ( .A(n16294), .B(n8149), .Z(n16297) );
  XNOR U18344 ( .A(n16290), .B(n16292), .Z(n8149) );
  NAND U18345 ( .A(n16298), .B(nreg[692]), .Z(n16292) );
  NAND U18346 ( .A(n12326), .B(nreg[692]), .Z(n16298) );
  XNOR U18347 ( .A(n16288), .B(n16299), .Z(n16290) );
  XOR U18348 ( .A(n16300), .B(n16301), .Z(n16288) );
  AND U18349 ( .A(n16302), .B(n16303), .Z(n16301) );
  XNOR U18350 ( .A(n16304), .B(n16300), .Z(n16303) );
  XOR U18351 ( .A(n16305), .B(nreg[692]), .Z(n16296) );
  IV U18352 ( .A(n16294), .Z(n16305) );
  XOR U18353 ( .A(n16306), .B(n16307), .Z(n16294) );
  AND U18354 ( .A(n16308), .B(n16309), .Z(n16307) );
  XNOR U18355 ( .A(n16306), .B(n8155), .Z(n16309) );
  XNOR U18356 ( .A(n16302), .B(n16304), .Z(n8155) );
  NAND U18357 ( .A(n16310), .B(nreg[691]), .Z(n16304) );
  NAND U18358 ( .A(n12326), .B(nreg[691]), .Z(n16310) );
  XNOR U18359 ( .A(n16300), .B(n16311), .Z(n16302) );
  XOR U18360 ( .A(n16312), .B(n16313), .Z(n16300) );
  AND U18361 ( .A(n16314), .B(n16315), .Z(n16313) );
  XNOR U18362 ( .A(n16316), .B(n16312), .Z(n16315) );
  XOR U18363 ( .A(n16317), .B(nreg[691]), .Z(n16308) );
  IV U18364 ( .A(n16306), .Z(n16317) );
  XOR U18365 ( .A(n16318), .B(n16319), .Z(n16306) );
  AND U18366 ( .A(n16320), .B(n16321), .Z(n16319) );
  XNOR U18367 ( .A(n16318), .B(n8161), .Z(n16321) );
  XNOR U18368 ( .A(n16314), .B(n16316), .Z(n8161) );
  NAND U18369 ( .A(n16322), .B(nreg[690]), .Z(n16316) );
  NAND U18370 ( .A(n12326), .B(nreg[690]), .Z(n16322) );
  XNOR U18371 ( .A(n16312), .B(n16323), .Z(n16314) );
  XOR U18372 ( .A(n16324), .B(n16325), .Z(n16312) );
  AND U18373 ( .A(n16326), .B(n16327), .Z(n16325) );
  XNOR U18374 ( .A(n16328), .B(n16324), .Z(n16327) );
  XOR U18375 ( .A(n16329), .B(nreg[690]), .Z(n16320) );
  IV U18376 ( .A(n16318), .Z(n16329) );
  XOR U18377 ( .A(n16330), .B(n16331), .Z(n16318) );
  AND U18378 ( .A(n16332), .B(n16333), .Z(n16331) );
  XNOR U18379 ( .A(n16330), .B(n8167), .Z(n16333) );
  XNOR U18380 ( .A(n16326), .B(n16328), .Z(n8167) );
  NAND U18381 ( .A(n16334), .B(nreg[689]), .Z(n16328) );
  NAND U18382 ( .A(n12326), .B(nreg[689]), .Z(n16334) );
  XNOR U18383 ( .A(n16324), .B(n16335), .Z(n16326) );
  XOR U18384 ( .A(n16336), .B(n16337), .Z(n16324) );
  AND U18385 ( .A(n16338), .B(n16339), .Z(n16337) );
  XNOR U18386 ( .A(n16340), .B(n16336), .Z(n16339) );
  XOR U18387 ( .A(n16341), .B(nreg[689]), .Z(n16332) );
  IV U18388 ( .A(n16330), .Z(n16341) );
  XOR U18389 ( .A(n16342), .B(n16343), .Z(n16330) );
  AND U18390 ( .A(n16344), .B(n16345), .Z(n16343) );
  XNOR U18391 ( .A(n16342), .B(n8173), .Z(n16345) );
  XNOR U18392 ( .A(n16338), .B(n16340), .Z(n8173) );
  NAND U18393 ( .A(n16346), .B(nreg[688]), .Z(n16340) );
  NAND U18394 ( .A(n12326), .B(nreg[688]), .Z(n16346) );
  XNOR U18395 ( .A(n16336), .B(n16347), .Z(n16338) );
  XOR U18396 ( .A(n16348), .B(n16349), .Z(n16336) );
  AND U18397 ( .A(n16350), .B(n16351), .Z(n16349) );
  XNOR U18398 ( .A(n16352), .B(n16348), .Z(n16351) );
  XOR U18399 ( .A(n16353), .B(nreg[688]), .Z(n16344) );
  IV U18400 ( .A(n16342), .Z(n16353) );
  XOR U18401 ( .A(n16354), .B(n16355), .Z(n16342) );
  AND U18402 ( .A(n16356), .B(n16357), .Z(n16355) );
  XNOR U18403 ( .A(n16354), .B(n8179), .Z(n16357) );
  XNOR U18404 ( .A(n16350), .B(n16352), .Z(n8179) );
  NAND U18405 ( .A(n16358), .B(nreg[687]), .Z(n16352) );
  NAND U18406 ( .A(n12326), .B(nreg[687]), .Z(n16358) );
  XNOR U18407 ( .A(n16348), .B(n16359), .Z(n16350) );
  XOR U18408 ( .A(n16360), .B(n16361), .Z(n16348) );
  AND U18409 ( .A(n16362), .B(n16363), .Z(n16361) );
  XNOR U18410 ( .A(n16364), .B(n16360), .Z(n16363) );
  XOR U18411 ( .A(n16365), .B(nreg[687]), .Z(n16356) );
  IV U18412 ( .A(n16354), .Z(n16365) );
  XOR U18413 ( .A(n16366), .B(n16367), .Z(n16354) );
  AND U18414 ( .A(n16368), .B(n16369), .Z(n16367) );
  XNOR U18415 ( .A(n16366), .B(n8185), .Z(n16369) );
  XNOR U18416 ( .A(n16362), .B(n16364), .Z(n8185) );
  NAND U18417 ( .A(n16370), .B(nreg[686]), .Z(n16364) );
  NAND U18418 ( .A(n12326), .B(nreg[686]), .Z(n16370) );
  XNOR U18419 ( .A(n16360), .B(n16371), .Z(n16362) );
  XOR U18420 ( .A(n16372), .B(n16373), .Z(n16360) );
  AND U18421 ( .A(n16374), .B(n16375), .Z(n16373) );
  XNOR U18422 ( .A(n16376), .B(n16372), .Z(n16375) );
  XOR U18423 ( .A(n16377), .B(nreg[686]), .Z(n16368) );
  IV U18424 ( .A(n16366), .Z(n16377) );
  XOR U18425 ( .A(n16378), .B(n16379), .Z(n16366) );
  AND U18426 ( .A(n16380), .B(n16381), .Z(n16379) );
  XNOR U18427 ( .A(n16378), .B(n8191), .Z(n16381) );
  XNOR U18428 ( .A(n16374), .B(n16376), .Z(n8191) );
  NAND U18429 ( .A(n16382), .B(nreg[685]), .Z(n16376) );
  NAND U18430 ( .A(n12326), .B(nreg[685]), .Z(n16382) );
  XNOR U18431 ( .A(n16372), .B(n16383), .Z(n16374) );
  XOR U18432 ( .A(n16384), .B(n16385), .Z(n16372) );
  AND U18433 ( .A(n16386), .B(n16387), .Z(n16385) );
  XNOR U18434 ( .A(n16388), .B(n16384), .Z(n16387) );
  XOR U18435 ( .A(n16389), .B(nreg[685]), .Z(n16380) );
  IV U18436 ( .A(n16378), .Z(n16389) );
  XOR U18437 ( .A(n16390), .B(n16391), .Z(n16378) );
  AND U18438 ( .A(n16392), .B(n16393), .Z(n16391) );
  XNOR U18439 ( .A(n16390), .B(n8197), .Z(n16393) );
  XNOR U18440 ( .A(n16386), .B(n16388), .Z(n8197) );
  NAND U18441 ( .A(n16394), .B(nreg[684]), .Z(n16388) );
  NAND U18442 ( .A(n12326), .B(nreg[684]), .Z(n16394) );
  XNOR U18443 ( .A(n16384), .B(n16395), .Z(n16386) );
  XOR U18444 ( .A(n16396), .B(n16397), .Z(n16384) );
  AND U18445 ( .A(n16398), .B(n16399), .Z(n16397) );
  XNOR U18446 ( .A(n16400), .B(n16396), .Z(n16399) );
  XOR U18447 ( .A(n16401), .B(nreg[684]), .Z(n16392) );
  IV U18448 ( .A(n16390), .Z(n16401) );
  XOR U18449 ( .A(n16402), .B(n16403), .Z(n16390) );
  AND U18450 ( .A(n16404), .B(n16405), .Z(n16403) );
  XNOR U18451 ( .A(n16402), .B(n8203), .Z(n16405) );
  XNOR U18452 ( .A(n16398), .B(n16400), .Z(n8203) );
  NAND U18453 ( .A(n16406), .B(nreg[683]), .Z(n16400) );
  NAND U18454 ( .A(n12326), .B(nreg[683]), .Z(n16406) );
  XNOR U18455 ( .A(n16396), .B(n16407), .Z(n16398) );
  XOR U18456 ( .A(n16408), .B(n16409), .Z(n16396) );
  AND U18457 ( .A(n16410), .B(n16411), .Z(n16409) );
  XNOR U18458 ( .A(n16412), .B(n16408), .Z(n16411) );
  XOR U18459 ( .A(n16413), .B(nreg[683]), .Z(n16404) );
  IV U18460 ( .A(n16402), .Z(n16413) );
  XOR U18461 ( .A(n16414), .B(n16415), .Z(n16402) );
  AND U18462 ( .A(n16416), .B(n16417), .Z(n16415) );
  XNOR U18463 ( .A(n16414), .B(n8209), .Z(n16417) );
  XNOR U18464 ( .A(n16410), .B(n16412), .Z(n8209) );
  NAND U18465 ( .A(n16418), .B(nreg[682]), .Z(n16412) );
  NAND U18466 ( .A(n12326), .B(nreg[682]), .Z(n16418) );
  XNOR U18467 ( .A(n16408), .B(n16419), .Z(n16410) );
  XOR U18468 ( .A(n16420), .B(n16421), .Z(n16408) );
  AND U18469 ( .A(n16422), .B(n16423), .Z(n16421) );
  XNOR U18470 ( .A(n16424), .B(n16420), .Z(n16423) );
  XOR U18471 ( .A(n16425), .B(nreg[682]), .Z(n16416) );
  IV U18472 ( .A(n16414), .Z(n16425) );
  XOR U18473 ( .A(n16426), .B(n16427), .Z(n16414) );
  AND U18474 ( .A(n16428), .B(n16429), .Z(n16427) );
  XNOR U18475 ( .A(n16426), .B(n8215), .Z(n16429) );
  XNOR U18476 ( .A(n16422), .B(n16424), .Z(n8215) );
  NAND U18477 ( .A(n16430), .B(nreg[681]), .Z(n16424) );
  NAND U18478 ( .A(n12326), .B(nreg[681]), .Z(n16430) );
  XNOR U18479 ( .A(n16420), .B(n16431), .Z(n16422) );
  XOR U18480 ( .A(n16432), .B(n16433), .Z(n16420) );
  AND U18481 ( .A(n16434), .B(n16435), .Z(n16433) );
  XNOR U18482 ( .A(n16436), .B(n16432), .Z(n16435) );
  XOR U18483 ( .A(n16437), .B(nreg[681]), .Z(n16428) );
  IV U18484 ( .A(n16426), .Z(n16437) );
  XOR U18485 ( .A(n16438), .B(n16439), .Z(n16426) );
  AND U18486 ( .A(n16440), .B(n16441), .Z(n16439) );
  XNOR U18487 ( .A(n16438), .B(n8221), .Z(n16441) );
  XNOR U18488 ( .A(n16434), .B(n16436), .Z(n8221) );
  NAND U18489 ( .A(n16442), .B(nreg[680]), .Z(n16436) );
  NAND U18490 ( .A(n12326), .B(nreg[680]), .Z(n16442) );
  XNOR U18491 ( .A(n16432), .B(n16443), .Z(n16434) );
  XOR U18492 ( .A(n16444), .B(n16445), .Z(n16432) );
  AND U18493 ( .A(n16446), .B(n16447), .Z(n16445) );
  XNOR U18494 ( .A(n16448), .B(n16444), .Z(n16447) );
  XOR U18495 ( .A(n16449), .B(nreg[680]), .Z(n16440) );
  IV U18496 ( .A(n16438), .Z(n16449) );
  XOR U18497 ( .A(n16450), .B(n16451), .Z(n16438) );
  AND U18498 ( .A(n16452), .B(n16453), .Z(n16451) );
  XNOR U18499 ( .A(n16450), .B(n8227), .Z(n16453) );
  XNOR U18500 ( .A(n16446), .B(n16448), .Z(n8227) );
  NAND U18501 ( .A(n16454), .B(nreg[679]), .Z(n16448) );
  NAND U18502 ( .A(n12326), .B(nreg[679]), .Z(n16454) );
  XNOR U18503 ( .A(n16444), .B(n16455), .Z(n16446) );
  XOR U18504 ( .A(n16456), .B(n16457), .Z(n16444) );
  AND U18505 ( .A(n16458), .B(n16459), .Z(n16457) );
  XNOR U18506 ( .A(n16460), .B(n16456), .Z(n16459) );
  XOR U18507 ( .A(n16461), .B(nreg[679]), .Z(n16452) );
  IV U18508 ( .A(n16450), .Z(n16461) );
  XOR U18509 ( .A(n16462), .B(n16463), .Z(n16450) );
  AND U18510 ( .A(n16464), .B(n16465), .Z(n16463) );
  XNOR U18511 ( .A(n16462), .B(n8233), .Z(n16465) );
  XNOR U18512 ( .A(n16458), .B(n16460), .Z(n8233) );
  NAND U18513 ( .A(n16466), .B(nreg[678]), .Z(n16460) );
  NAND U18514 ( .A(n12326), .B(nreg[678]), .Z(n16466) );
  XNOR U18515 ( .A(n16456), .B(n16467), .Z(n16458) );
  XOR U18516 ( .A(n16468), .B(n16469), .Z(n16456) );
  AND U18517 ( .A(n16470), .B(n16471), .Z(n16469) );
  XNOR U18518 ( .A(n16472), .B(n16468), .Z(n16471) );
  XOR U18519 ( .A(n16473), .B(nreg[678]), .Z(n16464) );
  IV U18520 ( .A(n16462), .Z(n16473) );
  XOR U18521 ( .A(n16474), .B(n16475), .Z(n16462) );
  AND U18522 ( .A(n16476), .B(n16477), .Z(n16475) );
  XNOR U18523 ( .A(n16474), .B(n8239), .Z(n16477) );
  XNOR U18524 ( .A(n16470), .B(n16472), .Z(n8239) );
  NAND U18525 ( .A(n16478), .B(nreg[677]), .Z(n16472) );
  NAND U18526 ( .A(n12326), .B(nreg[677]), .Z(n16478) );
  XNOR U18527 ( .A(n16468), .B(n16479), .Z(n16470) );
  XOR U18528 ( .A(n16480), .B(n16481), .Z(n16468) );
  AND U18529 ( .A(n16482), .B(n16483), .Z(n16481) );
  XNOR U18530 ( .A(n16484), .B(n16480), .Z(n16483) );
  XOR U18531 ( .A(n16485), .B(nreg[677]), .Z(n16476) );
  IV U18532 ( .A(n16474), .Z(n16485) );
  XOR U18533 ( .A(n16486), .B(n16487), .Z(n16474) );
  AND U18534 ( .A(n16488), .B(n16489), .Z(n16487) );
  XNOR U18535 ( .A(n16486), .B(n8245), .Z(n16489) );
  XNOR U18536 ( .A(n16482), .B(n16484), .Z(n8245) );
  NAND U18537 ( .A(n16490), .B(nreg[676]), .Z(n16484) );
  NAND U18538 ( .A(n12326), .B(nreg[676]), .Z(n16490) );
  XNOR U18539 ( .A(n16480), .B(n16491), .Z(n16482) );
  XOR U18540 ( .A(n16492), .B(n16493), .Z(n16480) );
  AND U18541 ( .A(n16494), .B(n16495), .Z(n16493) );
  XNOR U18542 ( .A(n16496), .B(n16492), .Z(n16495) );
  XOR U18543 ( .A(n16497), .B(nreg[676]), .Z(n16488) );
  IV U18544 ( .A(n16486), .Z(n16497) );
  XOR U18545 ( .A(n16498), .B(n16499), .Z(n16486) );
  AND U18546 ( .A(n16500), .B(n16501), .Z(n16499) );
  XNOR U18547 ( .A(n16498), .B(n8251), .Z(n16501) );
  XNOR U18548 ( .A(n16494), .B(n16496), .Z(n8251) );
  NAND U18549 ( .A(n16502), .B(nreg[675]), .Z(n16496) );
  NAND U18550 ( .A(n12326), .B(nreg[675]), .Z(n16502) );
  XNOR U18551 ( .A(n16492), .B(n16503), .Z(n16494) );
  XOR U18552 ( .A(n16504), .B(n16505), .Z(n16492) );
  AND U18553 ( .A(n16506), .B(n16507), .Z(n16505) );
  XNOR U18554 ( .A(n16508), .B(n16504), .Z(n16507) );
  XOR U18555 ( .A(n16509), .B(nreg[675]), .Z(n16500) );
  IV U18556 ( .A(n16498), .Z(n16509) );
  XOR U18557 ( .A(n16510), .B(n16511), .Z(n16498) );
  AND U18558 ( .A(n16512), .B(n16513), .Z(n16511) );
  XNOR U18559 ( .A(n16510), .B(n8257), .Z(n16513) );
  XNOR U18560 ( .A(n16506), .B(n16508), .Z(n8257) );
  NAND U18561 ( .A(n16514), .B(nreg[674]), .Z(n16508) );
  NAND U18562 ( .A(n12326), .B(nreg[674]), .Z(n16514) );
  XNOR U18563 ( .A(n16504), .B(n16515), .Z(n16506) );
  XOR U18564 ( .A(n16516), .B(n16517), .Z(n16504) );
  AND U18565 ( .A(n16518), .B(n16519), .Z(n16517) );
  XNOR U18566 ( .A(n16520), .B(n16516), .Z(n16519) );
  XOR U18567 ( .A(n16521), .B(nreg[674]), .Z(n16512) );
  IV U18568 ( .A(n16510), .Z(n16521) );
  XOR U18569 ( .A(n16522), .B(n16523), .Z(n16510) );
  AND U18570 ( .A(n16524), .B(n16525), .Z(n16523) );
  XNOR U18571 ( .A(n16522), .B(n8263), .Z(n16525) );
  XNOR U18572 ( .A(n16518), .B(n16520), .Z(n8263) );
  NAND U18573 ( .A(n16526), .B(nreg[673]), .Z(n16520) );
  NAND U18574 ( .A(n12326), .B(nreg[673]), .Z(n16526) );
  XNOR U18575 ( .A(n16516), .B(n16527), .Z(n16518) );
  XOR U18576 ( .A(n16528), .B(n16529), .Z(n16516) );
  AND U18577 ( .A(n16530), .B(n16531), .Z(n16529) );
  XNOR U18578 ( .A(n16532), .B(n16528), .Z(n16531) );
  XOR U18579 ( .A(n16533), .B(nreg[673]), .Z(n16524) );
  IV U18580 ( .A(n16522), .Z(n16533) );
  XOR U18581 ( .A(n16534), .B(n16535), .Z(n16522) );
  AND U18582 ( .A(n16536), .B(n16537), .Z(n16535) );
  XNOR U18583 ( .A(n16534), .B(n8269), .Z(n16537) );
  XNOR U18584 ( .A(n16530), .B(n16532), .Z(n8269) );
  NAND U18585 ( .A(n16538), .B(nreg[672]), .Z(n16532) );
  NAND U18586 ( .A(n12326), .B(nreg[672]), .Z(n16538) );
  XNOR U18587 ( .A(n16528), .B(n16539), .Z(n16530) );
  XOR U18588 ( .A(n16540), .B(n16541), .Z(n16528) );
  AND U18589 ( .A(n16542), .B(n16543), .Z(n16541) );
  XNOR U18590 ( .A(n16544), .B(n16540), .Z(n16543) );
  XOR U18591 ( .A(n16545), .B(nreg[672]), .Z(n16536) );
  IV U18592 ( .A(n16534), .Z(n16545) );
  XOR U18593 ( .A(n16546), .B(n16547), .Z(n16534) );
  AND U18594 ( .A(n16548), .B(n16549), .Z(n16547) );
  XNOR U18595 ( .A(n16546), .B(n8275), .Z(n16549) );
  XNOR U18596 ( .A(n16542), .B(n16544), .Z(n8275) );
  NAND U18597 ( .A(n16550), .B(nreg[671]), .Z(n16544) );
  NAND U18598 ( .A(n12326), .B(nreg[671]), .Z(n16550) );
  XNOR U18599 ( .A(n16540), .B(n16551), .Z(n16542) );
  XOR U18600 ( .A(n16552), .B(n16553), .Z(n16540) );
  AND U18601 ( .A(n16554), .B(n16555), .Z(n16553) );
  XNOR U18602 ( .A(n16556), .B(n16552), .Z(n16555) );
  XOR U18603 ( .A(n16557), .B(nreg[671]), .Z(n16548) );
  IV U18604 ( .A(n16546), .Z(n16557) );
  XOR U18605 ( .A(n16558), .B(n16559), .Z(n16546) );
  AND U18606 ( .A(n16560), .B(n16561), .Z(n16559) );
  XNOR U18607 ( .A(n16558), .B(n8281), .Z(n16561) );
  XNOR U18608 ( .A(n16554), .B(n16556), .Z(n8281) );
  NAND U18609 ( .A(n16562), .B(nreg[670]), .Z(n16556) );
  NAND U18610 ( .A(n12326), .B(nreg[670]), .Z(n16562) );
  XNOR U18611 ( .A(n16552), .B(n16563), .Z(n16554) );
  XOR U18612 ( .A(n16564), .B(n16565), .Z(n16552) );
  AND U18613 ( .A(n16566), .B(n16567), .Z(n16565) );
  XNOR U18614 ( .A(n16568), .B(n16564), .Z(n16567) );
  XOR U18615 ( .A(n16569), .B(nreg[670]), .Z(n16560) );
  IV U18616 ( .A(n16558), .Z(n16569) );
  XOR U18617 ( .A(n16570), .B(n16571), .Z(n16558) );
  AND U18618 ( .A(n16572), .B(n16573), .Z(n16571) );
  XNOR U18619 ( .A(n16570), .B(n8287), .Z(n16573) );
  XNOR U18620 ( .A(n16566), .B(n16568), .Z(n8287) );
  NAND U18621 ( .A(n16574), .B(nreg[669]), .Z(n16568) );
  NAND U18622 ( .A(n12326), .B(nreg[669]), .Z(n16574) );
  XNOR U18623 ( .A(n16564), .B(n16575), .Z(n16566) );
  XOR U18624 ( .A(n16576), .B(n16577), .Z(n16564) );
  AND U18625 ( .A(n16578), .B(n16579), .Z(n16577) );
  XNOR U18626 ( .A(n16580), .B(n16576), .Z(n16579) );
  XOR U18627 ( .A(n16581), .B(nreg[669]), .Z(n16572) );
  IV U18628 ( .A(n16570), .Z(n16581) );
  XOR U18629 ( .A(n16582), .B(n16583), .Z(n16570) );
  AND U18630 ( .A(n16584), .B(n16585), .Z(n16583) );
  XNOR U18631 ( .A(n16582), .B(n8293), .Z(n16585) );
  XNOR U18632 ( .A(n16578), .B(n16580), .Z(n8293) );
  NAND U18633 ( .A(n16586), .B(nreg[668]), .Z(n16580) );
  NAND U18634 ( .A(n12326), .B(nreg[668]), .Z(n16586) );
  XNOR U18635 ( .A(n16576), .B(n16587), .Z(n16578) );
  XOR U18636 ( .A(n16588), .B(n16589), .Z(n16576) );
  AND U18637 ( .A(n16590), .B(n16591), .Z(n16589) );
  XNOR U18638 ( .A(n16592), .B(n16588), .Z(n16591) );
  XOR U18639 ( .A(n16593), .B(nreg[668]), .Z(n16584) );
  IV U18640 ( .A(n16582), .Z(n16593) );
  XOR U18641 ( .A(n16594), .B(n16595), .Z(n16582) );
  AND U18642 ( .A(n16596), .B(n16597), .Z(n16595) );
  XNOR U18643 ( .A(n16594), .B(n8299), .Z(n16597) );
  XNOR U18644 ( .A(n16590), .B(n16592), .Z(n8299) );
  NAND U18645 ( .A(n16598), .B(nreg[667]), .Z(n16592) );
  NAND U18646 ( .A(n12326), .B(nreg[667]), .Z(n16598) );
  XNOR U18647 ( .A(n16588), .B(n16599), .Z(n16590) );
  XOR U18648 ( .A(n16600), .B(n16601), .Z(n16588) );
  AND U18649 ( .A(n16602), .B(n16603), .Z(n16601) );
  XNOR U18650 ( .A(n16604), .B(n16600), .Z(n16603) );
  XOR U18651 ( .A(n16605), .B(nreg[667]), .Z(n16596) );
  IV U18652 ( .A(n16594), .Z(n16605) );
  XOR U18653 ( .A(n16606), .B(n16607), .Z(n16594) );
  AND U18654 ( .A(n16608), .B(n16609), .Z(n16607) );
  XNOR U18655 ( .A(n16606), .B(n8305), .Z(n16609) );
  XNOR U18656 ( .A(n16602), .B(n16604), .Z(n8305) );
  NAND U18657 ( .A(n16610), .B(nreg[666]), .Z(n16604) );
  NAND U18658 ( .A(n12326), .B(nreg[666]), .Z(n16610) );
  XNOR U18659 ( .A(n16600), .B(n16611), .Z(n16602) );
  XOR U18660 ( .A(n16612), .B(n16613), .Z(n16600) );
  AND U18661 ( .A(n16614), .B(n16615), .Z(n16613) );
  XNOR U18662 ( .A(n16616), .B(n16612), .Z(n16615) );
  XOR U18663 ( .A(n16617), .B(nreg[666]), .Z(n16608) );
  IV U18664 ( .A(n16606), .Z(n16617) );
  XOR U18665 ( .A(n16618), .B(n16619), .Z(n16606) );
  AND U18666 ( .A(n16620), .B(n16621), .Z(n16619) );
  XNOR U18667 ( .A(n16618), .B(n8311), .Z(n16621) );
  XNOR U18668 ( .A(n16614), .B(n16616), .Z(n8311) );
  NAND U18669 ( .A(n16622), .B(nreg[665]), .Z(n16616) );
  NAND U18670 ( .A(n12326), .B(nreg[665]), .Z(n16622) );
  XNOR U18671 ( .A(n16612), .B(n16623), .Z(n16614) );
  XOR U18672 ( .A(n16624), .B(n16625), .Z(n16612) );
  AND U18673 ( .A(n16626), .B(n16627), .Z(n16625) );
  XNOR U18674 ( .A(n16628), .B(n16624), .Z(n16627) );
  XOR U18675 ( .A(n16629), .B(nreg[665]), .Z(n16620) );
  IV U18676 ( .A(n16618), .Z(n16629) );
  XOR U18677 ( .A(n16630), .B(n16631), .Z(n16618) );
  AND U18678 ( .A(n16632), .B(n16633), .Z(n16631) );
  XNOR U18679 ( .A(n16630), .B(n8317), .Z(n16633) );
  XNOR U18680 ( .A(n16626), .B(n16628), .Z(n8317) );
  NAND U18681 ( .A(n16634), .B(nreg[664]), .Z(n16628) );
  NAND U18682 ( .A(n12326), .B(nreg[664]), .Z(n16634) );
  XNOR U18683 ( .A(n16624), .B(n16635), .Z(n16626) );
  XOR U18684 ( .A(n16636), .B(n16637), .Z(n16624) );
  AND U18685 ( .A(n16638), .B(n16639), .Z(n16637) );
  XNOR U18686 ( .A(n16640), .B(n16636), .Z(n16639) );
  XOR U18687 ( .A(n16641), .B(nreg[664]), .Z(n16632) );
  IV U18688 ( .A(n16630), .Z(n16641) );
  XOR U18689 ( .A(n16642), .B(n16643), .Z(n16630) );
  AND U18690 ( .A(n16644), .B(n16645), .Z(n16643) );
  XNOR U18691 ( .A(n16642), .B(n8323), .Z(n16645) );
  XNOR U18692 ( .A(n16638), .B(n16640), .Z(n8323) );
  NAND U18693 ( .A(n16646), .B(nreg[663]), .Z(n16640) );
  NAND U18694 ( .A(n12326), .B(nreg[663]), .Z(n16646) );
  XNOR U18695 ( .A(n16636), .B(n16647), .Z(n16638) );
  XOR U18696 ( .A(n16648), .B(n16649), .Z(n16636) );
  AND U18697 ( .A(n16650), .B(n16651), .Z(n16649) );
  XNOR U18698 ( .A(n16652), .B(n16648), .Z(n16651) );
  XOR U18699 ( .A(n16653), .B(nreg[663]), .Z(n16644) );
  IV U18700 ( .A(n16642), .Z(n16653) );
  XOR U18701 ( .A(n16654), .B(n16655), .Z(n16642) );
  AND U18702 ( .A(n16656), .B(n16657), .Z(n16655) );
  XNOR U18703 ( .A(n16654), .B(n8329), .Z(n16657) );
  XNOR U18704 ( .A(n16650), .B(n16652), .Z(n8329) );
  NAND U18705 ( .A(n16658), .B(nreg[662]), .Z(n16652) );
  NAND U18706 ( .A(n12326), .B(nreg[662]), .Z(n16658) );
  XNOR U18707 ( .A(n16648), .B(n16659), .Z(n16650) );
  XOR U18708 ( .A(n16660), .B(n16661), .Z(n16648) );
  AND U18709 ( .A(n16662), .B(n16663), .Z(n16661) );
  XNOR U18710 ( .A(n16664), .B(n16660), .Z(n16663) );
  XOR U18711 ( .A(n16665), .B(nreg[662]), .Z(n16656) );
  IV U18712 ( .A(n16654), .Z(n16665) );
  XOR U18713 ( .A(n16666), .B(n16667), .Z(n16654) );
  AND U18714 ( .A(n16668), .B(n16669), .Z(n16667) );
  XNOR U18715 ( .A(n16666), .B(n8335), .Z(n16669) );
  XNOR U18716 ( .A(n16662), .B(n16664), .Z(n8335) );
  NAND U18717 ( .A(n16670), .B(nreg[661]), .Z(n16664) );
  NAND U18718 ( .A(n12326), .B(nreg[661]), .Z(n16670) );
  XNOR U18719 ( .A(n16660), .B(n16671), .Z(n16662) );
  XOR U18720 ( .A(n16672), .B(n16673), .Z(n16660) );
  AND U18721 ( .A(n16674), .B(n16675), .Z(n16673) );
  XNOR U18722 ( .A(n16676), .B(n16672), .Z(n16675) );
  XOR U18723 ( .A(n16677), .B(nreg[661]), .Z(n16668) );
  IV U18724 ( .A(n16666), .Z(n16677) );
  XOR U18725 ( .A(n16678), .B(n16679), .Z(n16666) );
  AND U18726 ( .A(n16680), .B(n16681), .Z(n16679) );
  XNOR U18727 ( .A(n16678), .B(n8341), .Z(n16681) );
  XNOR U18728 ( .A(n16674), .B(n16676), .Z(n8341) );
  NAND U18729 ( .A(n16682), .B(nreg[660]), .Z(n16676) );
  NAND U18730 ( .A(n12326), .B(nreg[660]), .Z(n16682) );
  XNOR U18731 ( .A(n16672), .B(n16683), .Z(n16674) );
  XOR U18732 ( .A(n16684), .B(n16685), .Z(n16672) );
  AND U18733 ( .A(n16686), .B(n16687), .Z(n16685) );
  XNOR U18734 ( .A(n16688), .B(n16684), .Z(n16687) );
  XOR U18735 ( .A(n16689), .B(nreg[660]), .Z(n16680) );
  IV U18736 ( .A(n16678), .Z(n16689) );
  XOR U18737 ( .A(n16690), .B(n16691), .Z(n16678) );
  AND U18738 ( .A(n16692), .B(n16693), .Z(n16691) );
  XNOR U18739 ( .A(n16690), .B(n8347), .Z(n16693) );
  XNOR U18740 ( .A(n16686), .B(n16688), .Z(n8347) );
  NAND U18741 ( .A(n16694), .B(nreg[659]), .Z(n16688) );
  NAND U18742 ( .A(n12326), .B(nreg[659]), .Z(n16694) );
  XNOR U18743 ( .A(n16684), .B(n16695), .Z(n16686) );
  XOR U18744 ( .A(n16696), .B(n16697), .Z(n16684) );
  AND U18745 ( .A(n16698), .B(n16699), .Z(n16697) );
  XNOR U18746 ( .A(n16700), .B(n16696), .Z(n16699) );
  XOR U18747 ( .A(n16701), .B(nreg[659]), .Z(n16692) );
  IV U18748 ( .A(n16690), .Z(n16701) );
  XOR U18749 ( .A(n16702), .B(n16703), .Z(n16690) );
  AND U18750 ( .A(n16704), .B(n16705), .Z(n16703) );
  XNOR U18751 ( .A(n16702), .B(n8353), .Z(n16705) );
  XNOR U18752 ( .A(n16698), .B(n16700), .Z(n8353) );
  NAND U18753 ( .A(n16706), .B(nreg[658]), .Z(n16700) );
  NAND U18754 ( .A(n12326), .B(nreg[658]), .Z(n16706) );
  XNOR U18755 ( .A(n16696), .B(n16707), .Z(n16698) );
  XOR U18756 ( .A(n16708), .B(n16709), .Z(n16696) );
  AND U18757 ( .A(n16710), .B(n16711), .Z(n16709) );
  XNOR U18758 ( .A(n16712), .B(n16708), .Z(n16711) );
  XOR U18759 ( .A(n16713), .B(nreg[658]), .Z(n16704) );
  IV U18760 ( .A(n16702), .Z(n16713) );
  XOR U18761 ( .A(n16714), .B(n16715), .Z(n16702) );
  AND U18762 ( .A(n16716), .B(n16717), .Z(n16715) );
  XNOR U18763 ( .A(n16714), .B(n8359), .Z(n16717) );
  XNOR U18764 ( .A(n16710), .B(n16712), .Z(n8359) );
  NAND U18765 ( .A(n16718), .B(nreg[657]), .Z(n16712) );
  NAND U18766 ( .A(n12326), .B(nreg[657]), .Z(n16718) );
  XNOR U18767 ( .A(n16708), .B(n16719), .Z(n16710) );
  XOR U18768 ( .A(n16720), .B(n16721), .Z(n16708) );
  AND U18769 ( .A(n16722), .B(n16723), .Z(n16721) );
  XNOR U18770 ( .A(n16724), .B(n16720), .Z(n16723) );
  XOR U18771 ( .A(n16725), .B(nreg[657]), .Z(n16716) );
  IV U18772 ( .A(n16714), .Z(n16725) );
  XOR U18773 ( .A(n16726), .B(n16727), .Z(n16714) );
  AND U18774 ( .A(n16728), .B(n16729), .Z(n16727) );
  XNOR U18775 ( .A(n16726), .B(n8365), .Z(n16729) );
  XNOR U18776 ( .A(n16722), .B(n16724), .Z(n8365) );
  NAND U18777 ( .A(n16730), .B(nreg[656]), .Z(n16724) );
  NAND U18778 ( .A(n12326), .B(nreg[656]), .Z(n16730) );
  XNOR U18779 ( .A(n16720), .B(n16731), .Z(n16722) );
  XOR U18780 ( .A(n16732), .B(n16733), .Z(n16720) );
  AND U18781 ( .A(n16734), .B(n16735), .Z(n16733) );
  XNOR U18782 ( .A(n16736), .B(n16732), .Z(n16735) );
  XOR U18783 ( .A(n16737), .B(nreg[656]), .Z(n16728) );
  IV U18784 ( .A(n16726), .Z(n16737) );
  XOR U18785 ( .A(n16738), .B(n16739), .Z(n16726) );
  AND U18786 ( .A(n16740), .B(n16741), .Z(n16739) );
  XNOR U18787 ( .A(n16738), .B(n8371), .Z(n16741) );
  XNOR U18788 ( .A(n16734), .B(n16736), .Z(n8371) );
  NAND U18789 ( .A(n16742), .B(nreg[655]), .Z(n16736) );
  NAND U18790 ( .A(n12326), .B(nreg[655]), .Z(n16742) );
  XNOR U18791 ( .A(n16732), .B(n16743), .Z(n16734) );
  XOR U18792 ( .A(n16744), .B(n16745), .Z(n16732) );
  AND U18793 ( .A(n16746), .B(n16747), .Z(n16745) );
  XNOR U18794 ( .A(n16748), .B(n16744), .Z(n16747) );
  XOR U18795 ( .A(n16749), .B(nreg[655]), .Z(n16740) );
  IV U18796 ( .A(n16738), .Z(n16749) );
  XOR U18797 ( .A(n16750), .B(n16751), .Z(n16738) );
  AND U18798 ( .A(n16752), .B(n16753), .Z(n16751) );
  XNOR U18799 ( .A(n16750), .B(n8377), .Z(n16753) );
  XNOR U18800 ( .A(n16746), .B(n16748), .Z(n8377) );
  NAND U18801 ( .A(n16754), .B(nreg[654]), .Z(n16748) );
  NAND U18802 ( .A(n12326), .B(nreg[654]), .Z(n16754) );
  XNOR U18803 ( .A(n16744), .B(n16755), .Z(n16746) );
  XOR U18804 ( .A(n16756), .B(n16757), .Z(n16744) );
  AND U18805 ( .A(n16758), .B(n16759), .Z(n16757) );
  XNOR U18806 ( .A(n16760), .B(n16756), .Z(n16759) );
  XOR U18807 ( .A(n16761), .B(nreg[654]), .Z(n16752) );
  IV U18808 ( .A(n16750), .Z(n16761) );
  XOR U18809 ( .A(n16762), .B(n16763), .Z(n16750) );
  AND U18810 ( .A(n16764), .B(n16765), .Z(n16763) );
  XNOR U18811 ( .A(n16762), .B(n8383), .Z(n16765) );
  XNOR U18812 ( .A(n16758), .B(n16760), .Z(n8383) );
  NAND U18813 ( .A(n16766), .B(nreg[653]), .Z(n16760) );
  NAND U18814 ( .A(n12326), .B(nreg[653]), .Z(n16766) );
  XNOR U18815 ( .A(n16756), .B(n16767), .Z(n16758) );
  XOR U18816 ( .A(n16768), .B(n16769), .Z(n16756) );
  AND U18817 ( .A(n16770), .B(n16771), .Z(n16769) );
  XNOR U18818 ( .A(n16772), .B(n16768), .Z(n16771) );
  XOR U18819 ( .A(n16773), .B(nreg[653]), .Z(n16764) );
  IV U18820 ( .A(n16762), .Z(n16773) );
  XOR U18821 ( .A(n16774), .B(n16775), .Z(n16762) );
  AND U18822 ( .A(n16776), .B(n16777), .Z(n16775) );
  XNOR U18823 ( .A(n16774), .B(n8389), .Z(n16777) );
  XNOR U18824 ( .A(n16770), .B(n16772), .Z(n8389) );
  NAND U18825 ( .A(n16778), .B(nreg[652]), .Z(n16772) );
  NAND U18826 ( .A(n12326), .B(nreg[652]), .Z(n16778) );
  XNOR U18827 ( .A(n16768), .B(n16779), .Z(n16770) );
  XOR U18828 ( .A(n16780), .B(n16781), .Z(n16768) );
  AND U18829 ( .A(n16782), .B(n16783), .Z(n16781) );
  XNOR U18830 ( .A(n16784), .B(n16780), .Z(n16783) );
  XOR U18831 ( .A(n16785), .B(nreg[652]), .Z(n16776) );
  IV U18832 ( .A(n16774), .Z(n16785) );
  XOR U18833 ( .A(n16786), .B(n16787), .Z(n16774) );
  AND U18834 ( .A(n16788), .B(n16789), .Z(n16787) );
  XNOR U18835 ( .A(n16786), .B(n8395), .Z(n16789) );
  XNOR U18836 ( .A(n16782), .B(n16784), .Z(n8395) );
  NAND U18837 ( .A(n16790), .B(nreg[651]), .Z(n16784) );
  NAND U18838 ( .A(n12326), .B(nreg[651]), .Z(n16790) );
  XNOR U18839 ( .A(n16780), .B(n16791), .Z(n16782) );
  XOR U18840 ( .A(n16792), .B(n16793), .Z(n16780) );
  AND U18841 ( .A(n16794), .B(n16795), .Z(n16793) );
  XNOR U18842 ( .A(n16796), .B(n16792), .Z(n16795) );
  XOR U18843 ( .A(n16797), .B(nreg[651]), .Z(n16788) );
  IV U18844 ( .A(n16786), .Z(n16797) );
  XOR U18845 ( .A(n16798), .B(n16799), .Z(n16786) );
  AND U18846 ( .A(n16800), .B(n16801), .Z(n16799) );
  XNOR U18847 ( .A(n16798), .B(n8401), .Z(n16801) );
  XNOR U18848 ( .A(n16794), .B(n16796), .Z(n8401) );
  NAND U18849 ( .A(n16802), .B(nreg[650]), .Z(n16796) );
  NAND U18850 ( .A(n12326), .B(nreg[650]), .Z(n16802) );
  XNOR U18851 ( .A(n16792), .B(n16803), .Z(n16794) );
  XOR U18852 ( .A(n16804), .B(n16805), .Z(n16792) );
  AND U18853 ( .A(n16806), .B(n16807), .Z(n16805) );
  XNOR U18854 ( .A(n16808), .B(n16804), .Z(n16807) );
  XOR U18855 ( .A(n16809), .B(nreg[650]), .Z(n16800) );
  IV U18856 ( .A(n16798), .Z(n16809) );
  XOR U18857 ( .A(n16810), .B(n16811), .Z(n16798) );
  AND U18858 ( .A(n16812), .B(n16813), .Z(n16811) );
  XNOR U18859 ( .A(n16810), .B(n8407), .Z(n16813) );
  XNOR U18860 ( .A(n16806), .B(n16808), .Z(n8407) );
  NAND U18861 ( .A(n16814), .B(nreg[649]), .Z(n16808) );
  NAND U18862 ( .A(n12326), .B(nreg[649]), .Z(n16814) );
  XNOR U18863 ( .A(n16804), .B(n16815), .Z(n16806) );
  XOR U18864 ( .A(n16816), .B(n16817), .Z(n16804) );
  AND U18865 ( .A(n16818), .B(n16819), .Z(n16817) );
  XNOR U18866 ( .A(n16820), .B(n16816), .Z(n16819) );
  XOR U18867 ( .A(n16821), .B(nreg[649]), .Z(n16812) );
  IV U18868 ( .A(n16810), .Z(n16821) );
  XOR U18869 ( .A(n16822), .B(n16823), .Z(n16810) );
  AND U18870 ( .A(n16824), .B(n16825), .Z(n16823) );
  XNOR U18871 ( .A(n16822), .B(n8413), .Z(n16825) );
  XNOR U18872 ( .A(n16818), .B(n16820), .Z(n8413) );
  NAND U18873 ( .A(n16826), .B(nreg[648]), .Z(n16820) );
  NAND U18874 ( .A(n12326), .B(nreg[648]), .Z(n16826) );
  XNOR U18875 ( .A(n16816), .B(n16827), .Z(n16818) );
  XOR U18876 ( .A(n16828), .B(n16829), .Z(n16816) );
  AND U18877 ( .A(n16830), .B(n16831), .Z(n16829) );
  XNOR U18878 ( .A(n16832), .B(n16828), .Z(n16831) );
  XOR U18879 ( .A(n16833), .B(nreg[648]), .Z(n16824) );
  IV U18880 ( .A(n16822), .Z(n16833) );
  XOR U18881 ( .A(n16834), .B(n16835), .Z(n16822) );
  AND U18882 ( .A(n16836), .B(n16837), .Z(n16835) );
  XNOR U18883 ( .A(n16834), .B(n8419), .Z(n16837) );
  XNOR U18884 ( .A(n16830), .B(n16832), .Z(n8419) );
  NAND U18885 ( .A(n16838), .B(nreg[647]), .Z(n16832) );
  NAND U18886 ( .A(n12326), .B(nreg[647]), .Z(n16838) );
  XNOR U18887 ( .A(n16828), .B(n16839), .Z(n16830) );
  XOR U18888 ( .A(n16840), .B(n16841), .Z(n16828) );
  AND U18889 ( .A(n16842), .B(n16843), .Z(n16841) );
  XNOR U18890 ( .A(n16844), .B(n16840), .Z(n16843) );
  XOR U18891 ( .A(n16845), .B(nreg[647]), .Z(n16836) );
  IV U18892 ( .A(n16834), .Z(n16845) );
  XOR U18893 ( .A(n16846), .B(n16847), .Z(n16834) );
  AND U18894 ( .A(n16848), .B(n16849), .Z(n16847) );
  XNOR U18895 ( .A(n16846), .B(n8425), .Z(n16849) );
  XNOR U18896 ( .A(n16842), .B(n16844), .Z(n8425) );
  NAND U18897 ( .A(n16850), .B(nreg[646]), .Z(n16844) );
  NAND U18898 ( .A(n12326), .B(nreg[646]), .Z(n16850) );
  XNOR U18899 ( .A(n16840), .B(n16851), .Z(n16842) );
  XOR U18900 ( .A(n16852), .B(n16853), .Z(n16840) );
  AND U18901 ( .A(n16854), .B(n16855), .Z(n16853) );
  XNOR U18902 ( .A(n16856), .B(n16852), .Z(n16855) );
  XOR U18903 ( .A(n16857), .B(nreg[646]), .Z(n16848) );
  IV U18904 ( .A(n16846), .Z(n16857) );
  XOR U18905 ( .A(n16858), .B(n16859), .Z(n16846) );
  AND U18906 ( .A(n16860), .B(n16861), .Z(n16859) );
  XNOR U18907 ( .A(n16858), .B(n8431), .Z(n16861) );
  XNOR U18908 ( .A(n16854), .B(n16856), .Z(n8431) );
  NAND U18909 ( .A(n16862), .B(nreg[645]), .Z(n16856) );
  NAND U18910 ( .A(n12326), .B(nreg[645]), .Z(n16862) );
  XNOR U18911 ( .A(n16852), .B(n16863), .Z(n16854) );
  XOR U18912 ( .A(n16864), .B(n16865), .Z(n16852) );
  AND U18913 ( .A(n16866), .B(n16867), .Z(n16865) );
  XNOR U18914 ( .A(n16868), .B(n16864), .Z(n16867) );
  XOR U18915 ( .A(n16869), .B(nreg[645]), .Z(n16860) );
  IV U18916 ( .A(n16858), .Z(n16869) );
  XOR U18917 ( .A(n16870), .B(n16871), .Z(n16858) );
  AND U18918 ( .A(n16872), .B(n16873), .Z(n16871) );
  XNOR U18919 ( .A(n16870), .B(n8437), .Z(n16873) );
  XNOR U18920 ( .A(n16866), .B(n16868), .Z(n8437) );
  NAND U18921 ( .A(n16874), .B(nreg[644]), .Z(n16868) );
  NAND U18922 ( .A(n12326), .B(nreg[644]), .Z(n16874) );
  XNOR U18923 ( .A(n16864), .B(n16875), .Z(n16866) );
  XOR U18924 ( .A(n16876), .B(n16877), .Z(n16864) );
  AND U18925 ( .A(n16878), .B(n16879), .Z(n16877) );
  XNOR U18926 ( .A(n16880), .B(n16876), .Z(n16879) );
  XOR U18927 ( .A(n16881), .B(nreg[644]), .Z(n16872) );
  IV U18928 ( .A(n16870), .Z(n16881) );
  XOR U18929 ( .A(n16882), .B(n16883), .Z(n16870) );
  AND U18930 ( .A(n16884), .B(n16885), .Z(n16883) );
  XNOR U18931 ( .A(n16882), .B(n8443), .Z(n16885) );
  XNOR U18932 ( .A(n16878), .B(n16880), .Z(n8443) );
  NAND U18933 ( .A(n16886), .B(nreg[643]), .Z(n16880) );
  NAND U18934 ( .A(n12326), .B(nreg[643]), .Z(n16886) );
  XNOR U18935 ( .A(n16876), .B(n16887), .Z(n16878) );
  XOR U18936 ( .A(n16888), .B(n16889), .Z(n16876) );
  AND U18937 ( .A(n16890), .B(n16891), .Z(n16889) );
  XNOR U18938 ( .A(n16892), .B(n16888), .Z(n16891) );
  XOR U18939 ( .A(n16893), .B(nreg[643]), .Z(n16884) );
  IV U18940 ( .A(n16882), .Z(n16893) );
  XOR U18941 ( .A(n16894), .B(n16895), .Z(n16882) );
  AND U18942 ( .A(n16896), .B(n16897), .Z(n16895) );
  XNOR U18943 ( .A(n16894), .B(n8449), .Z(n16897) );
  XNOR U18944 ( .A(n16890), .B(n16892), .Z(n8449) );
  NAND U18945 ( .A(n16898), .B(nreg[642]), .Z(n16892) );
  NAND U18946 ( .A(n12326), .B(nreg[642]), .Z(n16898) );
  XNOR U18947 ( .A(n16888), .B(n16899), .Z(n16890) );
  XOR U18948 ( .A(n16900), .B(n16901), .Z(n16888) );
  AND U18949 ( .A(n16902), .B(n16903), .Z(n16901) );
  XNOR U18950 ( .A(n16904), .B(n16900), .Z(n16903) );
  XOR U18951 ( .A(n16905), .B(nreg[642]), .Z(n16896) );
  IV U18952 ( .A(n16894), .Z(n16905) );
  XOR U18953 ( .A(n16906), .B(n16907), .Z(n16894) );
  AND U18954 ( .A(n16908), .B(n16909), .Z(n16907) );
  XNOR U18955 ( .A(n16906), .B(n8455), .Z(n16909) );
  XNOR U18956 ( .A(n16902), .B(n16904), .Z(n8455) );
  NAND U18957 ( .A(n16910), .B(nreg[641]), .Z(n16904) );
  NAND U18958 ( .A(n12326), .B(nreg[641]), .Z(n16910) );
  XNOR U18959 ( .A(n16900), .B(n16911), .Z(n16902) );
  XOR U18960 ( .A(n16912), .B(n16913), .Z(n16900) );
  AND U18961 ( .A(n16914), .B(n16915), .Z(n16913) );
  XNOR U18962 ( .A(n16916), .B(n16912), .Z(n16915) );
  XOR U18963 ( .A(n16917), .B(nreg[641]), .Z(n16908) );
  IV U18964 ( .A(n16906), .Z(n16917) );
  XOR U18965 ( .A(n16918), .B(n16919), .Z(n16906) );
  AND U18966 ( .A(n16920), .B(n16921), .Z(n16919) );
  XNOR U18967 ( .A(n16918), .B(n8461), .Z(n16921) );
  XNOR U18968 ( .A(n16914), .B(n16916), .Z(n8461) );
  NAND U18969 ( .A(n16922), .B(nreg[640]), .Z(n16916) );
  NAND U18970 ( .A(n12326), .B(nreg[640]), .Z(n16922) );
  XNOR U18971 ( .A(n16912), .B(n16923), .Z(n16914) );
  XOR U18972 ( .A(n16924), .B(n16925), .Z(n16912) );
  AND U18973 ( .A(n16926), .B(n16927), .Z(n16925) );
  XNOR U18974 ( .A(n16928), .B(n16924), .Z(n16927) );
  XOR U18975 ( .A(n16929), .B(nreg[640]), .Z(n16920) );
  IV U18976 ( .A(n16918), .Z(n16929) );
  XOR U18977 ( .A(n16930), .B(n16931), .Z(n16918) );
  AND U18978 ( .A(n16932), .B(n16933), .Z(n16931) );
  XNOR U18979 ( .A(n16930), .B(n8467), .Z(n16933) );
  XNOR U18980 ( .A(n16926), .B(n16928), .Z(n8467) );
  NAND U18981 ( .A(n16934), .B(nreg[639]), .Z(n16928) );
  NAND U18982 ( .A(n12326), .B(nreg[639]), .Z(n16934) );
  XNOR U18983 ( .A(n16924), .B(n16935), .Z(n16926) );
  XOR U18984 ( .A(n16936), .B(n16937), .Z(n16924) );
  AND U18985 ( .A(n16938), .B(n16939), .Z(n16937) );
  XNOR U18986 ( .A(n16940), .B(n16936), .Z(n16939) );
  XOR U18987 ( .A(n16941), .B(nreg[639]), .Z(n16932) );
  IV U18988 ( .A(n16930), .Z(n16941) );
  XOR U18989 ( .A(n16942), .B(n16943), .Z(n16930) );
  AND U18990 ( .A(n16944), .B(n16945), .Z(n16943) );
  XNOR U18991 ( .A(n16942), .B(n8473), .Z(n16945) );
  XNOR U18992 ( .A(n16938), .B(n16940), .Z(n8473) );
  NAND U18993 ( .A(n16946), .B(nreg[638]), .Z(n16940) );
  NAND U18994 ( .A(n12326), .B(nreg[638]), .Z(n16946) );
  XNOR U18995 ( .A(n16936), .B(n16947), .Z(n16938) );
  XOR U18996 ( .A(n16948), .B(n16949), .Z(n16936) );
  AND U18997 ( .A(n16950), .B(n16951), .Z(n16949) );
  XNOR U18998 ( .A(n16952), .B(n16948), .Z(n16951) );
  XOR U18999 ( .A(n16953), .B(nreg[638]), .Z(n16944) );
  IV U19000 ( .A(n16942), .Z(n16953) );
  XOR U19001 ( .A(n16954), .B(n16955), .Z(n16942) );
  AND U19002 ( .A(n16956), .B(n16957), .Z(n16955) );
  XNOR U19003 ( .A(n16954), .B(n8479), .Z(n16957) );
  XNOR U19004 ( .A(n16950), .B(n16952), .Z(n8479) );
  NAND U19005 ( .A(n16958), .B(nreg[637]), .Z(n16952) );
  NAND U19006 ( .A(n12326), .B(nreg[637]), .Z(n16958) );
  XNOR U19007 ( .A(n16948), .B(n16959), .Z(n16950) );
  XOR U19008 ( .A(n16960), .B(n16961), .Z(n16948) );
  AND U19009 ( .A(n16962), .B(n16963), .Z(n16961) );
  XNOR U19010 ( .A(n16964), .B(n16960), .Z(n16963) );
  XOR U19011 ( .A(n16965), .B(nreg[637]), .Z(n16956) );
  IV U19012 ( .A(n16954), .Z(n16965) );
  XOR U19013 ( .A(n16966), .B(n16967), .Z(n16954) );
  AND U19014 ( .A(n16968), .B(n16969), .Z(n16967) );
  XNOR U19015 ( .A(n16966), .B(n8485), .Z(n16969) );
  XNOR U19016 ( .A(n16962), .B(n16964), .Z(n8485) );
  NAND U19017 ( .A(n16970), .B(nreg[636]), .Z(n16964) );
  NAND U19018 ( .A(n12326), .B(nreg[636]), .Z(n16970) );
  XNOR U19019 ( .A(n16960), .B(n16971), .Z(n16962) );
  XOR U19020 ( .A(n16972), .B(n16973), .Z(n16960) );
  AND U19021 ( .A(n16974), .B(n16975), .Z(n16973) );
  XNOR U19022 ( .A(n16976), .B(n16972), .Z(n16975) );
  XOR U19023 ( .A(n16977), .B(nreg[636]), .Z(n16968) );
  IV U19024 ( .A(n16966), .Z(n16977) );
  XOR U19025 ( .A(n16978), .B(n16979), .Z(n16966) );
  AND U19026 ( .A(n16980), .B(n16981), .Z(n16979) );
  XNOR U19027 ( .A(n16978), .B(n8491), .Z(n16981) );
  XNOR U19028 ( .A(n16974), .B(n16976), .Z(n8491) );
  NAND U19029 ( .A(n16982), .B(nreg[635]), .Z(n16976) );
  NAND U19030 ( .A(n12326), .B(nreg[635]), .Z(n16982) );
  XNOR U19031 ( .A(n16972), .B(n16983), .Z(n16974) );
  XOR U19032 ( .A(n16984), .B(n16985), .Z(n16972) );
  AND U19033 ( .A(n16986), .B(n16987), .Z(n16985) );
  XNOR U19034 ( .A(n16988), .B(n16984), .Z(n16987) );
  XOR U19035 ( .A(n16989), .B(nreg[635]), .Z(n16980) );
  IV U19036 ( .A(n16978), .Z(n16989) );
  XOR U19037 ( .A(n16990), .B(n16991), .Z(n16978) );
  AND U19038 ( .A(n16992), .B(n16993), .Z(n16991) );
  XNOR U19039 ( .A(n16990), .B(n8497), .Z(n16993) );
  XNOR U19040 ( .A(n16986), .B(n16988), .Z(n8497) );
  NAND U19041 ( .A(n16994), .B(nreg[634]), .Z(n16988) );
  NAND U19042 ( .A(n12326), .B(nreg[634]), .Z(n16994) );
  XNOR U19043 ( .A(n16984), .B(n16995), .Z(n16986) );
  XOR U19044 ( .A(n16996), .B(n16997), .Z(n16984) );
  AND U19045 ( .A(n16998), .B(n16999), .Z(n16997) );
  XNOR U19046 ( .A(n17000), .B(n16996), .Z(n16999) );
  XOR U19047 ( .A(n17001), .B(nreg[634]), .Z(n16992) );
  IV U19048 ( .A(n16990), .Z(n17001) );
  XOR U19049 ( .A(n17002), .B(n17003), .Z(n16990) );
  AND U19050 ( .A(n17004), .B(n17005), .Z(n17003) );
  XNOR U19051 ( .A(n17002), .B(n8503), .Z(n17005) );
  XNOR U19052 ( .A(n16998), .B(n17000), .Z(n8503) );
  NAND U19053 ( .A(n17006), .B(nreg[633]), .Z(n17000) );
  NAND U19054 ( .A(n12326), .B(nreg[633]), .Z(n17006) );
  XNOR U19055 ( .A(n16996), .B(n17007), .Z(n16998) );
  XOR U19056 ( .A(n17008), .B(n17009), .Z(n16996) );
  AND U19057 ( .A(n17010), .B(n17011), .Z(n17009) );
  XNOR U19058 ( .A(n17012), .B(n17008), .Z(n17011) );
  XOR U19059 ( .A(n17013), .B(nreg[633]), .Z(n17004) );
  IV U19060 ( .A(n17002), .Z(n17013) );
  XOR U19061 ( .A(n17014), .B(n17015), .Z(n17002) );
  AND U19062 ( .A(n17016), .B(n17017), .Z(n17015) );
  XNOR U19063 ( .A(n17014), .B(n8509), .Z(n17017) );
  XNOR U19064 ( .A(n17010), .B(n17012), .Z(n8509) );
  NAND U19065 ( .A(n17018), .B(nreg[632]), .Z(n17012) );
  NAND U19066 ( .A(n12326), .B(nreg[632]), .Z(n17018) );
  XNOR U19067 ( .A(n17008), .B(n17019), .Z(n17010) );
  XOR U19068 ( .A(n17020), .B(n17021), .Z(n17008) );
  AND U19069 ( .A(n17022), .B(n17023), .Z(n17021) );
  XNOR U19070 ( .A(n17024), .B(n17020), .Z(n17023) );
  XOR U19071 ( .A(n17025), .B(nreg[632]), .Z(n17016) );
  IV U19072 ( .A(n17014), .Z(n17025) );
  XOR U19073 ( .A(n17026), .B(n17027), .Z(n17014) );
  AND U19074 ( .A(n17028), .B(n17029), .Z(n17027) );
  XNOR U19075 ( .A(n17026), .B(n8515), .Z(n17029) );
  XNOR U19076 ( .A(n17022), .B(n17024), .Z(n8515) );
  NAND U19077 ( .A(n17030), .B(nreg[631]), .Z(n17024) );
  NAND U19078 ( .A(n12326), .B(nreg[631]), .Z(n17030) );
  XNOR U19079 ( .A(n17020), .B(n17031), .Z(n17022) );
  XOR U19080 ( .A(n17032), .B(n17033), .Z(n17020) );
  AND U19081 ( .A(n17034), .B(n17035), .Z(n17033) );
  XNOR U19082 ( .A(n17036), .B(n17032), .Z(n17035) );
  XOR U19083 ( .A(n17037), .B(nreg[631]), .Z(n17028) );
  IV U19084 ( .A(n17026), .Z(n17037) );
  XOR U19085 ( .A(n17038), .B(n17039), .Z(n17026) );
  AND U19086 ( .A(n17040), .B(n17041), .Z(n17039) );
  XNOR U19087 ( .A(n17038), .B(n8521), .Z(n17041) );
  XNOR U19088 ( .A(n17034), .B(n17036), .Z(n8521) );
  NAND U19089 ( .A(n17042), .B(nreg[630]), .Z(n17036) );
  NAND U19090 ( .A(n12326), .B(nreg[630]), .Z(n17042) );
  XNOR U19091 ( .A(n17032), .B(n17043), .Z(n17034) );
  XOR U19092 ( .A(n17044), .B(n17045), .Z(n17032) );
  AND U19093 ( .A(n17046), .B(n17047), .Z(n17045) );
  XNOR U19094 ( .A(n17048), .B(n17044), .Z(n17047) );
  XOR U19095 ( .A(n17049), .B(nreg[630]), .Z(n17040) );
  IV U19096 ( .A(n17038), .Z(n17049) );
  XOR U19097 ( .A(n17050), .B(n17051), .Z(n17038) );
  AND U19098 ( .A(n17052), .B(n17053), .Z(n17051) );
  XNOR U19099 ( .A(n17050), .B(n8527), .Z(n17053) );
  XNOR U19100 ( .A(n17046), .B(n17048), .Z(n8527) );
  NAND U19101 ( .A(n17054), .B(nreg[629]), .Z(n17048) );
  NAND U19102 ( .A(n12326), .B(nreg[629]), .Z(n17054) );
  XNOR U19103 ( .A(n17044), .B(n17055), .Z(n17046) );
  XOR U19104 ( .A(n17056), .B(n17057), .Z(n17044) );
  AND U19105 ( .A(n17058), .B(n17059), .Z(n17057) );
  XNOR U19106 ( .A(n17060), .B(n17056), .Z(n17059) );
  XOR U19107 ( .A(n17061), .B(nreg[629]), .Z(n17052) );
  IV U19108 ( .A(n17050), .Z(n17061) );
  XOR U19109 ( .A(n17062), .B(n17063), .Z(n17050) );
  AND U19110 ( .A(n17064), .B(n17065), .Z(n17063) );
  XNOR U19111 ( .A(n17062), .B(n8533), .Z(n17065) );
  XNOR U19112 ( .A(n17058), .B(n17060), .Z(n8533) );
  NAND U19113 ( .A(n17066), .B(nreg[628]), .Z(n17060) );
  NAND U19114 ( .A(n12326), .B(nreg[628]), .Z(n17066) );
  XNOR U19115 ( .A(n17056), .B(n17067), .Z(n17058) );
  XOR U19116 ( .A(n17068), .B(n17069), .Z(n17056) );
  AND U19117 ( .A(n17070), .B(n17071), .Z(n17069) );
  XNOR U19118 ( .A(n17072), .B(n17068), .Z(n17071) );
  XOR U19119 ( .A(n17073), .B(nreg[628]), .Z(n17064) );
  IV U19120 ( .A(n17062), .Z(n17073) );
  XOR U19121 ( .A(n17074), .B(n17075), .Z(n17062) );
  AND U19122 ( .A(n17076), .B(n17077), .Z(n17075) );
  XNOR U19123 ( .A(n17074), .B(n8539), .Z(n17077) );
  XNOR U19124 ( .A(n17070), .B(n17072), .Z(n8539) );
  NAND U19125 ( .A(n17078), .B(nreg[627]), .Z(n17072) );
  NAND U19126 ( .A(n12326), .B(nreg[627]), .Z(n17078) );
  XNOR U19127 ( .A(n17068), .B(n17079), .Z(n17070) );
  XOR U19128 ( .A(n17080), .B(n17081), .Z(n17068) );
  AND U19129 ( .A(n17082), .B(n17083), .Z(n17081) );
  XNOR U19130 ( .A(n17084), .B(n17080), .Z(n17083) );
  XOR U19131 ( .A(n17085), .B(nreg[627]), .Z(n17076) );
  IV U19132 ( .A(n17074), .Z(n17085) );
  XOR U19133 ( .A(n17086), .B(n17087), .Z(n17074) );
  AND U19134 ( .A(n17088), .B(n17089), .Z(n17087) );
  XNOR U19135 ( .A(n17086), .B(n8545), .Z(n17089) );
  XNOR U19136 ( .A(n17082), .B(n17084), .Z(n8545) );
  NAND U19137 ( .A(n17090), .B(nreg[626]), .Z(n17084) );
  NAND U19138 ( .A(n12326), .B(nreg[626]), .Z(n17090) );
  XNOR U19139 ( .A(n17080), .B(n17091), .Z(n17082) );
  XOR U19140 ( .A(n17092), .B(n17093), .Z(n17080) );
  AND U19141 ( .A(n17094), .B(n17095), .Z(n17093) );
  XNOR U19142 ( .A(n17096), .B(n17092), .Z(n17095) );
  XOR U19143 ( .A(n17097), .B(nreg[626]), .Z(n17088) );
  IV U19144 ( .A(n17086), .Z(n17097) );
  XOR U19145 ( .A(n17098), .B(n17099), .Z(n17086) );
  AND U19146 ( .A(n17100), .B(n17101), .Z(n17099) );
  XNOR U19147 ( .A(n17098), .B(n8551), .Z(n17101) );
  XNOR U19148 ( .A(n17094), .B(n17096), .Z(n8551) );
  NAND U19149 ( .A(n17102), .B(nreg[625]), .Z(n17096) );
  NAND U19150 ( .A(n12326), .B(nreg[625]), .Z(n17102) );
  XNOR U19151 ( .A(n17092), .B(n17103), .Z(n17094) );
  XOR U19152 ( .A(n17104), .B(n17105), .Z(n17092) );
  AND U19153 ( .A(n17106), .B(n17107), .Z(n17105) );
  XNOR U19154 ( .A(n17108), .B(n17104), .Z(n17107) );
  XOR U19155 ( .A(n17109), .B(nreg[625]), .Z(n17100) );
  IV U19156 ( .A(n17098), .Z(n17109) );
  XOR U19157 ( .A(n17110), .B(n17111), .Z(n17098) );
  AND U19158 ( .A(n17112), .B(n17113), .Z(n17111) );
  XNOR U19159 ( .A(n17110), .B(n8557), .Z(n17113) );
  XNOR U19160 ( .A(n17106), .B(n17108), .Z(n8557) );
  NAND U19161 ( .A(n17114), .B(nreg[624]), .Z(n17108) );
  NAND U19162 ( .A(n12326), .B(nreg[624]), .Z(n17114) );
  XNOR U19163 ( .A(n17104), .B(n17115), .Z(n17106) );
  XOR U19164 ( .A(n17116), .B(n17117), .Z(n17104) );
  AND U19165 ( .A(n17118), .B(n17119), .Z(n17117) );
  XNOR U19166 ( .A(n17120), .B(n17116), .Z(n17119) );
  XOR U19167 ( .A(n17121), .B(nreg[624]), .Z(n17112) );
  IV U19168 ( .A(n17110), .Z(n17121) );
  XOR U19169 ( .A(n17122), .B(n17123), .Z(n17110) );
  AND U19170 ( .A(n17124), .B(n17125), .Z(n17123) );
  XNOR U19171 ( .A(n17122), .B(n8563), .Z(n17125) );
  XNOR U19172 ( .A(n17118), .B(n17120), .Z(n8563) );
  NAND U19173 ( .A(n17126), .B(nreg[623]), .Z(n17120) );
  NAND U19174 ( .A(n12326), .B(nreg[623]), .Z(n17126) );
  XNOR U19175 ( .A(n17116), .B(n17127), .Z(n17118) );
  XOR U19176 ( .A(n17128), .B(n17129), .Z(n17116) );
  AND U19177 ( .A(n17130), .B(n17131), .Z(n17129) );
  XNOR U19178 ( .A(n17132), .B(n17128), .Z(n17131) );
  XOR U19179 ( .A(n17133), .B(nreg[623]), .Z(n17124) );
  IV U19180 ( .A(n17122), .Z(n17133) );
  XOR U19181 ( .A(n17134), .B(n17135), .Z(n17122) );
  AND U19182 ( .A(n17136), .B(n17137), .Z(n17135) );
  XNOR U19183 ( .A(n17134), .B(n8569), .Z(n17137) );
  XNOR U19184 ( .A(n17130), .B(n17132), .Z(n8569) );
  NAND U19185 ( .A(n17138), .B(nreg[622]), .Z(n17132) );
  NAND U19186 ( .A(n12326), .B(nreg[622]), .Z(n17138) );
  XNOR U19187 ( .A(n17128), .B(n17139), .Z(n17130) );
  XOR U19188 ( .A(n17140), .B(n17141), .Z(n17128) );
  AND U19189 ( .A(n17142), .B(n17143), .Z(n17141) );
  XNOR U19190 ( .A(n17144), .B(n17140), .Z(n17143) );
  XOR U19191 ( .A(n17145), .B(nreg[622]), .Z(n17136) );
  IV U19192 ( .A(n17134), .Z(n17145) );
  XOR U19193 ( .A(n17146), .B(n17147), .Z(n17134) );
  AND U19194 ( .A(n17148), .B(n17149), .Z(n17147) );
  XNOR U19195 ( .A(n17146), .B(n8575), .Z(n17149) );
  XNOR U19196 ( .A(n17142), .B(n17144), .Z(n8575) );
  NAND U19197 ( .A(n17150), .B(nreg[621]), .Z(n17144) );
  NAND U19198 ( .A(n12326), .B(nreg[621]), .Z(n17150) );
  XNOR U19199 ( .A(n17140), .B(n17151), .Z(n17142) );
  XOR U19200 ( .A(n17152), .B(n17153), .Z(n17140) );
  AND U19201 ( .A(n17154), .B(n17155), .Z(n17153) );
  XNOR U19202 ( .A(n17156), .B(n17152), .Z(n17155) );
  XOR U19203 ( .A(n17157), .B(nreg[621]), .Z(n17148) );
  IV U19204 ( .A(n17146), .Z(n17157) );
  XOR U19205 ( .A(n17158), .B(n17159), .Z(n17146) );
  AND U19206 ( .A(n17160), .B(n17161), .Z(n17159) );
  XNOR U19207 ( .A(n17158), .B(n8581), .Z(n17161) );
  XNOR U19208 ( .A(n17154), .B(n17156), .Z(n8581) );
  NAND U19209 ( .A(n17162), .B(nreg[620]), .Z(n17156) );
  NAND U19210 ( .A(n12326), .B(nreg[620]), .Z(n17162) );
  XNOR U19211 ( .A(n17152), .B(n17163), .Z(n17154) );
  XOR U19212 ( .A(n17164), .B(n17165), .Z(n17152) );
  AND U19213 ( .A(n17166), .B(n17167), .Z(n17165) );
  XNOR U19214 ( .A(n17168), .B(n17164), .Z(n17167) );
  XOR U19215 ( .A(n17169), .B(nreg[620]), .Z(n17160) );
  IV U19216 ( .A(n17158), .Z(n17169) );
  XOR U19217 ( .A(n17170), .B(n17171), .Z(n17158) );
  AND U19218 ( .A(n17172), .B(n17173), .Z(n17171) );
  XNOR U19219 ( .A(n17170), .B(n8587), .Z(n17173) );
  XNOR U19220 ( .A(n17166), .B(n17168), .Z(n8587) );
  NAND U19221 ( .A(n17174), .B(nreg[619]), .Z(n17168) );
  NAND U19222 ( .A(n12326), .B(nreg[619]), .Z(n17174) );
  XNOR U19223 ( .A(n17164), .B(n17175), .Z(n17166) );
  XOR U19224 ( .A(n17176), .B(n17177), .Z(n17164) );
  AND U19225 ( .A(n17178), .B(n17179), .Z(n17177) );
  XNOR U19226 ( .A(n17180), .B(n17176), .Z(n17179) );
  XOR U19227 ( .A(n17181), .B(nreg[619]), .Z(n17172) );
  IV U19228 ( .A(n17170), .Z(n17181) );
  XOR U19229 ( .A(n17182), .B(n17183), .Z(n17170) );
  AND U19230 ( .A(n17184), .B(n17185), .Z(n17183) );
  XNOR U19231 ( .A(n17182), .B(n8593), .Z(n17185) );
  XNOR U19232 ( .A(n17178), .B(n17180), .Z(n8593) );
  NAND U19233 ( .A(n17186), .B(nreg[618]), .Z(n17180) );
  NAND U19234 ( .A(n12326), .B(nreg[618]), .Z(n17186) );
  XNOR U19235 ( .A(n17176), .B(n17187), .Z(n17178) );
  XOR U19236 ( .A(n17188), .B(n17189), .Z(n17176) );
  AND U19237 ( .A(n17190), .B(n17191), .Z(n17189) );
  XNOR U19238 ( .A(n17192), .B(n17188), .Z(n17191) );
  XOR U19239 ( .A(n17193), .B(nreg[618]), .Z(n17184) );
  IV U19240 ( .A(n17182), .Z(n17193) );
  XOR U19241 ( .A(n17194), .B(n17195), .Z(n17182) );
  AND U19242 ( .A(n17196), .B(n17197), .Z(n17195) );
  XNOR U19243 ( .A(n17194), .B(n8599), .Z(n17197) );
  XNOR U19244 ( .A(n17190), .B(n17192), .Z(n8599) );
  NAND U19245 ( .A(n17198), .B(nreg[617]), .Z(n17192) );
  NAND U19246 ( .A(n12326), .B(nreg[617]), .Z(n17198) );
  XNOR U19247 ( .A(n17188), .B(n17199), .Z(n17190) );
  XOR U19248 ( .A(n17200), .B(n17201), .Z(n17188) );
  AND U19249 ( .A(n17202), .B(n17203), .Z(n17201) );
  XNOR U19250 ( .A(n17204), .B(n17200), .Z(n17203) );
  XOR U19251 ( .A(n17205), .B(nreg[617]), .Z(n17196) );
  IV U19252 ( .A(n17194), .Z(n17205) );
  XOR U19253 ( .A(n17206), .B(n17207), .Z(n17194) );
  AND U19254 ( .A(n17208), .B(n17209), .Z(n17207) );
  XNOR U19255 ( .A(n17206), .B(n8605), .Z(n17209) );
  XNOR U19256 ( .A(n17202), .B(n17204), .Z(n8605) );
  NAND U19257 ( .A(n17210), .B(nreg[616]), .Z(n17204) );
  NAND U19258 ( .A(n12326), .B(nreg[616]), .Z(n17210) );
  XNOR U19259 ( .A(n17200), .B(n17211), .Z(n17202) );
  XOR U19260 ( .A(n17212), .B(n17213), .Z(n17200) );
  AND U19261 ( .A(n17214), .B(n17215), .Z(n17213) );
  XNOR U19262 ( .A(n17216), .B(n17212), .Z(n17215) );
  XOR U19263 ( .A(n17217), .B(nreg[616]), .Z(n17208) );
  IV U19264 ( .A(n17206), .Z(n17217) );
  XOR U19265 ( .A(n17218), .B(n17219), .Z(n17206) );
  AND U19266 ( .A(n17220), .B(n17221), .Z(n17219) );
  XNOR U19267 ( .A(n17218), .B(n8611), .Z(n17221) );
  XNOR U19268 ( .A(n17214), .B(n17216), .Z(n8611) );
  NAND U19269 ( .A(n17222), .B(nreg[615]), .Z(n17216) );
  NAND U19270 ( .A(n12326), .B(nreg[615]), .Z(n17222) );
  XNOR U19271 ( .A(n17212), .B(n17223), .Z(n17214) );
  XOR U19272 ( .A(n17224), .B(n17225), .Z(n17212) );
  AND U19273 ( .A(n17226), .B(n17227), .Z(n17225) );
  XNOR U19274 ( .A(n17228), .B(n17224), .Z(n17227) );
  XOR U19275 ( .A(n17229), .B(nreg[615]), .Z(n17220) );
  IV U19276 ( .A(n17218), .Z(n17229) );
  XOR U19277 ( .A(n17230), .B(n17231), .Z(n17218) );
  AND U19278 ( .A(n17232), .B(n17233), .Z(n17231) );
  XNOR U19279 ( .A(n17230), .B(n8617), .Z(n17233) );
  XNOR U19280 ( .A(n17226), .B(n17228), .Z(n8617) );
  NAND U19281 ( .A(n17234), .B(nreg[614]), .Z(n17228) );
  NAND U19282 ( .A(n12326), .B(nreg[614]), .Z(n17234) );
  XNOR U19283 ( .A(n17224), .B(n17235), .Z(n17226) );
  XOR U19284 ( .A(n17236), .B(n17237), .Z(n17224) );
  AND U19285 ( .A(n17238), .B(n17239), .Z(n17237) );
  XNOR U19286 ( .A(n17240), .B(n17236), .Z(n17239) );
  XOR U19287 ( .A(n17241), .B(nreg[614]), .Z(n17232) );
  IV U19288 ( .A(n17230), .Z(n17241) );
  XOR U19289 ( .A(n17242), .B(n17243), .Z(n17230) );
  AND U19290 ( .A(n17244), .B(n17245), .Z(n17243) );
  XNOR U19291 ( .A(n17242), .B(n8623), .Z(n17245) );
  XNOR U19292 ( .A(n17238), .B(n17240), .Z(n8623) );
  NAND U19293 ( .A(n17246), .B(nreg[613]), .Z(n17240) );
  NAND U19294 ( .A(n12326), .B(nreg[613]), .Z(n17246) );
  XNOR U19295 ( .A(n17236), .B(n17247), .Z(n17238) );
  XOR U19296 ( .A(n17248), .B(n17249), .Z(n17236) );
  AND U19297 ( .A(n17250), .B(n17251), .Z(n17249) );
  XNOR U19298 ( .A(n17252), .B(n17248), .Z(n17251) );
  XOR U19299 ( .A(n17253), .B(nreg[613]), .Z(n17244) );
  IV U19300 ( .A(n17242), .Z(n17253) );
  XOR U19301 ( .A(n17254), .B(n17255), .Z(n17242) );
  AND U19302 ( .A(n17256), .B(n17257), .Z(n17255) );
  XNOR U19303 ( .A(n17254), .B(n8629), .Z(n17257) );
  XNOR U19304 ( .A(n17250), .B(n17252), .Z(n8629) );
  NAND U19305 ( .A(n17258), .B(nreg[612]), .Z(n17252) );
  NAND U19306 ( .A(n12326), .B(nreg[612]), .Z(n17258) );
  XNOR U19307 ( .A(n17248), .B(n17259), .Z(n17250) );
  XOR U19308 ( .A(n17260), .B(n17261), .Z(n17248) );
  AND U19309 ( .A(n17262), .B(n17263), .Z(n17261) );
  XNOR U19310 ( .A(n17264), .B(n17260), .Z(n17263) );
  XOR U19311 ( .A(n17265), .B(nreg[612]), .Z(n17256) );
  IV U19312 ( .A(n17254), .Z(n17265) );
  XOR U19313 ( .A(n17266), .B(n17267), .Z(n17254) );
  AND U19314 ( .A(n17268), .B(n17269), .Z(n17267) );
  XNOR U19315 ( .A(n17266), .B(n8635), .Z(n17269) );
  XNOR U19316 ( .A(n17262), .B(n17264), .Z(n8635) );
  NAND U19317 ( .A(n17270), .B(nreg[611]), .Z(n17264) );
  NAND U19318 ( .A(n12326), .B(nreg[611]), .Z(n17270) );
  XNOR U19319 ( .A(n17260), .B(n17271), .Z(n17262) );
  XOR U19320 ( .A(n17272), .B(n17273), .Z(n17260) );
  AND U19321 ( .A(n17274), .B(n17275), .Z(n17273) );
  XNOR U19322 ( .A(n17276), .B(n17272), .Z(n17275) );
  XOR U19323 ( .A(n17277), .B(nreg[611]), .Z(n17268) );
  IV U19324 ( .A(n17266), .Z(n17277) );
  XOR U19325 ( .A(n17278), .B(n17279), .Z(n17266) );
  AND U19326 ( .A(n17280), .B(n17281), .Z(n17279) );
  XNOR U19327 ( .A(n17278), .B(n8641), .Z(n17281) );
  XNOR U19328 ( .A(n17274), .B(n17276), .Z(n8641) );
  NAND U19329 ( .A(n17282), .B(nreg[610]), .Z(n17276) );
  NAND U19330 ( .A(n12326), .B(nreg[610]), .Z(n17282) );
  XNOR U19331 ( .A(n17272), .B(n17283), .Z(n17274) );
  XOR U19332 ( .A(n17284), .B(n17285), .Z(n17272) );
  AND U19333 ( .A(n17286), .B(n17287), .Z(n17285) );
  XNOR U19334 ( .A(n17288), .B(n17284), .Z(n17287) );
  XOR U19335 ( .A(n17289), .B(nreg[610]), .Z(n17280) );
  IV U19336 ( .A(n17278), .Z(n17289) );
  XOR U19337 ( .A(n17290), .B(n17291), .Z(n17278) );
  AND U19338 ( .A(n17292), .B(n17293), .Z(n17291) );
  XNOR U19339 ( .A(n17290), .B(n8647), .Z(n17293) );
  XNOR U19340 ( .A(n17286), .B(n17288), .Z(n8647) );
  NAND U19341 ( .A(n17294), .B(nreg[609]), .Z(n17288) );
  NAND U19342 ( .A(n12326), .B(nreg[609]), .Z(n17294) );
  XNOR U19343 ( .A(n17284), .B(n17295), .Z(n17286) );
  XOR U19344 ( .A(n17296), .B(n17297), .Z(n17284) );
  AND U19345 ( .A(n17298), .B(n17299), .Z(n17297) );
  XNOR U19346 ( .A(n17300), .B(n17296), .Z(n17299) );
  XOR U19347 ( .A(n17301), .B(nreg[609]), .Z(n17292) );
  IV U19348 ( .A(n17290), .Z(n17301) );
  XOR U19349 ( .A(n17302), .B(n17303), .Z(n17290) );
  AND U19350 ( .A(n17304), .B(n17305), .Z(n17303) );
  XNOR U19351 ( .A(n17302), .B(n8653), .Z(n17305) );
  XNOR U19352 ( .A(n17298), .B(n17300), .Z(n8653) );
  NAND U19353 ( .A(n17306), .B(nreg[608]), .Z(n17300) );
  NAND U19354 ( .A(n12326), .B(nreg[608]), .Z(n17306) );
  XNOR U19355 ( .A(n17296), .B(n17307), .Z(n17298) );
  XOR U19356 ( .A(n17308), .B(n17309), .Z(n17296) );
  AND U19357 ( .A(n17310), .B(n17311), .Z(n17309) );
  XNOR U19358 ( .A(n17312), .B(n17308), .Z(n17311) );
  XOR U19359 ( .A(n17313), .B(nreg[608]), .Z(n17304) );
  IV U19360 ( .A(n17302), .Z(n17313) );
  XOR U19361 ( .A(n17314), .B(n17315), .Z(n17302) );
  AND U19362 ( .A(n17316), .B(n17317), .Z(n17315) );
  XNOR U19363 ( .A(n17314), .B(n8659), .Z(n17317) );
  XNOR U19364 ( .A(n17310), .B(n17312), .Z(n8659) );
  NAND U19365 ( .A(n17318), .B(nreg[607]), .Z(n17312) );
  NAND U19366 ( .A(n12326), .B(nreg[607]), .Z(n17318) );
  XNOR U19367 ( .A(n17308), .B(n17319), .Z(n17310) );
  XOR U19368 ( .A(n17320), .B(n17321), .Z(n17308) );
  AND U19369 ( .A(n17322), .B(n17323), .Z(n17321) );
  XNOR U19370 ( .A(n17324), .B(n17320), .Z(n17323) );
  XOR U19371 ( .A(n17325), .B(nreg[607]), .Z(n17316) );
  IV U19372 ( .A(n17314), .Z(n17325) );
  XOR U19373 ( .A(n17326), .B(n17327), .Z(n17314) );
  AND U19374 ( .A(n17328), .B(n17329), .Z(n17327) );
  XNOR U19375 ( .A(n17326), .B(n8665), .Z(n17329) );
  XNOR U19376 ( .A(n17322), .B(n17324), .Z(n8665) );
  NAND U19377 ( .A(n17330), .B(nreg[606]), .Z(n17324) );
  NAND U19378 ( .A(n12326), .B(nreg[606]), .Z(n17330) );
  XNOR U19379 ( .A(n17320), .B(n17331), .Z(n17322) );
  XOR U19380 ( .A(n17332), .B(n17333), .Z(n17320) );
  AND U19381 ( .A(n17334), .B(n17335), .Z(n17333) );
  XNOR U19382 ( .A(n17336), .B(n17332), .Z(n17335) );
  XOR U19383 ( .A(n17337), .B(nreg[606]), .Z(n17328) );
  IV U19384 ( .A(n17326), .Z(n17337) );
  XOR U19385 ( .A(n17338), .B(n17339), .Z(n17326) );
  AND U19386 ( .A(n17340), .B(n17341), .Z(n17339) );
  XNOR U19387 ( .A(n17338), .B(n8671), .Z(n17341) );
  XNOR U19388 ( .A(n17334), .B(n17336), .Z(n8671) );
  NAND U19389 ( .A(n17342), .B(nreg[605]), .Z(n17336) );
  NAND U19390 ( .A(n12326), .B(nreg[605]), .Z(n17342) );
  XNOR U19391 ( .A(n17332), .B(n17343), .Z(n17334) );
  XOR U19392 ( .A(n17344), .B(n17345), .Z(n17332) );
  AND U19393 ( .A(n17346), .B(n17347), .Z(n17345) );
  XNOR U19394 ( .A(n17348), .B(n17344), .Z(n17347) );
  XOR U19395 ( .A(n17349), .B(nreg[605]), .Z(n17340) );
  IV U19396 ( .A(n17338), .Z(n17349) );
  XOR U19397 ( .A(n17350), .B(n17351), .Z(n17338) );
  AND U19398 ( .A(n17352), .B(n17353), .Z(n17351) );
  XNOR U19399 ( .A(n17350), .B(n8677), .Z(n17353) );
  XNOR U19400 ( .A(n17346), .B(n17348), .Z(n8677) );
  NAND U19401 ( .A(n17354), .B(nreg[604]), .Z(n17348) );
  NAND U19402 ( .A(n12326), .B(nreg[604]), .Z(n17354) );
  XNOR U19403 ( .A(n17344), .B(n17355), .Z(n17346) );
  XOR U19404 ( .A(n17356), .B(n17357), .Z(n17344) );
  AND U19405 ( .A(n17358), .B(n17359), .Z(n17357) );
  XNOR U19406 ( .A(n17360), .B(n17356), .Z(n17359) );
  XOR U19407 ( .A(n17361), .B(nreg[604]), .Z(n17352) );
  IV U19408 ( .A(n17350), .Z(n17361) );
  XOR U19409 ( .A(n17362), .B(n17363), .Z(n17350) );
  AND U19410 ( .A(n17364), .B(n17365), .Z(n17363) );
  XNOR U19411 ( .A(n17362), .B(n8683), .Z(n17365) );
  XNOR U19412 ( .A(n17358), .B(n17360), .Z(n8683) );
  NAND U19413 ( .A(n17366), .B(nreg[603]), .Z(n17360) );
  NAND U19414 ( .A(n12326), .B(nreg[603]), .Z(n17366) );
  XNOR U19415 ( .A(n17356), .B(n17367), .Z(n17358) );
  XOR U19416 ( .A(n17368), .B(n17369), .Z(n17356) );
  AND U19417 ( .A(n17370), .B(n17371), .Z(n17369) );
  XNOR U19418 ( .A(n17372), .B(n17368), .Z(n17371) );
  XOR U19419 ( .A(n17373), .B(nreg[603]), .Z(n17364) );
  IV U19420 ( .A(n17362), .Z(n17373) );
  XOR U19421 ( .A(n17374), .B(n17375), .Z(n17362) );
  AND U19422 ( .A(n17376), .B(n17377), .Z(n17375) );
  XNOR U19423 ( .A(n17374), .B(n8689), .Z(n17377) );
  XNOR U19424 ( .A(n17370), .B(n17372), .Z(n8689) );
  NAND U19425 ( .A(n17378), .B(nreg[602]), .Z(n17372) );
  NAND U19426 ( .A(n12326), .B(nreg[602]), .Z(n17378) );
  XNOR U19427 ( .A(n17368), .B(n17379), .Z(n17370) );
  XOR U19428 ( .A(n17380), .B(n17381), .Z(n17368) );
  AND U19429 ( .A(n17382), .B(n17383), .Z(n17381) );
  XNOR U19430 ( .A(n17384), .B(n17380), .Z(n17383) );
  XOR U19431 ( .A(n17385), .B(nreg[602]), .Z(n17376) );
  IV U19432 ( .A(n17374), .Z(n17385) );
  XOR U19433 ( .A(n17386), .B(n17387), .Z(n17374) );
  AND U19434 ( .A(n17388), .B(n17389), .Z(n17387) );
  XNOR U19435 ( .A(n17386), .B(n8695), .Z(n17389) );
  XNOR U19436 ( .A(n17382), .B(n17384), .Z(n8695) );
  NAND U19437 ( .A(n17390), .B(nreg[601]), .Z(n17384) );
  NAND U19438 ( .A(n12326), .B(nreg[601]), .Z(n17390) );
  XNOR U19439 ( .A(n17380), .B(n17391), .Z(n17382) );
  XOR U19440 ( .A(n17392), .B(n17393), .Z(n17380) );
  AND U19441 ( .A(n17394), .B(n17395), .Z(n17393) );
  XNOR U19442 ( .A(n17396), .B(n17392), .Z(n17395) );
  XOR U19443 ( .A(n17397), .B(nreg[601]), .Z(n17388) );
  IV U19444 ( .A(n17386), .Z(n17397) );
  XOR U19445 ( .A(n17398), .B(n17399), .Z(n17386) );
  AND U19446 ( .A(n17400), .B(n17401), .Z(n17399) );
  XNOR U19447 ( .A(n17398), .B(n8701), .Z(n17401) );
  XNOR U19448 ( .A(n17394), .B(n17396), .Z(n8701) );
  NAND U19449 ( .A(n17402), .B(nreg[600]), .Z(n17396) );
  NAND U19450 ( .A(n12326), .B(nreg[600]), .Z(n17402) );
  XNOR U19451 ( .A(n17392), .B(n17403), .Z(n17394) );
  XOR U19452 ( .A(n17404), .B(n17405), .Z(n17392) );
  AND U19453 ( .A(n17406), .B(n17407), .Z(n17405) );
  XNOR U19454 ( .A(n17408), .B(n17404), .Z(n17407) );
  XOR U19455 ( .A(n17409), .B(nreg[600]), .Z(n17400) );
  IV U19456 ( .A(n17398), .Z(n17409) );
  XOR U19457 ( .A(n17410), .B(n17411), .Z(n17398) );
  AND U19458 ( .A(n17412), .B(n17413), .Z(n17411) );
  XNOR U19459 ( .A(n17410), .B(n8707), .Z(n17413) );
  XNOR U19460 ( .A(n17406), .B(n17408), .Z(n8707) );
  NAND U19461 ( .A(n17414), .B(nreg[599]), .Z(n17408) );
  NAND U19462 ( .A(n12326), .B(nreg[599]), .Z(n17414) );
  XNOR U19463 ( .A(n17404), .B(n17415), .Z(n17406) );
  XOR U19464 ( .A(n17416), .B(n17417), .Z(n17404) );
  AND U19465 ( .A(n17418), .B(n17419), .Z(n17417) );
  XNOR U19466 ( .A(n17420), .B(n17416), .Z(n17419) );
  XOR U19467 ( .A(n17421), .B(nreg[599]), .Z(n17412) );
  IV U19468 ( .A(n17410), .Z(n17421) );
  XOR U19469 ( .A(n17422), .B(n17423), .Z(n17410) );
  AND U19470 ( .A(n17424), .B(n17425), .Z(n17423) );
  XNOR U19471 ( .A(n17422), .B(n8713), .Z(n17425) );
  XNOR U19472 ( .A(n17418), .B(n17420), .Z(n8713) );
  NAND U19473 ( .A(n17426), .B(nreg[598]), .Z(n17420) );
  NAND U19474 ( .A(n12326), .B(nreg[598]), .Z(n17426) );
  XNOR U19475 ( .A(n17416), .B(n17427), .Z(n17418) );
  XOR U19476 ( .A(n17428), .B(n17429), .Z(n17416) );
  AND U19477 ( .A(n17430), .B(n17431), .Z(n17429) );
  XNOR U19478 ( .A(n17432), .B(n17428), .Z(n17431) );
  XOR U19479 ( .A(n17433), .B(nreg[598]), .Z(n17424) );
  IV U19480 ( .A(n17422), .Z(n17433) );
  XOR U19481 ( .A(n17434), .B(n17435), .Z(n17422) );
  AND U19482 ( .A(n17436), .B(n17437), .Z(n17435) );
  XNOR U19483 ( .A(n17434), .B(n8719), .Z(n17437) );
  XNOR U19484 ( .A(n17430), .B(n17432), .Z(n8719) );
  NAND U19485 ( .A(n17438), .B(nreg[597]), .Z(n17432) );
  NAND U19486 ( .A(n12326), .B(nreg[597]), .Z(n17438) );
  XNOR U19487 ( .A(n17428), .B(n17439), .Z(n17430) );
  XOR U19488 ( .A(n17440), .B(n17441), .Z(n17428) );
  AND U19489 ( .A(n17442), .B(n17443), .Z(n17441) );
  XNOR U19490 ( .A(n17444), .B(n17440), .Z(n17443) );
  XOR U19491 ( .A(n17445), .B(nreg[597]), .Z(n17436) );
  IV U19492 ( .A(n17434), .Z(n17445) );
  XOR U19493 ( .A(n17446), .B(n17447), .Z(n17434) );
  AND U19494 ( .A(n17448), .B(n17449), .Z(n17447) );
  XNOR U19495 ( .A(n17446), .B(n8725), .Z(n17449) );
  XNOR U19496 ( .A(n17442), .B(n17444), .Z(n8725) );
  NAND U19497 ( .A(n17450), .B(nreg[596]), .Z(n17444) );
  NAND U19498 ( .A(n12326), .B(nreg[596]), .Z(n17450) );
  XNOR U19499 ( .A(n17440), .B(n17451), .Z(n17442) );
  XOR U19500 ( .A(n17452), .B(n17453), .Z(n17440) );
  AND U19501 ( .A(n17454), .B(n17455), .Z(n17453) );
  XNOR U19502 ( .A(n17456), .B(n17452), .Z(n17455) );
  XOR U19503 ( .A(n17457), .B(nreg[596]), .Z(n17448) );
  IV U19504 ( .A(n17446), .Z(n17457) );
  XOR U19505 ( .A(n17458), .B(n17459), .Z(n17446) );
  AND U19506 ( .A(n17460), .B(n17461), .Z(n17459) );
  XNOR U19507 ( .A(n17458), .B(n8731), .Z(n17461) );
  XNOR U19508 ( .A(n17454), .B(n17456), .Z(n8731) );
  NAND U19509 ( .A(n17462), .B(nreg[595]), .Z(n17456) );
  NAND U19510 ( .A(n12326), .B(nreg[595]), .Z(n17462) );
  XNOR U19511 ( .A(n17452), .B(n17463), .Z(n17454) );
  XOR U19512 ( .A(n17464), .B(n17465), .Z(n17452) );
  AND U19513 ( .A(n17466), .B(n17467), .Z(n17465) );
  XNOR U19514 ( .A(n17468), .B(n17464), .Z(n17467) );
  XOR U19515 ( .A(n17469), .B(nreg[595]), .Z(n17460) );
  IV U19516 ( .A(n17458), .Z(n17469) );
  XOR U19517 ( .A(n17470), .B(n17471), .Z(n17458) );
  AND U19518 ( .A(n17472), .B(n17473), .Z(n17471) );
  XNOR U19519 ( .A(n17470), .B(n8737), .Z(n17473) );
  XNOR U19520 ( .A(n17466), .B(n17468), .Z(n8737) );
  NAND U19521 ( .A(n17474), .B(nreg[594]), .Z(n17468) );
  NAND U19522 ( .A(n12326), .B(nreg[594]), .Z(n17474) );
  XNOR U19523 ( .A(n17464), .B(n17475), .Z(n17466) );
  XOR U19524 ( .A(n17476), .B(n17477), .Z(n17464) );
  AND U19525 ( .A(n17478), .B(n17479), .Z(n17477) );
  XNOR U19526 ( .A(n17480), .B(n17476), .Z(n17479) );
  XOR U19527 ( .A(n17481), .B(nreg[594]), .Z(n17472) );
  IV U19528 ( .A(n17470), .Z(n17481) );
  XOR U19529 ( .A(n17482), .B(n17483), .Z(n17470) );
  AND U19530 ( .A(n17484), .B(n17485), .Z(n17483) );
  XNOR U19531 ( .A(n17482), .B(n8743), .Z(n17485) );
  XNOR U19532 ( .A(n17478), .B(n17480), .Z(n8743) );
  NAND U19533 ( .A(n17486), .B(nreg[593]), .Z(n17480) );
  NAND U19534 ( .A(n12326), .B(nreg[593]), .Z(n17486) );
  XNOR U19535 ( .A(n17476), .B(n17487), .Z(n17478) );
  XOR U19536 ( .A(n17488), .B(n17489), .Z(n17476) );
  AND U19537 ( .A(n17490), .B(n17491), .Z(n17489) );
  XNOR U19538 ( .A(n17492), .B(n17488), .Z(n17491) );
  XOR U19539 ( .A(n17493), .B(nreg[593]), .Z(n17484) );
  IV U19540 ( .A(n17482), .Z(n17493) );
  XOR U19541 ( .A(n17494), .B(n17495), .Z(n17482) );
  AND U19542 ( .A(n17496), .B(n17497), .Z(n17495) );
  XNOR U19543 ( .A(n17494), .B(n8749), .Z(n17497) );
  XNOR U19544 ( .A(n17490), .B(n17492), .Z(n8749) );
  NAND U19545 ( .A(n17498), .B(nreg[592]), .Z(n17492) );
  NAND U19546 ( .A(n12326), .B(nreg[592]), .Z(n17498) );
  XNOR U19547 ( .A(n17488), .B(n17499), .Z(n17490) );
  XOR U19548 ( .A(n17500), .B(n17501), .Z(n17488) );
  AND U19549 ( .A(n17502), .B(n17503), .Z(n17501) );
  XNOR U19550 ( .A(n17504), .B(n17500), .Z(n17503) );
  XOR U19551 ( .A(n17505), .B(nreg[592]), .Z(n17496) );
  IV U19552 ( .A(n17494), .Z(n17505) );
  XOR U19553 ( .A(n17506), .B(n17507), .Z(n17494) );
  AND U19554 ( .A(n17508), .B(n17509), .Z(n17507) );
  XNOR U19555 ( .A(n17506), .B(n8755), .Z(n17509) );
  XNOR U19556 ( .A(n17502), .B(n17504), .Z(n8755) );
  NAND U19557 ( .A(n17510), .B(nreg[591]), .Z(n17504) );
  NAND U19558 ( .A(n12326), .B(nreg[591]), .Z(n17510) );
  XNOR U19559 ( .A(n17500), .B(n17511), .Z(n17502) );
  XOR U19560 ( .A(n17512), .B(n17513), .Z(n17500) );
  AND U19561 ( .A(n17514), .B(n17515), .Z(n17513) );
  XNOR U19562 ( .A(n17516), .B(n17512), .Z(n17515) );
  XOR U19563 ( .A(n17517), .B(nreg[591]), .Z(n17508) );
  IV U19564 ( .A(n17506), .Z(n17517) );
  XOR U19565 ( .A(n17518), .B(n17519), .Z(n17506) );
  AND U19566 ( .A(n17520), .B(n17521), .Z(n17519) );
  XNOR U19567 ( .A(n17518), .B(n8761), .Z(n17521) );
  XNOR U19568 ( .A(n17514), .B(n17516), .Z(n8761) );
  NAND U19569 ( .A(n17522), .B(nreg[590]), .Z(n17516) );
  NAND U19570 ( .A(n12326), .B(nreg[590]), .Z(n17522) );
  XNOR U19571 ( .A(n17512), .B(n17523), .Z(n17514) );
  XOR U19572 ( .A(n17524), .B(n17525), .Z(n17512) );
  AND U19573 ( .A(n17526), .B(n17527), .Z(n17525) );
  XNOR U19574 ( .A(n17528), .B(n17524), .Z(n17527) );
  XOR U19575 ( .A(n17529), .B(nreg[590]), .Z(n17520) );
  IV U19576 ( .A(n17518), .Z(n17529) );
  XOR U19577 ( .A(n17530), .B(n17531), .Z(n17518) );
  AND U19578 ( .A(n17532), .B(n17533), .Z(n17531) );
  XNOR U19579 ( .A(n17530), .B(n8767), .Z(n17533) );
  XNOR U19580 ( .A(n17526), .B(n17528), .Z(n8767) );
  NAND U19581 ( .A(n17534), .B(nreg[589]), .Z(n17528) );
  NAND U19582 ( .A(n12326), .B(nreg[589]), .Z(n17534) );
  XNOR U19583 ( .A(n17524), .B(n17535), .Z(n17526) );
  XOR U19584 ( .A(n17536), .B(n17537), .Z(n17524) );
  AND U19585 ( .A(n17538), .B(n17539), .Z(n17537) );
  XNOR U19586 ( .A(n17540), .B(n17536), .Z(n17539) );
  XOR U19587 ( .A(n17541), .B(nreg[589]), .Z(n17532) );
  IV U19588 ( .A(n17530), .Z(n17541) );
  XOR U19589 ( .A(n17542), .B(n17543), .Z(n17530) );
  AND U19590 ( .A(n17544), .B(n17545), .Z(n17543) );
  XNOR U19591 ( .A(n17542), .B(n8773), .Z(n17545) );
  XNOR U19592 ( .A(n17538), .B(n17540), .Z(n8773) );
  NAND U19593 ( .A(n17546), .B(nreg[588]), .Z(n17540) );
  NAND U19594 ( .A(n12326), .B(nreg[588]), .Z(n17546) );
  XNOR U19595 ( .A(n17536), .B(n17547), .Z(n17538) );
  XOR U19596 ( .A(n17548), .B(n17549), .Z(n17536) );
  AND U19597 ( .A(n17550), .B(n17551), .Z(n17549) );
  XNOR U19598 ( .A(n17552), .B(n17548), .Z(n17551) );
  XOR U19599 ( .A(n17553), .B(nreg[588]), .Z(n17544) );
  IV U19600 ( .A(n17542), .Z(n17553) );
  XOR U19601 ( .A(n17554), .B(n17555), .Z(n17542) );
  AND U19602 ( .A(n17556), .B(n17557), .Z(n17555) );
  XNOR U19603 ( .A(n17554), .B(n8779), .Z(n17557) );
  XNOR U19604 ( .A(n17550), .B(n17552), .Z(n8779) );
  NAND U19605 ( .A(n17558), .B(nreg[587]), .Z(n17552) );
  NAND U19606 ( .A(n12326), .B(nreg[587]), .Z(n17558) );
  XNOR U19607 ( .A(n17548), .B(n17559), .Z(n17550) );
  XOR U19608 ( .A(n17560), .B(n17561), .Z(n17548) );
  AND U19609 ( .A(n17562), .B(n17563), .Z(n17561) );
  XNOR U19610 ( .A(n17564), .B(n17560), .Z(n17563) );
  XOR U19611 ( .A(n17565), .B(nreg[587]), .Z(n17556) );
  IV U19612 ( .A(n17554), .Z(n17565) );
  XOR U19613 ( .A(n17566), .B(n17567), .Z(n17554) );
  AND U19614 ( .A(n17568), .B(n17569), .Z(n17567) );
  XNOR U19615 ( .A(n17566), .B(n8785), .Z(n17569) );
  XNOR U19616 ( .A(n17562), .B(n17564), .Z(n8785) );
  NAND U19617 ( .A(n17570), .B(nreg[586]), .Z(n17564) );
  NAND U19618 ( .A(n12326), .B(nreg[586]), .Z(n17570) );
  XNOR U19619 ( .A(n17560), .B(n17571), .Z(n17562) );
  XOR U19620 ( .A(n17572), .B(n17573), .Z(n17560) );
  AND U19621 ( .A(n17574), .B(n17575), .Z(n17573) );
  XNOR U19622 ( .A(n17576), .B(n17572), .Z(n17575) );
  XOR U19623 ( .A(n17577), .B(nreg[586]), .Z(n17568) );
  IV U19624 ( .A(n17566), .Z(n17577) );
  XOR U19625 ( .A(n17578), .B(n17579), .Z(n17566) );
  AND U19626 ( .A(n17580), .B(n17581), .Z(n17579) );
  XNOR U19627 ( .A(n17578), .B(n8791), .Z(n17581) );
  XNOR U19628 ( .A(n17574), .B(n17576), .Z(n8791) );
  NAND U19629 ( .A(n17582), .B(nreg[585]), .Z(n17576) );
  NAND U19630 ( .A(n12326), .B(nreg[585]), .Z(n17582) );
  XNOR U19631 ( .A(n17572), .B(n17583), .Z(n17574) );
  XOR U19632 ( .A(n17584), .B(n17585), .Z(n17572) );
  AND U19633 ( .A(n17586), .B(n17587), .Z(n17585) );
  XNOR U19634 ( .A(n17588), .B(n17584), .Z(n17587) );
  XOR U19635 ( .A(n17589), .B(nreg[585]), .Z(n17580) );
  IV U19636 ( .A(n17578), .Z(n17589) );
  XOR U19637 ( .A(n17590), .B(n17591), .Z(n17578) );
  AND U19638 ( .A(n17592), .B(n17593), .Z(n17591) );
  XNOR U19639 ( .A(n17590), .B(n8797), .Z(n17593) );
  XNOR U19640 ( .A(n17586), .B(n17588), .Z(n8797) );
  NAND U19641 ( .A(n17594), .B(nreg[584]), .Z(n17588) );
  NAND U19642 ( .A(n12326), .B(nreg[584]), .Z(n17594) );
  XNOR U19643 ( .A(n17584), .B(n17595), .Z(n17586) );
  XOR U19644 ( .A(n17596), .B(n17597), .Z(n17584) );
  AND U19645 ( .A(n17598), .B(n17599), .Z(n17597) );
  XNOR U19646 ( .A(n17600), .B(n17596), .Z(n17599) );
  XOR U19647 ( .A(n17601), .B(nreg[584]), .Z(n17592) );
  IV U19648 ( .A(n17590), .Z(n17601) );
  XOR U19649 ( .A(n17602), .B(n17603), .Z(n17590) );
  AND U19650 ( .A(n17604), .B(n17605), .Z(n17603) );
  XNOR U19651 ( .A(n17602), .B(n8803), .Z(n17605) );
  XNOR U19652 ( .A(n17598), .B(n17600), .Z(n8803) );
  NAND U19653 ( .A(n17606), .B(nreg[583]), .Z(n17600) );
  NAND U19654 ( .A(n12326), .B(nreg[583]), .Z(n17606) );
  XNOR U19655 ( .A(n17596), .B(n17607), .Z(n17598) );
  XOR U19656 ( .A(n17608), .B(n17609), .Z(n17596) );
  AND U19657 ( .A(n17610), .B(n17611), .Z(n17609) );
  XNOR U19658 ( .A(n17612), .B(n17608), .Z(n17611) );
  XOR U19659 ( .A(n17613), .B(nreg[583]), .Z(n17604) );
  IV U19660 ( .A(n17602), .Z(n17613) );
  XOR U19661 ( .A(n17614), .B(n17615), .Z(n17602) );
  AND U19662 ( .A(n17616), .B(n17617), .Z(n17615) );
  XNOR U19663 ( .A(n17614), .B(n8809), .Z(n17617) );
  XNOR U19664 ( .A(n17610), .B(n17612), .Z(n8809) );
  NAND U19665 ( .A(n17618), .B(nreg[582]), .Z(n17612) );
  NAND U19666 ( .A(n12326), .B(nreg[582]), .Z(n17618) );
  XNOR U19667 ( .A(n17608), .B(n17619), .Z(n17610) );
  XOR U19668 ( .A(n17620), .B(n17621), .Z(n17608) );
  AND U19669 ( .A(n17622), .B(n17623), .Z(n17621) );
  XNOR U19670 ( .A(n17624), .B(n17620), .Z(n17623) );
  XOR U19671 ( .A(n17625), .B(nreg[582]), .Z(n17616) );
  IV U19672 ( .A(n17614), .Z(n17625) );
  XOR U19673 ( .A(n17626), .B(n17627), .Z(n17614) );
  AND U19674 ( .A(n17628), .B(n17629), .Z(n17627) );
  XNOR U19675 ( .A(n17626), .B(n8815), .Z(n17629) );
  XNOR U19676 ( .A(n17622), .B(n17624), .Z(n8815) );
  NAND U19677 ( .A(n17630), .B(nreg[581]), .Z(n17624) );
  NAND U19678 ( .A(n12326), .B(nreg[581]), .Z(n17630) );
  XNOR U19679 ( .A(n17620), .B(n17631), .Z(n17622) );
  XOR U19680 ( .A(n17632), .B(n17633), .Z(n17620) );
  AND U19681 ( .A(n17634), .B(n17635), .Z(n17633) );
  XNOR U19682 ( .A(n17636), .B(n17632), .Z(n17635) );
  XOR U19683 ( .A(n17637), .B(nreg[581]), .Z(n17628) );
  IV U19684 ( .A(n17626), .Z(n17637) );
  XOR U19685 ( .A(n17638), .B(n17639), .Z(n17626) );
  AND U19686 ( .A(n17640), .B(n17641), .Z(n17639) );
  XNOR U19687 ( .A(n17638), .B(n8821), .Z(n17641) );
  XNOR U19688 ( .A(n17634), .B(n17636), .Z(n8821) );
  NAND U19689 ( .A(n17642), .B(nreg[580]), .Z(n17636) );
  NAND U19690 ( .A(n12326), .B(nreg[580]), .Z(n17642) );
  XNOR U19691 ( .A(n17632), .B(n17643), .Z(n17634) );
  XOR U19692 ( .A(n17644), .B(n17645), .Z(n17632) );
  AND U19693 ( .A(n17646), .B(n17647), .Z(n17645) );
  XNOR U19694 ( .A(n17648), .B(n17644), .Z(n17647) );
  XOR U19695 ( .A(n17649), .B(nreg[580]), .Z(n17640) );
  IV U19696 ( .A(n17638), .Z(n17649) );
  XOR U19697 ( .A(n17650), .B(n17651), .Z(n17638) );
  AND U19698 ( .A(n17652), .B(n17653), .Z(n17651) );
  XNOR U19699 ( .A(n17650), .B(n8827), .Z(n17653) );
  XNOR U19700 ( .A(n17646), .B(n17648), .Z(n8827) );
  NAND U19701 ( .A(n17654), .B(nreg[579]), .Z(n17648) );
  NAND U19702 ( .A(n12326), .B(nreg[579]), .Z(n17654) );
  XNOR U19703 ( .A(n17644), .B(n17655), .Z(n17646) );
  XOR U19704 ( .A(n17656), .B(n17657), .Z(n17644) );
  AND U19705 ( .A(n17658), .B(n17659), .Z(n17657) );
  XNOR U19706 ( .A(n17660), .B(n17656), .Z(n17659) );
  XOR U19707 ( .A(n17661), .B(nreg[579]), .Z(n17652) );
  IV U19708 ( .A(n17650), .Z(n17661) );
  XOR U19709 ( .A(n17662), .B(n17663), .Z(n17650) );
  AND U19710 ( .A(n17664), .B(n17665), .Z(n17663) );
  XNOR U19711 ( .A(n17662), .B(n8833), .Z(n17665) );
  XNOR U19712 ( .A(n17658), .B(n17660), .Z(n8833) );
  NAND U19713 ( .A(n17666), .B(nreg[578]), .Z(n17660) );
  NAND U19714 ( .A(n12326), .B(nreg[578]), .Z(n17666) );
  XNOR U19715 ( .A(n17656), .B(n17667), .Z(n17658) );
  XOR U19716 ( .A(n17668), .B(n17669), .Z(n17656) );
  AND U19717 ( .A(n17670), .B(n17671), .Z(n17669) );
  XNOR U19718 ( .A(n17672), .B(n17668), .Z(n17671) );
  XOR U19719 ( .A(n17673), .B(nreg[578]), .Z(n17664) );
  IV U19720 ( .A(n17662), .Z(n17673) );
  XOR U19721 ( .A(n17674), .B(n17675), .Z(n17662) );
  AND U19722 ( .A(n17676), .B(n17677), .Z(n17675) );
  XNOR U19723 ( .A(n17674), .B(n8839), .Z(n17677) );
  XNOR U19724 ( .A(n17670), .B(n17672), .Z(n8839) );
  NAND U19725 ( .A(n17678), .B(nreg[577]), .Z(n17672) );
  NAND U19726 ( .A(n12326), .B(nreg[577]), .Z(n17678) );
  XNOR U19727 ( .A(n17668), .B(n17679), .Z(n17670) );
  XOR U19728 ( .A(n17680), .B(n17681), .Z(n17668) );
  AND U19729 ( .A(n17682), .B(n17683), .Z(n17681) );
  XNOR U19730 ( .A(n17684), .B(n17680), .Z(n17683) );
  XOR U19731 ( .A(n17685), .B(nreg[577]), .Z(n17676) );
  IV U19732 ( .A(n17674), .Z(n17685) );
  XOR U19733 ( .A(n17686), .B(n17687), .Z(n17674) );
  AND U19734 ( .A(n17688), .B(n17689), .Z(n17687) );
  XNOR U19735 ( .A(n17686), .B(n8845), .Z(n17689) );
  XNOR U19736 ( .A(n17682), .B(n17684), .Z(n8845) );
  NAND U19737 ( .A(n17690), .B(nreg[576]), .Z(n17684) );
  NAND U19738 ( .A(n12326), .B(nreg[576]), .Z(n17690) );
  XNOR U19739 ( .A(n17680), .B(n17691), .Z(n17682) );
  XOR U19740 ( .A(n17692), .B(n17693), .Z(n17680) );
  AND U19741 ( .A(n17694), .B(n17695), .Z(n17693) );
  XNOR U19742 ( .A(n17696), .B(n17692), .Z(n17695) );
  XOR U19743 ( .A(n17697), .B(nreg[576]), .Z(n17688) );
  IV U19744 ( .A(n17686), .Z(n17697) );
  XOR U19745 ( .A(n17698), .B(n17699), .Z(n17686) );
  AND U19746 ( .A(n17700), .B(n17701), .Z(n17699) );
  XNOR U19747 ( .A(n17698), .B(n8851), .Z(n17701) );
  XNOR U19748 ( .A(n17694), .B(n17696), .Z(n8851) );
  NAND U19749 ( .A(n17702), .B(nreg[575]), .Z(n17696) );
  NAND U19750 ( .A(n12326), .B(nreg[575]), .Z(n17702) );
  XNOR U19751 ( .A(n17692), .B(n17703), .Z(n17694) );
  XOR U19752 ( .A(n17704), .B(n17705), .Z(n17692) );
  AND U19753 ( .A(n17706), .B(n17707), .Z(n17705) );
  XNOR U19754 ( .A(n17708), .B(n17704), .Z(n17707) );
  XOR U19755 ( .A(n17709), .B(nreg[575]), .Z(n17700) );
  IV U19756 ( .A(n17698), .Z(n17709) );
  XOR U19757 ( .A(n17710), .B(n17711), .Z(n17698) );
  AND U19758 ( .A(n17712), .B(n17713), .Z(n17711) );
  XNOR U19759 ( .A(n17710), .B(n8857), .Z(n17713) );
  XNOR U19760 ( .A(n17706), .B(n17708), .Z(n8857) );
  NAND U19761 ( .A(n17714), .B(nreg[574]), .Z(n17708) );
  NAND U19762 ( .A(n12326), .B(nreg[574]), .Z(n17714) );
  XNOR U19763 ( .A(n17704), .B(n17715), .Z(n17706) );
  XOR U19764 ( .A(n17716), .B(n17717), .Z(n17704) );
  AND U19765 ( .A(n17718), .B(n17719), .Z(n17717) );
  XNOR U19766 ( .A(n17720), .B(n17716), .Z(n17719) );
  XOR U19767 ( .A(n17721), .B(nreg[574]), .Z(n17712) );
  IV U19768 ( .A(n17710), .Z(n17721) );
  XOR U19769 ( .A(n17722), .B(n17723), .Z(n17710) );
  AND U19770 ( .A(n17724), .B(n17725), .Z(n17723) );
  XNOR U19771 ( .A(n17722), .B(n8863), .Z(n17725) );
  XNOR U19772 ( .A(n17718), .B(n17720), .Z(n8863) );
  NAND U19773 ( .A(n17726), .B(nreg[573]), .Z(n17720) );
  NAND U19774 ( .A(n12326), .B(nreg[573]), .Z(n17726) );
  XNOR U19775 ( .A(n17716), .B(n17727), .Z(n17718) );
  XOR U19776 ( .A(n17728), .B(n17729), .Z(n17716) );
  AND U19777 ( .A(n17730), .B(n17731), .Z(n17729) );
  XNOR U19778 ( .A(n17732), .B(n17728), .Z(n17731) );
  XOR U19779 ( .A(n17733), .B(nreg[573]), .Z(n17724) );
  IV U19780 ( .A(n17722), .Z(n17733) );
  XOR U19781 ( .A(n17734), .B(n17735), .Z(n17722) );
  AND U19782 ( .A(n17736), .B(n17737), .Z(n17735) );
  XNOR U19783 ( .A(n17734), .B(n8869), .Z(n17737) );
  XNOR U19784 ( .A(n17730), .B(n17732), .Z(n8869) );
  NAND U19785 ( .A(n17738), .B(nreg[572]), .Z(n17732) );
  NAND U19786 ( .A(n12326), .B(nreg[572]), .Z(n17738) );
  XNOR U19787 ( .A(n17728), .B(n17739), .Z(n17730) );
  XOR U19788 ( .A(n17740), .B(n17741), .Z(n17728) );
  AND U19789 ( .A(n17742), .B(n17743), .Z(n17741) );
  XNOR U19790 ( .A(n17744), .B(n17740), .Z(n17743) );
  XOR U19791 ( .A(n17745), .B(nreg[572]), .Z(n17736) );
  IV U19792 ( .A(n17734), .Z(n17745) );
  XOR U19793 ( .A(n17746), .B(n17747), .Z(n17734) );
  AND U19794 ( .A(n17748), .B(n17749), .Z(n17747) );
  XNOR U19795 ( .A(n17746), .B(n8875), .Z(n17749) );
  XNOR U19796 ( .A(n17742), .B(n17744), .Z(n8875) );
  NAND U19797 ( .A(n17750), .B(nreg[571]), .Z(n17744) );
  NAND U19798 ( .A(n12326), .B(nreg[571]), .Z(n17750) );
  XNOR U19799 ( .A(n17740), .B(n17751), .Z(n17742) );
  XOR U19800 ( .A(n17752), .B(n17753), .Z(n17740) );
  AND U19801 ( .A(n17754), .B(n17755), .Z(n17753) );
  XNOR U19802 ( .A(n17756), .B(n17752), .Z(n17755) );
  XOR U19803 ( .A(n17757), .B(nreg[571]), .Z(n17748) );
  IV U19804 ( .A(n17746), .Z(n17757) );
  XOR U19805 ( .A(n17758), .B(n17759), .Z(n17746) );
  AND U19806 ( .A(n17760), .B(n17761), .Z(n17759) );
  XNOR U19807 ( .A(n17758), .B(n8881), .Z(n17761) );
  XNOR U19808 ( .A(n17754), .B(n17756), .Z(n8881) );
  NAND U19809 ( .A(n17762), .B(nreg[570]), .Z(n17756) );
  NAND U19810 ( .A(n12326), .B(nreg[570]), .Z(n17762) );
  XNOR U19811 ( .A(n17752), .B(n17763), .Z(n17754) );
  XOR U19812 ( .A(n17764), .B(n17765), .Z(n17752) );
  AND U19813 ( .A(n17766), .B(n17767), .Z(n17765) );
  XNOR U19814 ( .A(n17768), .B(n17764), .Z(n17767) );
  XOR U19815 ( .A(n17769), .B(nreg[570]), .Z(n17760) );
  IV U19816 ( .A(n17758), .Z(n17769) );
  XOR U19817 ( .A(n17770), .B(n17771), .Z(n17758) );
  AND U19818 ( .A(n17772), .B(n17773), .Z(n17771) );
  XNOR U19819 ( .A(n17770), .B(n8887), .Z(n17773) );
  XNOR U19820 ( .A(n17766), .B(n17768), .Z(n8887) );
  NAND U19821 ( .A(n17774), .B(nreg[569]), .Z(n17768) );
  NAND U19822 ( .A(n12326), .B(nreg[569]), .Z(n17774) );
  XNOR U19823 ( .A(n17764), .B(n17775), .Z(n17766) );
  XOR U19824 ( .A(n17776), .B(n17777), .Z(n17764) );
  AND U19825 ( .A(n17778), .B(n17779), .Z(n17777) );
  XNOR U19826 ( .A(n17780), .B(n17776), .Z(n17779) );
  XOR U19827 ( .A(n17781), .B(nreg[569]), .Z(n17772) );
  IV U19828 ( .A(n17770), .Z(n17781) );
  XOR U19829 ( .A(n17782), .B(n17783), .Z(n17770) );
  AND U19830 ( .A(n17784), .B(n17785), .Z(n17783) );
  XNOR U19831 ( .A(n17782), .B(n8893), .Z(n17785) );
  XNOR U19832 ( .A(n17778), .B(n17780), .Z(n8893) );
  NAND U19833 ( .A(n17786), .B(nreg[568]), .Z(n17780) );
  NAND U19834 ( .A(n12326), .B(nreg[568]), .Z(n17786) );
  XNOR U19835 ( .A(n17776), .B(n17787), .Z(n17778) );
  XOR U19836 ( .A(n17788), .B(n17789), .Z(n17776) );
  AND U19837 ( .A(n17790), .B(n17791), .Z(n17789) );
  XNOR U19838 ( .A(n17792), .B(n17788), .Z(n17791) );
  XOR U19839 ( .A(n17793), .B(nreg[568]), .Z(n17784) );
  IV U19840 ( .A(n17782), .Z(n17793) );
  XOR U19841 ( .A(n17794), .B(n17795), .Z(n17782) );
  AND U19842 ( .A(n17796), .B(n17797), .Z(n17795) );
  XNOR U19843 ( .A(n17794), .B(n8899), .Z(n17797) );
  XNOR U19844 ( .A(n17790), .B(n17792), .Z(n8899) );
  NAND U19845 ( .A(n17798), .B(nreg[567]), .Z(n17792) );
  NAND U19846 ( .A(n12326), .B(nreg[567]), .Z(n17798) );
  XNOR U19847 ( .A(n17788), .B(n17799), .Z(n17790) );
  XOR U19848 ( .A(n17800), .B(n17801), .Z(n17788) );
  AND U19849 ( .A(n17802), .B(n17803), .Z(n17801) );
  XNOR U19850 ( .A(n17804), .B(n17800), .Z(n17803) );
  XOR U19851 ( .A(n17805), .B(nreg[567]), .Z(n17796) );
  IV U19852 ( .A(n17794), .Z(n17805) );
  XOR U19853 ( .A(n17806), .B(n17807), .Z(n17794) );
  AND U19854 ( .A(n17808), .B(n17809), .Z(n17807) );
  XNOR U19855 ( .A(n17806), .B(n8905), .Z(n17809) );
  XNOR U19856 ( .A(n17802), .B(n17804), .Z(n8905) );
  NAND U19857 ( .A(n17810), .B(nreg[566]), .Z(n17804) );
  NAND U19858 ( .A(n12326), .B(nreg[566]), .Z(n17810) );
  XNOR U19859 ( .A(n17800), .B(n17811), .Z(n17802) );
  XOR U19860 ( .A(n17812), .B(n17813), .Z(n17800) );
  AND U19861 ( .A(n17814), .B(n17815), .Z(n17813) );
  XNOR U19862 ( .A(n17816), .B(n17812), .Z(n17815) );
  XOR U19863 ( .A(n17817), .B(nreg[566]), .Z(n17808) );
  IV U19864 ( .A(n17806), .Z(n17817) );
  XOR U19865 ( .A(n17818), .B(n17819), .Z(n17806) );
  AND U19866 ( .A(n17820), .B(n17821), .Z(n17819) );
  XNOR U19867 ( .A(n17818), .B(n8911), .Z(n17821) );
  XNOR U19868 ( .A(n17814), .B(n17816), .Z(n8911) );
  NAND U19869 ( .A(n17822), .B(nreg[565]), .Z(n17816) );
  NAND U19870 ( .A(n12326), .B(nreg[565]), .Z(n17822) );
  XNOR U19871 ( .A(n17812), .B(n17823), .Z(n17814) );
  XOR U19872 ( .A(n17824), .B(n17825), .Z(n17812) );
  AND U19873 ( .A(n17826), .B(n17827), .Z(n17825) );
  XNOR U19874 ( .A(n17828), .B(n17824), .Z(n17827) );
  XOR U19875 ( .A(n17829), .B(nreg[565]), .Z(n17820) );
  IV U19876 ( .A(n17818), .Z(n17829) );
  XOR U19877 ( .A(n17830), .B(n17831), .Z(n17818) );
  AND U19878 ( .A(n17832), .B(n17833), .Z(n17831) );
  XNOR U19879 ( .A(n17830), .B(n8917), .Z(n17833) );
  XNOR U19880 ( .A(n17826), .B(n17828), .Z(n8917) );
  NAND U19881 ( .A(n17834), .B(nreg[564]), .Z(n17828) );
  NAND U19882 ( .A(n12326), .B(nreg[564]), .Z(n17834) );
  XNOR U19883 ( .A(n17824), .B(n17835), .Z(n17826) );
  XOR U19884 ( .A(n17836), .B(n17837), .Z(n17824) );
  AND U19885 ( .A(n17838), .B(n17839), .Z(n17837) );
  XNOR U19886 ( .A(n17840), .B(n17836), .Z(n17839) );
  XOR U19887 ( .A(n17841), .B(nreg[564]), .Z(n17832) );
  IV U19888 ( .A(n17830), .Z(n17841) );
  XOR U19889 ( .A(n17842), .B(n17843), .Z(n17830) );
  AND U19890 ( .A(n17844), .B(n17845), .Z(n17843) );
  XNOR U19891 ( .A(n17842), .B(n8923), .Z(n17845) );
  XNOR U19892 ( .A(n17838), .B(n17840), .Z(n8923) );
  NAND U19893 ( .A(n17846), .B(nreg[563]), .Z(n17840) );
  NAND U19894 ( .A(n12326), .B(nreg[563]), .Z(n17846) );
  XNOR U19895 ( .A(n17836), .B(n17847), .Z(n17838) );
  XOR U19896 ( .A(n17848), .B(n17849), .Z(n17836) );
  AND U19897 ( .A(n17850), .B(n17851), .Z(n17849) );
  XNOR U19898 ( .A(n17852), .B(n17848), .Z(n17851) );
  XOR U19899 ( .A(n17853), .B(nreg[563]), .Z(n17844) );
  IV U19900 ( .A(n17842), .Z(n17853) );
  XOR U19901 ( .A(n17854), .B(n17855), .Z(n17842) );
  AND U19902 ( .A(n17856), .B(n17857), .Z(n17855) );
  XNOR U19903 ( .A(n17854), .B(n8929), .Z(n17857) );
  XNOR U19904 ( .A(n17850), .B(n17852), .Z(n8929) );
  NAND U19905 ( .A(n17858), .B(nreg[562]), .Z(n17852) );
  NAND U19906 ( .A(n12326), .B(nreg[562]), .Z(n17858) );
  XNOR U19907 ( .A(n17848), .B(n17859), .Z(n17850) );
  XOR U19908 ( .A(n17860), .B(n17861), .Z(n17848) );
  AND U19909 ( .A(n17862), .B(n17863), .Z(n17861) );
  XNOR U19910 ( .A(n17864), .B(n17860), .Z(n17863) );
  XOR U19911 ( .A(n17865), .B(nreg[562]), .Z(n17856) );
  IV U19912 ( .A(n17854), .Z(n17865) );
  XOR U19913 ( .A(n17866), .B(n17867), .Z(n17854) );
  AND U19914 ( .A(n17868), .B(n17869), .Z(n17867) );
  XNOR U19915 ( .A(n17866), .B(n8935), .Z(n17869) );
  XNOR U19916 ( .A(n17862), .B(n17864), .Z(n8935) );
  NAND U19917 ( .A(n17870), .B(nreg[561]), .Z(n17864) );
  NAND U19918 ( .A(n12326), .B(nreg[561]), .Z(n17870) );
  XNOR U19919 ( .A(n17860), .B(n17871), .Z(n17862) );
  XOR U19920 ( .A(n17872), .B(n17873), .Z(n17860) );
  AND U19921 ( .A(n17874), .B(n17875), .Z(n17873) );
  XNOR U19922 ( .A(n17876), .B(n17872), .Z(n17875) );
  XOR U19923 ( .A(n17877), .B(nreg[561]), .Z(n17868) );
  IV U19924 ( .A(n17866), .Z(n17877) );
  XOR U19925 ( .A(n17878), .B(n17879), .Z(n17866) );
  AND U19926 ( .A(n17880), .B(n17881), .Z(n17879) );
  XNOR U19927 ( .A(n17878), .B(n8941), .Z(n17881) );
  XNOR U19928 ( .A(n17874), .B(n17876), .Z(n8941) );
  NAND U19929 ( .A(n17882), .B(nreg[560]), .Z(n17876) );
  NAND U19930 ( .A(n12326), .B(nreg[560]), .Z(n17882) );
  XNOR U19931 ( .A(n17872), .B(n17883), .Z(n17874) );
  XOR U19932 ( .A(n17884), .B(n17885), .Z(n17872) );
  AND U19933 ( .A(n17886), .B(n17887), .Z(n17885) );
  XNOR U19934 ( .A(n17888), .B(n17884), .Z(n17887) );
  XOR U19935 ( .A(n17889), .B(nreg[560]), .Z(n17880) );
  IV U19936 ( .A(n17878), .Z(n17889) );
  XOR U19937 ( .A(n17890), .B(n17891), .Z(n17878) );
  AND U19938 ( .A(n17892), .B(n17893), .Z(n17891) );
  XNOR U19939 ( .A(n17890), .B(n8947), .Z(n17893) );
  XNOR U19940 ( .A(n17886), .B(n17888), .Z(n8947) );
  NAND U19941 ( .A(n17894), .B(nreg[559]), .Z(n17888) );
  NAND U19942 ( .A(n12326), .B(nreg[559]), .Z(n17894) );
  XNOR U19943 ( .A(n17884), .B(n17895), .Z(n17886) );
  XOR U19944 ( .A(n17896), .B(n17897), .Z(n17884) );
  AND U19945 ( .A(n17898), .B(n17899), .Z(n17897) );
  XNOR U19946 ( .A(n17900), .B(n17896), .Z(n17899) );
  XOR U19947 ( .A(n17901), .B(nreg[559]), .Z(n17892) );
  IV U19948 ( .A(n17890), .Z(n17901) );
  XOR U19949 ( .A(n17902), .B(n17903), .Z(n17890) );
  AND U19950 ( .A(n17904), .B(n17905), .Z(n17903) );
  XNOR U19951 ( .A(n17902), .B(n8953), .Z(n17905) );
  XNOR U19952 ( .A(n17898), .B(n17900), .Z(n8953) );
  NAND U19953 ( .A(n17906), .B(nreg[558]), .Z(n17900) );
  NAND U19954 ( .A(n12326), .B(nreg[558]), .Z(n17906) );
  XNOR U19955 ( .A(n17896), .B(n17907), .Z(n17898) );
  XOR U19956 ( .A(n17908), .B(n17909), .Z(n17896) );
  AND U19957 ( .A(n17910), .B(n17911), .Z(n17909) );
  XNOR U19958 ( .A(n17912), .B(n17908), .Z(n17911) );
  XOR U19959 ( .A(n17913), .B(nreg[558]), .Z(n17904) );
  IV U19960 ( .A(n17902), .Z(n17913) );
  XOR U19961 ( .A(n17914), .B(n17915), .Z(n17902) );
  AND U19962 ( .A(n17916), .B(n17917), .Z(n17915) );
  XNOR U19963 ( .A(n17914), .B(n8959), .Z(n17917) );
  XNOR U19964 ( .A(n17910), .B(n17912), .Z(n8959) );
  NAND U19965 ( .A(n17918), .B(nreg[557]), .Z(n17912) );
  NAND U19966 ( .A(n12326), .B(nreg[557]), .Z(n17918) );
  XNOR U19967 ( .A(n17908), .B(n17919), .Z(n17910) );
  XOR U19968 ( .A(n17920), .B(n17921), .Z(n17908) );
  AND U19969 ( .A(n17922), .B(n17923), .Z(n17921) );
  XNOR U19970 ( .A(n17924), .B(n17920), .Z(n17923) );
  XOR U19971 ( .A(n17925), .B(nreg[557]), .Z(n17916) );
  IV U19972 ( .A(n17914), .Z(n17925) );
  XOR U19973 ( .A(n17926), .B(n17927), .Z(n17914) );
  AND U19974 ( .A(n17928), .B(n17929), .Z(n17927) );
  XNOR U19975 ( .A(n17926), .B(n8965), .Z(n17929) );
  XNOR U19976 ( .A(n17922), .B(n17924), .Z(n8965) );
  NAND U19977 ( .A(n17930), .B(nreg[556]), .Z(n17924) );
  NAND U19978 ( .A(n12326), .B(nreg[556]), .Z(n17930) );
  XNOR U19979 ( .A(n17920), .B(n17931), .Z(n17922) );
  XOR U19980 ( .A(n17932), .B(n17933), .Z(n17920) );
  AND U19981 ( .A(n17934), .B(n17935), .Z(n17933) );
  XNOR U19982 ( .A(n17936), .B(n17932), .Z(n17935) );
  XOR U19983 ( .A(n17937), .B(nreg[556]), .Z(n17928) );
  IV U19984 ( .A(n17926), .Z(n17937) );
  XOR U19985 ( .A(n17938), .B(n17939), .Z(n17926) );
  AND U19986 ( .A(n17940), .B(n17941), .Z(n17939) );
  XNOR U19987 ( .A(n17938), .B(n8971), .Z(n17941) );
  XNOR U19988 ( .A(n17934), .B(n17936), .Z(n8971) );
  NAND U19989 ( .A(n17942), .B(nreg[555]), .Z(n17936) );
  NAND U19990 ( .A(n12326), .B(nreg[555]), .Z(n17942) );
  XNOR U19991 ( .A(n17932), .B(n17943), .Z(n17934) );
  XOR U19992 ( .A(n17944), .B(n17945), .Z(n17932) );
  AND U19993 ( .A(n17946), .B(n17947), .Z(n17945) );
  XNOR U19994 ( .A(n17948), .B(n17944), .Z(n17947) );
  XOR U19995 ( .A(n17949), .B(nreg[555]), .Z(n17940) );
  IV U19996 ( .A(n17938), .Z(n17949) );
  XOR U19997 ( .A(n17950), .B(n17951), .Z(n17938) );
  AND U19998 ( .A(n17952), .B(n17953), .Z(n17951) );
  XNOR U19999 ( .A(n17950), .B(n8977), .Z(n17953) );
  XNOR U20000 ( .A(n17946), .B(n17948), .Z(n8977) );
  NAND U20001 ( .A(n17954), .B(nreg[554]), .Z(n17948) );
  NAND U20002 ( .A(n12326), .B(nreg[554]), .Z(n17954) );
  XNOR U20003 ( .A(n17944), .B(n17955), .Z(n17946) );
  XOR U20004 ( .A(n17956), .B(n17957), .Z(n17944) );
  AND U20005 ( .A(n17958), .B(n17959), .Z(n17957) );
  XNOR U20006 ( .A(n17960), .B(n17956), .Z(n17959) );
  XOR U20007 ( .A(n17961), .B(nreg[554]), .Z(n17952) );
  IV U20008 ( .A(n17950), .Z(n17961) );
  XOR U20009 ( .A(n17962), .B(n17963), .Z(n17950) );
  AND U20010 ( .A(n17964), .B(n17965), .Z(n17963) );
  XNOR U20011 ( .A(n17962), .B(n8983), .Z(n17965) );
  XNOR U20012 ( .A(n17958), .B(n17960), .Z(n8983) );
  NAND U20013 ( .A(n17966), .B(nreg[553]), .Z(n17960) );
  NAND U20014 ( .A(n12326), .B(nreg[553]), .Z(n17966) );
  XNOR U20015 ( .A(n17956), .B(n17967), .Z(n17958) );
  XOR U20016 ( .A(n17968), .B(n17969), .Z(n17956) );
  AND U20017 ( .A(n17970), .B(n17971), .Z(n17969) );
  XNOR U20018 ( .A(n17972), .B(n17968), .Z(n17971) );
  XOR U20019 ( .A(n17973), .B(nreg[553]), .Z(n17964) );
  IV U20020 ( .A(n17962), .Z(n17973) );
  XOR U20021 ( .A(n17974), .B(n17975), .Z(n17962) );
  AND U20022 ( .A(n17976), .B(n17977), .Z(n17975) );
  XNOR U20023 ( .A(n17974), .B(n8989), .Z(n17977) );
  XNOR U20024 ( .A(n17970), .B(n17972), .Z(n8989) );
  NAND U20025 ( .A(n17978), .B(nreg[552]), .Z(n17972) );
  NAND U20026 ( .A(n12326), .B(nreg[552]), .Z(n17978) );
  XNOR U20027 ( .A(n17968), .B(n17979), .Z(n17970) );
  XOR U20028 ( .A(n17980), .B(n17981), .Z(n17968) );
  AND U20029 ( .A(n17982), .B(n17983), .Z(n17981) );
  XNOR U20030 ( .A(n17984), .B(n17980), .Z(n17983) );
  XOR U20031 ( .A(n17985), .B(nreg[552]), .Z(n17976) );
  IV U20032 ( .A(n17974), .Z(n17985) );
  XOR U20033 ( .A(n17986), .B(n17987), .Z(n17974) );
  AND U20034 ( .A(n17988), .B(n17989), .Z(n17987) );
  XNOR U20035 ( .A(n17986), .B(n8995), .Z(n17989) );
  XNOR U20036 ( .A(n17982), .B(n17984), .Z(n8995) );
  NAND U20037 ( .A(n17990), .B(nreg[551]), .Z(n17984) );
  NAND U20038 ( .A(n12326), .B(nreg[551]), .Z(n17990) );
  XNOR U20039 ( .A(n17980), .B(n17991), .Z(n17982) );
  XOR U20040 ( .A(n17992), .B(n17993), .Z(n17980) );
  AND U20041 ( .A(n17994), .B(n17995), .Z(n17993) );
  XNOR U20042 ( .A(n17996), .B(n17992), .Z(n17995) );
  XOR U20043 ( .A(n17997), .B(nreg[551]), .Z(n17988) );
  IV U20044 ( .A(n17986), .Z(n17997) );
  XOR U20045 ( .A(n17998), .B(n17999), .Z(n17986) );
  AND U20046 ( .A(n18000), .B(n18001), .Z(n17999) );
  XNOR U20047 ( .A(n17998), .B(n9001), .Z(n18001) );
  XNOR U20048 ( .A(n17994), .B(n17996), .Z(n9001) );
  NAND U20049 ( .A(n18002), .B(nreg[550]), .Z(n17996) );
  NAND U20050 ( .A(n12326), .B(nreg[550]), .Z(n18002) );
  XNOR U20051 ( .A(n17992), .B(n18003), .Z(n17994) );
  XOR U20052 ( .A(n18004), .B(n18005), .Z(n17992) );
  AND U20053 ( .A(n18006), .B(n18007), .Z(n18005) );
  XNOR U20054 ( .A(n18008), .B(n18004), .Z(n18007) );
  XOR U20055 ( .A(n18009), .B(nreg[550]), .Z(n18000) );
  IV U20056 ( .A(n17998), .Z(n18009) );
  XOR U20057 ( .A(n18010), .B(n18011), .Z(n17998) );
  AND U20058 ( .A(n18012), .B(n18013), .Z(n18011) );
  XNOR U20059 ( .A(n18010), .B(n9007), .Z(n18013) );
  XNOR U20060 ( .A(n18006), .B(n18008), .Z(n9007) );
  NAND U20061 ( .A(n18014), .B(nreg[549]), .Z(n18008) );
  NAND U20062 ( .A(n12326), .B(nreg[549]), .Z(n18014) );
  XNOR U20063 ( .A(n18004), .B(n18015), .Z(n18006) );
  XOR U20064 ( .A(n18016), .B(n18017), .Z(n18004) );
  AND U20065 ( .A(n18018), .B(n18019), .Z(n18017) );
  XNOR U20066 ( .A(n18020), .B(n18016), .Z(n18019) );
  XOR U20067 ( .A(n18021), .B(nreg[549]), .Z(n18012) );
  IV U20068 ( .A(n18010), .Z(n18021) );
  XOR U20069 ( .A(n18022), .B(n18023), .Z(n18010) );
  AND U20070 ( .A(n18024), .B(n18025), .Z(n18023) );
  XNOR U20071 ( .A(n18022), .B(n9013), .Z(n18025) );
  XNOR U20072 ( .A(n18018), .B(n18020), .Z(n9013) );
  NAND U20073 ( .A(n18026), .B(nreg[548]), .Z(n18020) );
  NAND U20074 ( .A(n12326), .B(nreg[548]), .Z(n18026) );
  XNOR U20075 ( .A(n18016), .B(n18027), .Z(n18018) );
  XOR U20076 ( .A(n18028), .B(n18029), .Z(n18016) );
  AND U20077 ( .A(n18030), .B(n18031), .Z(n18029) );
  XNOR U20078 ( .A(n18032), .B(n18028), .Z(n18031) );
  XOR U20079 ( .A(n18033), .B(nreg[548]), .Z(n18024) );
  IV U20080 ( .A(n18022), .Z(n18033) );
  XOR U20081 ( .A(n18034), .B(n18035), .Z(n18022) );
  AND U20082 ( .A(n18036), .B(n18037), .Z(n18035) );
  XNOR U20083 ( .A(n18034), .B(n9019), .Z(n18037) );
  XNOR U20084 ( .A(n18030), .B(n18032), .Z(n9019) );
  NAND U20085 ( .A(n18038), .B(nreg[547]), .Z(n18032) );
  NAND U20086 ( .A(n12326), .B(nreg[547]), .Z(n18038) );
  XNOR U20087 ( .A(n18028), .B(n18039), .Z(n18030) );
  XOR U20088 ( .A(n18040), .B(n18041), .Z(n18028) );
  AND U20089 ( .A(n18042), .B(n18043), .Z(n18041) );
  XNOR U20090 ( .A(n18044), .B(n18040), .Z(n18043) );
  XOR U20091 ( .A(n18045), .B(nreg[547]), .Z(n18036) );
  IV U20092 ( .A(n18034), .Z(n18045) );
  XOR U20093 ( .A(n18046), .B(n18047), .Z(n18034) );
  AND U20094 ( .A(n18048), .B(n18049), .Z(n18047) );
  XNOR U20095 ( .A(n18046), .B(n9025), .Z(n18049) );
  XNOR U20096 ( .A(n18042), .B(n18044), .Z(n9025) );
  NAND U20097 ( .A(n18050), .B(nreg[546]), .Z(n18044) );
  NAND U20098 ( .A(n12326), .B(nreg[546]), .Z(n18050) );
  XNOR U20099 ( .A(n18040), .B(n18051), .Z(n18042) );
  XOR U20100 ( .A(n18052), .B(n18053), .Z(n18040) );
  AND U20101 ( .A(n18054), .B(n18055), .Z(n18053) );
  XNOR U20102 ( .A(n18056), .B(n18052), .Z(n18055) );
  XOR U20103 ( .A(n18057), .B(nreg[546]), .Z(n18048) );
  IV U20104 ( .A(n18046), .Z(n18057) );
  XOR U20105 ( .A(n18058), .B(n18059), .Z(n18046) );
  AND U20106 ( .A(n18060), .B(n18061), .Z(n18059) );
  XNOR U20107 ( .A(n18058), .B(n9031), .Z(n18061) );
  XNOR U20108 ( .A(n18054), .B(n18056), .Z(n9031) );
  NAND U20109 ( .A(n18062), .B(nreg[545]), .Z(n18056) );
  NAND U20110 ( .A(n12326), .B(nreg[545]), .Z(n18062) );
  XNOR U20111 ( .A(n18052), .B(n18063), .Z(n18054) );
  XOR U20112 ( .A(n18064), .B(n18065), .Z(n18052) );
  AND U20113 ( .A(n18066), .B(n18067), .Z(n18065) );
  XNOR U20114 ( .A(n18068), .B(n18064), .Z(n18067) );
  XOR U20115 ( .A(n18069), .B(nreg[545]), .Z(n18060) );
  IV U20116 ( .A(n18058), .Z(n18069) );
  XOR U20117 ( .A(n18070), .B(n18071), .Z(n18058) );
  AND U20118 ( .A(n18072), .B(n18073), .Z(n18071) );
  XNOR U20119 ( .A(n18070), .B(n9037), .Z(n18073) );
  XNOR U20120 ( .A(n18066), .B(n18068), .Z(n9037) );
  NAND U20121 ( .A(n18074), .B(nreg[544]), .Z(n18068) );
  NAND U20122 ( .A(n12326), .B(nreg[544]), .Z(n18074) );
  XNOR U20123 ( .A(n18064), .B(n18075), .Z(n18066) );
  XOR U20124 ( .A(n18076), .B(n18077), .Z(n18064) );
  AND U20125 ( .A(n18078), .B(n18079), .Z(n18077) );
  XNOR U20126 ( .A(n18080), .B(n18076), .Z(n18079) );
  XOR U20127 ( .A(n18081), .B(nreg[544]), .Z(n18072) );
  IV U20128 ( .A(n18070), .Z(n18081) );
  XOR U20129 ( .A(n18082), .B(n18083), .Z(n18070) );
  AND U20130 ( .A(n18084), .B(n18085), .Z(n18083) );
  XNOR U20131 ( .A(n18082), .B(n9043), .Z(n18085) );
  XNOR U20132 ( .A(n18078), .B(n18080), .Z(n9043) );
  NAND U20133 ( .A(n18086), .B(nreg[543]), .Z(n18080) );
  NAND U20134 ( .A(n12326), .B(nreg[543]), .Z(n18086) );
  XNOR U20135 ( .A(n18076), .B(n18087), .Z(n18078) );
  XOR U20136 ( .A(n18088), .B(n18089), .Z(n18076) );
  AND U20137 ( .A(n18090), .B(n18091), .Z(n18089) );
  XNOR U20138 ( .A(n18092), .B(n18088), .Z(n18091) );
  XOR U20139 ( .A(n18093), .B(nreg[543]), .Z(n18084) );
  IV U20140 ( .A(n18082), .Z(n18093) );
  XOR U20141 ( .A(n18094), .B(n18095), .Z(n18082) );
  AND U20142 ( .A(n18096), .B(n18097), .Z(n18095) );
  XNOR U20143 ( .A(n18094), .B(n9049), .Z(n18097) );
  XNOR U20144 ( .A(n18090), .B(n18092), .Z(n9049) );
  NAND U20145 ( .A(n18098), .B(nreg[542]), .Z(n18092) );
  NAND U20146 ( .A(n12326), .B(nreg[542]), .Z(n18098) );
  XNOR U20147 ( .A(n18088), .B(n18099), .Z(n18090) );
  XOR U20148 ( .A(n18100), .B(n18101), .Z(n18088) );
  AND U20149 ( .A(n18102), .B(n18103), .Z(n18101) );
  XNOR U20150 ( .A(n18104), .B(n18100), .Z(n18103) );
  XOR U20151 ( .A(n18105), .B(nreg[542]), .Z(n18096) );
  IV U20152 ( .A(n18094), .Z(n18105) );
  XOR U20153 ( .A(n18106), .B(n18107), .Z(n18094) );
  AND U20154 ( .A(n18108), .B(n18109), .Z(n18107) );
  XNOR U20155 ( .A(n18106), .B(n9055), .Z(n18109) );
  XNOR U20156 ( .A(n18102), .B(n18104), .Z(n9055) );
  NAND U20157 ( .A(n18110), .B(nreg[541]), .Z(n18104) );
  NAND U20158 ( .A(n12326), .B(nreg[541]), .Z(n18110) );
  XNOR U20159 ( .A(n18100), .B(n18111), .Z(n18102) );
  XOR U20160 ( .A(n18112), .B(n18113), .Z(n18100) );
  AND U20161 ( .A(n18114), .B(n18115), .Z(n18113) );
  XNOR U20162 ( .A(n18116), .B(n18112), .Z(n18115) );
  XOR U20163 ( .A(n18117), .B(nreg[541]), .Z(n18108) );
  IV U20164 ( .A(n18106), .Z(n18117) );
  XOR U20165 ( .A(n18118), .B(n18119), .Z(n18106) );
  AND U20166 ( .A(n18120), .B(n18121), .Z(n18119) );
  XNOR U20167 ( .A(n18118), .B(n9061), .Z(n18121) );
  XNOR U20168 ( .A(n18114), .B(n18116), .Z(n9061) );
  NAND U20169 ( .A(n18122), .B(nreg[540]), .Z(n18116) );
  NAND U20170 ( .A(n12326), .B(nreg[540]), .Z(n18122) );
  XNOR U20171 ( .A(n18112), .B(n18123), .Z(n18114) );
  XOR U20172 ( .A(n18124), .B(n18125), .Z(n18112) );
  AND U20173 ( .A(n18126), .B(n18127), .Z(n18125) );
  XNOR U20174 ( .A(n18128), .B(n18124), .Z(n18127) );
  XOR U20175 ( .A(n18129), .B(nreg[540]), .Z(n18120) );
  IV U20176 ( .A(n18118), .Z(n18129) );
  XOR U20177 ( .A(n18130), .B(n18131), .Z(n18118) );
  AND U20178 ( .A(n18132), .B(n18133), .Z(n18131) );
  XNOR U20179 ( .A(n18130), .B(n9067), .Z(n18133) );
  XNOR U20180 ( .A(n18126), .B(n18128), .Z(n9067) );
  NAND U20181 ( .A(n18134), .B(nreg[539]), .Z(n18128) );
  NAND U20182 ( .A(n12326), .B(nreg[539]), .Z(n18134) );
  XNOR U20183 ( .A(n18124), .B(n18135), .Z(n18126) );
  XOR U20184 ( .A(n18136), .B(n18137), .Z(n18124) );
  AND U20185 ( .A(n18138), .B(n18139), .Z(n18137) );
  XNOR U20186 ( .A(n18140), .B(n18136), .Z(n18139) );
  XOR U20187 ( .A(n18141), .B(nreg[539]), .Z(n18132) );
  IV U20188 ( .A(n18130), .Z(n18141) );
  XOR U20189 ( .A(n18142), .B(n18143), .Z(n18130) );
  AND U20190 ( .A(n18144), .B(n18145), .Z(n18143) );
  XNOR U20191 ( .A(n18142), .B(n9073), .Z(n18145) );
  XNOR U20192 ( .A(n18138), .B(n18140), .Z(n9073) );
  NAND U20193 ( .A(n18146), .B(nreg[538]), .Z(n18140) );
  NAND U20194 ( .A(n12326), .B(nreg[538]), .Z(n18146) );
  XNOR U20195 ( .A(n18136), .B(n18147), .Z(n18138) );
  XOR U20196 ( .A(n18148), .B(n18149), .Z(n18136) );
  AND U20197 ( .A(n18150), .B(n18151), .Z(n18149) );
  XNOR U20198 ( .A(n18152), .B(n18148), .Z(n18151) );
  XOR U20199 ( .A(n18153), .B(nreg[538]), .Z(n18144) );
  IV U20200 ( .A(n18142), .Z(n18153) );
  XOR U20201 ( .A(n18154), .B(n18155), .Z(n18142) );
  AND U20202 ( .A(n18156), .B(n18157), .Z(n18155) );
  XNOR U20203 ( .A(n18154), .B(n9079), .Z(n18157) );
  XNOR U20204 ( .A(n18150), .B(n18152), .Z(n9079) );
  NAND U20205 ( .A(n18158), .B(nreg[537]), .Z(n18152) );
  NAND U20206 ( .A(n12326), .B(nreg[537]), .Z(n18158) );
  XNOR U20207 ( .A(n18148), .B(n18159), .Z(n18150) );
  XOR U20208 ( .A(n18160), .B(n18161), .Z(n18148) );
  AND U20209 ( .A(n18162), .B(n18163), .Z(n18161) );
  XNOR U20210 ( .A(n18164), .B(n18160), .Z(n18163) );
  XOR U20211 ( .A(n18165), .B(nreg[537]), .Z(n18156) );
  IV U20212 ( .A(n18154), .Z(n18165) );
  XOR U20213 ( .A(n18166), .B(n18167), .Z(n18154) );
  AND U20214 ( .A(n18168), .B(n18169), .Z(n18167) );
  XNOR U20215 ( .A(n18166), .B(n9085), .Z(n18169) );
  XNOR U20216 ( .A(n18162), .B(n18164), .Z(n9085) );
  NAND U20217 ( .A(n18170), .B(nreg[536]), .Z(n18164) );
  NAND U20218 ( .A(n12326), .B(nreg[536]), .Z(n18170) );
  XNOR U20219 ( .A(n18160), .B(n18171), .Z(n18162) );
  XOR U20220 ( .A(n18172), .B(n18173), .Z(n18160) );
  AND U20221 ( .A(n18174), .B(n18175), .Z(n18173) );
  XNOR U20222 ( .A(n18176), .B(n18172), .Z(n18175) );
  XOR U20223 ( .A(n18177), .B(nreg[536]), .Z(n18168) );
  IV U20224 ( .A(n18166), .Z(n18177) );
  XOR U20225 ( .A(n18178), .B(n18179), .Z(n18166) );
  AND U20226 ( .A(n18180), .B(n18181), .Z(n18179) );
  XNOR U20227 ( .A(n18178), .B(n9091), .Z(n18181) );
  XNOR U20228 ( .A(n18174), .B(n18176), .Z(n9091) );
  NAND U20229 ( .A(n18182), .B(nreg[535]), .Z(n18176) );
  NAND U20230 ( .A(n12326), .B(nreg[535]), .Z(n18182) );
  XNOR U20231 ( .A(n18172), .B(n18183), .Z(n18174) );
  XOR U20232 ( .A(n18184), .B(n18185), .Z(n18172) );
  AND U20233 ( .A(n18186), .B(n18187), .Z(n18185) );
  XNOR U20234 ( .A(n18188), .B(n18184), .Z(n18187) );
  XOR U20235 ( .A(n18189), .B(nreg[535]), .Z(n18180) );
  IV U20236 ( .A(n18178), .Z(n18189) );
  XOR U20237 ( .A(n18190), .B(n18191), .Z(n18178) );
  AND U20238 ( .A(n18192), .B(n18193), .Z(n18191) );
  XNOR U20239 ( .A(n18190), .B(n9097), .Z(n18193) );
  XNOR U20240 ( .A(n18186), .B(n18188), .Z(n9097) );
  NAND U20241 ( .A(n18194), .B(nreg[534]), .Z(n18188) );
  NAND U20242 ( .A(n12326), .B(nreg[534]), .Z(n18194) );
  XNOR U20243 ( .A(n18184), .B(n18195), .Z(n18186) );
  XOR U20244 ( .A(n18196), .B(n18197), .Z(n18184) );
  AND U20245 ( .A(n18198), .B(n18199), .Z(n18197) );
  XNOR U20246 ( .A(n18200), .B(n18196), .Z(n18199) );
  XOR U20247 ( .A(n18201), .B(nreg[534]), .Z(n18192) );
  IV U20248 ( .A(n18190), .Z(n18201) );
  XOR U20249 ( .A(n18202), .B(n18203), .Z(n18190) );
  AND U20250 ( .A(n18204), .B(n18205), .Z(n18203) );
  XNOR U20251 ( .A(n18202), .B(n9103), .Z(n18205) );
  XNOR U20252 ( .A(n18198), .B(n18200), .Z(n9103) );
  NAND U20253 ( .A(n18206), .B(nreg[533]), .Z(n18200) );
  NAND U20254 ( .A(n12326), .B(nreg[533]), .Z(n18206) );
  XNOR U20255 ( .A(n18196), .B(n18207), .Z(n18198) );
  XOR U20256 ( .A(n18208), .B(n18209), .Z(n18196) );
  AND U20257 ( .A(n18210), .B(n18211), .Z(n18209) );
  XNOR U20258 ( .A(n18212), .B(n18208), .Z(n18211) );
  XOR U20259 ( .A(n18213), .B(nreg[533]), .Z(n18204) );
  IV U20260 ( .A(n18202), .Z(n18213) );
  XOR U20261 ( .A(n18214), .B(n18215), .Z(n18202) );
  AND U20262 ( .A(n18216), .B(n18217), .Z(n18215) );
  XNOR U20263 ( .A(n18214), .B(n9109), .Z(n18217) );
  XNOR U20264 ( .A(n18210), .B(n18212), .Z(n9109) );
  NAND U20265 ( .A(n18218), .B(nreg[532]), .Z(n18212) );
  NAND U20266 ( .A(n12326), .B(nreg[532]), .Z(n18218) );
  XNOR U20267 ( .A(n18208), .B(n18219), .Z(n18210) );
  XOR U20268 ( .A(n18220), .B(n18221), .Z(n18208) );
  AND U20269 ( .A(n18222), .B(n18223), .Z(n18221) );
  XNOR U20270 ( .A(n18224), .B(n18220), .Z(n18223) );
  XOR U20271 ( .A(n18225), .B(nreg[532]), .Z(n18216) );
  IV U20272 ( .A(n18214), .Z(n18225) );
  XOR U20273 ( .A(n18226), .B(n18227), .Z(n18214) );
  AND U20274 ( .A(n18228), .B(n18229), .Z(n18227) );
  XNOR U20275 ( .A(n18226), .B(n9115), .Z(n18229) );
  XNOR U20276 ( .A(n18222), .B(n18224), .Z(n9115) );
  NAND U20277 ( .A(n18230), .B(nreg[531]), .Z(n18224) );
  NAND U20278 ( .A(n12326), .B(nreg[531]), .Z(n18230) );
  XNOR U20279 ( .A(n18220), .B(n18231), .Z(n18222) );
  XOR U20280 ( .A(n18232), .B(n18233), .Z(n18220) );
  AND U20281 ( .A(n18234), .B(n18235), .Z(n18233) );
  XNOR U20282 ( .A(n18236), .B(n18232), .Z(n18235) );
  XOR U20283 ( .A(n18237), .B(nreg[531]), .Z(n18228) );
  IV U20284 ( .A(n18226), .Z(n18237) );
  XOR U20285 ( .A(n18238), .B(n18239), .Z(n18226) );
  AND U20286 ( .A(n18240), .B(n18241), .Z(n18239) );
  XNOR U20287 ( .A(n18238), .B(n9121), .Z(n18241) );
  XNOR U20288 ( .A(n18234), .B(n18236), .Z(n9121) );
  NAND U20289 ( .A(n18242), .B(nreg[530]), .Z(n18236) );
  NAND U20290 ( .A(n12326), .B(nreg[530]), .Z(n18242) );
  XNOR U20291 ( .A(n18232), .B(n18243), .Z(n18234) );
  XOR U20292 ( .A(n18244), .B(n18245), .Z(n18232) );
  AND U20293 ( .A(n18246), .B(n18247), .Z(n18245) );
  XNOR U20294 ( .A(n18248), .B(n18244), .Z(n18247) );
  XOR U20295 ( .A(n18249), .B(nreg[530]), .Z(n18240) );
  IV U20296 ( .A(n18238), .Z(n18249) );
  XOR U20297 ( .A(n18250), .B(n18251), .Z(n18238) );
  AND U20298 ( .A(n18252), .B(n18253), .Z(n18251) );
  XNOR U20299 ( .A(n18250), .B(n9127), .Z(n18253) );
  XNOR U20300 ( .A(n18246), .B(n18248), .Z(n9127) );
  NAND U20301 ( .A(n18254), .B(nreg[529]), .Z(n18248) );
  NAND U20302 ( .A(n12326), .B(nreg[529]), .Z(n18254) );
  XNOR U20303 ( .A(n18244), .B(n18255), .Z(n18246) );
  XOR U20304 ( .A(n18256), .B(n18257), .Z(n18244) );
  AND U20305 ( .A(n18258), .B(n18259), .Z(n18257) );
  XNOR U20306 ( .A(n18260), .B(n18256), .Z(n18259) );
  XOR U20307 ( .A(n18261), .B(nreg[529]), .Z(n18252) );
  IV U20308 ( .A(n18250), .Z(n18261) );
  XOR U20309 ( .A(n18262), .B(n18263), .Z(n18250) );
  AND U20310 ( .A(n18264), .B(n18265), .Z(n18263) );
  XNOR U20311 ( .A(n18262), .B(n9133), .Z(n18265) );
  XNOR U20312 ( .A(n18258), .B(n18260), .Z(n9133) );
  NAND U20313 ( .A(n18266), .B(nreg[528]), .Z(n18260) );
  NAND U20314 ( .A(n12326), .B(nreg[528]), .Z(n18266) );
  XNOR U20315 ( .A(n18256), .B(n18267), .Z(n18258) );
  XOR U20316 ( .A(n18268), .B(n18269), .Z(n18256) );
  AND U20317 ( .A(n18270), .B(n18271), .Z(n18269) );
  XNOR U20318 ( .A(n18272), .B(n18268), .Z(n18271) );
  XOR U20319 ( .A(n18273), .B(nreg[528]), .Z(n18264) );
  IV U20320 ( .A(n18262), .Z(n18273) );
  XOR U20321 ( .A(n18274), .B(n18275), .Z(n18262) );
  AND U20322 ( .A(n18276), .B(n18277), .Z(n18275) );
  XNOR U20323 ( .A(n18274), .B(n9139), .Z(n18277) );
  XNOR U20324 ( .A(n18270), .B(n18272), .Z(n9139) );
  NAND U20325 ( .A(n18278), .B(nreg[527]), .Z(n18272) );
  NAND U20326 ( .A(n12326), .B(nreg[527]), .Z(n18278) );
  XNOR U20327 ( .A(n18268), .B(n18279), .Z(n18270) );
  XOR U20328 ( .A(n18280), .B(n18281), .Z(n18268) );
  AND U20329 ( .A(n18282), .B(n18283), .Z(n18281) );
  XNOR U20330 ( .A(n18284), .B(n18280), .Z(n18283) );
  XOR U20331 ( .A(n18285), .B(nreg[527]), .Z(n18276) );
  IV U20332 ( .A(n18274), .Z(n18285) );
  XOR U20333 ( .A(n18286), .B(n18287), .Z(n18274) );
  AND U20334 ( .A(n18288), .B(n18289), .Z(n18287) );
  XNOR U20335 ( .A(n18286), .B(n9145), .Z(n18289) );
  XNOR U20336 ( .A(n18282), .B(n18284), .Z(n9145) );
  NAND U20337 ( .A(n18290), .B(nreg[526]), .Z(n18284) );
  NAND U20338 ( .A(n12326), .B(nreg[526]), .Z(n18290) );
  XNOR U20339 ( .A(n18280), .B(n18291), .Z(n18282) );
  XOR U20340 ( .A(n18292), .B(n18293), .Z(n18280) );
  AND U20341 ( .A(n18294), .B(n18295), .Z(n18293) );
  XNOR U20342 ( .A(n18296), .B(n18292), .Z(n18295) );
  XOR U20343 ( .A(n18297), .B(nreg[526]), .Z(n18288) );
  IV U20344 ( .A(n18286), .Z(n18297) );
  XOR U20345 ( .A(n18298), .B(n18299), .Z(n18286) );
  AND U20346 ( .A(n18300), .B(n18301), .Z(n18299) );
  XNOR U20347 ( .A(n18298), .B(n9151), .Z(n18301) );
  XNOR U20348 ( .A(n18294), .B(n18296), .Z(n9151) );
  NAND U20349 ( .A(n18302), .B(nreg[525]), .Z(n18296) );
  NAND U20350 ( .A(n12326), .B(nreg[525]), .Z(n18302) );
  XNOR U20351 ( .A(n18292), .B(n18303), .Z(n18294) );
  XOR U20352 ( .A(n18304), .B(n18305), .Z(n18292) );
  AND U20353 ( .A(n18306), .B(n18307), .Z(n18305) );
  XNOR U20354 ( .A(n18308), .B(n18304), .Z(n18307) );
  XOR U20355 ( .A(n18309), .B(nreg[525]), .Z(n18300) );
  IV U20356 ( .A(n18298), .Z(n18309) );
  XOR U20357 ( .A(n18310), .B(n18311), .Z(n18298) );
  AND U20358 ( .A(n18312), .B(n18313), .Z(n18311) );
  XNOR U20359 ( .A(n18310), .B(n9157), .Z(n18313) );
  XNOR U20360 ( .A(n18306), .B(n18308), .Z(n9157) );
  NAND U20361 ( .A(n18314), .B(nreg[524]), .Z(n18308) );
  NAND U20362 ( .A(n12326), .B(nreg[524]), .Z(n18314) );
  XNOR U20363 ( .A(n18304), .B(n18315), .Z(n18306) );
  XOR U20364 ( .A(n18316), .B(n18317), .Z(n18304) );
  AND U20365 ( .A(n18318), .B(n18319), .Z(n18317) );
  XNOR U20366 ( .A(n18320), .B(n18316), .Z(n18319) );
  XOR U20367 ( .A(n18321), .B(nreg[524]), .Z(n18312) );
  IV U20368 ( .A(n18310), .Z(n18321) );
  XOR U20369 ( .A(n18322), .B(n18323), .Z(n18310) );
  AND U20370 ( .A(n18324), .B(n18325), .Z(n18323) );
  XNOR U20371 ( .A(n18322), .B(n9163), .Z(n18325) );
  XNOR U20372 ( .A(n18318), .B(n18320), .Z(n9163) );
  NAND U20373 ( .A(n18326), .B(nreg[523]), .Z(n18320) );
  NAND U20374 ( .A(n12326), .B(nreg[523]), .Z(n18326) );
  XNOR U20375 ( .A(n18316), .B(n18327), .Z(n18318) );
  XOR U20376 ( .A(n18328), .B(n18329), .Z(n18316) );
  AND U20377 ( .A(n18330), .B(n18331), .Z(n18329) );
  XNOR U20378 ( .A(n18332), .B(n18328), .Z(n18331) );
  XOR U20379 ( .A(n18333), .B(nreg[523]), .Z(n18324) );
  IV U20380 ( .A(n18322), .Z(n18333) );
  XOR U20381 ( .A(n18334), .B(n18335), .Z(n18322) );
  AND U20382 ( .A(n18336), .B(n18337), .Z(n18335) );
  XNOR U20383 ( .A(n18334), .B(n9169), .Z(n18337) );
  XNOR U20384 ( .A(n18330), .B(n18332), .Z(n9169) );
  NAND U20385 ( .A(n18338), .B(nreg[522]), .Z(n18332) );
  NAND U20386 ( .A(n12326), .B(nreg[522]), .Z(n18338) );
  XNOR U20387 ( .A(n18328), .B(n18339), .Z(n18330) );
  XOR U20388 ( .A(n18340), .B(n18341), .Z(n18328) );
  AND U20389 ( .A(n18342), .B(n18343), .Z(n18341) );
  XNOR U20390 ( .A(n18344), .B(n18340), .Z(n18343) );
  XOR U20391 ( .A(n18345), .B(nreg[522]), .Z(n18336) );
  IV U20392 ( .A(n18334), .Z(n18345) );
  XOR U20393 ( .A(n18346), .B(n18347), .Z(n18334) );
  AND U20394 ( .A(n18348), .B(n18349), .Z(n18347) );
  XNOR U20395 ( .A(n18346), .B(n9175), .Z(n18349) );
  XNOR U20396 ( .A(n18342), .B(n18344), .Z(n9175) );
  NAND U20397 ( .A(n18350), .B(nreg[521]), .Z(n18344) );
  NAND U20398 ( .A(n12326), .B(nreg[521]), .Z(n18350) );
  XNOR U20399 ( .A(n18340), .B(n18351), .Z(n18342) );
  XOR U20400 ( .A(n18352), .B(n18353), .Z(n18340) );
  AND U20401 ( .A(n18354), .B(n18355), .Z(n18353) );
  XNOR U20402 ( .A(n18356), .B(n18352), .Z(n18355) );
  XOR U20403 ( .A(n18357), .B(nreg[521]), .Z(n18348) );
  IV U20404 ( .A(n18346), .Z(n18357) );
  XOR U20405 ( .A(n18358), .B(n18359), .Z(n18346) );
  AND U20406 ( .A(n18360), .B(n18361), .Z(n18359) );
  XNOR U20407 ( .A(n18358), .B(n9181), .Z(n18361) );
  XNOR U20408 ( .A(n18354), .B(n18356), .Z(n9181) );
  NAND U20409 ( .A(n18362), .B(nreg[520]), .Z(n18356) );
  NAND U20410 ( .A(n12326), .B(nreg[520]), .Z(n18362) );
  XNOR U20411 ( .A(n18352), .B(n18363), .Z(n18354) );
  XOR U20412 ( .A(n18364), .B(n18365), .Z(n18352) );
  AND U20413 ( .A(n18366), .B(n18367), .Z(n18365) );
  XNOR U20414 ( .A(n18368), .B(n18364), .Z(n18367) );
  XOR U20415 ( .A(n18369), .B(nreg[520]), .Z(n18360) );
  IV U20416 ( .A(n18358), .Z(n18369) );
  XOR U20417 ( .A(n18370), .B(n18371), .Z(n18358) );
  AND U20418 ( .A(n18372), .B(n18373), .Z(n18371) );
  XNOR U20419 ( .A(n18370), .B(n9187), .Z(n18373) );
  XNOR U20420 ( .A(n18366), .B(n18368), .Z(n9187) );
  NAND U20421 ( .A(n18374), .B(nreg[519]), .Z(n18368) );
  NAND U20422 ( .A(n12326), .B(nreg[519]), .Z(n18374) );
  XNOR U20423 ( .A(n18364), .B(n18375), .Z(n18366) );
  XOR U20424 ( .A(n18376), .B(n18377), .Z(n18364) );
  AND U20425 ( .A(n18378), .B(n18379), .Z(n18377) );
  XNOR U20426 ( .A(n18380), .B(n18376), .Z(n18379) );
  XOR U20427 ( .A(n18381), .B(nreg[519]), .Z(n18372) );
  IV U20428 ( .A(n18370), .Z(n18381) );
  XOR U20429 ( .A(n18382), .B(n18383), .Z(n18370) );
  AND U20430 ( .A(n18384), .B(n18385), .Z(n18383) );
  XNOR U20431 ( .A(n18382), .B(n9193), .Z(n18385) );
  XNOR U20432 ( .A(n18378), .B(n18380), .Z(n9193) );
  NAND U20433 ( .A(n18386), .B(nreg[518]), .Z(n18380) );
  NAND U20434 ( .A(n12326), .B(nreg[518]), .Z(n18386) );
  XNOR U20435 ( .A(n18376), .B(n18387), .Z(n18378) );
  XOR U20436 ( .A(n18388), .B(n18389), .Z(n18376) );
  AND U20437 ( .A(n18390), .B(n18391), .Z(n18389) );
  XNOR U20438 ( .A(n18392), .B(n18388), .Z(n18391) );
  XOR U20439 ( .A(n18393), .B(nreg[518]), .Z(n18384) );
  IV U20440 ( .A(n18382), .Z(n18393) );
  XOR U20441 ( .A(n18394), .B(n18395), .Z(n18382) );
  AND U20442 ( .A(n18396), .B(n18397), .Z(n18395) );
  XNOR U20443 ( .A(n18394), .B(n9199), .Z(n18397) );
  XNOR U20444 ( .A(n18390), .B(n18392), .Z(n9199) );
  NAND U20445 ( .A(n18398), .B(nreg[517]), .Z(n18392) );
  NAND U20446 ( .A(n12326), .B(nreg[517]), .Z(n18398) );
  XNOR U20447 ( .A(n18388), .B(n18399), .Z(n18390) );
  XOR U20448 ( .A(n18400), .B(n18401), .Z(n18388) );
  AND U20449 ( .A(n18402), .B(n18403), .Z(n18401) );
  XNOR U20450 ( .A(n18404), .B(n18400), .Z(n18403) );
  XOR U20451 ( .A(n18405), .B(nreg[517]), .Z(n18396) );
  IV U20452 ( .A(n18394), .Z(n18405) );
  XOR U20453 ( .A(n18406), .B(n18407), .Z(n18394) );
  AND U20454 ( .A(n18408), .B(n18409), .Z(n18407) );
  XNOR U20455 ( .A(n18406), .B(n9205), .Z(n18409) );
  XNOR U20456 ( .A(n18402), .B(n18404), .Z(n9205) );
  NAND U20457 ( .A(n18410), .B(nreg[516]), .Z(n18404) );
  NAND U20458 ( .A(n12326), .B(nreg[516]), .Z(n18410) );
  XNOR U20459 ( .A(n18400), .B(n18411), .Z(n18402) );
  XOR U20460 ( .A(n18412), .B(n18413), .Z(n18400) );
  AND U20461 ( .A(n18414), .B(n18415), .Z(n18413) );
  XNOR U20462 ( .A(n18416), .B(n18412), .Z(n18415) );
  XOR U20463 ( .A(n18417), .B(nreg[516]), .Z(n18408) );
  IV U20464 ( .A(n18406), .Z(n18417) );
  XOR U20465 ( .A(n18418), .B(n18419), .Z(n18406) );
  AND U20466 ( .A(n18420), .B(n18421), .Z(n18419) );
  XNOR U20467 ( .A(n18418), .B(n9211), .Z(n18421) );
  XNOR U20468 ( .A(n18414), .B(n18416), .Z(n9211) );
  NAND U20469 ( .A(n18422), .B(nreg[515]), .Z(n18416) );
  NAND U20470 ( .A(n12326), .B(nreg[515]), .Z(n18422) );
  XNOR U20471 ( .A(n18412), .B(n18423), .Z(n18414) );
  XOR U20472 ( .A(n18424), .B(n18425), .Z(n18412) );
  AND U20473 ( .A(n18426), .B(n18427), .Z(n18425) );
  XNOR U20474 ( .A(n18428), .B(n18424), .Z(n18427) );
  XOR U20475 ( .A(n18429), .B(nreg[515]), .Z(n18420) );
  IV U20476 ( .A(n18418), .Z(n18429) );
  XOR U20477 ( .A(n18430), .B(n18431), .Z(n18418) );
  AND U20478 ( .A(n18432), .B(n18433), .Z(n18431) );
  XNOR U20479 ( .A(n18430), .B(n9217), .Z(n18433) );
  XNOR U20480 ( .A(n18426), .B(n18428), .Z(n9217) );
  NAND U20481 ( .A(n18434), .B(nreg[514]), .Z(n18428) );
  NAND U20482 ( .A(n12326), .B(nreg[514]), .Z(n18434) );
  XNOR U20483 ( .A(n18424), .B(n18435), .Z(n18426) );
  XOR U20484 ( .A(n18436), .B(n18437), .Z(n18424) );
  AND U20485 ( .A(n18438), .B(n18439), .Z(n18437) );
  XNOR U20486 ( .A(n18440), .B(n18436), .Z(n18439) );
  XOR U20487 ( .A(n18441), .B(nreg[514]), .Z(n18432) );
  IV U20488 ( .A(n18430), .Z(n18441) );
  XOR U20489 ( .A(n18442), .B(n18443), .Z(n18430) );
  AND U20490 ( .A(n18444), .B(n18445), .Z(n18443) );
  XNOR U20491 ( .A(n18442), .B(n9223), .Z(n18445) );
  XNOR U20492 ( .A(n18438), .B(n18440), .Z(n9223) );
  NAND U20493 ( .A(n18446), .B(nreg[513]), .Z(n18440) );
  NAND U20494 ( .A(n12326), .B(nreg[513]), .Z(n18446) );
  XNOR U20495 ( .A(n18436), .B(n18447), .Z(n18438) );
  XOR U20496 ( .A(n18448), .B(n18449), .Z(n18436) );
  AND U20497 ( .A(n18450), .B(n18451), .Z(n18449) );
  XNOR U20498 ( .A(n18452), .B(n18448), .Z(n18451) );
  XOR U20499 ( .A(n18453), .B(nreg[513]), .Z(n18444) );
  IV U20500 ( .A(n18442), .Z(n18453) );
  XOR U20501 ( .A(n18454), .B(n18455), .Z(n18442) );
  AND U20502 ( .A(n18456), .B(n18457), .Z(n18455) );
  XNOR U20503 ( .A(n18454), .B(n9229), .Z(n18457) );
  XNOR U20504 ( .A(n18450), .B(n18452), .Z(n9229) );
  NAND U20505 ( .A(n18458), .B(nreg[512]), .Z(n18452) );
  NAND U20506 ( .A(n12326), .B(nreg[512]), .Z(n18458) );
  XNOR U20507 ( .A(n18448), .B(n18459), .Z(n18450) );
  XOR U20508 ( .A(n18460), .B(n18461), .Z(n18448) );
  AND U20509 ( .A(n18462), .B(n18463), .Z(n18461) );
  XNOR U20510 ( .A(n18464), .B(n18460), .Z(n18463) );
  XOR U20511 ( .A(n18465), .B(nreg[512]), .Z(n18456) );
  IV U20512 ( .A(n18454), .Z(n18465) );
  XOR U20513 ( .A(n18466), .B(n18467), .Z(n18454) );
  AND U20514 ( .A(n18468), .B(n18469), .Z(n18467) );
  XNOR U20515 ( .A(n18466), .B(n9235), .Z(n18469) );
  XNOR U20516 ( .A(n18462), .B(n18464), .Z(n9235) );
  NAND U20517 ( .A(n18470), .B(nreg[511]), .Z(n18464) );
  NAND U20518 ( .A(n12326), .B(nreg[511]), .Z(n18470) );
  XNOR U20519 ( .A(n18460), .B(n18471), .Z(n18462) );
  XOR U20520 ( .A(n18472), .B(n18473), .Z(n18460) );
  AND U20521 ( .A(n18474), .B(n18475), .Z(n18473) );
  XNOR U20522 ( .A(n18476), .B(n18472), .Z(n18475) );
  XOR U20523 ( .A(n18477), .B(nreg[511]), .Z(n18468) );
  IV U20524 ( .A(n18466), .Z(n18477) );
  XOR U20525 ( .A(n18478), .B(n18479), .Z(n18466) );
  AND U20526 ( .A(n18480), .B(n18481), .Z(n18479) );
  XNOR U20527 ( .A(n18478), .B(n9241), .Z(n18481) );
  XNOR U20528 ( .A(n18474), .B(n18476), .Z(n9241) );
  NAND U20529 ( .A(n18482), .B(nreg[510]), .Z(n18476) );
  NAND U20530 ( .A(n12326), .B(nreg[510]), .Z(n18482) );
  XNOR U20531 ( .A(n18472), .B(n18483), .Z(n18474) );
  XOR U20532 ( .A(n18484), .B(n18485), .Z(n18472) );
  AND U20533 ( .A(n18486), .B(n18487), .Z(n18485) );
  XNOR U20534 ( .A(n18488), .B(n18484), .Z(n18487) );
  XOR U20535 ( .A(n18489), .B(nreg[510]), .Z(n18480) );
  IV U20536 ( .A(n18478), .Z(n18489) );
  XOR U20537 ( .A(n18490), .B(n18491), .Z(n18478) );
  AND U20538 ( .A(n18492), .B(n18493), .Z(n18491) );
  XNOR U20539 ( .A(n18490), .B(n9247), .Z(n18493) );
  XNOR U20540 ( .A(n18486), .B(n18488), .Z(n9247) );
  NAND U20541 ( .A(n18494), .B(nreg[509]), .Z(n18488) );
  NAND U20542 ( .A(n12326), .B(nreg[509]), .Z(n18494) );
  XNOR U20543 ( .A(n18484), .B(n18495), .Z(n18486) );
  XOR U20544 ( .A(n18496), .B(n18497), .Z(n18484) );
  AND U20545 ( .A(n18498), .B(n18499), .Z(n18497) );
  XNOR U20546 ( .A(n18500), .B(n18496), .Z(n18499) );
  XOR U20547 ( .A(n18501), .B(nreg[509]), .Z(n18492) );
  IV U20548 ( .A(n18490), .Z(n18501) );
  XOR U20549 ( .A(n18502), .B(n18503), .Z(n18490) );
  AND U20550 ( .A(n18504), .B(n18505), .Z(n18503) );
  XNOR U20551 ( .A(n18502), .B(n9253), .Z(n18505) );
  XNOR U20552 ( .A(n18498), .B(n18500), .Z(n9253) );
  NAND U20553 ( .A(n18506), .B(nreg[508]), .Z(n18500) );
  NAND U20554 ( .A(n12326), .B(nreg[508]), .Z(n18506) );
  XNOR U20555 ( .A(n18496), .B(n18507), .Z(n18498) );
  XOR U20556 ( .A(n18508), .B(n18509), .Z(n18496) );
  AND U20557 ( .A(n18510), .B(n18511), .Z(n18509) );
  XNOR U20558 ( .A(n18512), .B(n18508), .Z(n18511) );
  XOR U20559 ( .A(n18513), .B(nreg[508]), .Z(n18504) );
  IV U20560 ( .A(n18502), .Z(n18513) );
  XOR U20561 ( .A(n18514), .B(n18515), .Z(n18502) );
  AND U20562 ( .A(n18516), .B(n18517), .Z(n18515) );
  XNOR U20563 ( .A(n18514), .B(n9259), .Z(n18517) );
  XNOR U20564 ( .A(n18510), .B(n18512), .Z(n9259) );
  NAND U20565 ( .A(n18518), .B(nreg[507]), .Z(n18512) );
  NAND U20566 ( .A(n12326), .B(nreg[507]), .Z(n18518) );
  XNOR U20567 ( .A(n18508), .B(n18519), .Z(n18510) );
  XOR U20568 ( .A(n18520), .B(n18521), .Z(n18508) );
  AND U20569 ( .A(n18522), .B(n18523), .Z(n18521) );
  XNOR U20570 ( .A(n18524), .B(n18520), .Z(n18523) );
  XOR U20571 ( .A(n18525), .B(nreg[507]), .Z(n18516) );
  IV U20572 ( .A(n18514), .Z(n18525) );
  XOR U20573 ( .A(n18526), .B(n18527), .Z(n18514) );
  AND U20574 ( .A(n18528), .B(n18529), .Z(n18527) );
  XNOR U20575 ( .A(n18526), .B(n9265), .Z(n18529) );
  XNOR U20576 ( .A(n18522), .B(n18524), .Z(n9265) );
  NAND U20577 ( .A(n18530), .B(nreg[506]), .Z(n18524) );
  NAND U20578 ( .A(n12326), .B(nreg[506]), .Z(n18530) );
  XNOR U20579 ( .A(n18520), .B(n18531), .Z(n18522) );
  XOR U20580 ( .A(n18532), .B(n18533), .Z(n18520) );
  AND U20581 ( .A(n18534), .B(n18535), .Z(n18533) );
  XNOR U20582 ( .A(n18536), .B(n18532), .Z(n18535) );
  XOR U20583 ( .A(n18537), .B(nreg[506]), .Z(n18528) );
  IV U20584 ( .A(n18526), .Z(n18537) );
  XOR U20585 ( .A(n18538), .B(n18539), .Z(n18526) );
  AND U20586 ( .A(n18540), .B(n18541), .Z(n18539) );
  XNOR U20587 ( .A(n18538), .B(n9271), .Z(n18541) );
  XNOR U20588 ( .A(n18534), .B(n18536), .Z(n9271) );
  NAND U20589 ( .A(n18542), .B(nreg[505]), .Z(n18536) );
  NAND U20590 ( .A(n12326), .B(nreg[505]), .Z(n18542) );
  XNOR U20591 ( .A(n18532), .B(n18543), .Z(n18534) );
  XOR U20592 ( .A(n18544), .B(n18545), .Z(n18532) );
  AND U20593 ( .A(n18546), .B(n18547), .Z(n18545) );
  XNOR U20594 ( .A(n18548), .B(n18544), .Z(n18547) );
  XOR U20595 ( .A(n18549), .B(nreg[505]), .Z(n18540) );
  IV U20596 ( .A(n18538), .Z(n18549) );
  XOR U20597 ( .A(n18550), .B(n18551), .Z(n18538) );
  AND U20598 ( .A(n18552), .B(n18553), .Z(n18551) );
  XNOR U20599 ( .A(n18550), .B(n9277), .Z(n18553) );
  XNOR U20600 ( .A(n18546), .B(n18548), .Z(n9277) );
  NAND U20601 ( .A(n18554), .B(nreg[504]), .Z(n18548) );
  NAND U20602 ( .A(n12326), .B(nreg[504]), .Z(n18554) );
  XNOR U20603 ( .A(n18544), .B(n18555), .Z(n18546) );
  XOR U20604 ( .A(n18556), .B(n18557), .Z(n18544) );
  AND U20605 ( .A(n18558), .B(n18559), .Z(n18557) );
  XNOR U20606 ( .A(n18560), .B(n18556), .Z(n18559) );
  XOR U20607 ( .A(n18561), .B(nreg[504]), .Z(n18552) );
  IV U20608 ( .A(n18550), .Z(n18561) );
  XOR U20609 ( .A(n18562), .B(n18563), .Z(n18550) );
  AND U20610 ( .A(n18564), .B(n18565), .Z(n18563) );
  XNOR U20611 ( .A(n18562), .B(n9283), .Z(n18565) );
  XNOR U20612 ( .A(n18558), .B(n18560), .Z(n9283) );
  NAND U20613 ( .A(n18566), .B(nreg[503]), .Z(n18560) );
  NAND U20614 ( .A(n12326), .B(nreg[503]), .Z(n18566) );
  XNOR U20615 ( .A(n18556), .B(n18567), .Z(n18558) );
  XOR U20616 ( .A(n18568), .B(n18569), .Z(n18556) );
  AND U20617 ( .A(n18570), .B(n18571), .Z(n18569) );
  XNOR U20618 ( .A(n18572), .B(n18568), .Z(n18571) );
  XOR U20619 ( .A(n18573), .B(nreg[503]), .Z(n18564) );
  IV U20620 ( .A(n18562), .Z(n18573) );
  XOR U20621 ( .A(n18574), .B(n18575), .Z(n18562) );
  AND U20622 ( .A(n18576), .B(n18577), .Z(n18575) );
  XNOR U20623 ( .A(n18574), .B(n9289), .Z(n18577) );
  XNOR U20624 ( .A(n18570), .B(n18572), .Z(n9289) );
  NAND U20625 ( .A(n18578), .B(nreg[502]), .Z(n18572) );
  NAND U20626 ( .A(n12326), .B(nreg[502]), .Z(n18578) );
  XNOR U20627 ( .A(n18568), .B(n18579), .Z(n18570) );
  XOR U20628 ( .A(n18580), .B(n18581), .Z(n18568) );
  AND U20629 ( .A(n18582), .B(n18583), .Z(n18581) );
  XNOR U20630 ( .A(n18584), .B(n18580), .Z(n18583) );
  XOR U20631 ( .A(n18585), .B(nreg[502]), .Z(n18576) );
  IV U20632 ( .A(n18574), .Z(n18585) );
  XOR U20633 ( .A(n18586), .B(n18587), .Z(n18574) );
  AND U20634 ( .A(n18588), .B(n18589), .Z(n18587) );
  XNOR U20635 ( .A(n18586), .B(n9295), .Z(n18589) );
  XNOR U20636 ( .A(n18582), .B(n18584), .Z(n9295) );
  NAND U20637 ( .A(n18590), .B(nreg[501]), .Z(n18584) );
  NAND U20638 ( .A(n12326), .B(nreg[501]), .Z(n18590) );
  XNOR U20639 ( .A(n18580), .B(n18591), .Z(n18582) );
  XOR U20640 ( .A(n18592), .B(n18593), .Z(n18580) );
  AND U20641 ( .A(n18594), .B(n18595), .Z(n18593) );
  XNOR U20642 ( .A(n18596), .B(n18592), .Z(n18595) );
  XOR U20643 ( .A(n18597), .B(nreg[501]), .Z(n18588) );
  IV U20644 ( .A(n18586), .Z(n18597) );
  XOR U20645 ( .A(n18598), .B(n18599), .Z(n18586) );
  AND U20646 ( .A(n18600), .B(n18601), .Z(n18599) );
  XNOR U20647 ( .A(n18598), .B(n9301), .Z(n18601) );
  XNOR U20648 ( .A(n18594), .B(n18596), .Z(n9301) );
  NAND U20649 ( .A(n18602), .B(nreg[500]), .Z(n18596) );
  NAND U20650 ( .A(n12326), .B(nreg[500]), .Z(n18602) );
  XNOR U20651 ( .A(n18592), .B(n18603), .Z(n18594) );
  XOR U20652 ( .A(n18604), .B(n18605), .Z(n18592) );
  AND U20653 ( .A(n18606), .B(n18607), .Z(n18605) );
  XNOR U20654 ( .A(n18608), .B(n18604), .Z(n18607) );
  XOR U20655 ( .A(n18609), .B(nreg[500]), .Z(n18600) );
  IV U20656 ( .A(n18598), .Z(n18609) );
  XOR U20657 ( .A(n18610), .B(n18611), .Z(n18598) );
  AND U20658 ( .A(n18612), .B(n18613), .Z(n18611) );
  XNOR U20659 ( .A(n18610), .B(n9307), .Z(n18613) );
  XNOR U20660 ( .A(n18606), .B(n18608), .Z(n9307) );
  NAND U20661 ( .A(n18614), .B(nreg[499]), .Z(n18608) );
  NAND U20662 ( .A(n12326), .B(nreg[499]), .Z(n18614) );
  XNOR U20663 ( .A(n18604), .B(n18615), .Z(n18606) );
  XOR U20664 ( .A(n18616), .B(n18617), .Z(n18604) );
  AND U20665 ( .A(n18618), .B(n18619), .Z(n18617) );
  XNOR U20666 ( .A(n18620), .B(n18616), .Z(n18619) );
  XOR U20667 ( .A(n18621), .B(nreg[499]), .Z(n18612) );
  IV U20668 ( .A(n18610), .Z(n18621) );
  XOR U20669 ( .A(n18622), .B(n18623), .Z(n18610) );
  AND U20670 ( .A(n18624), .B(n18625), .Z(n18623) );
  XNOR U20671 ( .A(n18622), .B(n9313), .Z(n18625) );
  XNOR U20672 ( .A(n18618), .B(n18620), .Z(n9313) );
  NAND U20673 ( .A(n18626), .B(nreg[498]), .Z(n18620) );
  NAND U20674 ( .A(n12326), .B(nreg[498]), .Z(n18626) );
  XNOR U20675 ( .A(n18616), .B(n18627), .Z(n18618) );
  XOR U20676 ( .A(n18628), .B(n18629), .Z(n18616) );
  AND U20677 ( .A(n18630), .B(n18631), .Z(n18629) );
  XNOR U20678 ( .A(n18632), .B(n18628), .Z(n18631) );
  XOR U20679 ( .A(n18633), .B(nreg[498]), .Z(n18624) );
  IV U20680 ( .A(n18622), .Z(n18633) );
  XOR U20681 ( .A(n18634), .B(n18635), .Z(n18622) );
  AND U20682 ( .A(n18636), .B(n18637), .Z(n18635) );
  XNOR U20683 ( .A(n18634), .B(n9319), .Z(n18637) );
  XNOR U20684 ( .A(n18630), .B(n18632), .Z(n9319) );
  NAND U20685 ( .A(n18638), .B(nreg[497]), .Z(n18632) );
  NAND U20686 ( .A(n12326), .B(nreg[497]), .Z(n18638) );
  XNOR U20687 ( .A(n18628), .B(n18639), .Z(n18630) );
  XOR U20688 ( .A(n18640), .B(n18641), .Z(n18628) );
  AND U20689 ( .A(n18642), .B(n18643), .Z(n18641) );
  XNOR U20690 ( .A(n18644), .B(n18640), .Z(n18643) );
  XOR U20691 ( .A(n18645), .B(nreg[497]), .Z(n18636) );
  IV U20692 ( .A(n18634), .Z(n18645) );
  XOR U20693 ( .A(n18646), .B(n18647), .Z(n18634) );
  AND U20694 ( .A(n18648), .B(n18649), .Z(n18647) );
  XNOR U20695 ( .A(n18646), .B(n9325), .Z(n18649) );
  XNOR U20696 ( .A(n18642), .B(n18644), .Z(n9325) );
  NAND U20697 ( .A(n18650), .B(nreg[496]), .Z(n18644) );
  NAND U20698 ( .A(n12326), .B(nreg[496]), .Z(n18650) );
  XNOR U20699 ( .A(n18640), .B(n18651), .Z(n18642) );
  XOR U20700 ( .A(n18652), .B(n18653), .Z(n18640) );
  AND U20701 ( .A(n18654), .B(n18655), .Z(n18653) );
  XNOR U20702 ( .A(n18656), .B(n18652), .Z(n18655) );
  XOR U20703 ( .A(n18657), .B(nreg[496]), .Z(n18648) );
  IV U20704 ( .A(n18646), .Z(n18657) );
  XOR U20705 ( .A(n18658), .B(n18659), .Z(n18646) );
  AND U20706 ( .A(n18660), .B(n18661), .Z(n18659) );
  XNOR U20707 ( .A(n18658), .B(n9331), .Z(n18661) );
  XNOR U20708 ( .A(n18654), .B(n18656), .Z(n9331) );
  NAND U20709 ( .A(n18662), .B(nreg[495]), .Z(n18656) );
  NAND U20710 ( .A(n12326), .B(nreg[495]), .Z(n18662) );
  XNOR U20711 ( .A(n18652), .B(n18663), .Z(n18654) );
  XOR U20712 ( .A(n18664), .B(n18665), .Z(n18652) );
  AND U20713 ( .A(n18666), .B(n18667), .Z(n18665) );
  XNOR U20714 ( .A(n18668), .B(n18664), .Z(n18667) );
  XOR U20715 ( .A(n18669), .B(nreg[495]), .Z(n18660) );
  IV U20716 ( .A(n18658), .Z(n18669) );
  XOR U20717 ( .A(n18670), .B(n18671), .Z(n18658) );
  AND U20718 ( .A(n18672), .B(n18673), .Z(n18671) );
  XNOR U20719 ( .A(n18670), .B(n9337), .Z(n18673) );
  XNOR U20720 ( .A(n18666), .B(n18668), .Z(n9337) );
  NAND U20721 ( .A(n18674), .B(nreg[494]), .Z(n18668) );
  NAND U20722 ( .A(n12326), .B(nreg[494]), .Z(n18674) );
  XNOR U20723 ( .A(n18664), .B(n18675), .Z(n18666) );
  XOR U20724 ( .A(n18676), .B(n18677), .Z(n18664) );
  AND U20725 ( .A(n18678), .B(n18679), .Z(n18677) );
  XNOR U20726 ( .A(n18680), .B(n18676), .Z(n18679) );
  XOR U20727 ( .A(n18681), .B(nreg[494]), .Z(n18672) );
  IV U20728 ( .A(n18670), .Z(n18681) );
  XOR U20729 ( .A(n18682), .B(n18683), .Z(n18670) );
  AND U20730 ( .A(n18684), .B(n18685), .Z(n18683) );
  XNOR U20731 ( .A(n18682), .B(n9343), .Z(n18685) );
  XNOR U20732 ( .A(n18678), .B(n18680), .Z(n9343) );
  NAND U20733 ( .A(n18686), .B(nreg[493]), .Z(n18680) );
  NAND U20734 ( .A(n12326), .B(nreg[493]), .Z(n18686) );
  XNOR U20735 ( .A(n18676), .B(n18687), .Z(n18678) );
  XOR U20736 ( .A(n18688), .B(n18689), .Z(n18676) );
  AND U20737 ( .A(n18690), .B(n18691), .Z(n18689) );
  XNOR U20738 ( .A(n18692), .B(n18688), .Z(n18691) );
  XOR U20739 ( .A(n18693), .B(nreg[493]), .Z(n18684) );
  IV U20740 ( .A(n18682), .Z(n18693) );
  XOR U20741 ( .A(n18694), .B(n18695), .Z(n18682) );
  AND U20742 ( .A(n18696), .B(n18697), .Z(n18695) );
  XNOR U20743 ( .A(n18694), .B(n9349), .Z(n18697) );
  XNOR U20744 ( .A(n18690), .B(n18692), .Z(n9349) );
  NAND U20745 ( .A(n18698), .B(nreg[492]), .Z(n18692) );
  NAND U20746 ( .A(n12326), .B(nreg[492]), .Z(n18698) );
  XNOR U20747 ( .A(n18688), .B(n18699), .Z(n18690) );
  XOR U20748 ( .A(n18700), .B(n18701), .Z(n18688) );
  AND U20749 ( .A(n18702), .B(n18703), .Z(n18701) );
  XNOR U20750 ( .A(n18704), .B(n18700), .Z(n18703) );
  XOR U20751 ( .A(n18705), .B(nreg[492]), .Z(n18696) );
  IV U20752 ( .A(n18694), .Z(n18705) );
  XOR U20753 ( .A(n18706), .B(n18707), .Z(n18694) );
  AND U20754 ( .A(n18708), .B(n18709), .Z(n18707) );
  XNOR U20755 ( .A(n18706), .B(n9355), .Z(n18709) );
  XNOR U20756 ( .A(n18702), .B(n18704), .Z(n9355) );
  NAND U20757 ( .A(n18710), .B(nreg[491]), .Z(n18704) );
  NAND U20758 ( .A(n12326), .B(nreg[491]), .Z(n18710) );
  XNOR U20759 ( .A(n18700), .B(n18711), .Z(n18702) );
  XOR U20760 ( .A(n18712), .B(n18713), .Z(n18700) );
  AND U20761 ( .A(n18714), .B(n18715), .Z(n18713) );
  XNOR U20762 ( .A(n18716), .B(n18712), .Z(n18715) );
  XOR U20763 ( .A(n18717), .B(nreg[491]), .Z(n18708) );
  IV U20764 ( .A(n18706), .Z(n18717) );
  XOR U20765 ( .A(n18718), .B(n18719), .Z(n18706) );
  AND U20766 ( .A(n18720), .B(n18721), .Z(n18719) );
  XNOR U20767 ( .A(n18718), .B(n9361), .Z(n18721) );
  XNOR U20768 ( .A(n18714), .B(n18716), .Z(n9361) );
  NAND U20769 ( .A(n18722), .B(nreg[490]), .Z(n18716) );
  NAND U20770 ( .A(n12326), .B(nreg[490]), .Z(n18722) );
  XNOR U20771 ( .A(n18712), .B(n18723), .Z(n18714) );
  XOR U20772 ( .A(n18724), .B(n18725), .Z(n18712) );
  AND U20773 ( .A(n18726), .B(n18727), .Z(n18725) );
  XNOR U20774 ( .A(n18728), .B(n18724), .Z(n18727) );
  XOR U20775 ( .A(n18729), .B(nreg[490]), .Z(n18720) );
  IV U20776 ( .A(n18718), .Z(n18729) );
  XOR U20777 ( .A(n18730), .B(n18731), .Z(n18718) );
  AND U20778 ( .A(n18732), .B(n18733), .Z(n18731) );
  XNOR U20779 ( .A(n18730), .B(n9367), .Z(n18733) );
  XNOR U20780 ( .A(n18726), .B(n18728), .Z(n9367) );
  NAND U20781 ( .A(n18734), .B(nreg[489]), .Z(n18728) );
  NAND U20782 ( .A(n12326), .B(nreg[489]), .Z(n18734) );
  XNOR U20783 ( .A(n18724), .B(n18735), .Z(n18726) );
  XOR U20784 ( .A(n18736), .B(n18737), .Z(n18724) );
  AND U20785 ( .A(n18738), .B(n18739), .Z(n18737) );
  XNOR U20786 ( .A(n18740), .B(n18736), .Z(n18739) );
  XOR U20787 ( .A(n18741), .B(nreg[489]), .Z(n18732) );
  IV U20788 ( .A(n18730), .Z(n18741) );
  XOR U20789 ( .A(n18742), .B(n18743), .Z(n18730) );
  AND U20790 ( .A(n18744), .B(n18745), .Z(n18743) );
  XNOR U20791 ( .A(n18742), .B(n9373), .Z(n18745) );
  XNOR U20792 ( .A(n18738), .B(n18740), .Z(n9373) );
  NAND U20793 ( .A(n18746), .B(nreg[488]), .Z(n18740) );
  NAND U20794 ( .A(n12326), .B(nreg[488]), .Z(n18746) );
  XNOR U20795 ( .A(n18736), .B(n18747), .Z(n18738) );
  XOR U20796 ( .A(n18748), .B(n18749), .Z(n18736) );
  AND U20797 ( .A(n18750), .B(n18751), .Z(n18749) );
  XNOR U20798 ( .A(n18752), .B(n18748), .Z(n18751) );
  XOR U20799 ( .A(n18753), .B(nreg[488]), .Z(n18744) );
  IV U20800 ( .A(n18742), .Z(n18753) );
  XOR U20801 ( .A(n18754), .B(n18755), .Z(n18742) );
  AND U20802 ( .A(n18756), .B(n18757), .Z(n18755) );
  XNOR U20803 ( .A(n18754), .B(n9379), .Z(n18757) );
  XNOR U20804 ( .A(n18750), .B(n18752), .Z(n9379) );
  NAND U20805 ( .A(n18758), .B(nreg[487]), .Z(n18752) );
  NAND U20806 ( .A(n12326), .B(nreg[487]), .Z(n18758) );
  XNOR U20807 ( .A(n18748), .B(n18759), .Z(n18750) );
  XOR U20808 ( .A(n18760), .B(n18761), .Z(n18748) );
  AND U20809 ( .A(n18762), .B(n18763), .Z(n18761) );
  XNOR U20810 ( .A(n18764), .B(n18760), .Z(n18763) );
  XOR U20811 ( .A(n18765), .B(nreg[487]), .Z(n18756) );
  IV U20812 ( .A(n18754), .Z(n18765) );
  XOR U20813 ( .A(n18766), .B(n18767), .Z(n18754) );
  AND U20814 ( .A(n18768), .B(n18769), .Z(n18767) );
  XNOR U20815 ( .A(n18766), .B(n9385), .Z(n18769) );
  XNOR U20816 ( .A(n18762), .B(n18764), .Z(n9385) );
  NAND U20817 ( .A(n18770), .B(nreg[486]), .Z(n18764) );
  NAND U20818 ( .A(n12326), .B(nreg[486]), .Z(n18770) );
  XNOR U20819 ( .A(n18760), .B(n18771), .Z(n18762) );
  XOR U20820 ( .A(n18772), .B(n18773), .Z(n18760) );
  AND U20821 ( .A(n18774), .B(n18775), .Z(n18773) );
  XNOR U20822 ( .A(n18776), .B(n18772), .Z(n18775) );
  XOR U20823 ( .A(n18777), .B(nreg[486]), .Z(n18768) );
  IV U20824 ( .A(n18766), .Z(n18777) );
  XOR U20825 ( .A(n18778), .B(n18779), .Z(n18766) );
  AND U20826 ( .A(n18780), .B(n18781), .Z(n18779) );
  XNOR U20827 ( .A(n18778), .B(n9391), .Z(n18781) );
  XNOR U20828 ( .A(n18774), .B(n18776), .Z(n9391) );
  NAND U20829 ( .A(n18782), .B(nreg[485]), .Z(n18776) );
  NAND U20830 ( .A(n12326), .B(nreg[485]), .Z(n18782) );
  XNOR U20831 ( .A(n18772), .B(n18783), .Z(n18774) );
  XOR U20832 ( .A(n18784), .B(n18785), .Z(n18772) );
  AND U20833 ( .A(n18786), .B(n18787), .Z(n18785) );
  XNOR U20834 ( .A(n18788), .B(n18784), .Z(n18787) );
  XOR U20835 ( .A(n18789), .B(nreg[485]), .Z(n18780) );
  IV U20836 ( .A(n18778), .Z(n18789) );
  XOR U20837 ( .A(n18790), .B(n18791), .Z(n18778) );
  AND U20838 ( .A(n18792), .B(n18793), .Z(n18791) );
  XNOR U20839 ( .A(n18790), .B(n9397), .Z(n18793) );
  XNOR U20840 ( .A(n18786), .B(n18788), .Z(n9397) );
  NAND U20841 ( .A(n18794), .B(nreg[484]), .Z(n18788) );
  NAND U20842 ( .A(n12326), .B(nreg[484]), .Z(n18794) );
  XNOR U20843 ( .A(n18784), .B(n18795), .Z(n18786) );
  XOR U20844 ( .A(n18796), .B(n18797), .Z(n18784) );
  AND U20845 ( .A(n18798), .B(n18799), .Z(n18797) );
  XNOR U20846 ( .A(n18800), .B(n18796), .Z(n18799) );
  XOR U20847 ( .A(n18801), .B(nreg[484]), .Z(n18792) );
  IV U20848 ( .A(n18790), .Z(n18801) );
  XOR U20849 ( .A(n18802), .B(n18803), .Z(n18790) );
  AND U20850 ( .A(n18804), .B(n18805), .Z(n18803) );
  XNOR U20851 ( .A(n18802), .B(n9403), .Z(n18805) );
  XNOR U20852 ( .A(n18798), .B(n18800), .Z(n9403) );
  NAND U20853 ( .A(n18806), .B(nreg[483]), .Z(n18800) );
  NAND U20854 ( .A(n12326), .B(nreg[483]), .Z(n18806) );
  XNOR U20855 ( .A(n18796), .B(n18807), .Z(n18798) );
  XOR U20856 ( .A(n18808), .B(n18809), .Z(n18796) );
  AND U20857 ( .A(n18810), .B(n18811), .Z(n18809) );
  XNOR U20858 ( .A(n18812), .B(n18808), .Z(n18811) );
  XOR U20859 ( .A(n18813), .B(nreg[483]), .Z(n18804) );
  IV U20860 ( .A(n18802), .Z(n18813) );
  XOR U20861 ( .A(n18814), .B(n18815), .Z(n18802) );
  AND U20862 ( .A(n18816), .B(n18817), .Z(n18815) );
  XNOR U20863 ( .A(n18814), .B(n9409), .Z(n18817) );
  XNOR U20864 ( .A(n18810), .B(n18812), .Z(n9409) );
  NAND U20865 ( .A(n18818), .B(nreg[482]), .Z(n18812) );
  NAND U20866 ( .A(n12326), .B(nreg[482]), .Z(n18818) );
  XNOR U20867 ( .A(n18808), .B(n18819), .Z(n18810) );
  XOR U20868 ( .A(n18820), .B(n18821), .Z(n18808) );
  AND U20869 ( .A(n18822), .B(n18823), .Z(n18821) );
  XNOR U20870 ( .A(n18824), .B(n18820), .Z(n18823) );
  XOR U20871 ( .A(n18825), .B(nreg[482]), .Z(n18816) );
  IV U20872 ( .A(n18814), .Z(n18825) );
  XOR U20873 ( .A(n18826), .B(n18827), .Z(n18814) );
  AND U20874 ( .A(n18828), .B(n18829), .Z(n18827) );
  XNOR U20875 ( .A(n18826), .B(n9415), .Z(n18829) );
  XNOR U20876 ( .A(n18822), .B(n18824), .Z(n9415) );
  NAND U20877 ( .A(n18830), .B(nreg[481]), .Z(n18824) );
  NAND U20878 ( .A(n12326), .B(nreg[481]), .Z(n18830) );
  XNOR U20879 ( .A(n18820), .B(n18831), .Z(n18822) );
  XOR U20880 ( .A(n18832), .B(n18833), .Z(n18820) );
  AND U20881 ( .A(n18834), .B(n18835), .Z(n18833) );
  XNOR U20882 ( .A(n18836), .B(n18832), .Z(n18835) );
  XOR U20883 ( .A(n18837), .B(nreg[481]), .Z(n18828) );
  IV U20884 ( .A(n18826), .Z(n18837) );
  XOR U20885 ( .A(n18838), .B(n18839), .Z(n18826) );
  AND U20886 ( .A(n18840), .B(n18841), .Z(n18839) );
  XNOR U20887 ( .A(n18838), .B(n9421), .Z(n18841) );
  XNOR U20888 ( .A(n18834), .B(n18836), .Z(n9421) );
  NAND U20889 ( .A(n18842), .B(nreg[480]), .Z(n18836) );
  NAND U20890 ( .A(n12326), .B(nreg[480]), .Z(n18842) );
  XNOR U20891 ( .A(n18832), .B(n18843), .Z(n18834) );
  XOR U20892 ( .A(n18844), .B(n18845), .Z(n18832) );
  AND U20893 ( .A(n18846), .B(n18847), .Z(n18845) );
  XNOR U20894 ( .A(n18848), .B(n18844), .Z(n18847) );
  XOR U20895 ( .A(n18849), .B(nreg[480]), .Z(n18840) );
  IV U20896 ( .A(n18838), .Z(n18849) );
  XOR U20897 ( .A(n18850), .B(n18851), .Z(n18838) );
  AND U20898 ( .A(n18852), .B(n18853), .Z(n18851) );
  XNOR U20899 ( .A(n18850), .B(n9427), .Z(n18853) );
  XNOR U20900 ( .A(n18846), .B(n18848), .Z(n9427) );
  NAND U20901 ( .A(n18854), .B(nreg[479]), .Z(n18848) );
  NAND U20902 ( .A(n12326), .B(nreg[479]), .Z(n18854) );
  XNOR U20903 ( .A(n18844), .B(n18855), .Z(n18846) );
  XOR U20904 ( .A(n18856), .B(n18857), .Z(n18844) );
  AND U20905 ( .A(n18858), .B(n18859), .Z(n18857) );
  XNOR U20906 ( .A(n18860), .B(n18856), .Z(n18859) );
  XOR U20907 ( .A(n18861), .B(nreg[479]), .Z(n18852) );
  IV U20908 ( .A(n18850), .Z(n18861) );
  XOR U20909 ( .A(n18862), .B(n18863), .Z(n18850) );
  AND U20910 ( .A(n18864), .B(n18865), .Z(n18863) );
  XNOR U20911 ( .A(n18862), .B(n9433), .Z(n18865) );
  XNOR U20912 ( .A(n18858), .B(n18860), .Z(n9433) );
  NAND U20913 ( .A(n18866), .B(nreg[478]), .Z(n18860) );
  NAND U20914 ( .A(n12326), .B(nreg[478]), .Z(n18866) );
  XNOR U20915 ( .A(n18856), .B(n18867), .Z(n18858) );
  XOR U20916 ( .A(n18868), .B(n18869), .Z(n18856) );
  AND U20917 ( .A(n18870), .B(n18871), .Z(n18869) );
  XNOR U20918 ( .A(n18872), .B(n18868), .Z(n18871) );
  XOR U20919 ( .A(n18873), .B(nreg[478]), .Z(n18864) );
  IV U20920 ( .A(n18862), .Z(n18873) );
  XOR U20921 ( .A(n18874), .B(n18875), .Z(n18862) );
  AND U20922 ( .A(n18876), .B(n18877), .Z(n18875) );
  XNOR U20923 ( .A(n18874), .B(n9439), .Z(n18877) );
  XNOR U20924 ( .A(n18870), .B(n18872), .Z(n9439) );
  NAND U20925 ( .A(n18878), .B(nreg[477]), .Z(n18872) );
  NAND U20926 ( .A(n12326), .B(nreg[477]), .Z(n18878) );
  XNOR U20927 ( .A(n18868), .B(n18879), .Z(n18870) );
  XOR U20928 ( .A(n18880), .B(n18881), .Z(n18868) );
  AND U20929 ( .A(n18882), .B(n18883), .Z(n18881) );
  XNOR U20930 ( .A(n18884), .B(n18880), .Z(n18883) );
  XOR U20931 ( .A(n18885), .B(nreg[477]), .Z(n18876) );
  IV U20932 ( .A(n18874), .Z(n18885) );
  XOR U20933 ( .A(n18886), .B(n18887), .Z(n18874) );
  AND U20934 ( .A(n18888), .B(n18889), .Z(n18887) );
  XNOR U20935 ( .A(n18886), .B(n9445), .Z(n18889) );
  XNOR U20936 ( .A(n18882), .B(n18884), .Z(n9445) );
  NAND U20937 ( .A(n18890), .B(nreg[476]), .Z(n18884) );
  NAND U20938 ( .A(n12326), .B(nreg[476]), .Z(n18890) );
  XNOR U20939 ( .A(n18880), .B(n18891), .Z(n18882) );
  XOR U20940 ( .A(n18892), .B(n18893), .Z(n18880) );
  AND U20941 ( .A(n18894), .B(n18895), .Z(n18893) );
  XNOR U20942 ( .A(n18896), .B(n18892), .Z(n18895) );
  XOR U20943 ( .A(n18897), .B(nreg[476]), .Z(n18888) );
  IV U20944 ( .A(n18886), .Z(n18897) );
  XOR U20945 ( .A(n18898), .B(n18899), .Z(n18886) );
  AND U20946 ( .A(n18900), .B(n18901), .Z(n18899) );
  XNOR U20947 ( .A(n18898), .B(n9451), .Z(n18901) );
  XNOR U20948 ( .A(n18894), .B(n18896), .Z(n9451) );
  NAND U20949 ( .A(n18902), .B(nreg[475]), .Z(n18896) );
  NAND U20950 ( .A(n12326), .B(nreg[475]), .Z(n18902) );
  XNOR U20951 ( .A(n18892), .B(n18903), .Z(n18894) );
  XOR U20952 ( .A(n18904), .B(n18905), .Z(n18892) );
  AND U20953 ( .A(n18906), .B(n18907), .Z(n18905) );
  XNOR U20954 ( .A(n18908), .B(n18904), .Z(n18907) );
  XOR U20955 ( .A(n18909), .B(nreg[475]), .Z(n18900) );
  IV U20956 ( .A(n18898), .Z(n18909) );
  XOR U20957 ( .A(n18910), .B(n18911), .Z(n18898) );
  AND U20958 ( .A(n18912), .B(n18913), .Z(n18911) );
  XNOR U20959 ( .A(n18910), .B(n9457), .Z(n18913) );
  XNOR U20960 ( .A(n18906), .B(n18908), .Z(n9457) );
  NAND U20961 ( .A(n18914), .B(nreg[474]), .Z(n18908) );
  NAND U20962 ( .A(n12326), .B(nreg[474]), .Z(n18914) );
  XNOR U20963 ( .A(n18904), .B(n18915), .Z(n18906) );
  XOR U20964 ( .A(n18916), .B(n18917), .Z(n18904) );
  AND U20965 ( .A(n18918), .B(n18919), .Z(n18917) );
  XNOR U20966 ( .A(n18920), .B(n18916), .Z(n18919) );
  XOR U20967 ( .A(n18921), .B(nreg[474]), .Z(n18912) );
  IV U20968 ( .A(n18910), .Z(n18921) );
  XOR U20969 ( .A(n18922), .B(n18923), .Z(n18910) );
  AND U20970 ( .A(n18924), .B(n18925), .Z(n18923) );
  XNOR U20971 ( .A(n18922), .B(n9463), .Z(n18925) );
  XNOR U20972 ( .A(n18918), .B(n18920), .Z(n9463) );
  NAND U20973 ( .A(n18926), .B(nreg[473]), .Z(n18920) );
  NAND U20974 ( .A(n12326), .B(nreg[473]), .Z(n18926) );
  XNOR U20975 ( .A(n18916), .B(n18927), .Z(n18918) );
  XOR U20976 ( .A(n18928), .B(n18929), .Z(n18916) );
  AND U20977 ( .A(n18930), .B(n18931), .Z(n18929) );
  XNOR U20978 ( .A(n18932), .B(n18928), .Z(n18931) );
  XOR U20979 ( .A(n18933), .B(nreg[473]), .Z(n18924) );
  IV U20980 ( .A(n18922), .Z(n18933) );
  XOR U20981 ( .A(n18934), .B(n18935), .Z(n18922) );
  AND U20982 ( .A(n18936), .B(n18937), .Z(n18935) );
  XNOR U20983 ( .A(n18934), .B(n9469), .Z(n18937) );
  XNOR U20984 ( .A(n18930), .B(n18932), .Z(n9469) );
  NAND U20985 ( .A(n18938), .B(nreg[472]), .Z(n18932) );
  NAND U20986 ( .A(n12326), .B(nreg[472]), .Z(n18938) );
  XNOR U20987 ( .A(n18928), .B(n18939), .Z(n18930) );
  XOR U20988 ( .A(n18940), .B(n18941), .Z(n18928) );
  AND U20989 ( .A(n18942), .B(n18943), .Z(n18941) );
  XNOR U20990 ( .A(n18944), .B(n18940), .Z(n18943) );
  XOR U20991 ( .A(n18945), .B(nreg[472]), .Z(n18936) );
  IV U20992 ( .A(n18934), .Z(n18945) );
  XOR U20993 ( .A(n18946), .B(n18947), .Z(n18934) );
  AND U20994 ( .A(n18948), .B(n18949), .Z(n18947) );
  XNOR U20995 ( .A(n18946), .B(n9475), .Z(n18949) );
  XNOR U20996 ( .A(n18942), .B(n18944), .Z(n9475) );
  NAND U20997 ( .A(n18950), .B(nreg[471]), .Z(n18944) );
  NAND U20998 ( .A(n12326), .B(nreg[471]), .Z(n18950) );
  XNOR U20999 ( .A(n18940), .B(n18951), .Z(n18942) );
  XOR U21000 ( .A(n18952), .B(n18953), .Z(n18940) );
  AND U21001 ( .A(n18954), .B(n18955), .Z(n18953) );
  XNOR U21002 ( .A(n18956), .B(n18952), .Z(n18955) );
  XOR U21003 ( .A(n18957), .B(nreg[471]), .Z(n18948) );
  IV U21004 ( .A(n18946), .Z(n18957) );
  XOR U21005 ( .A(n18958), .B(n18959), .Z(n18946) );
  AND U21006 ( .A(n18960), .B(n18961), .Z(n18959) );
  XNOR U21007 ( .A(n18958), .B(n9481), .Z(n18961) );
  XNOR U21008 ( .A(n18954), .B(n18956), .Z(n9481) );
  NAND U21009 ( .A(n18962), .B(nreg[470]), .Z(n18956) );
  NAND U21010 ( .A(n12326), .B(nreg[470]), .Z(n18962) );
  XNOR U21011 ( .A(n18952), .B(n18963), .Z(n18954) );
  XOR U21012 ( .A(n18964), .B(n18965), .Z(n18952) );
  AND U21013 ( .A(n18966), .B(n18967), .Z(n18965) );
  XNOR U21014 ( .A(n18968), .B(n18964), .Z(n18967) );
  XOR U21015 ( .A(n18969), .B(nreg[470]), .Z(n18960) );
  IV U21016 ( .A(n18958), .Z(n18969) );
  XOR U21017 ( .A(n18970), .B(n18971), .Z(n18958) );
  AND U21018 ( .A(n18972), .B(n18973), .Z(n18971) );
  XNOR U21019 ( .A(n18970), .B(n9487), .Z(n18973) );
  XNOR U21020 ( .A(n18966), .B(n18968), .Z(n9487) );
  NAND U21021 ( .A(n18974), .B(nreg[469]), .Z(n18968) );
  NAND U21022 ( .A(n12326), .B(nreg[469]), .Z(n18974) );
  XNOR U21023 ( .A(n18964), .B(n18975), .Z(n18966) );
  XOR U21024 ( .A(n18976), .B(n18977), .Z(n18964) );
  AND U21025 ( .A(n18978), .B(n18979), .Z(n18977) );
  XNOR U21026 ( .A(n18980), .B(n18976), .Z(n18979) );
  XOR U21027 ( .A(n18981), .B(nreg[469]), .Z(n18972) );
  IV U21028 ( .A(n18970), .Z(n18981) );
  XOR U21029 ( .A(n18982), .B(n18983), .Z(n18970) );
  AND U21030 ( .A(n18984), .B(n18985), .Z(n18983) );
  XNOR U21031 ( .A(n18982), .B(n9493), .Z(n18985) );
  XNOR U21032 ( .A(n18978), .B(n18980), .Z(n9493) );
  NAND U21033 ( .A(n18986), .B(nreg[468]), .Z(n18980) );
  NAND U21034 ( .A(n12326), .B(nreg[468]), .Z(n18986) );
  XNOR U21035 ( .A(n18976), .B(n18987), .Z(n18978) );
  XOR U21036 ( .A(n18988), .B(n18989), .Z(n18976) );
  AND U21037 ( .A(n18990), .B(n18991), .Z(n18989) );
  XNOR U21038 ( .A(n18992), .B(n18988), .Z(n18991) );
  XOR U21039 ( .A(n18993), .B(nreg[468]), .Z(n18984) );
  IV U21040 ( .A(n18982), .Z(n18993) );
  XOR U21041 ( .A(n18994), .B(n18995), .Z(n18982) );
  AND U21042 ( .A(n18996), .B(n18997), .Z(n18995) );
  XNOR U21043 ( .A(n18994), .B(n9499), .Z(n18997) );
  XNOR U21044 ( .A(n18990), .B(n18992), .Z(n9499) );
  NAND U21045 ( .A(n18998), .B(nreg[467]), .Z(n18992) );
  NAND U21046 ( .A(n12326), .B(nreg[467]), .Z(n18998) );
  XNOR U21047 ( .A(n18988), .B(n18999), .Z(n18990) );
  XOR U21048 ( .A(n19000), .B(n19001), .Z(n18988) );
  AND U21049 ( .A(n19002), .B(n19003), .Z(n19001) );
  XNOR U21050 ( .A(n19004), .B(n19000), .Z(n19003) );
  XOR U21051 ( .A(n19005), .B(nreg[467]), .Z(n18996) );
  IV U21052 ( .A(n18994), .Z(n19005) );
  XOR U21053 ( .A(n19006), .B(n19007), .Z(n18994) );
  AND U21054 ( .A(n19008), .B(n19009), .Z(n19007) );
  XNOR U21055 ( .A(n19006), .B(n9505), .Z(n19009) );
  XNOR U21056 ( .A(n19002), .B(n19004), .Z(n9505) );
  NAND U21057 ( .A(n19010), .B(nreg[466]), .Z(n19004) );
  NAND U21058 ( .A(n12326), .B(nreg[466]), .Z(n19010) );
  XNOR U21059 ( .A(n19000), .B(n19011), .Z(n19002) );
  XOR U21060 ( .A(n19012), .B(n19013), .Z(n19000) );
  AND U21061 ( .A(n19014), .B(n19015), .Z(n19013) );
  XNOR U21062 ( .A(n19016), .B(n19012), .Z(n19015) );
  XOR U21063 ( .A(n19017), .B(nreg[466]), .Z(n19008) );
  IV U21064 ( .A(n19006), .Z(n19017) );
  XOR U21065 ( .A(n19018), .B(n19019), .Z(n19006) );
  AND U21066 ( .A(n19020), .B(n19021), .Z(n19019) );
  XNOR U21067 ( .A(n19018), .B(n9511), .Z(n19021) );
  XNOR U21068 ( .A(n19014), .B(n19016), .Z(n9511) );
  NAND U21069 ( .A(n19022), .B(nreg[465]), .Z(n19016) );
  NAND U21070 ( .A(n12326), .B(nreg[465]), .Z(n19022) );
  XNOR U21071 ( .A(n19012), .B(n19023), .Z(n19014) );
  XOR U21072 ( .A(n19024), .B(n19025), .Z(n19012) );
  AND U21073 ( .A(n19026), .B(n19027), .Z(n19025) );
  XNOR U21074 ( .A(n19028), .B(n19024), .Z(n19027) );
  XOR U21075 ( .A(n19029), .B(nreg[465]), .Z(n19020) );
  IV U21076 ( .A(n19018), .Z(n19029) );
  XOR U21077 ( .A(n19030), .B(n19031), .Z(n19018) );
  AND U21078 ( .A(n19032), .B(n19033), .Z(n19031) );
  XNOR U21079 ( .A(n19030), .B(n9517), .Z(n19033) );
  XNOR U21080 ( .A(n19026), .B(n19028), .Z(n9517) );
  NAND U21081 ( .A(n19034), .B(nreg[464]), .Z(n19028) );
  NAND U21082 ( .A(n12326), .B(nreg[464]), .Z(n19034) );
  XNOR U21083 ( .A(n19024), .B(n19035), .Z(n19026) );
  XOR U21084 ( .A(n19036), .B(n19037), .Z(n19024) );
  AND U21085 ( .A(n19038), .B(n19039), .Z(n19037) );
  XNOR U21086 ( .A(n19040), .B(n19036), .Z(n19039) );
  XOR U21087 ( .A(n19041), .B(nreg[464]), .Z(n19032) );
  IV U21088 ( .A(n19030), .Z(n19041) );
  XOR U21089 ( .A(n19042), .B(n19043), .Z(n19030) );
  AND U21090 ( .A(n19044), .B(n19045), .Z(n19043) );
  XNOR U21091 ( .A(n19042), .B(n9523), .Z(n19045) );
  XNOR U21092 ( .A(n19038), .B(n19040), .Z(n9523) );
  NAND U21093 ( .A(n19046), .B(nreg[463]), .Z(n19040) );
  NAND U21094 ( .A(n12326), .B(nreg[463]), .Z(n19046) );
  XNOR U21095 ( .A(n19036), .B(n19047), .Z(n19038) );
  XOR U21096 ( .A(n19048), .B(n19049), .Z(n19036) );
  AND U21097 ( .A(n19050), .B(n19051), .Z(n19049) );
  XNOR U21098 ( .A(n19052), .B(n19048), .Z(n19051) );
  XOR U21099 ( .A(n19053), .B(nreg[463]), .Z(n19044) );
  IV U21100 ( .A(n19042), .Z(n19053) );
  XOR U21101 ( .A(n19054), .B(n19055), .Z(n19042) );
  AND U21102 ( .A(n19056), .B(n19057), .Z(n19055) );
  XNOR U21103 ( .A(n19054), .B(n9529), .Z(n19057) );
  XNOR U21104 ( .A(n19050), .B(n19052), .Z(n9529) );
  NAND U21105 ( .A(n19058), .B(nreg[462]), .Z(n19052) );
  NAND U21106 ( .A(n12326), .B(nreg[462]), .Z(n19058) );
  XNOR U21107 ( .A(n19048), .B(n19059), .Z(n19050) );
  XOR U21108 ( .A(n19060), .B(n19061), .Z(n19048) );
  AND U21109 ( .A(n19062), .B(n19063), .Z(n19061) );
  XNOR U21110 ( .A(n19064), .B(n19060), .Z(n19063) );
  XOR U21111 ( .A(n19065), .B(nreg[462]), .Z(n19056) );
  IV U21112 ( .A(n19054), .Z(n19065) );
  XOR U21113 ( .A(n19066), .B(n19067), .Z(n19054) );
  AND U21114 ( .A(n19068), .B(n19069), .Z(n19067) );
  XNOR U21115 ( .A(n19066), .B(n9535), .Z(n19069) );
  XNOR U21116 ( .A(n19062), .B(n19064), .Z(n9535) );
  NAND U21117 ( .A(n19070), .B(nreg[461]), .Z(n19064) );
  NAND U21118 ( .A(n12326), .B(nreg[461]), .Z(n19070) );
  XNOR U21119 ( .A(n19060), .B(n19071), .Z(n19062) );
  XOR U21120 ( .A(n19072), .B(n19073), .Z(n19060) );
  AND U21121 ( .A(n19074), .B(n19075), .Z(n19073) );
  XNOR U21122 ( .A(n19076), .B(n19072), .Z(n19075) );
  XOR U21123 ( .A(n19077), .B(nreg[461]), .Z(n19068) );
  IV U21124 ( .A(n19066), .Z(n19077) );
  XOR U21125 ( .A(n19078), .B(n19079), .Z(n19066) );
  AND U21126 ( .A(n19080), .B(n19081), .Z(n19079) );
  XNOR U21127 ( .A(n19078), .B(n9541), .Z(n19081) );
  XNOR U21128 ( .A(n19074), .B(n19076), .Z(n9541) );
  NAND U21129 ( .A(n19082), .B(nreg[460]), .Z(n19076) );
  NAND U21130 ( .A(n12326), .B(nreg[460]), .Z(n19082) );
  XNOR U21131 ( .A(n19072), .B(n19083), .Z(n19074) );
  XOR U21132 ( .A(n19084), .B(n19085), .Z(n19072) );
  AND U21133 ( .A(n19086), .B(n19087), .Z(n19085) );
  XNOR U21134 ( .A(n19088), .B(n19084), .Z(n19087) );
  XOR U21135 ( .A(n19089), .B(nreg[460]), .Z(n19080) );
  IV U21136 ( .A(n19078), .Z(n19089) );
  XOR U21137 ( .A(n19090), .B(n19091), .Z(n19078) );
  AND U21138 ( .A(n19092), .B(n19093), .Z(n19091) );
  XNOR U21139 ( .A(n19090), .B(n9547), .Z(n19093) );
  XNOR U21140 ( .A(n19086), .B(n19088), .Z(n9547) );
  NAND U21141 ( .A(n19094), .B(nreg[459]), .Z(n19088) );
  NAND U21142 ( .A(n12326), .B(nreg[459]), .Z(n19094) );
  XNOR U21143 ( .A(n19084), .B(n19095), .Z(n19086) );
  XOR U21144 ( .A(n19096), .B(n19097), .Z(n19084) );
  AND U21145 ( .A(n19098), .B(n19099), .Z(n19097) );
  XNOR U21146 ( .A(n19100), .B(n19096), .Z(n19099) );
  XOR U21147 ( .A(n19101), .B(nreg[459]), .Z(n19092) );
  IV U21148 ( .A(n19090), .Z(n19101) );
  XOR U21149 ( .A(n19102), .B(n19103), .Z(n19090) );
  AND U21150 ( .A(n19104), .B(n19105), .Z(n19103) );
  XNOR U21151 ( .A(n19102), .B(n9553), .Z(n19105) );
  XNOR U21152 ( .A(n19098), .B(n19100), .Z(n9553) );
  NAND U21153 ( .A(n19106), .B(nreg[458]), .Z(n19100) );
  NAND U21154 ( .A(n12326), .B(nreg[458]), .Z(n19106) );
  XNOR U21155 ( .A(n19096), .B(n19107), .Z(n19098) );
  XOR U21156 ( .A(n19108), .B(n19109), .Z(n19096) );
  AND U21157 ( .A(n19110), .B(n19111), .Z(n19109) );
  XNOR U21158 ( .A(n19112), .B(n19108), .Z(n19111) );
  XOR U21159 ( .A(n19113), .B(nreg[458]), .Z(n19104) );
  IV U21160 ( .A(n19102), .Z(n19113) );
  XOR U21161 ( .A(n19114), .B(n19115), .Z(n19102) );
  AND U21162 ( .A(n19116), .B(n19117), .Z(n19115) );
  XNOR U21163 ( .A(n19114), .B(n9559), .Z(n19117) );
  XNOR U21164 ( .A(n19110), .B(n19112), .Z(n9559) );
  NAND U21165 ( .A(n19118), .B(nreg[457]), .Z(n19112) );
  NAND U21166 ( .A(n12326), .B(nreg[457]), .Z(n19118) );
  XNOR U21167 ( .A(n19108), .B(n19119), .Z(n19110) );
  XOR U21168 ( .A(n19120), .B(n19121), .Z(n19108) );
  AND U21169 ( .A(n19122), .B(n19123), .Z(n19121) );
  XNOR U21170 ( .A(n19124), .B(n19120), .Z(n19123) );
  XOR U21171 ( .A(n19125), .B(nreg[457]), .Z(n19116) );
  IV U21172 ( .A(n19114), .Z(n19125) );
  XOR U21173 ( .A(n19126), .B(n19127), .Z(n19114) );
  AND U21174 ( .A(n19128), .B(n19129), .Z(n19127) );
  XNOR U21175 ( .A(n19126), .B(n9565), .Z(n19129) );
  XNOR U21176 ( .A(n19122), .B(n19124), .Z(n9565) );
  NAND U21177 ( .A(n19130), .B(nreg[456]), .Z(n19124) );
  NAND U21178 ( .A(n12326), .B(nreg[456]), .Z(n19130) );
  XNOR U21179 ( .A(n19120), .B(n19131), .Z(n19122) );
  XOR U21180 ( .A(n19132), .B(n19133), .Z(n19120) );
  AND U21181 ( .A(n19134), .B(n19135), .Z(n19133) );
  XNOR U21182 ( .A(n19136), .B(n19132), .Z(n19135) );
  XOR U21183 ( .A(n19137), .B(nreg[456]), .Z(n19128) );
  IV U21184 ( .A(n19126), .Z(n19137) );
  XOR U21185 ( .A(n19138), .B(n19139), .Z(n19126) );
  AND U21186 ( .A(n19140), .B(n19141), .Z(n19139) );
  XNOR U21187 ( .A(n19138), .B(n9571), .Z(n19141) );
  XNOR U21188 ( .A(n19134), .B(n19136), .Z(n9571) );
  NAND U21189 ( .A(n19142), .B(nreg[455]), .Z(n19136) );
  NAND U21190 ( .A(n12326), .B(nreg[455]), .Z(n19142) );
  XNOR U21191 ( .A(n19132), .B(n19143), .Z(n19134) );
  XOR U21192 ( .A(n19144), .B(n19145), .Z(n19132) );
  AND U21193 ( .A(n19146), .B(n19147), .Z(n19145) );
  XNOR U21194 ( .A(n19148), .B(n19144), .Z(n19147) );
  XOR U21195 ( .A(n19149), .B(nreg[455]), .Z(n19140) );
  IV U21196 ( .A(n19138), .Z(n19149) );
  XOR U21197 ( .A(n19150), .B(n19151), .Z(n19138) );
  AND U21198 ( .A(n19152), .B(n19153), .Z(n19151) );
  XNOR U21199 ( .A(n19150), .B(n9577), .Z(n19153) );
  XNOR U21200 ( .A(n19146), .B(n19148), .Z(n9577) );
  NAND U21201 ( .A(n19154), .B(nreg[454]), .Z(n19148) );
  NAND U21202 ( .A(n12326), .B(nreg[454]), .Z(n19154) );
  XNOR U21203 ( .A(n19144), .B(n19155), .Z(n19146) );
  XOR U21204 ( .A(n19156), .B(n19157), .Z(n19144) );
  AND U21205 ( .A(n19158), .B(n19159), .Z(n19157) );
  XNOR U21206 ( .A(n19160), .B(n19156), .Z(n19159) );
  XOR U21207 ( .A(n19161), .B(nreg[454]), .Z(n19152) );
  IV U21208 ( .A(n19150), .Z(n19161) );
  XOR U21209 ( .A(n19162), .B(n19163), .Z(n19150) );
  AND U21210 ( .A(n19164), .B(n19165), .Z(n19163) );
  XNOR U21211 ( .A(n19162), .B(n9583), .Z(n19165) );
  XNOR U21212 ( .A(n19158), .B(n19160), .Z(n9583) );
  NAND U21213 ( .A(n19166), .B(nreg[453]), .Z(n19160) );
  NAND U21214 ( .A(n12326), .B(nreg[453]), .Z(n19166) );
  XNOR U21215 ( .A(n19156), .B(n19167), .Z(n19158) );
  XOR U21216 ( .A(n19168), .B(n19169), .Z(n19156) );
  AND U21217 ( .A(n19170), .B(n19171), .Z(n19169) );
  XNOR U21218 ( .A(n19172), .B(n19168), .Z(n19171) );
  XOR U21219 ( .A(n19173), .B(nreg[453]), .Z(n19164) );
  IV U21220 ( .A(n19162), .Z(n19173) );
  XOR U21221 ( .A(n19174), .B(n19175), .Z(n19162) );
  AND U21222 ( .A(n19176), .B(n19177), .Z(n19175) );
  XNOR U21223 ( .A(n19174), .B(n9589), .Z(n19177) );
  XNOR U21224 ( .A(n19170), .B(n19172), .Z(n9589) );
  NAND U21225 ( .A(n19178), .B(nreg[452]), .Z(n19172) );
  NAND U21226 ( .A(n12326), .B(nreg[452]), .Z(n19178) );
  XNOR U21227 ( .A(n19168), .B(n19179), .Z(n19170) );
  XOR U21228 ( .A(n19180), .B(n19181), .Z(n19168) );
  AND U21229 ( .A(n19182), .B(n19183), .Z(n19181) );
  XNOR U21230 ( .A(n19184), .B(n19180), .Z(n19183) );
  XOR U21231 ( .A(n19185), .B(nreg[452]), .Z(n19176) );
  IV U21232 ( .A(n19174), .Z(n19185) );
  XOR U21233 ( .A(n19186), .B(n19187), .Z(n19174) );
  AND U21234 ( .A(n19188), .B(n19189), .Z(n19187) );
  XNOR U21235 ( .A(n19186), .B(n9595), .Z(n19189) );
  XNOR U21236 ( .A(n19182), .B(n19184), .Z(n9595) );
  NAND U21237 ( .A(n19190), .B(nreg[451]), .Z(n19184) );
  NAND U21238 ( .A(n12326), .B(nreg[451]), .Z(n19190) );
  XNOR U21239 ( .A(n19180), .B(n19191), .Z(n19182) );
  XOR U21240 ( .A(n19192), .B(n19193), .Z(n19180) );
  AND U21241 ( .A(n19194), .B(n19195), .Z(n19193) );
  XNOR U21242 ( .A(n19196), .B(n19192), .Z(n19195) );
  XOR U21243 ( .A(n19197), .B(nreg[451]), .Z(n19188) );
  IV U21244 ( .A(n19186), .Z(n19197) );
  XOR U21245 ( .A(n19198), .B(n19199), .Z(n19186) );
  AND U21246 ( .A(n19200), .B(n19201), .Z(n19199) );
  XNOR U21247 ( .A(n19198), .B(n9601), .Z(n19201) );
  XNOR U21248 ( .A(n19194), .B(n19196), .Z(n9601) );
  NAND U21249 ( .A(n19202), .B(nreg[450]), .Z(n19196) );
  NAND U21250 ( .A(n12326), .B(nreg[450]), .Z(n19202) );
  XNOR U21251 ( .A(n19192), .B(n19203), .Z(n19194) );
  XOR U21252 ( .A(n19204), .B(n19205), .Z(n19192) );
  AND U21253 ( .A(n19206), .B(n19207), .Z(n19205) );
  XNOR U21254 ( .A(n19208), .B(n19204), .Z(n19207) );
  XOR U21255 ( .A(n19209), .B(nreg[450]), .Z(n19200) );
  IV U21256 ( .A(n19198), .Z(n19209) );
  XOR U21257 ( .A(n19210), .B(n19211), .Z(n19198) );
  AND U21258 ( .A(n19212), .B(n19213), .Z(n19211) );
  XNOR U21259 ( .A(n19210), .B(n9607), .Z(n19213) );
  XNOR U21260 ( .A(n19206), .B(n19208), .Z(n9607) );
  NAND U21261 ( .A(n19214), .B(nreg[449]), .Z(n19208) );
  NAND U21262 ( .A(n12326), .B(nreg[449]), .Z(n19214) );
  XNOR U21263 ( .A(n19204), .B(n19215), .Z(n19206) );
  XOR U21264 ( .A(n19216), .B(n19217), .Z(n19204) );
  AND U21265 ( .A(n19218), .B(n19219), .Z(n19217) );
  XNOR U21266 ( .A(n19220), .B(n19216), .Z(n19219) );
  XOR U21267 ( .A(n19221), .B(nreg[449]), .Z(n19212) );
  IV U21268 ( .A(n19210), .Z(n19221) );
  XOR U21269 ( .A(n19222), .B(n19223), .Z(n19210) );
  AND U21270 ( .A(n19224), .B(n19225), .Z(n19223) );
  XNOR U21271 ( .A(n19222), .B(n9613), .Z(n19225) );
  XNOR U21272 ( .A(n19218), .B(n19220), .Z(n9613) );
  NAND U21273 ( .A(n19226), .B(nreg[448]), .Z(n19220) );
  NAND U21274 ( .A(n12326), .B(nreg[448]), .Z(n19226) );
  XNOR U21275 ( .A(n19216), .B(n19227), .Z(n19218) );
  XOR U21276 ( .A(n19228), .B(n19229), .Z(n19216) );
  AND U21277 ( .A(n19230), .B(n19231), .Z(n19229) );
  XNOR U21278 ( .A(n19232), .B(n19228), .Z(n19231) );
  XOR U21279 ( .A(n19233), .B(nreg[448]), .Z(n19224) );
  IV U21280 ( .A(n19222), .Z(n19233) );
  XOR U21281 ( .A(n19234), .B(n19235), .Z(n19222) );
  AND U21282 ( .A(n19236), .B(n19237), .Z(n19235) );
  XNOR U21283 ( .A(n19234), .B(n9619), .Z(n19237) );
  XNOR U21284 ( .A(n19230), .B(n19232), .Z(n9619) );
  NAND U21285 ( .A(n19238), .B(nreg[447]), .Z(n19232) );
  NAND U21286 ( .A(n12326), .B(nreg[447]), .Z(n19238) );
  XNOR U21287 ( .A(n19228), .B(n19239), .Z(n19230) );
  XOR U21288 ( .A(n19240), .B(n19241), .Z(n19228) );
  AND U21289 ( .A(n19242), .B(n19243), .Z(n19241) );
  XNOR U21290 ( .A(n19244), .B(n19240), .Z(n19243) );
  XOR U21291 ( .A(n19245), .B(nreg[447]), .Z(n19236) );
  IV U21292 ( .A(n19234), .Z(n19245) );
  XOR U21293 ( .A(n19246), .B(n19247), .Z(n19234) );
  AND U21294 ( .A(n19248), .B(n19249), .Z(n19247) );
  XNOR U21295 ( .A(n19246), .B(n9625), .Z(n19249) );
  XNOR U21296 ( .A(n19242), .B(n19244), .Z(n9625) );
  NAND U21297 ( .A(n19250), .B(nreg[446]), .Z(n19244) );
  NAND U21298 ( .A(n12326), .B(nreg[446]), .Z(n19250) );
  XNOR U21299 ( .A(n19240), .B(n19251), .Z(n19242) );
  XOR U21300 ( .A(n19252), .B(n19253), .Z(n19240) );
  AND U21301 ( .A(n19254), .B(n19255), .Z(n19253) );
  XNOR U21302 ( .A(n19256), .B(n19252), .Z(n19255) );
  XOR U21303 ( .A(n19257), .B(nreg[446]), .Z(n19248) );
  IV U21304 ( .A(n19246), .Z(n19257) );
  XOR U21305 ( .A(n19258), .B(n19259), .Z(n19246) );
  AND U21306 ( .A(n19260), .B(n19261), .Z(n19259) );
  XNOR U21307 ( .A(n19258), .B(n9631), .Z(n19261) );
  XNOR U21308 ( .A(n19254), .B(n19256), .Z(n9631) );
  NAND U21309 ( .A(n19262), .B(nreg[445]), .Z(n19256) );
  NAND U21310 ( .A(n12326), .B(nreg[445]), .Z(n19262) );
  XNOR U21311 ( .A(n19252), .B(n19263), .Z(n19254) );
  XOR U21312 ( .A(n19264), .B(n19265), .Z(n19252) );
  AND U21313 ( .A(n19266), .B(n19267), .Z(n19265) );
  XNOR U21314 ( .A(n19268), .B(n19264), .Z(n19267) );
  XOR U21315 ( .A(n19269), .B(nreg[445]), .Z(n19260) );
  IV U21316 ( .A(n19258), .Z(n19269) );
  XOR U21317 ( .A(n19270), .B(n19271), .Z(n19258) );
  AND U21318 ( .A(n19272), .B(n19273), .Z(n19271) );
  XNOR U21319 ( .A(n19270), .B(n9637), .Z(n19273) );
  XNOR U21320 ( .A(n19266), .B(n19268), .Z(n9637) );
  NAND U21321 ( .A(n19274), .B(nreg[444]), .Z(n19268) );
  NAND U21322 ( .A(n12326), .B(nreg[444]), .Z(n19274) );
  XNOR U21323 ( .A(n19264), .B(n19275), .Z(n19266) );
  XOR U21324 ( .A(n19276), .B(n19277), .Z(n19264) );
  AND U21325 ( .A(n19278), .B(n19279), .Z(n19277) );
  XNOR U21326 ( .A(n19280), .B(n19276), .Z(n19279) );
  XOR U21327 ( .A(n19281), .B(nreg[444]), .Z(n19272) );
  IV U21328 ( .A(n19270), .Z(n19281) );
  XOR U21329 ( .A(n19282), .B(n19283), .Z(n19270) );
  AND U21330 ( .A(n19284), .B(n19285), .Z(n19283) );
  XNOR U21331 ( .A(n19282), .B(n9643), .Z(n19285) );
  XNOR U21332 ( .A(n19278), .B(n19280), .Z(n9643) );
  NAND U21333 ( .A(n19286), .B(nreg[443]), .Z(n19280) );
  NAND U21334 ( .A(n12326), .B(nreg[443]), .Z(n19286) );
  XNOR U21335 ( .A(n19276), .B(n19287), .Z(n19278) );
  XOR U21336 ( .A(n19288), .B(n19289), .Z(n19276) );
  AND U21337 ( .A(n19290), .B(n19291), .Z(n19289) );
  XNOR U21338 ( .A(n19292), .B(n19288), .Z(n19291) );
  XOR U21339 ( .A(n19293), .B(nreg[443]), .Z(n19284) );
  IV U21340 ( .A(n19282), .Z(n19293) );
  XOR U21341 ( .A(n19294), .B(n19295), .Z(n19282) );
  AND U21342 ( .A(n19296), .B(n19297), .Z(n19295) );
  XNOR U21343 ( .A(n19294), .B(n9649), .Z(n19297) );
  XNOR U21344 ( .A(n19290), .B(n19292), .Z(n9649) );
  NAND U21345 ( .A(n19298), .B(nreg[442]), .Z(n19292) );
  NAND U21346 ( .A(n12326), .B(nreg[442]), .Z(n19298) );
  XNOR U21347 ( .A(n19288), .B(n19299), .Z(n19290) );
  XOR U21348 ( .A(n19300), .B(n19301), .Z(n19288) );
  AND U21349 ( .A(n19302), .B(n19303), .Z(n19301) );
  XNOR U21350 ( .A(n19304), .B(n19300), .Z(n19303) );
  XOR U21351 ( .A(n19305), .B(nreg[442]), .Z(n19296) );
  IV U21352 ( .A(n19294), .Z(n19305) );
  XOR U21353 ( .A(n19306), .B(n19307), .Z(n19294) );
  AND U21354 ( .A(n19308), .B(n19309), .Z(n19307) );
  XNOR U21355 ( .A(n19306), .B(n9655), .Z(n19309) );
  XNOR U21356 ( .A(n19302), .B(n19304), .Z(n9655) );
  NAND U21357 ( .A(n19310), .B(nreg[441]), .Z(n19304) );
  NAND U21358 ( .A(n12326), .B(nreg[441]), .Z(n19310) );
  XNOR U21359 ( .A(n19300), .B(n19311), .Z(n19302) );
  XOR U21360 ( .A(n19312), .B(n19313), .Z(n19300) );
  AND U21361 ( .A(n19314), .B(n19315), .Z(n19313) );
  XNOR U21362 ( .A(n19316), .B(n19312), .Z(n19315) );
  XOR U21363 ( .A(n19317), .B(nreg[441]), .Z(n19308) );
  IV U21364 ( .A(n19306), .Z(n19317) );
  XOR U21365 ( .A(n19318), .B(n19319), .Z(n19306) );
  AND U21366 ( .A(n19320), .B(n19321), .Z(n19319) );
  XNOR U21367 ( .A(n19318), .B(n9661), .Z(n19321) );
  XNOR U21368 ( .A(n19314), .B(n19316), .Z(n9661) );
  NAND U21369 ( .A(n19322), .B(nreg[440]), .Z(n19316) );
  NAND U21370 ( .A(n12326), .B(nreg[440]), .Z(n19322) );
  XNOR U21371 ( .A(n19312), .B(n19323), .Z(n19314) );
  XOR U21372 ( .A(n19324), .B(n19325), .Z(n19312) );
  AND U21373 ( .A(n19326), .B(n19327), .Z(n19325) );
  XNOR U21374 ( .A(n19328), .B(n19324), .Z(n19327) );
  XOR U21375 ( .A(n19329), .B(nreg[440]), .Z(n19320) );
  IV U21376 ( .A(n19318), .Z(n19329) );
  XOR U21377 ( .A(n19330), .B(n19331), .Z(n19318) );
  AND U21378 ( .A(n19332), .B(n19333), .Z(n19331) );
  XNOR U21379 ( .A(n19330), .B(n9667), .Z(n19333) );
  XNOR U21380 ( .A(n19326), .B(n19328), .Z(n9667) );
  NAND U21381 ( .A(n19334), .B(nreg[439]), .Z(n19328) );
  NAND U21382 ( .A(n12326), .B(nreg[439]), .Z(n19334) );
  XNOR U21383 ( .A(n19324), .B(n19335), .Z(n19326) );
  XOR U21384 ( .A(n19336), .B(n19337), .Z(n19324) );
  AND U21385 ( .A(n19338), .B(n19339), .Z(n19337) );
  XNOR U21386 ( .A(n19340), .B(n19336), .Z(n19339) );
  XOR U21387 ( .A(n19341), .B(nreg[439]), .Z(n19332) );
  IV U21388 ( .A(n19330), .Z(n19341) );
  XOR U21389 ( .A(n19342), .B(n19343), .Z(n19330) );
  AND U21390 ( .A(n19344), .B(n19345), .Z(n19343) );
  XNOR U21391 ( .A(n19342), .B(n9673), .Z(n19345) );
  XNOR U21392 ( .A(n19338), .B(n19340), .Z(n9673) );
  NAND U21393 ( .A(n19346), .B(nreg[438]), .Z(n19340) );
  NAND U21394 ( .A(n12326), .B(nreg[438]), .Z(n19346) );
  XNOR U21395 ( .A(n19336), .B(n19347), .Z(n19338) );
  XOR U21396 ( .A(n19348), .B(n19349), .Z(n19336) );
  AND U21397 ( .A(n19350), .B(n19351), .Z(n19349) );
  XNOR U21398 ( .A(n19352), .B(n19348), .Z(n19351) );
  XOR U21399 ( .A(n19353), .B(nreg[438]), .Z(n19344) );
  IV U21400 ( .A(n19342), .Z(n19353) );
  XOR U21401 ( .A(n19354), .B(n19355), .Z(n19342) );
  AND U21402 ( .A(n19356), .B(n19357), .Z(n19355) );
  XNOR U21403 ( .A(n19354), .B(n9679), .Z(n19357) );
  XNOR U21404 ( .A(n19350), .B(n19352), .Z(n9679) );
  NAND U21405 ( .A(n19358), .B(nreg[437]), .Z(n19352) );
  NAND U21406 ( .A(n12326), .B(nreg[437]), .Z(n19358) );
  XNOR U21407 ( .A(n19348), .B(n19359), .Z(n19350) );
  XOR U21408 ( .A(n19360), .B(n19361), .Z(n19348) );
  AND U21409 ( .A(n19362), .B(n19363), .Z(n19361) );
  XNOR U21410 ( .A(n19364), .B(n19360), .Z(n19363) );
  XOR U21411 ( .A(n19365), .B(nreg[437]), .Z(n19356) );
  IV U21412 ( .A(n19354), .Z(n19365) );
  XOR U21413 ( .A(n19366), .B(n19367), .Z(n19354) );
  AND U21414 ( .A(n19368), .B(n19369), .Z(n19367) );
  XNOR U21415 ( .A(n19366), .B(n9685), .Z(n19369) );
  XNOR U21416 ( .A(n19362), .B(n19364), .Z(n9685) );
  NAND U21417 ( .A(n19370), .B(nreg[436]), .Z(n19364) );
  NAND U21418 ( .A(n12326), .B(nreg[436]), .Z(n19370) );
  XNOR U21419 ( .A(n19360), .B(n19371), .Z(n19362) );
  XOR U21420 ( .A(n19372), .B(n19373), .Z(n19360) );
  AND U21421 ( .A(n19374), .B(n19375), .Z(n19373) );
  XNOR U21422 ( .A(n19376), .B(n19372), .Z(n19375) );
  XOR U21423 ( .A(n19377), .B(nreg[436]), .Z(n19368) );
  IV U21424 ( .A(n19366), .Z(n19377) );
  XOR U21425 ( .A(n19378), .B(n19379), .Z(n19366) );
  AND U21426 ( .A(n19380), .B(n19381), .Z(n19379) );
  XNOR U21427 ( .A(n19378), .B(n9691), .Z(n19381) );
  XNOR U21428 ( .A(n19374), .B(n19376), .Z(n9691) );
  NAND U21429 ( .A(n19382), .B(nreg[435]), .Z(n19376) );
  NAND U21430 ( .A(n12326), .B(nreg[435]), .Z(n19382) );
  XNOR U21431 ( .A(n19372), .B(n19383), .Z(n19374) );
  XOR U21432 ( .A(n19384), .B(n19385), .Z(n19372) );
  AND U21433 ( .A(n19386), .B(n19387), .Z(n19385) );
  XNOR U21434 ( .A(n19388), .B(n19384), .Z(n19387) );
  XOR U21435 ( .A(n19389), .B(nreg[435]), .Z(n19380) );
  IV U21436 ( .A(n19378), .Z(n19389) );
  XOR U21437 ( .A(n19390), .B(n19391), .Z(n19378) );
  AND U21438 ( .A(n19392), .B(n19393), .Z(n19391) );
  XNOR U21439 ( .A(n19390), .B(n9697), .Z(n19393) );
  XNOR U21440 ( .A(n19386), .B(n19388), .Z(n9697) );
  NAND U21441 ( .A(n19394), .B(nreg[434]), .Z(n19388) );
  NAND U21442 ( .A(n12326), .B(nreg[434]), .Z(n19394) );
  XNOR U21443 ( .A(n19384), .B(n19395), .Z(n19386) );
  XOR U21444 ( .A(n19396), .B(n19397), .Z(n19384) );
  AND U21445 ( .A(n19398), .B(n19399), .Z(n19397) );
  XNOR U21446 ( .A(n19400), .B(n19396), .Z(n19399) );
  XOR U21447 ( .A(n19401), .B(nreg[434]), .Z(n19392) );
  IV U21448 ( .A(n19390), .Z(n19401) );
  XOR U21449 ( .A(n19402), .B(n19403), .Z(n19390) );
  AND U21450 ( .A(n19404), .B(n19405), .Z(n19403) );
  XNOR U21451 ( .A(n19402), .B(n9703), .Z(n19405) );
  XNOR U21452 ( .A(n19398), .B(n19400), .Z(n9703) );
  NAND U21453 ( .A(n19406), .B(nreg[433]), .Z(n19400) );
  NAND U21454 ( .A(n12326), .B(nreg[433]), .Z(n19406) );
  XNOR U21455 ( .A(n19396), .B(n19407), .Z(n19398) );
  XOR U21456 ( .A(n19408), .B(n19409), .Z(n19396) );
  AND U21457 ( .A(n19410), .B(n19411), .Z(n19409) );
  XNOR U21458 ( .A(n19412), .B(n19408), .Z(n19411) );
  XOR U21459 ( .A(n19413), .B(nreg[433]), .Z(n19404) );
  IV U21460 ( .A(n19402), .Z(n19413) );
  XOR U21461 ( .A(n19414), .B(n19415), .Z(n19402) );
  AND U21462 ( .A(n19416), .B(n19417), .Z(n19415) );
  XNOR U21463 ( .A(n19414), .B(n9709), .Z(n19417) );
  XNOR U21464 ( .A(n19410), .B(n19412), .Z(n9709) );
  NAND U21465 ( .A(n19418), .B(nreg[432]), .Z(n19412) );
  NAND U21466 ( .A(n12326), .B(nreg[432]), .Z(n19418) );
  XNOR U21467 ( .A(n19408), .B(n19419), .Z(n19410) );
  XOR U21468 ( .A(n19420), .B(n19421), .Z(n19408) );
  AND U21469 ( .A(n19422), .B(n19423), .Z(n19421) );
  XNOR U21470 ( .A(n19424), .B(n19420), .Z(n19423) );
  XOR U21471 ( .A(n19425), .B(nreg[432]), .Z(n19416) );
  IV U21472 ( .A(n19414), .Z(n19425) );
  XOR U21473 ( .A(n19426), .B(n19427), .Z(n19414) );
  AND U21474 ( .A(n19428), .B(n19429), .Z(n19427) );
  XNOR U21475 ( .A(n19426), .B(n9715), .Z(n19429) );
  XNOR U21476 ( .A(n19422), .B(n19424), .Z(n9715) );
  NAND U21477 ( .A(n19430), .B(nreg[431]), .Z(n19424) );
  NAND U21478 ( .A(n12326), .B(nreg[431]), .Z(n19430) );
  XNOR U21479 ( .A(n19420), .B(n19431), .Z(n19422) );
  XOR U21480 ( .A(n19432), .B(n19433), .Z(n19420) );
  AND U21481 ( .A(n19434), .B(n19435), .Z(n19433) );
  XNOR U21482 ( .A(n19436), .B(n19432), .Z(n19435) );
  XOR U21483 ( .A(n19437), .B(nreg[431]), .Z(n19428) );
  IV U21484 ( .A(n19426), .Z(n19437) );
  XOR U21485 ( .A(n19438), .B(n19439), .Z(n19426) );
  AND U21486 ( .A(n19440), .B(n19441), .Z(n19439) );
  XNOR U21487 ( .A(n19438), .B(n9721), .Z(n19441) );
  XNOR U21488 ( .A(n19434), .B(n19436), .Z(n9721) );
  NAND U21489 ( .A(n19442), .B(nreg[430]), .Z(n19436) );
  NAND U21490 ( .A(n12326), .B(nreg[430]), .Z(n19442) );
  XNOR U21491 ( .A(n19432), .B(n19443), .Z(n19434) );
  XOR U21492 ( .A(n19444), .B(n19445), .Z(n19432) );
  AND U21493 ( .A(n19446), .B(n19447), .Z(n19445) );
  XNOR U21494 ( .A(n19448), .B(n19444), .Z(n19447) );
  XOR U21495 ( .A(n19449), .B(nreg[430]), .Z(n19440) );
  IV U21496 ( .A(n19438), .Z(n19449) );
  XOR U21497 ( .A(n19450), .B(n19451), .Z(n19438) );
  AND U21498 ( .A(n19452), .B(n19453), .Z(n19451) );
  XNOR U21499 ( .A(n19450), .B(n9727), .Z(n19453) );
  XNOR U21500 ( .A(n19446), .B(n19448), .Z(n9727) );
  NAND U21501 ( .A(n19454), .B(nreg[429]), .Z(n19448) );
  NAND U21502 ( .A(n12326), .B(nreg[429]), .Z(n19454) );
  XNOR U21503 ( .A(n19444), .B(n19455), .Z(n19446) );
  XOR U21504 ( .A(n19456), .B(n19457), .Z(n19444) );
  AND U21505 ( .A(n19458), .B(n19459), .Z(n19457) );
  XNOR U21506 ( .A(n19460), .B(n19456), .Z(n19459) );
  XOR U21507 ( .A(n19461), .B(nreg[429]), .Z(n19452) );
  IV U21508 ( .A(n19450), .Z(n19461) );
  XOR U21509 ( .A(n19462), .B(n19463), .Z(n19450) );
  AND U21510 ( .A(n19464), .B(n19465), .Z(n19463) );
  XNOR U21511 ( .A(n19462), .B(n9733), .Z(n19465) );
  XNOR U21512 ( .A(n19458), .B(n19460), .Z(n9733) );
  NAND U21513 ( .A(n19466), .B(nreg[428]), .Z(n19460) );
  NAND U21514 ( .A(n12326), .B(nreg[428]), .Z(n19466) );
  XNOR U21515 ( .A(n19456), .B(n19467), .Z(n19458) );
  XOR U21516 ( .A(n19468), .B(n19469), .Z(n19456) );
  AND U21517 ( .A(n19470), .B(n19471), .Z(n19469) );
  XNOR U21518 ( .A(n19472), .B(n19468), .Z(n19471) );
  XOR U21519 ( .A(n19473), .B(nreg[428]), .Z(n19464) );
  IV U21520 ( .A(n19462), .Z(n19473) );
  XOR U21521 ( .A(n19474), .B(n19475), .Z(n19462) );
  AND U21522 ( .A(n19476), .B(n19477), .Z(n19475) );
  XNOR U21523 ( .A(n19474), .B(n9739), .Z(n19477) );
  XNOR U21524 ( .A(n19470), .B(n19472), .Z(n9739) );
  NAND U21525 ( .A(n19478), .B(nreg[427]), .Z(n19472) );
  NAND U21526 ( .A(n12326), .B(nreg[427]), .Z(n19478) );
  XNOR U21527 ( .A(n19468), .B(n19479), .Z(n19470) );
  XOR U21528 ( .A(n19480), .B(n19481), .Z(n19468) );
  AND U21529 ( .A(n19482), .B(n19483), .Z(n19481) );
  XNOR U21530 ( .A(n19484), .B(n19480), .Z(n19483) );
  XOR U21531 ( .A(n19485), .B(nreg[427]), .Z(n19476) );
  IV U21532 ( .A(n19474), .Z(n19485) );
  XOR U21533 ( .A(n19486), .B(n19487), .Z(n19474) );
  AND U21534 ( .A(n19488), .B(n19489), .Z(n19487) );
  XNOR U21535 ( .A(n19486), .B(n9745), .Z(n19489) );
  XNOR U21536 ( .A(n19482), .B(n19484), .Z(n9745) );
  NAND U21537 ( .A(n19490), .B(nreg[426]), .Z(n19484) );
  NAND U21538 ( .A(n12326), .B(nreg[426]), .Z(n19490) );
  XNOR U21539 ( .A(n19480), .B(n19491), .Z(n19482) );
  XOR U21540 ( .A(n19492), .B(n19493), .Z(n19480) );
  AND U21541 ( .A(n19494), .B(n19495), .Z(n19493) );
  XNOR U21542 ( .A(n19496), .B(n19492), .Z(n19495) );
  XOR U21543 ( .A(n19497), .B(nreg[426]), .Z(n19488) );
  IV U21544 ( .A(n19486), .Z(n19497) );
  XOR U21545 ( .A(n19498), .B(n19499), .Z(n19486) );
  AND U21546 ( .A(n19500), .B(n19501), .Z(n19499) );
  XNOR U21547 ( .A(n19498), .B(n9751), .Z(n19501) );
  XNOR U21548 ( .A(n19494), .B(n19496), .Z(n9751) );
  NAND U21549 ( .A(n19502), .B(nreg[425]), .Z(n19496) );
  NAND U21550 ( .A(n12326), .B(nreg[425]), .Z(n19502) );
  XNOR U21551 ( .A(n19492), .B(n19503), .Z(n19494) );
  XOR U21552 ( .A(n19504), .B(n19505), .Z(n19492) );
  AND U21553 ( .A(n19506), .B(n19507), .Z(n19505) );
  XNOR U21554 ( .A(n19508), .B(n19504), .Z(n19507) );
  XOR U21555 ( .A(n19509), .B(nreg[425]), .Z(n19500) );
  IV U21556 ( .A(n19498), .Z(n19509) );
  XOR U21557 ( .A(n19510), .B(n19511), .Z(n19498) );
  AND U21558 ( .A(n19512), .B(n19513), .Z(n19511) );
  XNOR U21559 ( .A(n19510), .B(n9757), .Z(n19513) );
  XNOR U21560 ( .A(n19506), .B(n19508), .Z(n9757) );
  NAND U21561 ( .A(n19514), .B(nreg[424]), .Z(n19508) );
  NAND U21562 ( .A(n12326), .B(nreg[424]), .Z(n19514) );
  XNOR U21563 ( .A(n19504), .B(n19515), .Z(n19506) );
  XOR U21564 ( .A(n19516), .B(n19517), .Z(n19504) );
  AND U21565 ( .A(n19518), .B(n19519), .Z(n19517) );
  XNOR U21566 ( .A(n19520), .B(n19516), .Z(n19519) );
  XOR U21567 ( .A(n19521), .B(nreg[424]), .Z(n19512) );
  IV U21568 ( .A(n19510), .Z(n19521) );
  XOR U21569 ( .A(n19522), .B(n19523), .Z(n19510) );
  AND U21570 ( .A(n19524), .B(n19525), .Z(n19523) );
  XNOR U21571 ( .A(n19522), .B(n9763), .Z(n19525) );
  XNOR U21572 ( .A(n19518), .B(n19520), .Z(n9763) );
  NAND U21573 ( .A(n19526), .B(nreg[423]), .Z(n19520) );
  NAND U21574 ( .A(n12326), .B(nreg[423]), .Z(n19526) );
  XNOR U21575 ( .A(n19516), .B(n19527), .Z(n19518) );
  XOR U21576 ( .A(n19528), .B(n19529), .Z(n19516) );
  AND U21577 ( .A(n19530), .B(n19531), .Z(n19529) );
  XNOR U21578 ( .A(n19532), .B(n19528), .Z(n19531) );
  XOR U21579 ( .A(n19533), .B(nreg[423]), .Z(n19524) );
  IV U21580 ( .A(n19522), .Z(n19533) );
  XOR U21581 ( .A(n19534), .B(n19535), .Z(n19522) );
  AND U21582 ( .A(n19536), .B(n19537), .Z(n19535) );
  XNOR U21583 ( .A(n19534), .B(n9769), .Z(n19537) );
  XNOR U21584 ( .A(n19530), .B(n19532), .Z(n9769) );
  NAND U21585 ( .A(n19538), .B(nreg[422]), .Z(n19532) );
  NAND U21586 ( .A(n12326), .B(nreg[422]), .Z(n19538) );
  XNOR U21587 ( .A(n19528), .B(n19539), .Z(n19530) );
  XOR U21588 ( .A(n19540), .B(n19541), .Z(n19528) );
  AND U21589 ( .A(n19542), .B(n19543), .Z(n19541) );
  XNOR U21590 ( .A(n19544), .B(n19540), .Z(n19543) );
  XOR U21591 ( .A(n19545), .B(nreg[422]), .Z(n19536) );
  IV U21592 ( .A(n19534), .Z(n19545) );
  XOR U21593 ( .A(n19546), .B(n19547), .Z(n19534) );
  AND U21594 ( .A(n19548), .B(n19549), .Z(n19547) );
  XNOR U21595 ( .A(n19546), .B(n9775), .Z(n19549) );
  XNOR U21596 ( .A(n19542), .B(n19544), .Z(n9775) );
  NAND U21597 ( .A(n19550), .B(nreg[421]), .Z(n19544) );
  NAND U21598 ( .A(n12326), .B(nreg[421]), .Z(n19550) );
  XNOR U21599 ( .A(n19540), .B(n19551), .Z(n19542) );
  XOR U21600 ( .A(n19552), .B(n19553), .Z(n19540) );
  AND U21601 ( .A(n19554), .B(n19555), .Z(n19553) );
  XNOR U21602 ( .A(n19556), .B(n19552), .Z(n19555) );
  XOR U21603 ( .A(n19557), .B(nreg[421]), .Z(n19548) );
  IV U21604 ( .A(n19546), .Z(n19557) );
  XOR U21605 ( .A(n19558), .B(n19559), .Z(n19546) );
  AND U21606 ( .A(n19560), .B(n19561), .Z(n19559) );
  XNOR U21607 ( .A(n19558), .B(n9781), .Z(n19561) );
  XNOR U21608 ( .A(n19554), .B(n19556), .Z(n9781) );
  NAND U21609 ( .A(n19562), .B(nreg[420]), .Z(n19556) );
  NAND U21610 ( .A(n12326), .B(nreg[420]), .Z(n19562) );
  XNOR U21611 ( .A(n19552), .B(n19563), .Z(n19554) );
  XOR U21612 ( .A(n19564), .B(n19565), .Z(n19552) );
  AND U21613 ( .A(n19566), .B(n19567), .Z(n19565) );
  XNOR U21614 ( .A(n19568), .B(n19564), .Z(n19567) );
  XOR U21615 ( .A(n19569), .B(nreg[420]), .Z(n19560) );
  IV U21616 ( .A(n19558), .Z(n19569) );
  XOR U21617 ( .A(n19570), .B(n19571), .Z(n19558) );
  AND U21618 ( .A(n19572), .B(n19573), .Z(n19571) );
  XNOR U21619 ( .A(n19570), .B(n9787), .Z(n19573) );
  XNOR U21620 ( .A(n19566), .B(n19568), .Z(n9787) );
  NAND U21621 ( .A(n19574), .B(nreg[419]), .Z(n19568) );
  NAND U21622 ( .A(n12326), .B(nreg[419]), .Z(n19574) );
  XNOR U21623 ( .A(n19564), .B(n19575), .Z(n19566) );
  XOR U21624 ( .A(n19576), .B(n19577), .Z(n19564) );
  AND U21625 ( .A(n19578), .B(n19579), .Z(n19577) );
  XNOR U21626 ( .A(n19580), .B(n19576), .Z(n19579) );
  XOR U21627 ( .A(n19581), .B(nreg[419]), .Z(n19572) );
  IV U21628 ( .A(n19570), .Z(n19581) );
  XOR U21629 ( .A(n19582), .B(n19583), .Z(n19570) );
  AND U21630 ( .A(n19584), .B(n19585), .Z(n19583) );
  XNOR U21631 ( .A(n19582), .B(n9793), .Z(n19585) );
  XNOR U21632 ( .A(n19578), .B(n19580), .Z(n9793) );
  NAND U21633 ( .A(n19586), .B(nreg[418]), .Z(n19580) );
  NAND U21634 ( .A(n12326), .B(nreg[418]), .Z(n19586) );
  XNOR U21635 ( .A(n19576), .B(n19587), .Z(n19578) );
  XOR U21636 ( .A(n19588), .B(n19589), .Z(n19576) );
  AND U21637 ( .A(n19590), .B(n19591), .Z(n19589) );
  XNOR U21638 ( .A(n19592), .B(n19588), .Z(n19591) );
  XOR U21639 ( .A(n19593), .B(nreg[418]), .Z(n19584) );
  IV U21640 ( .A(n19582), .Z(n19593) );
  XOR U21641 ( .A(n19594), .B(n19595), .Z(n19582) );
  AND U21642 ( .A(n19596), .B(n19597), .Z(n19595) );
  XNOR U21643 ( .A(n19594), .B(n9799), .Z(n19597) );
  XNOR U21644 ( .A(n19590), .B(n19592), .Z(n9799) );
  NAND U21645 ( .A(n19598), .B(nreg[417]), .Z(n19592) );
  NAND U21646 ( .A(n12326), .B(nreg[417]), .Z(n19598) );
  XNOR U21647 ( .A(n19588), .B(n19599), .Z(n19590) );
  XOR U21648 ( .A(n19600), .B(n19601), .Z(n19588) );
  AND U21649 ( .A(n19602), .B(n19603), .Z(n19601) );
  XNOR U21650 ( .A(n19604), .B(n19600), .Z(n19603) );
  XOR U21651 ( .A(n19605), .B(nreg[417]), .Z(n19596) );
  IV U21652 ( .A(n19594), .Z(n19605) );
  XOR U21653 ( .A(n19606), .B(n19607), .Z(n19594) );
  AND U21654 ( .A(n19608), .B(n19609), .Z(n19607) );
  XNOR U21655 ( .A(n19606), .B(n9805), .Z(n19609) );
  XNOR U21656 ( .A(n19602), .B(n19604), .Z(n9805) );
  NAND U21657 ( .A(n19610), .B(nreg[416]), .Z(n19604) );
  NAND U21658 ( .A(n12326), .B(nreg[416]), .Z(n19610) );
  XNOR U21659 ( .A(n19600), .B(n19611), .Z(n19602) );
  XOR U21660 ( .A(n19612), .B(n19613), .Z(n19600) );
  AND U21661 ( .A(n19614), .B(n19615), .Z(n19613) );
  XNOR U21662 ( .A(n19616), .B(n19612), .Z(n19615) );
  XOR U21663 ( .A(n19617), .B(nreg[416]), .Z(n19608) );
  IV U21664 ( .A(n19606), .Z(n19617) );
  XOR U21665 ( .A(n19618), .B(n19619), .Z(n19606) );
  AND U21666 ( .A(n19620), .B(n19621), .Z(n19619) );
  XNOR U21667 ( .A(n19618), .B(n9811), .Z(n19621) );
  XNOR U21668 ( .A(n19614), .B(n19616), .Z(n9811) );
  NAND U21669 ( .A(n19622), .B(nreg[415]), .Z(n19616) );
  NAND U21670 ( .A(n12326), .B(nreg[415]), .Z(n19622) );
  XNOR U21671 ( .A(n19612), .B(n19623), .Z(n19614) );
  XOR U21672 ( .A(n19624), .B(n19625), .Z(n19612) );
  AND U21673 ( .A(n19626), .B(n19627), .Z(n19625) );
  XNOR U21674 ( .A(n19628), .B(n19624), .Z(n19627) );
  XOR U21675 ( .A(n19629), .B(nreg[415]), .Z(n19620) );
  IV U21676 ( .A(n19618), .Z(n19629) );
  XOR U21677 ( .A(n19630), .B(n19631), .Z(n19618) );
  AND U21678 ( .A(n19632), .B(n19633), .Z(n19631) );
  XNOR U21679 ( .A(n19630), .B(n9817), .Z(n19633) );
  XNOR U21680 ( .A(n19626), .B(n19628), .Z(n9817) );
  NAND U21681 ( .A(n19634), .B(nreg[414]), .Z(n19628) );
  NAND U21682 ( .A(n12326), .B(nreg[414]), .Z(n19634) );
  XNOR U21683 ( .A(n19624), .B(n19635), .Z(n19626) );
  XOR U21684 ( .A(n19636), .B(n19637), .Z(n19624) );
  AND U21685 ( .A(n19638), .B(n19639), .Z(n19637) );
  XNOR U21686 ( .A(n19640), .B(n19636), .Z(n19639) );
  XOR U21687 ( .A(n19641), .B(nreg[414]), .Z(n19632) );
  IV U21688 ( .A(n19630), .Z(n19641) );
  XOR U21689 ( .A(n19642), .B(n19643), .Z(n19630) );
  AND U21690 ( .A(n19644), .B(n19645), .Z(n19643) );
  XNOR U21691 ( .A(n19642), .B(n9823), .Z(n19645) );
  XNOR U21692 ( .A(n19638), .B(n19640), .Z(n9823) );
  NAND U21693 ( .A(n19646), .B(nreg[413]), .Z(n19640) );
  NAND U21694 ( .A(n12326), .B(nreg[413]), .Z(n19646) );
  XNOR U21695 ( .A(n19636), .B(n19647), .Z(n19638) );
  XOR U21696 ( .A(n19648), .B(n19649), .Z(n19636) );
  AND U21697 ( .A(n19650), .B(n19651), .Z(n19649) );
  XNOR U21698 ( .A(n19652), .B(n19648), .Z(n19651) );
  XOR U21699 ( .A(n19653), .B(nreg[413]), .Z(n19644) );
  IV U21700 ( .A(n19642), .Z(n19653) );
  XOR U21701 ( .A(n19654), .B(n19655), .Z(n19642) );
  AND U21702 ( .A(n19656), .B(n19657), .Z(n19655) );
  XNOR U21703 ( .A(n19654), .B(n9829), .Z(n19657) );
  XNOR U21704 ( .A(n19650), .B(n19652), .Z(n9829) );
  NAND U21705 ( .A(n19658), .B(nreg[412]), .Z(n19652) );
  NAND U21706 ( .A(n12326), .B(nreg[412]), .Z(n19658) );
  XNOR U21707 ( .A(n19648), .B(n19659), .Z(n19650) );
  XOR U21708 ( .A(n19660), .B(n19661), .Z(n19648) );
  AND U21709 ( .A(n19662), .B(n19663), .Z(n19661) );
  XNOR U21710 ( .A(n19664), .B(n19660), .Z(n19663) );
  XOR U21711 ( .A(n19665), .B(nreg[412]), .Z(n19656) );
  IV U21712 ( .A(n19654), .Z(n19665) );
  XOR U21713 ( .A(n19666), .B(n19667), .Z(n19654) );
  AND U21714 ( .A(n19668), .B(n19669), .Z(n19667) );
  XNOR U21715 ( .A(n19666), .B(n9835), .Z(n19669) );
  XNOR U21716 ( .A(n19662), .B(n19664), .Z(n9835) );
  NAND U21717 ( .A(n19670), .B(nreg[411]), .Z(n19664) );
  NAND U21718 ( .A(n12326), .B(nreg[411]), .Z(n19670) );
  XNOR U21719 ( .A(n19660), .B(n19671), .Z(n19662) );
  XOR U21720 ( .A(n19672), .B(n19673), .Z(n19660) );
  AND U21721 ( .A(n19674), .B(n19675), .Z(n19673) );
  XNOR U21722 ( .A(n19676), .B(n19672), .Z(n19675) );
  XOR U21723 ( .A(n19677), .B(nreg[411]), .Z(n19668) );
  IV U21724 ( .A(n19666), .Z(n19677) );
  XOR U21725 ( .A(n19678), .B(n19679), .Z(n19666) );
  AND U21726 ( .A(n19680), .B(n19681), .Z(n19679) );
  XNOR U21727 ( .A(n19678), .B(n9841), .Z(n19681) );
  XNOR U21728 ( .A(n19674), .B(n19676), .Z(n9841) );
  NAND U21729 ( .A(n19682), .B(nreg[410]), .Z(n19676) );
  NAND U21730 ( .A(n12326), .B(nreg[410]), .Z(n19682) );
  XNOR U21731 ( .A(n19672), .B(n19683), .Z(n19674) );
  XOR U21732 ( .A(n19684), .B(n19685), .Z(n19672) );
  AND U21733 ( .A(n19686), .B(n19687), .Z(n19685) );
  XNOR U21734 ( .A(n19688), .B(n19684), .Z(n19687) );
  XOR U21735 ( .A(n19689), .B(nreg[410]), .Z(n19680) );
  IV U21736 ( .A(n19678), .Z(n19689) );
  XOR U21737 ( .A(n19690), .B(n19691), .Z(n19678) );
  AND U21738 ( .A(n19692), .B(n19693), .Z(n19691) );
  XNOR U21739 ( .A(n19690), .B(n9847), .Z(n19693) );
  XNOR U21740 ( .A(n19686), .B(n19688), .Z(n9847) );
  NAND U21741 ( .A(n19694), .B(nreg[409]), .Z(n19688) );
  NAND U21742 ( .A(n12326), .B(nreg[409]), .Z(n19694) );
  XNOR U21743 ( .A(n19684), .B(n19695), .Z(n19686) );
  XOR U21744 ( .A(n19696), .B(n19697), .Z(n19684) );
  AND U21745 ( .A(n19698), .B(n19699), .Z(n19697) );
  XNOR U21746 ( .A(n19700), .B(n19696), .Z(n19699) );
  XOR U21747 ( .A(n19701), .B(nreg[409]), .Z(n19692) );
  IV U21748 ( .A(n19690), .Z(n19701) );
  XOR U21749 ( .A(n19702), .B(n19703), .Z(n19690) );
  AND U21750 ( .A(n19704), .B(n19705), .Z(n19703) );
  XNOR U21751 ( .A(n19702), .B(n9853), .Z(n19705) );
  XNOR U21752 ( .A(n19698), .B(n19700), .Z(n9853) );
  NAND U21753 ( .A(n19706), .B(nreg[408]), .Z(n19700) );
  NAND U21754 ( .A(n12326), .B(nreg[408]), .Z(n19706) );
  XNOR U21755 ( .A(n19696), .B(n19707), .Z(n19698) );
  XOR U21756 ( .A(n19708), .B(n19709), .Z(n19696) );
  AND U21757 ( .A(n19710), .B(n19711), .Z(n19709) );
  XNOR U21758 ( .A(n19712), .B(n19708), .Z(n19711) );
  XOR U21759 ( .A(n19713), .B(nreg[408]), .Z(n19704) );
  IV U21760 ( .A(n19702), .Z(n19713) );
  XOR U21761 ( .A(n19714), .B(n19715), .Z(n19702) );
  AND U21762 ( .A(n19716), .B(n19717), .Z(n19715) );
  XNOR U21763 ( .A(n19714), .B(n9859), .Z(n19717) );
  XNOR U21764 ( .A(n19710), .B(n19712), .Z(n9859) );
  NAND U21765 ( .A(n19718), .B(nreg[407]), .Z(n19712) );
  NAND U21766 ( .A(n12326), .B(nreg[407]), .Z(n19718) );
  XNOR U21767 ( .A(n19708), .B(n19719), .Z(n19710) );
  XOR U21768 ( .A(n19720), .B(n19721), .Z(n19708) );
  AND U21769 ( .A(n19722), .B(n19723), .Z(n19721) );
  XNOR U21770 ( .A(n19724), .B(n19720), .Z(n19723) );
  XOR U21771 ( .A(n19725), .B(nreg[407]), .Z(n19716) );
  IV U21772 ( .A(n19714), .Z(n19725) );
  XOR U21773 ( .A(n19726), .B(n19727), .Z(n19714) );
  AND U21774 ( .A(n19728), .B(n19729), .Z(n19727) );
  XNOR U21775 ( .A(n19726), .B(n9865), .Z(n19729) );
  XNOR U21776 ( .A(n19722), .B(n19724), .Z(n9865) );
  NAND U21777 ( .A(n19730), .B(nreg[406]), .Z(n19724) );
  NAND U21778 ( .A(n12326), .B(nreg[406]), .Z(n19730) );
  XNOR U21779 ( .A(n19720), .B(n19731), .Z(n19722) );
  XOR U21780 ( .A(n19732), .B(n19733), .Z(n19720) );
  AND U21781 ( .A(n19734), .B(n19735), .Z(n19733) );
  XNOR U21782 ( .A(n19736), .B(n19732), .Z(n19735) );
  XOR U21783 ( .A(n19737), .B(nreg[406]), .Z(n19728) );
  IV U21784 ( .A(n19726), .Z(n19737) );
  XOR U21785 ( .A(n19738), .B(n19739), .Z(n19726) );
  AND U21786 ( .A(n19740), .B(n19741), .Z(n19739) );
  XNOR U21787 ( .A(n19738), .B(n9871), .Z(n19741) );
  XNOR U21788 ( .A(n19734), .B(n19736), .Z(n9871) );
  NAND U21789 ( .A(n19742), .B(nreg[405]), .Z(n19736) );
  NAND U21790 ( .A(n12326), .B(nreg[405]), .Z(n19742) );
  XNOR U21791 ( .A(n19732), .B(n19743), .Z(n19734) );
  XOR U21792 ( .A(n19744), .B(n19745), .Z(n19732) );
  AND U21793 ( .A(n19746), .B(n19747), .Z(n19745) );
  XNOR U21794 ( .A(n19748), .B(n19744), .Z(n19747) );
  XOR U21795 ( .A(n19749), .B(nreg[405]), .Z(n19740) );
  IV U21796 ( .A(n19738), .Z(n19749) );
  XOR U21797 ( .A(n19750), .B(n19751), .Z(n19738) );
  AND U21798 ( .A(n19752), .B(n19753), .Z(n19751) );
  XNOR U21799 ( .A(n19750), .B(n9877), .Z(n19753) );
  XNOR U21800 ( .A(n19746), .B(n19748), .Z(n9877) );
  NAND U21801 ( .A(n19754), .B(nreg[404]), .Z(n19748) );
  NAND U21802 ( .A(n12326), .B(nreg[404]), .Z(n19754) );
  XNOR U21803 ( .A(n19744), .B(n19755), .Z(n19746) );
  XOR U21804 ( .A(n19756), .B(n19757), .Z(n19744) );
  AND U21805 ( .A(n19758), .B(n19759), .Z(n19757) );
  XNOR U21806 ( .A(n19760), .B(n19756), .Z(n19759) );
  XOR U21807 ( .A(n19761), .B(nreg[404]), .Z(n19752) );
  IV U21808 ( .A(n19750), .Z(n19761) );
  XOR U21809 ( .A(n19762), .B(n19763), .Z(n19750) );
  AND U21810 ( .A(n19764), .B(n19765), .Z(n19763) );
  XNOR U21811 ( .A(n19762), .B(n9883), .Z(n19765) );
  XNOR U21812 ( .A(n19758), .B(n19760), .Z(n9883) );
  NAND U21813 ( .A(n19766), .B(nreg[403]), .Z(n19760) );
  NAND U21814 ( .A(n12326), .B(nreg[403]), .Z(n19766) );
  XNOR U21815 ( .A(n19756), .B(n19767), .Z(n19758) );
  XOR U21816 ( .A(n19768), .B(n19769), .Z(n19756) );
  AND U21817 ( .A(n19770), .B(n19771), .Z(n19769) );
  XNOR U21818 ( .A(n19772), .B(n19768), .Z(n19771) );
  XOR U21819 ( .A(n19773), .B(nreg[403]), .Z(n19764) );
  IV U21820 ( .A(n19762), .Z(n19773) );
  XOR U21821 ( .A(n19774), .B(n19775), .Z(n19762) );
  AND U21822 ( .A(n19776), .B(n19777), .Z(n19775) );
  XNOR U21823 ( .A(n19774), .B(n9889), .Z(n19777) );
  XNOR U21824 ( .A(n19770), .B(n19772), .Z(n9889) );
  NAND U21825 ( .A(n19778), .B(nreg[402]), .Z(n19772) );
  NAND U21826 ( .A(n12326), .B(nreg[402]), .Z(n19778) );
  XNOR U21827 ( .A(n19768), .B(n19779), .Z(n19770) );
  XOR U21828 ( .A(n19780), .B(n19781), .Z(n19768) );
  AND U21829 ( .A(n19782), .B(n19783), .Z(n19781) );
  XNOR U21830 ( .A(n19784), .B(n19780), .Z(n19783) );
  XOR U21831 ( .A(n19785), .B(nreg[402]), .Z(n19776) );
  IV U21832 ( .A(n19774), .Z(n19785) );
  XOR U21833 ( .A(n19786), .B(n19787), .Z(n19774) );
  AND U21834 ( .A(n19788), .B(n19789), .Z(n19787) );
  XNOR U21835 ( .A(n19786), .B(n9895), .Z(n19789) );
  XNOR U21836 ( .A(n19782), .B(n19784), .Z(n9895) );
  NAND U21837 ( .A(n19790), .B(nreg[401]), .Z(n19784) );
  NAND U21838 ( .A(n12326), .B(nreg[401]), .Z(n19790) );
  XNOR U21839 ( .A(n19780), .B(n19791), .Z(n19782) );
  XOR U21840 ( .A(n19792), .B(n19793), .Z(n19780) );
  AND U21841 ( .A(n19794), .B(n19795), .Z(n19793) );
  XNOR U21842 ( .A(n19796), .B(n19792), .Z(n19795) );
  XOR U21843 ( .A(n19797), .B(nreg[401]), .Z(n19788) );
  IV U21844 ( .A(n19786), .Z(n19797) );
  XOR U21845 ( .A(n19798), .B(n19799), .Z(n19786) );
  AND U21846 ( .A(n19800), .B(n19801), .Z(n19799) );
  XNOR U21847 ( .A(n19798), .B(n9901), .Z(n19801) );
  XNOR U21848 ( .A(n19794), .B(n19796), .Z(n9901) );
  NAND U21849 ( .A(n19802), .B(nreg[400]), .Z(n19796) );
  NAND U21850 ( .A(n12326), .B(nreg[400]), .Z(n19802) );
  XNOR U21851 ( .A(n19792), .B(n19803), .Z(n19794) );
  XOR U21852 ( .A(n19804), .B(n19805), .Z(n19792) );
  AND U21853 ( .A(n19806), .B(n19807), .Z(n19805) );
  XNOR U21854 ( .A(n19808), .B(n19804), .Z(n19807) );
  XOR U21855 ( .A(n19809), .B(nreg[400]), .Z(n19800) );
  IV U21856 ( .A(n19798), .Z(n19809) );
  XOR U21857 ( .A(n19810), .B(n19811), .Z(n19798) );
  AND U21858 ( .A(n19812), .B(n19813), .Z(n19811) );
  XNOR U21859 ( .A(n19810), .B(n9907), .Z(n19813) );
  XNOR U21860 ( .A(n19806), .B(n19808), .Z(n9907) );
  NAND U21861 ( .A(n19814), .B(nreg[399]), .Z(n19808) );
  NAND U21862 ( .A(n12326), .B(nreg[399]), .Z(n19814) );
  XNOR U21863 ( .A(n19804), .B(n19815), .Z(n19806) );
  XOR U21864 ( .A(n19816), .B(n19817), .Z(n19804) );
  AND U21865 ( .A(n19818), .B(n19819), .Z(n19817) );
  XNOR U21866 ( .A(n19820), .B(n19816), .Z(n19819) );
  XOR U21867 ( .A(n19821), .B(nreg[399]), .Z(n19812) );
  IV U21868 ( .A(n19810), .Z(n19821) );
  XOR U21869 ( .A(n19822), .B(n19823), .Z(n19810) );
  AND U21870 ( .A(n19824), .B(n19825), .Z(n19823) );
  XNOR U21871 ( .A(n19822), .B(n9913), .Z(n19825) );
  XNOR U21872 ( .A(n19818), .B(n19820), .Z(n9913) );
  NAND U21873 ( .A(n19826), .B(nreg[398]), .Z(n19820) );
  NAND U21874 ( .A(n12326), .B(nreg[398]), .Z(n19826) );
  XNOR U21875 ( .A(n19816), .B(n19827), .Z(n19818) );
  XOR U21876 ( .A(n19828), .B(n19829), .Z(n19816) );
  AND U21877 ( .A(n19830), .B(n19831), .Z(n19829) );
  XNOR U21878 ( .A(n19832), .B(n19828), .Z(n19831) );
  XOR U21879 ( .A(n19833), .B(nreg[398]), .Z(n19824) );
  IV U21880 ( .A(n19822), .Z(n19833) );
  XOR U21881 ( .A(n19834), .B(n19835), .Z(n19822) );
  AND U21882 ( .A(n19836), .B(n19837), .Z(n19835) );
  XNOR U21883 ( .A(n19834), .B(n9919), .Z(n19837) );
  XNOR U21884 ( .A(n19830), .B(n19832), .Z(n9919) );
  NAND U21885 ( .A(n19838), .B(nreg[397]), .Z(n19832) );
  NAND U21886 ( .A(n12326), .B(nreg[397]), .Z(n19838) );
  XNOR U21887 ( .A(n19828), .B(n19839), .Z(n19830) );
  XOR U21888 ( .A(n19840), .B(n19841), .Z(n19828) );
  AND U21889 ( .A(n19842), .B(n19843), .Z(n19841) );
  XNOR U21890 ( .A(n19844), .B(n19840), .Z(n19843) );
  XOR U21891 ( .A(n19845), .B(nreg[397]), .Z(n19836) );
  IV U21892 ( .A(n19834), .Z(n19845) );
  XOR U21893 ( .A(n19846), .B(n19847), .Z(n19834) );
  AND U21894 ( .A(n19848), .B(n19849), .Z(n19847) );
  XNOR U21895 ( .A(n19846), .B(n9925), .Z(n19849) );
  XNOR U21896 ( .A(n19842), .B(n19844), .Z(n9925) );
  NAND U21897 ( .A(n19850), .B(nreg[396]), .Z(n19844) );
  NAND U21898 ( .A(n12326), .B(nreg[396]), .Z(n19850) );
  XNOR U21899 ( .A(n19840), .B(n19851), .Z(n19842) );
  XOR U21900 ( .A(n19852), .B(n19853), .Z(n19840) );
  AND U21901 ( .A(n19854), .B(n19855), .Z(n19853) );
  XNOR U21902 ( .A(n19856), .B(n19852), .Z(n19855) );
  XOR U21903 ( .A(n19857), .B(nreg[396]), .Z(n19848) );
  IV U21904 ( .A(n19846), .Z(n19857) );
  XOR U21905 ( .A(n19858), .B(n19859), .Z(n19846) );
  AND U21906 ( .A(n19860), .B(n19861), .Z(n19859) );
  XNOR U21907 ( .A(n19858), .B(n9931), .Z(n19861) );
  XNOR U21908 ( .A(n19854), .B(n19856), .Z(n9931) );
  NAND U21909 ( .A(n19862), .B(nreg[395]), .Z(n19856) );
  NAND U21910 ( .A(n12326), .B(nreg[395]), .Z(n19862) );
  XNOR U21911 ( .A(n19852), .B(n19863), .Z(n19854) );
  XOR U21912 ( .A(n19864), .B(n19865), .Z(n19852) );
  AND U21913 ( .A(n19866), .B(n19867), .Z(n19865) );
  XNOR U21914 ( .A(n19868), .B(n19864), .Z(n19867) );
  XOR U21915 ( .A(n19869), .B(nreg[395]), .Z(n19860) );
  IV U21916 ( .A(n19858), .Z(n19869) );
  XOR U21917 ( .A(n19870), .B(n19871), .Z(n19858) );
  AND U21918 ( .A(n19872), .B(n19873), .Z(n19871) );
  XNOR U21919 ( .A(n19870), .B(n9937), .Z(n19873) );
  XNOR U21920 ( .A(n19866), .B(n19868), .Z(n9937) );
  NAND U21921 ( .A(n19874), .B(nreg[394]), .Z(n19868) );
  NAND U21922 ( .A(n12326), .B(nreg[394]), .Z(n19874) );
  XNOR U21923 ( .A(n19864), .B(n19875), .Z(n19866) );
  XOR U21924 ( .A(n19876), .B(n19877), .Z(n19864) );
  AND U21925 ( .A(n19878), .B(n19879), .Z(n19877) );
  XNOR U21926 ( .A(n19880), .B(n19876), .Z(n19879) );
  XOR U21927 ( .A(n19881), .B(nreg[394]), .Z(n19872) );
  IV U21928 ( .A(n19870), .Z(n19881) );
  XOR U21929 ( .A(n19882), .B(n19883), .Z(n19870) );
  AND U21930 ( .A(n19884), .B(n19885), .Z(n19883) );
  XNOR U21931 ( .A(n19882), .B(n9943), .Z(n19885) );
  XNOR U21932 ( .A(n19878), .B(n19880), .Z(n9943) );
  NAND U21933 ( .A(n19886), .B(nreg[393]), .Z(n19880) );
  NAND U21934 ( .A(n12326), .B(nreg[393]), .Z(n19886) );
  XNOR U21935 ( .A(n19876), .B(n19887), .Z(n19878) );
  XOR U21936 ( .A(n19888), .B(n19889), .Z(n19876) );
  AND U21937 ( .A(n19890), .B(n19891), .Z(n19889) );
  XNOR U21938 ( .A(n19892), .B(n19888), .Z(n19891) );
  XOR U21939 ( .A(n19893), .B(nreg[393]), .Z(n19884) );
  IV U21940 ( .A(n19882), .Z(n19893) );
  XOR U21941 ( .A(n19894), .B(n19895), .Z(n19882) );
  AND U21942 ( .A(n19896), .B(n19897), .Z(n19895) );
  XNOR U21943 ( .A(n19894), .B(n9949), .Z(n19897) );
  XNOR U21944 ( .A(n19890), .B(n19892), .Z(n9949) );
  NAND U21945 ( .A(n19898), .B(nreg[392]), .Z(n19892) );
  NAND U21946 ( .A(n12326), .B(nreg[392]), .Z(n19898) );
  XNOR U21947 ( .A(n19888), .B(n19899), .Z(n19890) );
  XOR U21948 ( .A(n19900), .B(n19901), .Z(n19888) );
  AND U21949 ( .A(n19902), .B(n19903), .Z(n19901) );
  XNOR U21950 ( .A(n19904), .B(n19900), .Z(n19903) );
  XOR U21951 ( .A(n19905), .B(nreg[392]), .Z(n19896) );
  IV U21952 ( .A(n19894), .Z(n19905) );
  XOR U21953 ( .A(n19906), .B(n19907), .Z(n19894) );
  AND U21954 ( .A(n19908), .B(n19909), .Z(n19907) );
  XNOR U21955 ( .A(n19906), .B(n9955), .Z(n19909) );
  XNOR U21956 ( .A(n19902), .B(n19904), .Z(n9955) );
  NAND U21957 ( .A(n19910), .B(nreg[391]), .Z(n19904) );
  NAND U21958 ( .A(n12326), .B(nreg[391]), .Z(n19910) );
  XNOR U21959 ( .A(n19900), .B(n19911), .Z(n19902) );
  XOR U21960 ( .A(n19912), .B(n19913), .Z(n19900) );
  AND U21961 ( .A(n19914), .B(n19915), .Z(n19913) );
  XNOR U21962 ( .A(n19916), .B(n19912), .Z(n19915) );
  XOR U21963 ( .A(n19917), .B(nreg[391]), .Z(n19908) );
  IV U21964 ( .A(n19906), .Z(n19917) );
  XOR U21965 ( .A(n19918), .B(n19919), .Z(n19906) );
  AND U21966 ( .A(n19920), .B(n19921), .Z(n19919) );
  XNOR U21967 ( .A(n19918), .B(n9961), .Z(n19921) );
  XNOR U21968 ( .A(n19914), .B(n19916), .Z(n9961) );
  NAND U21969 ( .A(n19922), .B(nreg[390]), .Z(n19916) );
  NAND U21970 ( .A(n12326), .B(nreg[390]), .Z(n19922) );
  XNOR U21971 ( .A(n19912), .B(n19923), .Z(n19914) );
  XOR U21972 ( .A(n19924), .B(n19925), .Z(n19912) );
  AND U21973 ( .A(n19926), .B(n19927), .Z(n19925) );
  XNOR U21974 ( .A(n19928), .B(n19924), .Z(n19927) );
  XOR U21975 ( .A(n19929), .B(nreg[390]), .Z(n19920) );
  IV U21976 ( .A(n19918), .Z(n19929) );
  XOR U21977 ( .A(n19930), .B(n19931), .Z(n19918) );
  AND U21978 ( .A(n19932), .B(n19933), .Z(n19931) );
  XNOR U21979 ( .A(n19930), .B(n9967), .Z(n19933) );
  XNOR U21980 ( .A(n19926), .B(n19928), .Z(n9967) );
  NAND U21981 ( .A(n19934), .B(nreg[389]), .Z(n19928) );
  NAND U21982 ( .A(n12326), .B(nreg[389]), .Z(n19934) );
  XNOR U21983 ( .A(n19924), .B(n19935), .Z(n19926) );
  XOR U21984 ( .A(n19936), .B(n19937), .Z(n19924) );
  AND U21985 ( .A(n19938), .B(n19939), .Z(n19937) );
  XNOR U21986 ( .A(n19940), .B(n19936), .Z(n19939) );
  XOR U21987 ( .A(n19941), .B(nreg[389]), .Z(n19932) );
  IV U21988 ( .A(n19930), .Z(n19941) );
  XOR U21989 ( .A(n19942), .B(n19943), .Z(n19930) );
  AND U21990 ( .A(n19944), .B(n19945), .Z(n19943) );
  XNOR U21991 ( .A(n19942), .B(n9973), .Z(n19945) );
  XNOR U21992 ( .A(n19938), .B(n19940), .Z(n9973) );
  NAND U21993 ( .A(n19946), .B(nreg[388]), .Z(n19940) );
  NAND U21994 ( .A(n12326), .B(nreg[388]), .Z(n19946) );
  XNOR U21995 ( .A(n19936), .B(n19947), .Z(n19938) );
  XOR U21996 ( .A(n19948), .B(n19949), .Z(n19936) );
  AND U21997 ( .A(n19950), .B(n19951), .Z(n19949) );
  XNOR U21998 ( .A(n19952), .B(n19948), .Z(n19951) );
  XOR U21999 ( .A(n19953), .B(nreg[388]), .Z(n19944) );
  IV U22000 ( .A(n19942), .Z(n19953) );
  XOR U22001 ( .A(n19954), .B(n19955), .Z(n19942) );
  AND U22002 ( .A(n19956), .B(n19957), .Z(n19955) );
  XNOR U22003 ( .A(n19954), .B(n9979), .Z(n19957) );
  XNOR U22004 ( .A(n19950), .B(n19952), .Z(n9979) );
  NAND U22005 ( .A(n19958), .B(nreg[387]), .Z(n19952) );
  NAND U22006 ( .A(n12326), .B(nreg[387]), .Z(n19958) );
  XNOR U22007 ( .A(n19948), .B(n19959), .Z(n19950) );
  XOR U22008 ( .A(n19960), .B(n19961), .Z(n19948) );
  AND U22009 ( .A(n19962), .B(n19963), .Z(n19961) );
  XNOR U22010 ( .A(n19964), .B(n19960), .Z(n19963) );
  XOR U22011 ( .A(n19965), .B(nreg[387]), .Z(n19956) );
  IV U22012 ( .A(n19954), .Z(n19965) );
  XOR U22013 ( .A(n19966), .B(n19967), .Z(n19954) );
  AND U22014 ( .A(n19968), .B(n19969), .Z(n19967) );
  XNOR U22015 ( .A(n19966), .B(n9985), .Z(n19969) );
  XNOR U22016 ( .A(n19962), .B(n19964), .Z(n9985) );
  NAND U22017 ( .A(n19970), .B(nreg[386]), .Z(n19964) );
  NAND U22018 ( .A(n12326), .B(nreg[386]), .Z(n19970) );
  XNOR U22019 ( .A(n19960), .B(n19971), .Z(n19962) );
  XOR U22020 ( .A(n19972), .B(n19973), .Z(n19960) );
  AND U22021 ( .A(n19974), .B(n19975), .Z(n19973) );
  XNOR U22022 ( .A(n19976), .B(n19972), .Z(n19975) );
  XOR U22023 ( .A(n19977), .B(nreg[386]), .Z(n19968) );
  IV U22024 ( .A(n19966), .Z(n19977) );
  XOR U22025 ( .A(n19978), .B(n19979), .Z(n19966) );
  AND U22026 ( .A(n19980), .B(n19981), .Z(n19979) );
  XNOR U22027 ( .A(n19978), .B(n9991), .Z(n19981) );
  XNOR U22028 ( .A(n19974), .B(n19976), .Z(n9991) );
  NAND U22029 ( .A(n19982), .B(nreg[385]), .Z(n19976) );
  NAND U22030 ( .A(n12326), .B(nreg[385]), .Z(n19982) );
  XNOR U22031 ( .A(n19972), .B(n19983), .Z(n19974) );
  XOR U22032 ( .A(n19984), .B(n19985), .Z(n19972) );
  AND U22033 ( .A(n19986), .B(n19987), .Z(n19985) );
  XNOR U22034 ( .A(n19988), .B(n19984), .Z(n19987) );
  XOR U22035 ( .A(n19989), .B(nreg[385]), .Z(n19980) );
  IV U22036 ( .A(n19978), .Z(n19989) );
  XOR U22037 ( .A(n19990), .B(n19991), .Z(n19978) );
  AND U22038 ( .A(n19992), .B(n19993), .Z(n19991) );
  XNOR U22039 ( .A(n19990), .B(n9997), .Z(n19993) );
  XNOR U22040 ( .A(n19986), .B(n19988), .Z(n9997) );
  NAND U22041 ( .A(n19994), .B(nreg[384]), .Z(n19988) );
  NAND U22042 ( .A(n12326), .B(nreg[384]), .Z(n19994) );
  XNOR U22043 ( .A(n19984), .B(n19995), .Z(n19986) );
  XOR U22044 ( .A(n19996), .B(n19997), .Z(n19984) );
  AND U22045 ( .A(n19998), .B(n19999), .Z(n19997) );
  XNOR U22046 ( .A(n20000), .B(n19996), .Z(n19999) );
  XOR U22047 ( .A(n20001), .B(nreg[384]), .Z(n19992) );
  IV U22048 ( .A(n19990), .Z(n20001) );
  XOR U22049 ( .A(n20002), .B(n20003), .Z(n19990) );
  AND U22050 ( .A(n20004), .B(n20005), .Z(n20003) );
  XNOR U22051 ( .A(n20002), .B(n10003), .Z(n20005) );
  XNOR U22052 ( .A(n19998), .B(n20000), .Z(n10003) );
  NAND U22053 ( .A(n20006), .B(nreg[383]), .Z(n20000) );
  NAND U22054 ( .A(n12326), .B(nreg[383]), .Z(n20006) );
  XNOR U22055 ( .A(n19996), .B(n20007), .Z(n19998) );
  XOR U22056 ( .A(n20008), .B(n20009), .Z(n19996) );
  AND U22057 ( .A(n20010), .B(n20011), .Z(n20009) );
  XNOR U22058 ( .A(n20012), .B(n20008), .Z(n20011) );
  XOR U22059 ( .A(n20013), .B(nreg[383]), .Z(n20004) );
  IV U22060 ( .A(n20002), .Z(n20013) );
  XOR U22061 ( .A(n20014), .B(n20015), .Z(n20002) );
  AND U22062 ( .A(n20016), .B(n20017), .Z(n20015) );
  XNOR U22063 ( .A(n20014), .B(n10009), .Z(n20017) );
  XNOR U22064 ( .A(n20010), .B(n20012), .Z(n10009) );
  NAND U22065 ( .A(n20018), .B(nreg[382]), .Z(n20012) );
  NAND U22066 ( .A(n12326), .B(nreg[382]), .Z(n20018) );
  XNOR U22067 ( .A(n20008), .B(n20019), .Z(n20010) );
  XOR U22068 ( .A(n20020), .B(n20021), .Z(n20008) );
  AND U22069 ( .A(n20022), .B(n20023), .Z(n20021) );
  XNOR U22070 ( .A(n20024), .B(n20020), .Z(n20023) );
  XOR U22071 ( .A(n20025), .B(nreg[382]), .Z(n20016) );
  IV U22072 ( .A(n20014), .Z(n20025) );
  XOR U22073 ( .A(n20026), .B(n20027), .Z(n20014) );
  AND U22074 ( .A(n20028), .B(n20029), .Z(n20027) );
  XNOR U22075 ( .A(n20026), .B(n10015), .Z(n20029) );
  XNOR U22076 ( .A(n20022), .B(n20024), .Z(n10015) );
  NAND U22077 ( .A(n20030), .B(nreg[381]), .Z(n20024) );
  NAND U22078 ( .A(n12326), .B(nreg[381]), .Z(n20030) );
  XNOR U22079 ( .A(n20020), .B(n20031), .Z(n20022) );
  XOR U22080 ( .A(n20032), .B(n20033), .Z(n20020) );
  AND U22081 ( .A(n20034), .B(n20035), .Z(n20033) );
  XNOR U22082 ( .A(n20036), .B(n20032), .Z(n20035) );
  XOR U22083 ( .A(n20037), .B(nreg[381]), .Z(n20028) );
  IV U22084 ( .A(n20026), .Z(n20037) );
  XOR U22085 ( .A(n20038), .B(n20039), .Z(n20026) );
  AND U22086 ( .A(n20040), .B(n20041), .Z(n20039) );
  XNOR U22087 ( .A(n20038), .B(n10021), .Z(n20041) );
  XNOR U22088 ( .A(n20034), .B(n20036), .Z(n10021) );
  NAND U22089 ( .A(n20042), .B(nreg[380]), .Z(n20036) );
  NAND U22090 ( .A(n12326), .B(nreg[380]), .Z(n20042) );
  XNOR U22091 ( .A(n20032), .B(n20043), .Z(n20034) );
  XOR U22092 ( .A(n20044), .B(n20045), .Z(n20032) );
  AND U22093 ( .A(n20046), .B(n20047), .Z(n20045) );
  XNOR U22094 ( .A(n20048), .B(n20044), .Z(n20047) );
  XOR U22095 ( .A(n20049), .B(nreg[380]), .Z(n20040) );
  IV U22096 ( .A(n20038), .Z(n20049) );
  XOR U22097 ( .A(n20050), .B(n20051), .Z(n20038) );
  AND U22098 ( .A(n20052), .B(n20053), .Z(n20051) );
  XNOR U22099 ( .A(n20050), .B(n10027), .Z(n20053) );
  XNOR U22100 ( .A(n20046), .B(n20048), .Z(n10027) );
  NAND U22101 ( .A(n20054), .B(nreg[379]), .Z(n20048) );
  NAND U22102 ( .A(n12326), .B(nreg[379]), .Z(n20054) );
  XNOR U22103 ( .A(n20044), .B(n20055), .Z(n20046) );
  XOR U22104 ( .A(n20056), .B(n20057), .Z(n20044) );
  AND U22105 ( .A(n20058), .B(n20059), .Z(n20057) );
  XNOR U22106 ( .A(n20060), .B(n20056), .Z(n20059) );
  XOR U22107 ( .A(n20061), .B(nreg[379]), .Z(n20052) );
  IV U22108 ( .A(n20050), .Z(n20061) );
  XOR U22109 ( .A(n20062), .B(n20063), .Z(n20050) );
  AND U22110 ( .A(n20064), .B(n20065), .Z(n20063) );
  XNOR U22111 ( .A(n20062), .B(n10033), .Z(n20065) );
  XNOR U22112 ( .A(n20058), .B(n20060), .Z(n10033) );
  NAND U22113 ( .A(n20066), .B(nreg[378]), .Z(n20060) );
  NAND U22114 ( .A(n12326), .B(nreg[378]), .Z(n20066) );
  XNOR U22115 ( .A(n20056), .B(n20067), .Z(n20058) );
  XOR U22116 ( .A(n20068), .B(n20069), .Z(n20056) );
  AND U22117 ( .A(n20070), .B(n20071), .Z(n20069) );
  XNOR U22118 ( .A(n20072), .B(n20068), .Z(n20071) );
  XOR U22119 ( .A(n20073), .B(nreg[378]), .Z(n20064) );
  IV U22120 ( .A(n20062), .Z(n20073) );
  XOR U22121 ( .A(n20074), .B(n20075), .Z(n20062) );
  AND U22122 ( .A(n20076), .B(n20077), .Z(n20075) );
  XNOR U22123 ( .A(n20074), .B(n10039), .Z(n20077) );
  XNOR U22124 ( .A(n20070), .B(n20072), .Z(n10039) );
  NAND U22125 ( .A(n20078), .B(nreg[377]), .Z(n20072) );
  NAND U22126 ( .A(n12326), .B(nreg[377]), .Z(n20078) );
  XNOR U22127 ( .A(n20068), .B(n20079), .Z(n20070) );
  XOR U22128 ( .A(n20080), .B(n20081), .Z(n20068) );
  AND U22129 ( .A(n20082), .B(n20083), .Z(n20081) );
  XNOR U22130 ( .A(n20084), .B(n20080), .Z(n20083) );
  XOR U22131 ( .A(n20085), .B(nreg[377]), .Z(n20076) );
  IV U22132 ( .A(n20074), .Z(n20085) );
  XOR U22133 ( .A(n20086), .B(n20087), .Z(n20074) );
  AND U22134 ( .A(n20088), .B(n20089), .Z(n20087) );
  XNOR U22135 ( .A(n20086), .B(n10045), .Z(n20089) );
  XNOR U22136 ( .A(n20082), .B(n20084), .Z(n10045) );
  NAND U22137 ( .A(n20090), .B(nreg[376]), .Z(n20084) );
  NAND U22138 ( .A(n12326), .B(nreg[376]), .Z(n20090) );
  XNOR U22139 ( .A(n20080), .B(n20091), .Z(n20082) );
  XOR U22140 ( .A(n20092), .B(n20093), .Z(n20080) );
  AND U22141 ( .A(n20094), .B(n20095), .Z(n20093) );
  XNOR U22142 ( .A(n20096), .B(n20092), .Z(n20095) );
  XOR U22143 ( .A(n20097), .B(nreg[376]), .Z(n20088) );
  IV U22144 ( .A(n20086), .Z(n20097) );
  XOR U22145 ( .A(n20098), .B(n20099), .Z(n20086) );
  AND U22146 ( .A(n20100), .B(n20101), .Z(n20099) );
  XNOR U22147 ( .A(n20098), .B(n10051), .Z(n20101) );
  XNOR U22148 ( .A(n20094), .B(n20096), .Z(n10051) );
  NAND U22149 ( .A(n20102), .B(nreg[375]), .Z(n20096) );
  NAND U22150 ( .A(n12326), .B(nreg[375]), .Z(n20102) );
  XNOR U22151 ( .A(n20092), .B(n20103), .Z(n20094) );
  XOR U22152 ( .A(n20104), .B(n20105), .Z(n20092) );
  AND U22153 ( .A(n20106), .B(n20107), .Z(n20105) );
  XNOR U22154 ( .A(n20108), .B(n20104), .Z(n20107) );
  XOR U22155 ( .A(n20109), .B(nreg[375]), .Z(n20100) );
  IV U22156 ( .A(n20098), .Z(n20109) );
  XOR U22157 ( .A(n20110), .B(n20111), .Z(n20098) );
  AND U22158 ( .A(n20112), .B(n20113), .Z(n20111) );
  XNOR U22159 ( .A(n20110), .B(n10057), .Z(n20113) );
  XNOR U22160 ( .A(n20106), .B(n20108), .Z(n10057) );
  NAND U22161 ( .A(n20114), .B(nreg[374]), .Z(n20108) );
  NAND U22162 ( .A(n12326), .B(nreg[374]), .Z(n20114) );
  XNOR U22163 ( .A(n20104), .B(n20115), .Z(n20106) );
  XOR U22164 ( .A(n20116), .B(n20117), .Z(n20104) );
  AND U22165 ( .A(n20118), .B(n20119), .Z(n20117) );
  XNOR U22166 ( .A(n20120), .B(n20116), .Z(n20119) );
  XOR U22167 ( .A(n20121), .B(nreg[374]), .Z(n20112) );
  IV U22168 ( .A(n20110), .Z(n20121) );
  XOR U22169 ( .A(n20122), .B(n20123), .Z(n20110) );
  AND U22170 ( .A(n20124), .B(n20125), .Z(n20123) );
  XNOR U22171 ( .A(n20122), .B(n10063), .Z(n20125) );
  XNOR U22172 ( .A(n20118), .B(n20120), .Z(n10063) );
  NAND U22173 ( .A(n20126), .B(nreg[373]), .Z(n20120) );
  NAND U22174 ( .A(n12326), .B(nreg[373]), .Z(n20126) );
  XNOR U22175 ( .A(n20116), .B(n20127), .Z(n20118) );
  XOR U22176 ( .A(n20128), .B(n20129), .Z(n20116) );
  AND U22177 ( .A(n20130), .B(n20131), .Z(n20129) );
  XNOR U22178 ( .A(n20132), .B(n20128), .Z(n20131) );
  XOR U22179 ( .A(n20133), .B(nreg[373]), .Z(n20124) );
  IV U22180 ( .A(n20122), .Z(n20133) );
  XOR U22181 ( .A(n20134), .B(n20135), .Z(n20122) );
  AND U22182 ( .A(n20136), .B(n20137), .Z(n20135) );
  XNOR U22183 ( .A(n20134), .B(n10069), .Z(n20137) );
  XNOR U22184 ( .A(n20130), .B(n20132), .Z(n10069) );
  NAND U22185 ( .A(n20138), .B(nreg[372]), .Z(n20132) );
  NAND U22186 ( .A(n12326), .B(nreg[372]), .Z(n20138) );
  XNOR U22187 ( .A(n20128), .B(n20139), .Z(n20130) );
  XOR U22188 ( .A(n20140), .B(n20141), .Z(n20128) );
  AND U22189 ( .A(n20142), .B(n20143), .Z(n20141) );
  XNOR U22190 ( .A(n20144), .B(n20140), .Z(n20143) );
  XOR U22191 ( .A(n20145), .B(nreg[372]), .Z(n20136) );
  IV U22192 ( .A(n20134), .Z(n20145) );
  XOR U22193 ( .A(n20146), .B(n20147), .Z(n20134) );
  AND U22194 ( .A(n20148), .B(n20149), .Z(n20147) );
  XNOR U22195 ( .A(n20146), .B(n10075), .Z(n20149) );
  XNOR U22196 ( .A(n20142), .B(n20144), .Z(n10075) );
  NAND U22197 ( .A(n20150), .B(nreg[371]), .Z(n20144) );
  NAND U22198 ( .A(n12326), .B(nreg[371]), .Z(n20150) );
  XNOR U22199 ( .A(n20140), .B(n20151), .Z(n20142) );
  XOR U22200 ( .A(n20152), .B(n20153), .Z(n20140) );
  AND U22201 ( .A(n20154), .B(n20155), .Z(n20153) );
  XNOR U22202 ( .A(n20156), .B(n20152), .Z(n20155) );
  XOR U22203 ( .A(n20157), .B(nreg[371]), .Z(n20148) );
  IV U22204 ( .A(n20146), .Z(n20157) );
  XOR U22205 ( .A(n20158), .B(n20159), .Z(n20146) );
  AND U22206 ( .A(n20160), .B(n20161), .Z(n20159) );
  XNOR U22207 ( .A(n20158), .B(n10081), .Z(n20161) );
  XNOR U22208 ( .A(n20154), .B(n20156), .Z(n10081) );
  NAND U22209 ( .A(n20162), .B(nreg[370]), .Z(n20156) );
  NAND U22210 ( .A(n12326), .B(nreg[370]), .Z(n20162) );
  XNOR U22211 ( .A(n20152), .B(n20163), .Z(n20154) );
  XOR U22212 ( .A(n20164), .B(n20165), .Z(n20152) );
  AND U22213 ( .A(n20166), .B(n20167), .Z(n20165) );
  XNOR U22214 ( .A(n20168), .B(n20164), .Z(n20167) );
  XOR U22215 ( .A(n20169), .B(nreg[370]), .Z(n20160) );
  IV U22216 ( .A(n20158), .Z(n20169) );
  XOR U22217 ( .A(n20170), .B(n20171), .Z(n20158) );
  AND U22218 ( .A(n20172), .B(n20173), .Z(n20171) );
  XNOR U22219 ( .A(n20170), .B(n10087), .Z(n20173) );
  XNOR U22220 ( .A(n20166), .B(n20168), .Z(n10087) );
  NAND U22221 ( .A(n20174), .B(nreg[369]), .Z(n20168) );
  NAND U22222 ( .A(n12326), .B(nreg[369]), .Z(n20174) );
  XNOR U22223 ( .A(n20164), .B(n20175), .Z(n20166) );
  XOR U22224 ( .A(n20176), .B(n20177), .Z(n20164) );
  AND U22225 ( .A(n20178), .B(n20179), .Z(n20177) );
  XNOR U22226 ( .A(n20180), .B(n20176), .Z(n20179) );
  XOR U22227 ( .A(n20181), .B(nreg[369]), .Z(n20172) );
  IV U22228 ( .A(n20170), .Z(n20181) );
  XOR U22229 ( .A(n20182), .B(n20183), .Z(n20170) );
  AND U22230 ( .A(n20184), .B(n20185), .Z(n20183) );
  XNOR U22231 ( .A(n20182), .B(n10093), .Z(n20185) );
  XNOR U22232 ( .A(n20178), .B(n20180), .Z(n10093) );
  NAND U22233 ( .A(n20186), .B(nreg[368]), .Z(n20180) );
  NAND U22234 ( .A(n12326), .B(nreg[368]), .Z(n20186) );
  XNOR U22235 ( .A(n20176), .B(n20187), .Z(n20178) );
  XOR U22236 ( .A(n20188), .B(n20189), .Z(n20176) );
  AND U22237 ( .A(n20190), .B(n20191), .Z(n20189) );
  XNOR U22238 ( .A(n20192), .B(n20188), .Z(n20191) );
  XOR U22239 ( .A(n20193), .B(nreg[368]), .Z(n20184) );
  IV U22240 ( .A(n20182), .Z(n20193) );
  XOR U22241 ( .A(n20194), .B(n20195), .Z(n20182) );
  AND U22242 ( .A(n20196), .B(n20197), .Z(n20195) );
  XNOR U22243 ( .A(n20194), .B(n10099), .Z(n20197) );
  XNOR U22244 ( .A(n20190), .B(n20192), .Z(n10099) );
  NAND U22245 ( .A(n20198), .B(nreg[367]), .Z(n20192) );
  NAND U22246 ( .A(n12326), .B(nreg[367]), .Z(n20198) );
  XNOR U22247 ( .A(n20188), .B(n20199), .Z(n20190) );
  XOR U22248 ( .A(n20200), .B(n20201), .Z(n20188) );
  AND U22249 ( .A(n20202), .B(n20203), .Z(n20201) );
  XNOR U22250 ( .A(n20204), .B(n20200), .Z(n20203) );
  XOR U22251 ( .A(n20205), .B(nreg[367]), .Z(n20196) );
  IV U22252 ( .A(n20194), .Z(n20205) );
  XOR U22253 ( .A(n20206), .B(n20207), .Z(n20194) );
  AND U22254 ( .A(n20208), .B(n20209), .Z(n20207) );
  XNOR U22255 ( .A(n20206), .B(n10105), .Z(n20209) );
  XNOR U22256 ( .A(n20202), .B(n20204), .Z(n10105) );
  NAND U22257 ( .A(n20210), .B(nreg[366]), .Z(n20204) );
  NAND U22258 ( .A(n12326), .B(nreg[366]), .Z(n20210) );
  XNOR U22259 ( .A(n20200), .B(n20211), .Z(n20202) );
  XOR U22260 ( .A(n20212), .B(n20213), .Z(n20200) );
  AND U22261 ( .A(n20214), .B(n20215), .Z(n20213) );
  XNOR U22262 ( .A(n20216), .B(n20212), .Z(n20215) );
  XOR U22263 ( .A(n20217), .B(nreg[366]), .Z(n20208) );
  IV U22264 ( .A(n20206), .Z(n20217) );
  XOR U22265 ( .A(n20218), .B(n20219), .Z(n20206) );
  AND U22266 ( .A(n20220), .B(n20221), .Z(n20219) );
  XNOR U22267 ( .A(n20218), .B(n10111), .Z(n20221) );
  XNOR U22268 ( .A(n20214), .B(n20216), .Z(n10111) );
  NAND U22269 ( .A(n20222), .B(nreg[365]), .Z(n20216) );
  NAND U22270 ( .A(n12326), .B(nreg[365]), .Z(n20222) );
  XNOR U22271 ( .A(n20212), .B(n20223), .Z(n20214) );
  XOR U22272 ( .A(n20224), .B(n20225), .Z(n20212) );
  AND U22273 ( .A(n20226), .B(n20227), .Z(n20225) );
  XNOR U22274 ( .A(n20228), .B(n20224), .Z(n20227) );
  XOR U22275 ( .A(n20229), .B(nreg[365]), .Z(n20220) );
  IV U22276 ( .A(n20218), .Z(n20229) );
  XOR U22277 ( .A(n20230), .B(n20231), .Z(n20218) );
  AND U22278 ( .A(n20232), .B(n20233), .Z(n20231) );
  XNOR U22279 ( .A(n20230), .B(n10117), .Z(n20233) );
  XNOR U22280 ( .A(n20226), .B(n20228), .Z(n10117) );
  NAND U22281 ( .A(n20234), .B(nreg[364]), .Z(n20228) );
  NAND U22282 ( .A(n12326), .B(nreg[364]), .Z(n20234) );
  XNOR U22283 ( .A(n20224), .B(n20235), .Z(n20226) );
  XOR U22284 ( .A(n20236), .B(n20237), .Z(n20224) );
  AND U22285 ( .A(n20238), .B(n20239), .Z(n20237) );
  XNOR U22286 ( .A(n20240), .B(n20236), .Z(n20239) );
  XOR U22287 ( .A(n20241), .B(nreg[364]), .Z(n20232) );
  IV U22288 ( .A(n20230), .Z(n20241) );
  XOR U22289 ( .A(n20242), .B(n20243), .Z(n20230) );
  AND U22290 ( .A(n20244), .B(n20245), .Z(n20243) );
  XNOR U22291 ( .A(n20242), .B(n10123), .Z(n20245) );
  XNOR U22292 ( .A(n20238), .B(n20240), .Z(n10123) );
  NAND U22293 ( .A(n20246), .B(nreg[363]), .Z(n20240) );
  NAND U22294 ( .A(n12326), .B(nreg[363]), .Z(n20246) );
  XNOR U22295 ( .A(n20236), .B(n20247), .Z(n20238) );
  XOR U22296 ( .A(n20248), .B(n20249), .Z(n20236) );
  AND U22297 ( .A(n20250), .B(n20251), .Z(n20249) );
  XNOR U22298 ( .A(n20252), .B(n20248), .Z(n20251) );
  XOR U22299 ( .A(n20253), .B(nreg[363]), .Z(n20244) );
  IV U22300 ( .A(n20242), .Z(n20253) );
  XOR U22301 ( .A(n20254), .B(n20255), .Z(n20242) );
  AND U22302 ( .A(n20256), .B(n20257), .Z(n20255) );
  XNOR U22303 ( .A(n20254), .B(n10129), .Z(n20257) );
  XNOR U22304 ( .A(n20250), .B(n20252), .Z(n10129) );
  NAND U22305 ( .A(n20258), .B(nreg[362]), .Z(n20252) );
  NAND U22306 ( .A(n12326), .B(nreg[362]), .Z(n20258) );
  XNOR U22307 ( .A(n20248), .B(n20259), .Z(n20250) );
  XOR U22308 ( .A(n20260), .B(n20261), .Z(n20248) );
  AND U22309 ( .A(n20262), .B(n20263), .Z(n20261) );
  XNOR U22310 ( .A(n20264), .B(n20260), .Z(n20263) );
  XOR U22311 ( .A(n20265), .B(nreg[362]), .Z(n20256) );
  IV U22312 ( .A(n20254), .Z(n20265) );
  XOR U22313 ( .A(n20266), .B(n20267), .Z(n20254) );
  AND U22314 ( .A(n20268), .B(n20269), .Z(n20267) );
  XNOR U22315 ( .A(n20266), .B(n10135), .Z(n20269) );
  XNOR U22316 ( .A(n20262), .B(n20264), .Z(n10135) );
  NAND U22317 ( .A(n20270), .B(nreg[361]), .Z(n20264) );
  NAND U22318 ( .A(n12326), .B(nreg[361]), .Z(n20270) );
  XNOR U22319 ( .A(n20260), .B(n20271), .Z(n20262) );
  XOR U22320 ( .A(n20272), .B(n20273), .Z(n20260) );
  AND U22321 ( .A(n20274), .B(n20275), .Z(n20273) );
  XNOR U22322 ( .A(n20276), .B(n20272), .Z(n20275) );
  XOR U22323 ( .A(n20277), .B(nreg[361]), .Z(n20268) );
  IV U22324 ( .A(n20266), .Z(n20277) );
  XOR U22325 ( .A(n20278), .B(n20279), .Z(n20266) );
  AND U22326 ( .A(n20280), .B(n20281), .Z(n20279) );
  XNOR U22327 ( .A(n20278), .B(n10141), .Z(n20281) );
  XNOR U22328 ( .A(n20274), .B(n20276), .Z(n10141) );
  NAND U22329 ( .A(n20282), .B(nreg[360]), .Z(n20276) );
  NAND U22330 ( .A(n12326), .B(nreg[360]), .Z(n20282) );
  XNOR U22331 ( .A(n20272), .B(n20283), .Z(n20274) );
  XOR U22332 ( .A(n20284), .B(n20285), .Z(n20272) );
  AND U22333 ( .A(n20286), .B(n20287), .Z(n20285) );
  XNOR U22334 ( .A(n20288), .B(n20284), .Z(n20287) );
  XOR U22335 ( .A(n20289), .B(nreg[360]), .Z(n20280) );
  IV U22336 ( .A(n20278), .Z(n20289) );
  XOR U22337 ( .A(n20290), .B(n20291), .Z(n20278) );
  AND U22338 ( .A(n20292), .B(n20293), .Z(n20291) );
  XNOR U22339 ( .A(n20290), .B(n10147), .Z(n20293) );
  XNOR U22340 ( .A(n20286), .B(n20288), .Z(n10147) );
  NAND U22341 ( .A(n20294), .B(nreg[359]), .Z(n20288) );
  NAND U22342 ( .A(n12326), .B(nreg[359]), .Z(n20294) );
  XNOR U22343 ( .A(n20284), .B(n20295), .Z(n20286) );
  XOR U22344 ( .A(n20296), .B(n20297), .Z(n20284) );
  AND U22345 ( .A(n20298), .B(n20299), .Z(n20297) );
  XNOR U22346 ( .A(n20300), .B(n20296), .Z(n20299) );
  XOR U22347 ( .A(n20301), .B(nreg[359]), .Z(n20292) );
  IV U22348 ( .A(n20290), .Z(n20301) );
  XOR U22349 ( .A(n20302), .B(n20303), .Z(n20290) );
  AND U22350 ( .A(n20304), .B(n20305), .Z(n20303) );
  XNOR U22351 ( .A(n20302), .B(n10153), .Z(n20305) );
  XNOR U22352 ( .A(n20298), .B(n20300), .Z(n10153) );
  NAND U22353 ( .A(n20306), .B(nreg[358]), .Z(n20300) );
  NAND U22354 ( .A(n12326), .B(nreg[358]), .Z(n20306) );
  XNOR U22355 ( .A(n20296), .B(n20307), .Z(n20298) );
  XOR U22356 ( .A(n20308), .B(n20309), .Z(n20296) );
  AND U22357 ( .A(n20310), .B(n20311), .Z(n20309) );
  XNOR U22358 ( .A(n20312), .B(n20308), .Z(n20311) );
  XOR U22359 ( .A(n20313), .B(nreg[358]), .Z(n20304) );
  IV U22360 ( .A(n20302), .Z(n20313) );
  XOR U22361 ( .A(n20314), .B(n20315), .Z(n20302) );
  AND U22362 ( .A(n20316), .B(n20317), .Z(n20315) );
  XNOR U22363 ( .A(n20314), .B(n10159), .Z(n20317) );
  XNOR U22364 ( .A(n20310), .B(n20312), .Z(n10159) );
  NAND U22365 ( .A(n20318), .B(nreg[357]), .Z(n20312) );
  NAND U22366 ( .A(n12326), .B(nreg[357]), .Z(n20318) );
  XNOR U22367 ( .A(n20308), .B(n20319), .Z(n20310) );
  XOR U22368 ( .A(n20320), .B(n20321), .Z(n20308) );
  AND U22369 ( .A(n20322), .B(n20323), .Z(n20321) );
  XNOR U22370 ( .A(n20324), .B(n20320), .Z(n20323) );
  XOR U22371 ( .A(n20325), .B(nreg[357]), .Z(n20316) );
  IV U22372 ( .A(n20314), .Z(n20325) );
  XOR U22373 ( .A(n20326), .B(n20327), .Z(n20314) );
  AND U22374 ( .A(n20328), .B(n20329), .Z(n20327) );
  XNOR U22375 ( .A(n20326), .B(n10165), .Z(n20329) );
  XNOR U22376 ( .A(n20322), .B(n20324), .Z(n10165) );
  NAND U22377 ( .A(n20330), .B(nreg[356]), .Z(n20324) );
  NAND U22378 ( .A(n12326), .B(nreg[356]), .Z(n20330) );
  XNOR U22379 ( .A(n20320), .B(n20331), .Z(n20322) );
  XOR U22380 ( .A(n20332), .B(n20333), .Z(n20320) );
  AND U22381 ( .A(n20334), .B(n20335), .Z(n20333) );
  XNOR U22382 ( .A(n20336), .B(n20332), .Z(n20335) );
  XOR U22383 ( .A(n20337), .B(nreg[356]), .Z(n20328) );
  IV U22384 ( .A(n20326), .Z(n20337) );
  XOR U22385 ( .A(n20338), .B(n20339), .Z(n20326) );
  AND U22386 ( .A(n20340), .B(n20341), .Z(n20339) );
  XNOR U22387 ( .A(n20338), .B(n10171), .Z(n20341) );
  XNOR U22388 ( .A(n20334), .B(n20336), .Z(n10171) );
  NAND U22389 ( .A(n20342), .B(nreg[355]), .Z(n20336) );
  NAND U22390 ( .A(n12326), .B(nreg[355]), .Z(n20342) );
  XNOR U22391 ( .A(n20332), .B(n20343), .Z(n20334) );
  XOR U22392 ( .A(n20344), .B(n20345), .Z(n20332) );
  AND U22393 ( .A(n20346), .B(n20347), .Z(n20345) );
  XNOR U22394 ( .A(n20348), .B(n20344), .Z(n20347) );
  XOR U22395 ( .A(n20349), .B(nreg[355]), .Z(n20340) );
  IV U22396 ( .A(n20338), .Z(n20349) );
  XOR U22397 ( .A(n20350), .B(n20351), .Z(n20338) );
  AND U22398 ( .A(n20352), .B(n20353), .Z(n20351) );
  XNOR U22399 ( .A(n20350), .B(n10177), .Z(n20353) );
  XNOR U22400 ( .A(n20346), .B(n20348), .Z(n10177) );
  NAND U22401 ( .A(n20354), .B(nreg[354]), .Z(n20348) );
  NAND U22402 ( .A(n12326), .B(nreg[354]), .Z(n20354) );
  XNOR U22403 ( .A(n20344), .B(n20355), .Z(n20346) );
  XOR U22404 ( .A(n20356), .B(n20357), .Z(n20344) );
  AND U22405 ( .A(n20358), .B(n20359), .Z(n20357) );
  XNOR U22406 ( .A(n20360), .B(n20356), .Z(n20359) );
  XOR U22407 ( .A(n20361), .B(nreg[354]), .Z(n20352) );
  IV U22408 ( .A(n20350), .Z(n20361) );
  XOR U22409 ( .A(n20362), .B(n20363), .Z(n20350) );
  AND U22410 ( .A(n20364), .B(n20365), .Z(n20363) );
  XNOR U22411 ( .A(n20362), .B(n10183), .Z(n20365) );
  XNOR U22412 ( .A(n20358), .B(n20360), .Z(n10183) );
  NAND U22413 ( .A(n20366), .B(nreg[353]), .Z(n20360) );
  NAND U22414 ( .A(n12326), .B(nreg[353]), .Z(n20366) );
  XNOR U22415 ( .A(n20356), .B(n20367), .Z(n20358) );
  XOR U22416 ( .A(n20368), .B(n20369), .Z(n20356) );
  AND U22417 ( .A(n20370), .B(n20371), .Z(n20369) );
  XNOR U22418 ( .A(n20372), .B(n20368), .Z(n20371) );
  XOR U22419 ( .A(n20373), .B(nreg[353]), .Z(n20364) );
  IV U22420 ( .A(n20362), .Z(n20373) );
  XOR U22421 ( .A(n20374), .B(n20375), .Z(n20362) );
  AND U22422 ( .A(n20376), .B(n20377), .Z(n20375) );
  XNOR U22423 ( .A(n20374), .B(n10189), .Z(n20377) );
  XNOR U22424 ( .A(n20370), .B(n20372), .Z(n10189) );
  NAND U22425 ( .A(n20378), .B(nreg[352]), .Z(n20372) );
  NAND U22426 ( .A(n12326), .B(nreg[352]), .Z(n20378) );
  XNOR U22427 ( .A(n20368), .B(n20379), .Z(n20370) );
  XOR U22428 ( .A(n20380), .B(n20381), .Z(n20368) );
  AND U22429 ( .A(n20382), .B(n20383), .Z(n20381) );
  XNOR U22430 ( .A(n20384), .B(n20380), .Z(n20383) );
  XOR U22431 ( .A(n20385), .B(nreg[352]), .Z(n20376) );
  IV U22432 ( .A(n20374), .Z(n20385) );
  XOR U22433 ( .A(n20386), .B(n20387), .Z(n20374) );
  AND U22434 ( .A(n20388), .B(n20389), .Z(n20387) );
  XNOR U22435 ( .A(n20386), .B(n10195), .Z(n20389) );
  XNOR U22436 ( .A(n20382), .B(n20384), .Z(n10195) );
  NAND U22437 ( .A(n20390), .B(nreg[351]), .Z(n20384) );
  NAND U22438 ( .A(n12326), .B(nreg[351]), .Z(n20390) );
  XNOR U22439 ( .A(n20380), .B(n20391), .Z(n20382) );
  XOR U22440 ( .A(n20392), .B(n20393), .Z(n20380) );
  AND U22441 ( .A(n20394), .B(n20395), .Z(n20393) );
  XNOR U22442 ( .A(n20396), .B(n20392), .Z(n20395) );
  XOR U22443 ( .A(n20397), .B(nreg[351]), .Z(n20388) );
  IV U22444 ( .A(n20386), .Z(n20397) );
  XOR U22445 ( .A(n20398), .B(n20399), .Z(n20386) );
  AND U22446 ( .A(n20400), .B(n20401), .Z(n20399) );
  XNOR U22447 ( .A(n20398), .B(n10201), .Z(n20401) );
  XNOR U22448 ( .A(n20394), .B(n20396), .Z(n10201) );
  NAND U22449 ( .A(n20402), .B(nreg[350]), .Z(n20396) );
  NAND U22450 ( .A(n12326), .B(nreg[350]), .Z(n20402) );
  XNOR U22451 ( .A(n20392), .B(n20403), .Z(n20394) );
  XOR U22452 ( .A(n20404), .B(n20405), .Z(n20392) );
  AND U22453 ( .A(n20406), .B(n20407), .Z(n20405) );
  XNOR U22454 ( .A(n20408), .B(n20404), .Z(n20407) );
  XOR U22455 ( .A(n20409), .B(nreg[350]), .Z(n20400) );
  IV U22456 ( .A(n20398), .Z(n20409) );
  XOR U22457 ( .A(n20410), .B(n20411), .Z(n20398) );
  AND U22458 ( .A(n20412), .B(n20413), .Z(n20411) );
  XNOR U22459 ( .A(n20410), .B(n10207), .Z(n20413) );
  XNOR U22460 ( .A(n20406), .B(n20408), .Z(n10207) );
  NAND U22461 ( .A(n20414), .B(nreg[349]), .Z(n20408) );
  NAND U22462 ( .A(n12326), .B(nreg[349]), .Z(n20414) );
  XNOR U22463 ( .A(n20404), .B(n20415), .Z(n20406) );
  XOR U22464 ( .A(n20416), .B(n20417), .Z(n20404) );
  AND U22465 ( .A(n20418), .B(n20419), .Z(n20417) );
  XNOR U22466 ( .A(n20420), .B(n20416), .Z(n20419) );
  XOR U22467 ( .A(n20421), .B(nreg[349]), .Z(n20412) );
  IV U22468 ( .A(n20410), .Z(n20421) );
  XOR U22469 ( .A(n20422), .B(n20423), .Z(n20410) );
  AND U22470 ( .A(n20424), .B(n20425), .Z(n20423) );
  XNOR U22471 ( .A(n20422), .B(n10213), .Z(n20425) );
  XNOR U22472 ( .A(n20418), .B(n20420), .Z(n10213) );
  NAND U22473 ( .A(n20426), .B(nreg[348]), .Z(n20420) );
  NAND U22474 ( .A(n12326), .B(nreg[348]), .Z(n20426) );
  XNOR U22475 ( .A(n20416), .B(n20427), .Z(n20418) );
  XOR U22476 ( .A(n20428), .B(n20429), .Z(n20416) );
  AND U22477 ( .A(n20430), .B(n20431), .Z(n20429) );
  XNOR U22478 ( .A(n20432), .B(n20428), .Z(n20431) );
  XOR U22479 ( .A(n20433), .B(nreg[348]), .Z(n20424) );
  IV U22480 ( .A(n20422), .Z(n20433) );
  XOR U22481 ( .A(n20434), .B(n20435), .Z(n20422) );
  AND U22482 ( .A(n20436), .B(n20437), .Z(n20435) );
  XNOR U22483 ( .A(n20434), .B(n10219), .Z(n20437) );
  XNOR U22484 ( .A(n20430), .B(n20432), .Z(n10219) );
  NAND U22485 ( .A(n20438), .B(nreg[347]), .Z(n20432) );
  NAND U22486 ( .A(n12326), .B(nreg[347]), .Z(n20438) );
  XNOR U22487 ( .A(n20428), .B(n20439), .Z(n20430) );
  XOR U22488 ( .A(n20440), .B(n20441), .Z(n20428) );
  AND U22489 ( .A(n20442), .B(n20443), .Z(n20441) );
  XNOR U22490 ( .A(n20444), .B(n20440), .Z(n20443) );
  XOR U22491 ( .A(n20445), .B(nreg[347]), .Z(n20436) );
  IV U22492 ( .A(n20434), .Z(n20445) );
  XOR U22493 ( .A(n20446), .B(n20447), .Z(n20434) );
  AND U22494 ( .A(n20448), .B(n20449), .Z(n20447) );
  XNOR U22495 ( .A(n20446), .B(n10225), .Z(n20449) );
  XNOR U22496 ( .A(n20442), .B(n20444), .Z(n10225) );
  NAND U22497 ( .A(n20450), .B(nreg[346]), .Z(n20444) );
  NAND U22498 ( .A(n12326), .B(nreg[346]), .Z(n20450) );
  XNOR U22499 ( .A(n20440), .B(n20451), .Z(n20442) );
  XOR U22500 ( .A(n20452), .B(n20453), .Z(n20440) );
  AND U22501 ( .A(n20454), .B(n20455), .Z(n20453) );
  XNOR U22502 ( .A(n20456), .B(n20452), .Z(n20455) );
  XOR U22503 ( .A(n20457), .B(nreg[346]), .Z(n20448) );
  IV U22504 ( .A(n20446), .Z(n20457) );
  XOR U22505 ( .A(n20458), .B(n20459), .Z(n20446) );
  AND U22506 ( .A(n20460), .B(n20461), .Z(n20459) );
  XNOR U22507 ( .A(n20458), .B(n10231), .Z(n20461) );
  XNOR U22508 ( .A(n20454), .B(n20456), .Z(n10231) );
  NAND U22509 ( .A(n20462), .B(nreg[345]), .Z(n20456) );
  NAND U22510 ( .A(n12326), .B(nreg[345]), .Z(n20462) );
  XNOR U22511 ( .A(n20452), .B(n20463), .Z(n20454) );
  XOR U22512 ( .A(n20464), .B(n20465), .Z(n20452) );
  AND U22513 ( .A(n20466), .B(n20467), .Z(n20465) );
  XNOR U22514 ( .A(n20468), .B(n20464), .Z(n20467) );
  XOR U22515 ( .A(n20469), .B(nreg[345]), .Z(n20460) );
  IV U22516 ( .A(n20458), .Z(n20469) );
  XOR U22517 ( .A(n20470), .B(n20471), .Z(n20458) );
  AND U22518 ( .A(n20472), .B(n20473), .Z(n20471) );
  XNOR U22519 ( .A(n20470), .B(n10237), .Z(n20473) );
  XNOR U22520 ( .A(n20466), .B(n20468), .Z(n10237) );
  NAND U22521 ( .A(n20474), .B(nreg[344]), .Z(n20468) );
  NAND U22522 ( .A(n12326), .B(nreg[344]), .Z(n20474) );
  XNOR U22523 ( .A(n20464), .B(n20475), .Z(n20466) );
  XOR U22524 ( .A(n20476), .B(n20477), .Z(n20464) );
  AND U22525 ( .A(n20478), .B(n20479), .Z(n20477) );
  XNOR U22526 ( .A(n20480), .B(n20476), .Z(n20479) );
  XOR U22527 ( .A(n20481), .B(nreg[344]), .Z(n20472) );
  IV U22528 ( .A(n20470), .Z(n20481) );
  XOR U22529 ( .A(n20482), .B(n20483), .Z(n20470) );
  AND U22530 ( .A(n20484), .B(n20485), .Z(n20483) );
  XNOR U22531 ( .A(n20482), .B(n10243), .Z(n20485) );
  XNOR U22532 ( .A(n20478), .B(n20480), .Z(n10243) );
  NAND U22533 ( .A(n20486), .B(nreg[343]), .Z(n20480) );
  NAND U22534 ( .A(n12326), .B(nreg[343]), .Z(n20486) );
  XNOR U22535 ( .A(n20476), .B(n20487), .Z(n20478) );
  XOR U22536 ( .A(n20488), .B(n20489), .Z(n20476) );
  AND U22537 ( .A(n20490), .B(n20491), .Z(n20489) );
  XNOR U22538 ( .A(n20492), .B(n20488), .Z(n20491) );
  XOR U22539 ( .A(n20493), .B(nreg[343]), .Z(n20484) );
  IV U22540 ( .A(n20482), .Z(n20493) );
  XOR U22541 ( .A(n20494), .B(n20495), .Z(n20482) );
  AND U22542 ( .A(n20496), .B(n20497), .Z(n20495) );
  XNOR U22543 ( .A(n20494), .B(n10249), .Z(n20497) );
  XNOR U22544 ( .A(n20490), .B(n20492), .Z(n10249) );
  NAND U22545 ( .A(n20498), .B(nreg[342]), .Z(n20492) );
  NAND U22546 ( .A(n12326), .B(nreg[342]), .Z(n20498) );
  XNOR U22547 ( .A(n20488), .B(n20499), .Z(n20490) );
  XOR U22548 ( .A(n20500), .B(n20501), .Z(n20488) );
  AND U22549 ( .A(n20502), .B(n20503), .Z(n20501) );
  XNOR U22550 ( .A(n20504), .B(n20500), .Z(n20503) );
  XOR U22551 ( .A(n20505), .B(nreg[342]), .Z(n20496) );
  IV U22552 ( .A(n20494), .Z(n20505) );
  XOR U22553 ( .A(n20506), .B(n20507), .Z(n20494) );
  AND U22554 ( .A(n20508), .B(n20509), .Z(n20507) );
  XNOR U22555 ( .A(n20506), .B(n10255), .Z(n20509) );
  XNOR U22556 ( .A(n20502), .B(n20504), .Z(n10255) );
  NAND U22557 ( .A(n20510), .B(nreg[341]), .Z(n20504) );
  NAND U22558 ( .A(n12326), .B(nreg[341]), .Z(n20510) );
  XNOR U22559 ( .A(n20500), .B(n20511), .Z(n20502) );
  XOR U22560 ( .A(n20512), .B(n20513), .Z(n20500) );
  AND U22561 ( .A(n20514), .B(n20515), .Z(n20513) );
  XNOR U22562 ( .A(n20516), .B(n20512), .Z(n20515) );
  XOR U22563 ( .A(n20517), .B(nreg[341]), .Z(n20508) );
  IV U22564 ( .A(n20506), .Z(n20517) );
  XOR U22565 ( .A(n20518), .B(n20519), .Z(n20506) );
  AND U22566 ( .A(n20520), .B(n20521), .Z(n20519) );
  XNOR U22567 ( .A(n20518), .B(n10261), .Z(n20521) );
  XNOR U22568 ( .A(n20514), .B(n20516), .Z(n10261) );
  NAND U22569 ( .A(n20522), .B(nreg[340]), .Z(n20516) );
  NAND U22570 ( .A(n12326), .B(nreg[340]), .Z(n20522) );
  XNOR U22571 ( .A(n20512), .B(n20523), .Z(n20514) );
  XOR U22572 ( .A(n20524), .B(n20525), .Z(n20512) );
  AND U22573 ( .A(n20526), .B(n20527), .Z(n20525) );
  XNOR U22574 ( .A(n20528), .B(n20524), .Z(n20527) );
  XOR U22575 ( .A(n20529), .B(nreg[340]), .Z(n20520) );
  IV U22576 ( .A(n20518), .Z(n20529) );
  XOR U22577 ( .A(n20530), .B(n20531), .Z(n20518) );
  AND U22578 ( .A(n20532), .B(n20533), .Z(n20531) );
  XNOR U22579 ( .A(n20530), .B(n10267), .Z(n20533) );
  XNOR U22580 ( .A(n20526), .B(n20528), .Z(n10267) );
  NAND U22581 ( .A(n20534), .B(nreg[339]), .Z(n20528) );
  NAND U22582 ( .A(n12326), .B(nreg[339]), .Z(n20534) );
  XNOR U22583 ( .A(n20524), .B(n20535), .Z(n20526) );
  XOR U22584 ( .A(n20536), .B(n20537), .Z(n20524) );
  AND U22585 ( .A(n20538), .B(n20539), .Z(n20537) );
  XNOR U22586 ( .A(n20540), .B(n20536), .Z(n20539) );
  XOR U22587 ( .A(n20541), .B(nreg[339]), .Z(n20532) );
  IV U22588 ( .A(n20530), .Z(n20541) );
  XOR U22589 ( .A(n20542), .B(n20543), .Z(n20530) );
  AND U22590 ( .A(n20544), .B(n20545), .Z(n20543) );
  XNOR U22591 ( .A(n20542), .B(n10273), .Z(n20545) );
  XNOR U22592 ( .A(n20538), .B(n20540), .Z(n10273) );
  NAND U22593 ( .A(n20546), .B(nreg[338]), .Z(n20540) );
  NAND U22594 ( .A(n12326), .B(nreg[338]), .Z(n20546) );
  XNOR U22595 ( .A(n20536), .B(n20547), .Z(n20538) );
  XOR U22596 ( .A(n20548), .B(n20549), .Z(n20536) );
  AND U22597 ( .A(n20550), .B(n20551), .Z(n20549) );
  XNOR U22598 ( .A(n20552), .B(n20548), .Z(n20551) );
  XOR U22599 ( .A(n20553), .B(nreg[338]), .Z(n20544) );
  IV U22600 ( .A(n20542), .Z(n20553) );
  XOR U22601 ( .A(n20554), .B(n20555), .Z(n20542) );
  AND U22602 ( .A(n20556), .B(n20557), .Z(n20555) );
  XNOR U22603 ( .A(n20554), .B(n10279), .Z(n20557) );
  XNOR U22604 ( .A(n20550), .B(n20552), .Z(n10279) );
  NAND U22605 ( .A(n20558), .B(nreg[337]), .Z(n20552) );
  NAND U22606 ( .A(n12326), .B(nreg[337]), .Z(n20558) );
  XNOR U22607 ( .A(n20548), .B(n20559), .Z(n20550) );
  XOR U22608 ( .A(n20560), .B(n20561), .Z(n20548) );
  AND U22609 ( .A(n20562), .B(n20563), .Z(n20561) );
  XNOR U22610 ( .A(n20564), .B(n20560), .Z(n20563) );
  XOR U22611 ( .A(n20565), .B(nreg[337]), .Z(n20556) );
  IV U22612 ( .A(n20554), .Z(n20565) );
  XOR U22613 ( .A(n20566), .B(n20567), .Z(n20554) );
  AND U22614 ( .A(n20568), .B(n20569), .Z(n20567) );
  XNOR U22615 ( .A(n20566), .B(n10285), .Z(n20569) );
  XNOR U22616 ( .A(n20562), .B(n20564), .Z(n10285) );
  NAND U22617 ( .A(n20570), .B(nreg[336]), .Z(n20564) );
  NAND U22618 ( .A(n12326), .B(nreg[336]), .Z(n20570) );
  XNOR U22619 ( .A(n20560), .B(n20571), .Z(n20562) );
  XOR U22620 ( .A(n20572), .B(n20573), .Z(n20560) );
  AND U22621 ( .A(n20574), .B(n20575), .Z(n20573) );
  XNOR U22622 ( .A(n20576), .B(n20572), .Z(n20575) );
  XOR U22623 ( .A(n20577), .B(nreg[336]), .Z(n20568) );
  IV U22624 ( .A(n20566), .Z(n20577) );
  XOR U22625 ( .A(n20578), .B(n20579), .Z(n20566) );
  AND U22626 ( .A(n20580), .B(n20581), .Z(n20579) );
  XNOR U22627 ( .A(n20578), .B(n10291), .Z(n20581) );
  XNOR U22628 ( .A(n20574), .B(n20576), .Z(n10291) );
  NAND U22629 ( .A(n20582), .B(nreg[335]), .Z(n20576) );
  NAND U22630 ( .A(n12326), .B(nreg[335]), .Z(n20582) );
  XNOR U22631 ( .A(n20572), .B(n20583), .Z(n20574) );
  XOR U22632 ( .A(n20584), .B(n20585), .Z(n20572) );
  AND U22633 ( .A(n20586), .B(n20587), .Z(n20585) );
  XNOR U22634 ( .A(n20588), .B(n20584), .Z(n20587) );
  XOR U22635 ( .A(n20589), .B(nreg[335]), .Z(n20580) );
  IV U22636 ( .A(n20578), .Z(n20589) );
  XOR U22637 ( .A(n20590), .B(n20591), .Z(n20578) );
  AND U22638 ( .A(n20592), .B(n20593), .Z(n20591) );
  XNOR U22639 ( .A(n20590), .B(n10297), .Z(n20593) );
  XNOR U22640 ( .A(n20586), .B(n20588), .Z(n10297) );
  NAND U22641 ( .A(n20594), .B(nreg[334]), .Z(n20588) );
  NAND U22642 ( .A(n12326), .B(nreg[334]), .Z(n20594) );
  XNOR U22643 ( .A(n20584), .B(n20595), .Z(n20586) );
  XOR U22644 ( .A(n20596), .B(n20597), .Z(n20584) );
  AND U22645 ( .A(n20598), .B(n20599), .Z(n20597) );
  XNOR U22646 ( .A(n20600), .B(n20596), .Z(n20599) );
  XOR U22647 ( .A(n20601), .B(nreg[334]), .Z(n20592) );
  IV U22648 ( .A(n20590), .Z(n20601) );
  XOR U22649 ( .A(n20602), .B(n20603), .Z(n20590) );
  AND U22650 ( .A(n20604), .B(n20605), .Z(n20603) );
  XNOR U22651 ( .A(n20602), .B(n10303), .Z(n20605) );
  XNOR U22652 ( .A(n20598), .B(n20600), .Z(n10303) );
  NAND U22653 ( .A(n20606), .B(nreg[333]), .Z(n20600) );
  NAND U22654 ( .A(n12326), .B(nreg[333]), .Z(n20606) );
  XNOR U22655 ( .A(n20596), .B(n20607), .Z(n20598) );
  XOR U22656 ( .A(n20608), .B(n20609), .Z(n20596) );
  AND U22657 ( .A(n20610), .B(n20611), .Z(n20609) );
  XNOR U22658 ( .A(n20612), .B(n20608), .Z(n20611) );
  XOR U22659 ( .A(n20613), .B(nreg[333]), .Z(n20604) );
  IV U22660 ( .A(n20602), .Z(n20613) );
  XOR U22661 ( .A(n20614), .B(n20615), .Z(n20602) );
  AND U22662 ( .A(n20616), .B(n20617), .Z(n20615) );
  XNOR U22663 ( .A(n20614), .B(n10309), .Z(n20617) );
  XNOR U22664 ( .A(n20610), .B(n20612), .Z(n10309) );
  NAND U22665 ( .A(n20618), .B(nreg[332]), .Z(n20612) );
  NAND U22666 ( .A(n12326), .B(nreg[332]), .Z(n20618) );
  XNOR U22667 ( .A(n20608), .B(n20619), .Z(n20610) );
  XOR U22668 ( .A(n20620), .B(n20621), .Z(n20608) );
  AND U22669 ( .A(n20622), .B(n20623), .Z(n20621) );
  XNOR U22670 ( .A(n20624), .B(n20620), .Z(n20623) );
  XOR U22671 ( .A(n20625), .B(nreg[332]), .Z(n20616) );
  IV U22672 ( .A(n20614), .Z(n20625) );
  XOR U22673 ( .A(n20626), .B(n20627), .Z(n20614) );
  AND U22674 ( .A(n20628), .B(n20629), .Z(n20627) );
  XNOR U22675 ( .A(n20626), .B(n10315), .Z(n20629) );
  XNOR U22676 ( .A(n20622), .B(n20624), .Z(n10315) );
  NAND U22677 ( .A(n20630), .B(nreg[331]), .Z(n20624) );
  NAND U22678 ( .A(n12326), .B(nreg[331]), .Z(n20630) );
  XNOR U22679 ( .A(n20620), .B(n20631), .Z(n20622) );
  XOR U22680 ( .A(n20632), .B(n20633), .Z(n20620) );
  AND U22681 ( .A(n20634), .B(n20635), .Z(n20633) );
  XNOR U22682 ( .A(n20636), .B(n20632), .Z(n20635) );
  XOR U22683 ( .A(n20637), .B(nreg[331]), .Z(n20628) );
  IV U22684 ( .A(n20626), .Z(n20637) );
  XOR U22685 ( .A(n20638), .B(n20639), .Z(n20626) );
  AND U22686 ( .A(n20640), .B(n20641), .Z(n20639) );
  XNOR U22687 ( .A(n20638), .B(n10321), .Z(n20641) );
  XNOR U22688 ( .A(n20634), .B(n20636), .Z(n10321) );
  NAND U22689 ( .A(n20642), .B(nreg[330]), .Z(n20636) );
  NAND U22690 ( .A(n12326), .B(nreg[330]), .Z(n20642) );
  XNOR U22691 ( .A(n20632), .B(n20643), .Z(n20634) );
  XOR U22692 ( .A(n20644), .B(n20645), .Z(n20632) );
  AND U22693 ( .A(n20646), .B(n20647), .Z(n20645) );
  XNOR U22694 ( .A(n20648), .B(n20644), .Z(n20647) );
  XOR U22695 ( .A(n20649), .B(nreg[330]), .Z(n20640) );
  IV U22696 ( .A(n20638), .Z(n20649) );
  XOR U22697 ( .A(n20650), .B(n20651), .Z(n20638) );
  AND U22698 ( .A(n20652), .B(n20653), .Z(n20651) );
  XNOR U22699 ( .A(n20650), .B(n10327), .Z(n20653) );
  XNOR U22700 ( .A(n20646), .B(n20648), .Z(n10327) );
  NAND U22701 ( .A(n20654), .B(nreg[329]), .Z(n20648) );
  NAND U22702 ( .A(n12326), .B(nreg[329]), .Z(n20654) );
  XNOR U22703 ( .A(n20644), .B(n20655), .Z(n20646) );
  XOR U22704 ( .A(n20656), .B(n20657), .Z(n20644) );
  AND U22705 ( .A(n20658), .B(n20659), .Z(n20657) );
  XNOR U22706 ( .A(n20660), .B(n20656), .Z(n20659) );
  XOR U22707 ( .A(n20661), .B(nreg[329]), .Z(n20652) );
  IV U22708 ( .A(n20650), .Z(n20661) );
  XOR U22709 ( .A(n20662), .B(n20663), .Z(n20650) );
  AND U22710 ( .A(n20664), .B(n20665), .Z(n20663) );
  XNOR U22711 ( .A(n20662), .B(n10333), .Z(n20665) );
  XNOR U22712 ( .A(n20658), .B(n20660), .Z(n10333) );
  NAND U22713 ( .A(n20666), .B(nreg[328]), .Z(n20660) );
  NAND U22714 ( .A(n12326), .B(nreg[328]), .Z(n20666) );
  XNOR U22715 ( .A(n20656), .B(n20667), .Z(n20658) );
  XOR U22716 ( .A(n20668), .B(n20669), .Z(n20656) );
  AND U22717 ( .A(n20670), .B(n20671), .Z(n20669) );
  XNOR U22718 ( .A(n20672), .B(n20668), .Z(n20671) );
  XOR U22719 ( .A(n20673), .B(nreg[328]), .Z(n20664) );
  IV U22720 ( .A(n20662), .Z(n20673) );
  XOR U22721 ( .A(n20674), .B(n20675), .Z(n20662) );
  AND U22722 ( .A(n20676), .B(n20677), .Z(n20675) );
  XNOR U22723 ( .A(n20674), .B(n10339), .Z(n20677) );
  XNOR U22724 ( .A(n20670), .B(n20672), .Z(n10339) );
  NAND U22725 ( .A(n20678), .B(nreg[327]), .Z(n20672) );
  NAND U22726 ( .A(n12326), .B(nreg[327]), .Z(n20678) );
  XNOR U22727 ( .A(n20668), .B(n20679), .Z(n20670) );
  XOR U22728 ( .A(n20680), .B(n20681), .Z(n20668) );
  AND U22729 ( .A(n20682), .B(n20683), .Z(n20681) );
  XNOR U22730 ( .A(n20684), .B(n20680), .Z(n20683) );
  XOR U22731 ( .A(n20685), .B(nreg[327]), .Z(n20676) );
  IV U22732 ( .A(n20674), .Z(n20685) );
  XOR U22733 ( .A(n20686), .B(n20687), .Z(n20674) );
  AND U22734 ( .A(n20688), .B(n20689), .Z(n20687) );
  XNOR U22735 ( .A(n20686), .B(n10345), .Z(n20689) );
  XNOR U22736 ( .A(n20682), .B(n20684), .Z(n10345) );
  NAND U22737 ( .A(n20690), .B(nreg[326]), .Z(n20684) );
  NAND U22738 ( .A(n12326), .B(nreg[326]), .Z(n20690) );
  XNOR U22739 ( .A(n20680), .B(n20691), .Z(n20682) );
  XOR U22740 ( .A(n20692), .B(n20693), .Z(n20680) );
  AND U22741 ( .A(n20694), .B(n20695), .Z(n20693) );
  XNOR U22742 ( .A(n20696), .B(n20692), .Z(n20695) );
  XOR U22743 ( .A(n20697), .B(nreg[326]), .Z(n20688) );
  IV U22744 ( .A(n20686), .Z(n20697) );
  XOR U22745 ( .A(n20698), .B(n20699), .Z(n20686) );
  AND U22746 ( .A(n20700), .B(n20701), .Z(n20699) );
  XNOR U22747 ( .A(n20698), .B(n10351), .Z(n20701) );
  XNOR U22748 ( .A(n20694), .B(n20696), .Z(n10351) );
  NAND U22749 ( .A(n20702), .B(nreg[325]), .Z(n20696) );
  NAND U22750 ( .A(n12326), .B(nreg[325]), .Z(n20702) );
  XNOR U22751 ( .A(n20692), .B(n20703), .Z(n20694) );
  XOR U22752 ( .A(n20704), .B(n20705), .Z(n20692) );
  AND U22753 ( .A(n20706), .B(n20707), .Z(n20705) );
  XNOR U22754 ( .A(n20708), .B(n20704), .Z(n20707) );
  XOR U22755 ( .A(n20709), .B(nreg[325]), .Z(n20700) );
  IV U22756 ( .A(n20698), .Z(n20709) );
  XOR U22757 ( .A(n20710), .B(n20711), .Z(n20698) );
  AND U22758 ( .A(n20712), .B(n20713), .Z(n20711) );
  XNOR U22759 ( .A(n20710), .B(n10357), .Z(n20713) );
  XNOR U22760 ( .A(n20706), .B(n20708), .Z(n10357) );
  NAND U22761 ( .A(n20714), .B(nreg[324]), .Z(n20708) );
  NAND U22762 ( .A(n12326), .B(nreg[324]), .Z(n20714) );
  XNOR U22763 ( .A(n20704), .B(n20715), .Z(n20706) );
  XOR U22764 ( .A(n20716), .B(n20717), .Z(n20704) );
  AND U22765 ( .A(n20718), .B(n20719), .Z(n20717) );
  XNOR U22766 ( .A(n20720), .B(n20716), .Z(n20719) );
  XOR U22767 ( .A(n20721), .B(nreg[324]), .Z(n20712) );
  IV U22768 ( .A(n20710), .Z(n20721) );
  XOR U22769 ( .A(n20722), .B(n20723), .Z(n20710) );
  AND U22770 ( .A(n20724), .B(n20725), .Z(n20723) );
  XNOR U22771 ( .A(n20722), .B(n10363), .Z(n20725) );
  XNOR U22772 ( .A(n20718), .B(n20720), .Z(n10363) );
  NAND U22773 ( .A(n20726), .B(nreg[323]), .Z(n20720) );
  NAND U22774 ( .A(n12326), .B(nreg[323]), .Z(n20726) );
  XNOR U22775 ( .A(n20716), .B(n20727), .Z(n20718) );
  XOR U22776 ( .A(n20728), .B(n20729), .Z(n20716) );
  AND U22777 ( .A(n20730), .B(n20731), .Z(n20729) );
  XNOR U22778 ( .A(n20732), .B(n20728), .Z(n20731) );
  XOR U22779 ( .A(n20733), .B(nreg[323]), .Z(n20724) );
  IV U22780 ( .A(n20722), .Z(n20733) );
  XOR U22781 ( .A(n20734), .B(n20735), .Z(n20722) );
  AND U22782 ( .A(n20736), .B(n20737), .Z(n20735) );
  XNOR U22783 ( .A(n20734), .B(n10369), .Z(n20737) );
  XNOR U22784 ( .A(n20730), .B(n20732), .Z(n10369) );
  NAND U22785 ( .A(n20738), .B(nreg[322]), .Z(n20732) );
  NAND U22786 ( .A(n12326), .B(nreg[322]), .Z(n20738) );
  XNOR U22787 ( .A(n20728), .B(n20739), .Z(n20730) );
  XOR U22788 ( .A(n20740), .B(n20741), .Z(n20728) );
  AND U22789 ( .A(n20742), .B(n20743), .Z(n20741) );
  XNOR U22790 ( .A(n20744), .B(n20740), .Z(n20743) );
  XOR U22791 ( .A(n20745), .B(nreg[322]), .Z(n20736) );
  IV U22792 ( .A(n20734), .Z(n20745) );
  XOR U22793 ( .A(n20746), .B(n20747), .Z(n20734) );
  AND U22794 ( .A(n20748), .B(n20749), .Z(n20747) );
  XNOR U22795 ( .A(n20746), .B(n10375), .Z(n20749) );
  XNOR U22796 ( .A(n20742), .B(n20744), .Z(n10375) );
  NAND U22797 ( .A(n20750), .B(nreg[321]), .Z(n20744) );
  NAND U22798 ( .A(n12326), .B(nreg[321]), .Z(n20750) );
  XNOR U22799 ( .A(n20740), .B(n20751), .Z(n20742) );
  XOR U22800 ( .A(n20752), .B(n20753), .Z(n20740) );
  AND U22801 ( .A(n20754), .B(n20755), .Z(n20753) );
  XNOR U22802 ( .A(n20756), .B(n20752), .Z(n20755) );
  XOR U22803 ( .A(n20757), .B(nreg[321]), .Z(n20748) );
  IV U22804 ( .A(n20746), .Z(n20757) );
  XOR U22805 ( .A(n20758), .B(n20759), .Z(n20746) );
  AND U22806 ( .A(n20760), .B(n20761), .Z(n20759) );
  XNOR U22807 ( .A(n20758), .B(n10381), .Z(n20761) );
  XNOR U22808 ( .A(n20754), .B(n20756), .Z(n10381) );
  NAND U22809 ( .A(n20762), .B(nreg[320]), .Z(n20756) );
  NAND U22810 ( .A(n12326), .B(nreg[320]), .Z(n20762) );
  XNOR U22811 ( .A(n20752), .B(n20763), .Z(n20754) );
  XOR U22812 ( .A(n20764), .B(n20765), .Z(n20752) );
  AND U22813 ( .A(n20766), .B(n20767), .Z(n20765) );
  XNOR U22814 ( .A(n20768), .B(n20764), .Z(n20767) );
  XOR U22815 ( .A(n20769), .B(nreg[320]), .Z(n20760) );
  IV U22816 ( .A(n20758), .Z(n20769) );
  XOR U22817 ( .A(n20770), .B(n20771), .Z(n20758) );
  AND U22818 ( .A(n20772), .B(n20773), .Z(n20771) );
  XNOR U22819 ( .A(n20770), .B(n10387), .Z(n20773) );
  XNOR U22820 ( .A(n20766), .B(n20768), .Z(n10387) );
  NAND U22821 ( .A(n20774), .B(nreg[319]), .Z(n20768) );
  NAND U22822 ( .A(n12326), .B(nreg[319]), .Z(n20774) );
  XNOR U22823 ( .A(n20764), .B(n20775), .Z(n20766) );
  XOR U22824 ( .A(n20776), .B(n20777), .Z(n20764) );
  AND U22825 ( .A(n20778), .B(n20779), .Z(n20777) );
  XNOR U22826 ( .A(n20780), .B(n20776), .Z(n20779) );
  XOR U22827 ( .A(n20781), .B(nreg[319]), .Z(n20772) );
  IV U22828 ( .A(n20770), .Z(n20781) );
  XOR U22829 ( .A(n20782), .B(n20783), .Z(n20770) );
  AND U22830 ( .A(n20784), .B(n20785), .Z(n20783) );
  XNOR U22831 ( .A(n20782), .B(n10393), .Z(n20785) );
  XNOR U22832 ( .A(n20778), .B(n20780), .Z(n10393) );
  NAND U22833 ( .A(n20786), .B(nreg[318]), .Z(n20780) );
  NAND U22834 ( .A(n12326), .B(nreg[318]), .Z(n20786) );
  XNOR U22835 ( .A(n20776), .B(n20787), .Z(n20778) );
  XOR U22836 ( .A(n20788), .B(n20789), .Z(n20776) );
  AND U22837 ( .A(n20790), .B(n20791), .Z(n20789) );
  XNOR U22838 ( .A(n20792), .B(n20788), .Z(n20791) );
  XOR U22839 ( .A(n20793), .B(nreg[318]), .Z(n20784) );
  IV U22840 ( .A(n20782), .Z(n20793) );
  XOR U22841 ( .A(n20794), .B(n20795), .Z(n20782) );
  AND U22842 ( .A(n20796), .B(n20797), .Z(n20795) );
  XNOR U22843 ( .A(n20794), .B(n10399), .Z(n20797) );
  XNOR U22844 ( .A(n20790), .B(n20792), .Z(n10399) );
  NAND U22845 ( .A(n20798), .B(nreg[317]), .Z(n20792) );
  NAND U22846 ( .A(n12326), .B(nreg[317]), .Z(n20798) );
  XNOR U22847 ( .A(n20788), .B(n20799), .Z(n20790) );
  XOR U22848 ( .A(n20800), .B(n20801), .Z(n20788) );
  AND U22849 ( .A(n20802), .B(n20803), .Z(n20801) );
  XNOR U22850 ( .A(n20804), .B(n20800), .Z(n20803) );
  XOR U22851 ( .A(n20805), .B(nreg[317]), .Z(n20796) );
  IV U22852 ( .A(n20794), .Z(n20805) );
  XOR U22853 ( .A(n20806), .B(n20807), .Z(n20794) );
  AND U22854 ( .A(n20808), .B(n20809), .Z(n20807) );
  XNOR U22855 ( .A(n20806), .B(n10405), .Z(n20809) );
  XNOR U22856 ( .A(n20802), .B(n20804), .Z(n10405) );
  NAND U22857 ( .A(n20810), .B(nreg[316]), .Z(n20804) );
  NAND U22858 ( .A(n12326), .B(nreg[316]), .Z(n20810) );
  XNOR U22859 ( .A(n20800), .B(n20811), .Z(n20802) );
  XOR U22860 ( .A(n20812), .B(n20813), .Z(n20800) );
  AND U22861 ( .A(n20814), .B(n20815), .Z(n20813) );
  XNOR U22862 ( .A(n20816), .B(n20812), .Z(n20815) );
  XOR U22863 ( .A(n20817), .B(nreg[316]), .Z(n20808) );
  IV U22864 ( .A(n20806), .Z(n20817) );
  XOR U22865 ( .A(n20818), .B(n20819), .Z(n20806) );
  AND U22866 ( .A(n20820), .B(n20821), .Z(n20819) );
  XNOR U22867 ( .A(n20818), .B(n10411), .Z(n20821) );
  XNOR U22868 ( .A(n20814), .B(n20816), .Z(n10411) );
  NAND U22869 ( .A(n20822), .B(nreg[315]), .Z(n20816) );
  NAND U22870 ( .A(n12326), .B(nreg[315]), .Z(n20822) );
  XNOR U22871 ( .A(n20812), .B(n20823), .Z(n20814) );
  XOR U22872 ( .A(n20824), .B(n20825), .Z(n20812) );
  AND U22873 ( .A(n20826), .B(n20827), .Z(n20825) );
  XNOR U22874 ( .A(n20828), .B(n20824), .Z(n20827) );
  XOR U22875 ( .A(n20829), .B(nreg[315]), .Z(n20820) );
  IV U22876 ( .A(n20818), .Z(n20829) );
  XOR U22877 ( .A(n20830), .B(n20831), .Z(n20818) );
  AND U22878 ( .A(n20832), .B(n20833), .Z(n20831) );
  XNOR U22879 ( .A(n20830), .B(n10417), .Z(n20833) );
  XNOR U22880 ( .A(n20826), .B(n20828), .Z(n10417) );
  NAND U22881 ( .A(n20834), .B(nreg[314]), .Z(n20828) );
  NAND U22882 ( .A(n12326), .B(nreg[314]), .Z(n20834) );
  XNOR U22883 ( .A(n20824), .B(n20835), .Z(n20826) );
  XOR U22884 ( .A(n20836), .B(n20837), .Z(n20824) );
  AND U22885 ( .A(n20838), .B(n20839), .Z(n20837) );
  XNOR U22886 ( .A(n20840), .B(n20836), .Z(n20839) );
  XOR U22887 ( .A(n20841), .B(nreg[314]), .Z(n20832) );
  IV U22888 ( .A(n20830), .Z(n20841) );
  XOR U22889 ( .A(n20842), .B(n20843), .Z(n20830) );
  AND U22890 ( .A(n20844), .B(n20845), .Z(n20843) );
  XNOR U22891 ( .A(n20842), .B(n10423), .Z(n20845) );
  XNOR U22892 ( .A(n20838), .B(n20840), .Z(n10423) );
  NAND U22893 ( .A(n20846), .B(nreg[313]), .Z(n20840) );
  NAND U22894 ( .A(n12326), .B(nreg[313]), .Z(n20846) );
  XNOR U22895 ( .A(n20836), .B(n20847), .Z(n20838) );
  XOR U22896 ( .A(n20848), .B(n20849), .Z(n20836) );
  AND U22897 ( .A(n20850), .B(n20851), .Z(n20849) );
  XNOR U22898 ( .A(n20852), .B(n20848), .Z(n20851) );
  XOR U22899 ( .A(n20853), .B(nreg[313]), .Z(n20844) );
  IV U22900 ( .A(n20842), .Z(n20853) );
  XOR U22901 ( .A(n20854), .B(n20855), .Z(n20842) );
  AND U22902 ( .A(n20856), .B(n20857), .Z(n20855) );
  XNOR U22903 ( .A(n20854), .B(n10429), .Z(n20857) );
  XNOR U22904 ( .A(n20850), .B(n20852), .Z(n10429) );
  NAND U22905 ( .A(n20858), .B(nreg[312]), .Z(n20852) );
  NAND U22906 ( .A(n12326), .B(nreg[312]), .Z(n20858) );
  XNOR U22907 ( .A(n20848), .B(n20859), .Z(n20850) );
  XOR U22908 ( .A(n20860), .B(n20861), .Z(n20848) );
  AND U22909 ( .A(n20862), .B(n20863), .Z(n20861) );
  XNOR U22910 ( .A(n20864), .B(n20860), .Z(n20863) );
  XOR U22911 ( .A(n20865), .B(nreg[312]), .Z(n20856) );
  IV U22912 ( .A(n20854), .Z(n20865) );
  XOR U22913 ( .A(n20866), .B(n20867), .Z(n20854) );
  AND U22914 ( .A(n20868), .B(n20869), .Z(n20867) );
  XNOR U22915 ( .A(n20866), .B(n10435), .Z(n20869) );
  XNOR U22916 ( .A(n20862), .B(n20864), .Z(n10435) );
  NAND U22917 ( .A(n20870), .B(nreg[311]), .Z(n20864) );
  NAND U22918 ( .A(n12326), .B(nreg[311]), .Z(n20870) );
  XNOR U22919 ( .A(n20860), .B(n20871), .Z(n20862) );
  XOR U22920 ( .A(n20872), .B(n20873), .Z(n20860) );
  AND U22921 ( .A(n20874), .B(n20875), .Z(n20873) );
  XNOR U22922 ( .A(n20876), .B(n20872), .Z(n20875) );
  XOR U22923 ( .A(n20877), .B(nreg[311]), .Z(n20868) );
  IV U22924 ( .A(n20866), .Z(n20877) );
  XOR U22925 ( .A(n20878), .B(n20879), .Z(n20866) );
  AND U22926 ( .A(n20880), .B(n20881), .Z(n20879) );
  XNOR U22927 ( .A(n20878), .B(n10441), .Z(n20881) );
  XNOR U22928 ( .A(n20874), .B(n20876), .Z(n10441) );
  NAND U22929 ( .A(n20882), .B(nreg[310]), .Z(n20876) );
  NAND U22930 ( .A(n12326), .B(nreg[310]), .Z(n20882) );
  XNOR U22931 ( .A(n20872), .B(n20883), .Z(n20874) );
  XOR U22932 ( .A(n20884), .B(n20885), .Z(n20872) );
  AND U22933 ( .A(n20886), .B(n20887), .Z(n20885) );
  XNOR U22934 ( .A(n20888), .B(n20884), .Z(n20887) );
  XOR U22935 ( .A(n20889), .B(nreg[310]), .Z(n20880) );
  IV U22936 ( .A(n20878), .Z(n20889) );
  XOR U22937 ( .A(n20890), .B(n20891), .Z(n20878) );
  AND U22938 ( .A(n20892), .B(n20893), .Z(n20891) );
  XNOR U22939 ( .A(n20890), .B(n10447), .Z(n20893) );
  XNOR U22940 ( .A(n20886), .B(n20888), .Z(n10447) );
  NAND U22941 ( .A(n20894), .B(nreg[309]), .Z(n20888) );
  NAND U22942 ( .A(n12326), .B(nreg[309]), .Z(n20894) );
  XNOR U22943 ( .A(n20884), .B(n20895), .Z(n20886) );
  XOR U22944 ( .A(n20896), .B(n20897), .Z(n20884) );
  AND U22945 ( .A(n20898), .B(n20899), .Z(n20897) );
  XNOR U22946 ( .A(n20900), .B(n20896), .Z(n20899) );
  XOR U22947 ( .A(n20901), .B(nreg[309]), .Z(n20892) );
  IV U22948 ( .A(n20890), .Z(n20901) );
  XOR U22949 ( .A(n20902), .B(n20903), .Z(n20890) );
  AND U22950 ( .A(n20904), .B(n20905), .Z(n20903) );
  XNOR U22951 ( .A(n20902), .B(n10453), .Z(n20905) );
  XNOR U22952 ( .A(n20898), .B(n20900), .Z(n10453) );
  NAND U22953 ( .A(n20906), .B(nreg[308]), .Z(n20900) );
  NAND U22954 ( .A(n12326), .B(nreg[308]), .Z(n20906) );
  XNOR U22955 ( .A(n20896), .B(n20907), .Z(n20898) );
  XOR U22956 ( .A(n20908), .B(n20909), .Z(n20896) );
  AND U22957 ( .A(n20910), .B(n20911), .Z(n20909) );
  XNOR U22958 ( .A(n20912), .B(n20908), .Z(n20911) );
  XOR U22959 ( .A(n20913), .B(nreg[308]), .Z(n20904) );
  IV U22960 ( .A(n20902), .Z(n20913) );
  XOR U22961 ( .A(n20914), .B(n20915), .Z(n20902) );
  AND U22962 ( .A(n20916), .B(n20917), .Z(n20915) );
  XNOR U22963 ( .A(n20914), .B(n10459), .Z(n20917) );
  XNOR U22964 ( .A(n20910), .B(n20912), .Z(n10459) );
  NAND U22965 ( .A(n20918), .B(nreg[307]), .Z(n20912) );
  NAND U22966 ( .A(n12326), .B(nreg[307]), .Z(n20918) );
  XNOR U22967 ( .A(n20908), .B(n20919), .Z(n20910) );
  XOR U22968 ( .A(n20920), .B(n20921), .Z(n20908) );
  AND U22969 ( .A(n20922), .B(n20923), .Z(n20921) );
  XNOR U22970 ( .A(n20924), .B(n20920), .Z(n20923) );
  XOR U22971 ( .A(n20925), .B(nreg[307]), .Z(n20916) );
  IV U22972 ( .A(n20914), .Z(n20925) );
  XOR U22973 ( .A(n20926), .B(n20927), .Z(n20914) );
  AND U22974 ( .A(n20928), .B(n20929), .Z(n20927) );
  XNOR U22975 ( .A(n20926), .B(n10465), .Z(n20929) );
  XNOR U22976 ( .A(n20922), .B(n20924), .Z(n10465) );
  NAND U22977 ( .A(n20930), .B(nreg[306]), .Z(n20924) );
  NAND U22978 ( .A(n12326), .B(nreg[306]), .Z(n20930) );
  XNOR U22979 ( .A(n20920), .B(n20931), .Z(n20922) );
  XOR U22980 ( .A(n20932), .B(n20933), .Z(n20920) );
  AND U22981 ( .A(n20934), .B(n20935), .Z(n20933) );
  XNOR U22982 ( .A(n20936), .B(n20932), .Z(n20935) );
  XOR U22983 ( .A(n20937), .B(nreg[306]), .Z(n20928) );
  IV U22984 ( .A(n20926), .Z(n20937) );
  XOR U22985 ( .A(n20938), .B(n20939), .Z(n20926) );
  AND U22986 ( .A(n20940), .B(n20941), .Z(n20939) );
  XNOR U22987 ( .A(n20938), .B(n10471), .Z(n20941) );
  XNOR U22988 ( .A(n20934), .B(n20936), .Z(n10471) );
  NAND U22989 ( .A(n20942), .B(nreg[305]), .Z(n20936) );
  NAND U22990 ( .A(n12326), .B(nreg[305]), .Z(n20942) );
  XNOR U22991 ( .A(n20932), .B(n20943), .Z(n20934) );
  XOR U22992 ( .A(n20944), .B(n20945), .Z(n20932) );
  AND U22993 ( .A(n20946), .B(n20947), .Z(n20945) );
  XNOR U22994 ( .A(n20948), .B(n20944), .Z(n20947) );
  XOR U22995 ( .A(n20949), .B(nreg[305]), .Z(n20940) );
  IV U22996 ( .A(n20938), .Z(n20949) );
  XOR U22997 ( .A(n20950), .B(n20951), .Z(n20938) );
  AND U22998 ( .A(n20952), .B(n20953), .Z(n20951) );
  XNOR U22999 ( .A(n20950), .B(n10477), .Z(n20953) );
  XNOR U23000 ( .A(n20946), .B(n20948), .Z(n10477) );
  NAND U23001 ( .A(n20954), .B(nreg[304]), .Z(n20948) );
  NAND U23002 ( .A(n12326), .B(nreg[304]), .Z(n20954) );
  XNOR U23003 ( .A(n20944), .B(n20955), .Z(n20946) );
  XOR U23004 ( .A(n20956), .B(n20957), .Z(n20944) );
  AND U23005 ( .A(n20958), .B(n20959), .Z(n20957) );
  XNOR U23006 ( .A(n20960), .B(n20956), .Z(n20959) );
  XOR U23007 ( .A(n20961), .B(nreg[304]), .Z(n20952) );
  IV U23008 ( .A(n20950), .Z(n20961) );
  XOR U23009 ( .A(n20962), .B(n20963), .Z(n20950) );
  AND U23010 ( .A(n20964), .B(n20965), .Z(n20963) );
  XNOR U23011 ( .A(n20962), .B(n10483), .Z(n20965) );
  XNOR U23012 ( .A(n20958), .B(n20960), .Z(n10483) );
  NAND U23013 ( .A(n20966), .B(nreg[303]), .Z(n20960) );
  NAND U23014 ( .A(n12326), .B(nreg[303]), .Z(n20966) );
  XNOR U23015 ( .A(n20956), .B(n20967), .Z(n20958) );
  XOR U23016 ( .A(n20968), .B(n20969), .Z(n20956) );
  AND U23017 ( .A(n20970), .B(n20971), .Z(n20969) );
  XNOR U23018 ( .A(n20972), .B(n20968), .Z(n20971) );
  XOR U23019 ( .A(n20973), .B(nreg[303]), .Z(n20964) );
  IV U23020 ( .A(n20962), .Z(n20973) );
  XOR U23021 ( .A(n20974), .B(n20975), .Z(n20962) );
  AND U23022 ( .A(n20976), .B(n20977), .Z(n20975) );
  XNOR U23023 ( .A(n20974), .B(n10489), .Z(n20977) );
  XNOR U23024 ( .A(n20970), .B(n20972), .Z(n10489) );
  NAND U23025 ( .A(n20978), .B(nreg[302]), .Z(n20972) );
  NAND U23026 ( .A(n12326), .B(nreg[302]), .Z(n20978) );
  XNOR U23027 ( .A(n20968), .B(n20979), .Z(n20970) );
  XOR U23028 ( .A(n20980), .B(n20981), .Z(n20968) );
  AND U23029 ( .A(n20982), .B(n20983), .Z(n20981) );
  XNOR U23030 ( .A(n20984), .B(n20980), .Z(n20983) );
  XOR U23031 ( .A(n20985), .B(nreg[302]), .Z(n20976) );
  IV U23032 ( .A(n20974), .Z(n20985) );
  XOR U23033 ( .A(n20986), .B(n20987), .Z(n20974) );
  AND U23034 ( .A(n20988), .B(n20989), .Z(n20987) );
  XNOR U23035 ( .A(n20986), .B(n10495), .Z(n20989) );
  XNOR U23036 ( .A(n20982), .B(n20984), .Z(n10495) );
  NAND U23037 ( .A(n20990), .B(nreg[301]), .Z(n20984) );
  NAND U23038 ( .A(n12326), .B(nreg[301]), .Z(n20990) );
  XNOR U23039 ( .A(n20980), .B(n20991), .Z(n20982) );
  XOR U23040 ( .A(n20992), .B(n20993), .Z(n20980) );
  AND U23041 ( .A(n20994), .B(n20995), .Z(n20993) );
  XNOR U23042 ( .A(n20996), .B(n20992), .Z(n20995) );
  XOR U23043 ( .A(n20997), .B(nreg[301]), .Z(n20988) );
  IV U23044 ( .A(n20986), .Z(n20997) );
  XOR U23045 ( .A(n20998), .B(n20999), .Z(n20986) );
  AND U23046 ( .A(n21000), .B(n21001), .Z(n20999) );
  XNOR U23047 ( .A(n20998), .B(n10501), .Z(n21001) );
  XNOR U23048 ( .A(n20994), .B(n20996), .Z(n10501) );
  NAND U23049 ( .A(n21002), .B(nreg[300]), .Z(n20996) );
  NAND U23050 ( .A(n12326), .B(nreg[300]), .Z(n21002) );
  XNOR U23051 ( .A(n20992), .B(n21003), .Z(n20994) );
  XOR U23052 ( .A(n21004), .B(n21005), .Z(n20992) );
  AND U23053 ( .A(n21006), .B(n21007), .Z(n21005) );
  XNOR U23054 ( .A(n21008), .B(n21004), .Z(n21007) );
  XOR U23055 ( .A(n21009), .B(nreg[300]), .Z(n21000) );
  IV U23056 ( .A(n20998), .Z(n21009) );
  XOR U23057 ( .A(n21010), .B(n21011), .Z(n20998) );
  AND U23058 ( .A(n21012), .B(n21013), .Z(n21011) );
  XNOR U23059 ( .A(n21010), .B(n10507), .Z(n21013) );
  XNOR U23060 ( .A(n21006), .B(n21008), .Z(n10507) );
  NAND U23061 ( .A(n21014), .B(nreg[299]), .Z(n21008) );
  NAND U23062 ( .A(n12326), .B(nreg[299]), .Z(n21014) );
  XNOR U23063 ( .A(n21004), .B(n21015), .Z(n21006) );
  XOR U23064 ( .A(n21016), .B(n21017), .Z(n21004) );
  AND U23065 ( .A(n21018), .B(n21019), .Z(n21017) );
  XNOR U23066 ( .A(n21020), .B(n21016), .Z(n21019) );
  XOR U23067 ( .A(n21021), .B(nreg[299]), .Z(n21012) );
  IV U23068 ( .A(n21010), .Z(n21021) );
  XOR U23069 ( .A(n21022), .B(n21023), .Z(n21010) );
  AND U23070 ( .A(n21024), .B(n21025), .Z(n21023) );
  XNOR U23071 ( .A(n21022), .B(n10513), .Z(n21025) );
  XNOR U23072 ( .A(n21018), .B(n21020), .Z(n10513) );
  NAND U23073 ( .A(n21026), .B(nreg[298]), .Z(n21020) );
  NAND U23074 ( .A(n12326), .B(nreg[298]), .Z(n21026) );
  XNOR U23075 ( .A(n21016), .B(n21027), .Z(n21018) );
  XOR U23076 ( .A(n21028), .B(n21029), .Z(n21016) );
  AND U23077 ( .A(n21030), .B(n21031), .Z(n21029) );
  XNOR U23078 ( .A(n21032), .B(n21028), .Z(n21031) );
  XOR U23079 ( .A(n21033), .B(nreg[298]), .Z(n21024) );
  IV U23080 ( .A(n21022), .Z(n21033) );
  XOR U23081 ( .A(n21034), .B(n21035), .Z(n21022) );
  AND U23082 ( .A(n21036), .B(n21037), .Z(n21035) );
  XNOR U23083 ( .A(n21034), .B(n10519), .Z(n21037) );
  XNOR U23084 ( .A(n21030), .B(n21032), .Z(n10519) );
  NAND U23085 ( .A(n21038), .B(nreg[297]), .Z(n21032) );
  NAND U23086 ( .A(n12326), .B(nreg[297]), .Z(n21038) );
  XNOR U23087 ( .A(n21028), .B(n21039), .Z(n21030) );
  XOR U23088 ( .A(n21040), .B(n21041), .Z(n21028) );
  AND U23089 ( .A(n21042), .B(n21043), .Z(n21041) );
  XNOR U23090 ( .A(n21044), .B(n21040), .Z(n21043) );
  XOR U23091 ( .A(n21045), .B(nreg[297]), .Z(n21036) );
  IV U23092 ( .A(n21034), .Z(n21045) );
  XOR U23093 ( .A(n21046), .B(n21047), .Z(n21034) );
  AND U23094 ( .A(n21048), .B(n21049), .Z(n21047) );
  XNOR U23095 ( .A(n21046), .B(n10525), .Z(n21049) );
  XNOR U23096 ( .A(n21042), .B(n21044), .Z(n10525) );
  NAND U23097 ( .A(n21050), .B(nreg[296]), .Z(n21044) );
  NAND U23098 ( .A(n12326), .B(nreg[296]), .Z(n21050) );
  XNOR U23099 ( .A(n21040), .B(n21051), .Z(n21042) );
  XOR U23100 ( .A(n21052), .B(n21053), .Z(n21040) );
  AND U23101 ( .A(n21054), .B(n21055), .Z(n21053) );
  XNOR U23102 ( .A(n21056), .B(n21052), .Z(n21055) );
  XOR U23103 ( .A(n21057), .B(nreg[296]), .Z(n21048) );
  IV U23104 ( .A(n21046), .Z(n21057) );
  XOR U23105 ( .A(n21058), .B(n21059), .Z(n21046) );
  AND U23106 ( .A(n21060), .B(n21061), .Z(n21059) );
  XNOR U23107 ( .A(n21058), .B(n10531), .Z(n21061) );
  XNOR U23108 ( .A(n21054), .B(n21056), .Z(n10531) );
  NAND U23109 ( .A(n21062), .B(nreg[295]), .Z(n21056) );
  NAND U23110 ( .A(n12326), .B(nreg[295]), .Z(n21062) );
  XNOR U23111 ( .A(n21052), .B(n21063), .Z(n21054) );
  XOR U23112 ( .A(n21064), .B(n21065), .Z(n21052) );
  AND U23113 ( .A(n21066), .B(n21067), .Z(n21065) );
  XNOR U23114 ( .A(n21068), .B(n21064), .Z(n21067) );
  XOR U23115 ( .A(n21069), .B(nreg[295]), .Z(n21060) );
  IV U23116 ( .A(n21058), .Z(n21069) );
  XOR U23117 ( .A(n21070), .B(n21071), .Z(n21058) );
  AND U23118 ( .A(n21072), .B(n21073), .Z(n21071) );
  XNOR U23119 ( .A(n21070), .B(n10537), .Z(n21073) );
  XNOR U23120 ( .A(n21066), .B(n21068), .Z(n10537) );
  NAND U23121 ( .A(n21074), .B(nreg[294]), .Z(n21068) );
  NAND U23122 ( .A(n12326), .B(nreg[294]), .Z(n21074) );
  XNOR U23123 ( .A(n21064), .B(n21075), .Z(n21066) );
  XOR U23124 ( .A(n21076), .B(n21077), .Z(n21064) );
  AND U23125 ( .A(n21078), .B(n21079), .Z(n21077) );
  XNOR U23126 ( .A(n21080), .B(n21076), .Z(n21079) );
  XOR U23127 ( .A(n21081), .B(nreg[294]), .Z(n21072) );
  IV U23128 ( .A(n21070), .Z(n21081) );
  XOR U23129 ( .A(n21082), .B(n21083), .Z(n21070) );
  AND U23130 ( .A(n21084), .B(n21085), .Z(n21083) );
  XNOR U23131 ( .A(n21082), .B(n10543), .Z(n21085) );
  XNOR U23132 ( .A(n21078), .B(n21080), .Z(n10543) );
  NAND U23133 ( .A(n21086), .B(nreg[293]), .Z(n21080) );
  NAND U23134 ( .A(n12326), .B(nreg[293]), .Z(n21086) );
  XNOR U23135 ( .A(n21076), .B(n21087), .Z(n21078) );
  XOR U23136 ( .A(n21088), .B(n21089), .Z(n21076) );
  AND U23137 ( .A(n21090), .B(n21091), .Z(n21089) );
  XNOR U23138 ( .A(n21092), .B(n21088), .Z(n21091) );
  XOR U23139 ( .A(n21093), .B(nreg[293]), .Z(n21084) );
  IV U23140 ( .A(n21082), .Z(n21093) );
  XOR U23141 ( .A(n21094), .B(n21095), .Z(n21082) );
  AND U23142 ( .A(n21096), .B(n21097), .Z(n21095) );
  XNOR U23143 ( .A(n21094), .B(n10549), .Z(n21097) );
  XNOR U23144 ( .A(n21090), .B(n21092), .Z(n10549) );
  NAND U23145 ( .A(n21098), .B(nreg[292]), .Z(n21092) );
  NAND U23146 ( .A(n12326), .B(nreg[292]), .Z(n21098) );
  XNOR U23147 ( .A(n21088), .B(n21099), .Z(n21090) );
  XOR U23148 ( .A(n21100), .B(n21101), .Z(n21088) );
  AND U23149 ( .A(n21102), .B(n21103), .Z(n21101) );
  XNOR U23150 ( .A(n21104), .B(n21100), .Z(n21103) );
  XOR U23151 ( .A(n21105), .B(nreg[292]), .Z(n21096) );
  IV U23152 ( .A(n21094), .Z(n21105) );
  XOR U23153 ( .A(n21106), .B(n21107), .Z(n21094) );
  AND U23154 ( .A(n21108), .B(n21109), .Z(n21107) );
  XNOR U23155 ( .A(n21106), .B(n10555), .Z(n21109) );
  XNOR U23156 ( .A(n21102), .B(n21104), .Z(n10555) );
  NAND U23157 ( .A(n21110), .B(nreg[291]), .Z(n21104) );
  NAND U23158 ( .A(n12326), .B(nreg[291]), .Z(n21110) );
  XNOR U23159 ( .A(n21100), .B(n21111), .Z(n21102) );
  XOR U23160 ( .A(n21112), .B(n21113), .Z(n21100) );
  AND U23161 ( .A(n21114), .B(n21115), .Z(n21113) );
  XNOR U23162 ( .A(n21116), .B(n21112), .Z(n21115) );
  XOR U23163 ( .A(n21117), .B(nreg[291]), .Z(n21108) );
  IV U23164 ( .A(n21106), .Z(n21117) );
  XOR U23165 ( .A(n21118), .B(n21119), .Z(n21106) );
  AND U23166 ( .A(n21120), .B(n21121), .Z(n21119) );
  XNOR U23167 ( .A(n21118), .B(n10561), .Z(n21121) );
  XNOR U23168 ( .A(n21114), .B(n21116), .Z(n10561) );
  NAND U23169 ( .A(n21122), .B(nreg[290]), .Z(n21116) );
  NAND U23170 ( .A(n12326), .B(nreg[290]), .Z(n21122) );
  XNOR U23171 ( .A(n21112), .B(n21123), .Z(n21114) );
  XOR U23172 ( .A(n21124), .B(n21125), .Z(n21112) );
  AND U23173 ( .A(n21126), .B(n21127), .Z(n21125) );
  XNOR U23174 ( .A(n21128), .B(n21124), .Z(n21127) );
  XOR U23175 ( .A(n21129), .B(nreg[290]), .Z(n21120) );
  IV U23176 ( .A(n21118), .Z(n21129) );
  XOR U23177 ( .A(n21130), .B(n21131), .Z(n21118) );
  AND U23178 ( .A(n21132), .B(n21133), .Z(n21131) );
  XNOR U23179 ( .A(n21130), .B(n10567), .Z(n21133) );
  XNOR U23180 ( .A(n21126), .B(n21128), .Z(n10567) );
  NAND U23181 ( .A(n21134), .B(nreg[289]), .Z(n21128) );
  NAND U23182 ( .A(n12326), .B(nreg[289]), .Z(n21134) );
  XNOR U23183 ( .A(n21124), .B(n21135), .Z(n21126) );
  XOR U23184 ( .A(n21136), .B(n21137), .Z(n21124) );
  AND U23185 ( .A(n21138), .B(n21139), .Z(n21137) );
  XNOR U23186 ( .A(n21140), .B(n21136), .Z(n21139) );
  XOR U23187 ( .A(n21141), .B(nreg[289]), .Z(n21132) );
  IV U23188 ( .A(n21130), .Z(n21141) );
  XOR U23189 ( .A(n21142), .B(n21143), .Z(n21130) );
  AND U23190 ( .A(n21144), .B(n21145), .Z(n21143) );
  XNOR U23191 ( .A(n21142), .B(n10573), .Z(n21145) );
  XNOR U23192 ( .A(n21138), .B(n21140), .Z(n10573) );
  NAND U23193 ( .A(n21146), .B(nreg[288]), .Z(n21140) );
  NAND U23194 ( .A(n12326), .B(nreg[288]), .Z(n21146) );
  XNOR U23195 ( .A(n21136), .B(n21147), .Z(n21138) );
  XOR U23196 ( .A(n21148), .B(n21149), .Z(n21136) );
  AND U23197 ( .A(n21150), .B(n21151), .Z(n21149) );
  XNOR U23198 ( .A(n21152), .B(n21148), .Z(n21151) );
  XOR U23199 ( .A(n21153), .B(nreg[288]), .Z(n21144) );
  IV U23200 ( .A(n21142), .Z(n21153) );
  XOR U23201 ( .A(n21154), .B(n21155), .Z(n21142) );
  AND U23202 ( .A(n21156), .B(n21157), .Z(n21155) );
  XNOR U23203 ( .A(n21154), .B(n10579), .Z(n21157) );
  XNOR U23204 ( .A(n21150), .B(n21152), .Z(n10579) );
  NAND U23205 ( .A(n21158), .B(nreg[287]), .Z(n21152) );
  NAND U23206 ( .A(n12326), .B(nreg[287]), .Z(n21158) );
  XNOR U23207 ( .A(n21148), .B(n21159), .Z(n21150) );
  XOR U23208 ( .A(n21160), .B(n21161), .Z(n21148) );
  AND U23209 ( .A(n21162), .B(n21163), .Z(n21161) );
  XNOR U23210 ( .A(n21164), .B(n21160), .Z(n21163) );
  XOR U23211 ( .A(n21165), .B(nreg[287]), .Z(n21156) );
  IV U23212 ( .A(n21154), .Z(n21165) );
  XOR U23213 ( .A(n21166), .B(n21167), .Z(n21154) );
  AND U23214 ( .A(n21168), .B(n21169), .Z(n21167) );
  XNOR U23215 ( .A(n21166), .B(n10585), .Z(n21169) );
  XNOR U23216 ( .A(n21162), .B(n21164), .Z(n10585) );
  NAND U23217 ( .A(n21170), .B(nreg[286]), .Z(n21164) );
  NAND U23218 ( .A(n12326), .B(nreg[286]), .Z(n21170) );
  XNOR U23219 ( .A(n21160), .B(n21171), .Z(n21162) );
  XOR U23220 ( .A(n21172), .B(n21173), .Z(n21160) );
  AND U23221 ( .A(n21174), .B(n21175), .Z(n21173) );
  XNOR U23222 ( .A(n21176), .B(n21172), .Z(n21175) );
  XOR U23223 ( .A(n21177), .B(nreg[286]), .Z(n21168) );
  IV U23224 ( .A(n21166), .Z(n21177) );
  XOR U23225 ( .A(n21178), .B(n21179), .Z(n21166) );
  AND U23226 ( .A(n21180), .B(n21181), .Z(n21179) );
  XNOR U23227 ( .A(n21178), .B(n10591), .Z(n21181) );
  XNOR U23228 ( .A(n21174), .B(n21176), .Z(n10591) );
  NAND U23229 ( .A(n21182), .B(nreg[285]), .Z(n21176) );
  NAND U23230 ( .A(n12326), .B(nreg[285]), .Z(n21182) );
  XNOR U23231 ( .A(n21172), .B(n21183), .Z(n21174) );
  XOR U23232 ( .A(n21184), .B(n21185), .Z(n21172) );
  AND U23233 ( .A(n21186), .B(n21187), .Z(n21185) );
  XNOR U23234 ( .A(n21188), .B(n21184), .Z(n21187) );
  XOR U23235 ( .A(n21189), .B(nreg[285]), .Z(n21180) );
  IV U23236 ( .A(n21178), .Z(n21189) );
  XOR U23237 ( .A(n21190), .B(n21191), .Z(n21178) );
  AND U23238 ( .A(n21192), .B(n21193), .Z(n21191) );
  XNOR U23239 ( .A(n21190), .B(n10597), .Z(n21193) );
  XNOR U23240 ( .A(n21186), .B(n21188), .Z(n10597) );
  NAND U23241 ( .A(n21194), .B(nreg[284]), .Z(n21188) );
  NAND U23242 ( .A(n12326), .B(nreg[284]), .Z(n21194) );
  XNOR U23243 ( .A(n21184), .B(n21195), .Z(n21186) );
  XOR U23244 ( .A(n21196), .B(n21197), .Z(n21184) );
  AND U23245 ( .A(n21198), .B(n21199), .Z(n21197) );
  XNOR U23246 ( .A(n21200), .B(n21196), .Z(n21199) );
  XOR U23247 ( .A(n21201), .B(nreg[284]), .Z(n21192) );
  IV U23248 ( .A(n21190), .Z(n21201) );
  XOR U23249 ( .A(n21202), .B(n21203), .Z(n21190) );
  AND U23250 ( .A(n21204), .B(n21205), .Z(n21203) );
  XNOR U23251 ( .A(n21202), .B(n10603), .Z(n21205) );
  XNOR U23252 ( .A(n21198), .B(n21200), .Z(n10603) );
  NAND U23253 ( .A(n21206), .B(nreg[283]), .Z(n21200) );
  NAND U23254 ( .A(n12326), .B(nreg[283]), .Z(n21206) );
  XNOR U23255 ( .A(n21196), .B(n21207), .Z(n21198) );
  XOR U23256 ( .A(n21208), .B(n21209), .Z(n21196) );
  AND U23257 ( .A(n21210), .B(n21211), .Z(n21209) );
  XNOR U23258 ( .A(n21212), .B(n21208), .Z(n21211) );
  XOR U23259 ( .A(n21213), .B(nreg[283]), .Z(n21204) );
  IV U23260 ( .A(n21202), .Z(n21213) );
  XOR U23261 ( .A(n21214), .B(n21215), .Z(n21202) );
  AND U23262 ( .A(n21216), .B(n21217), .Z(n21215) );
  XNOR U23263 ( .A(n21214), .B(n10609), .Z(n21217) );
  XNOR U23264 ( .A(n21210), .B(n21212), .Z(n10609) );
  NAND U23265 ( .A(n21218), .B(nreg[282]), .Z(n21212) );
  NAND U23266 ( .A(n12326), .B(nreg[282]), .Z(n21218) );
  XNOR U23267 ( .A(n21208), .B(n21219), .Z(n21210) );
  XOR U23268 ( .A(n21220), .B(n21221), .Z(n21208) );
  AND U23269 ( .A(n21222), .B(n21223), .Z(n21221) );
  XNOR U23270 ( .A(n21224), .B(n21220), .Z(n21223) );
  XOR U23271 ( .A(n21225), .B(nreg[282]), .Z(n21216) );
  IV U23272 ( .A(n21214), .Z(n21225) );
  XOR U23273 ( .A(n21226), .B(n21227), .Z(n21214) );
  AND U23274 ( .A(n21228), .B(n21229), .Z(n21227) );
  XNOR U23275 ( .A(n21226), .B(n10615), .Z(n21229) );
  XNOR U23276 ( .A(n21222), .B(n21224), .Z(n10615) );
  NAND U23277 ( .A(n21230), .B(nreg[281]), .Z(n21224) );
  NAND U23278 ( .A(n12326), .B(nreg[281]), .Z(n21230) );
  XNOR U23279 ( .A(n21220), .B(n21231), .Z(n21222) );
  XOR U23280 ( .A(n21232), .B(n21233), .Z(n21220) );
  AND U23281 ( .A(n21234), .B(n21235), .Z(n21233) );
  XNOR U23282 ( .A(n21236), .B(n21232), .Z(n21235) );
  XOR U23283 ( .A(n21237), .B(nreg[281]), .Z(n21228) );
  IV U23284 ( .A(n21226), .Z(n21237) );
  XOR U23285 ( .A(n21238), .B(n21239), .Z(n21226) );
  AND U23286 ( .A(n21240), .B(n21241), .Z(n21239) );
  XNOR U23287 ( .A(n21238), .B(n10621), .Z(n21241) );
  XNOR U23288 ( .A(n21234), .B(n21236), .Z(n10621) );
  NAND U23289 ( .A(n21242), .B(nreg[280]), .Z(n21236) );
  NAND U23290 ( .A(n12326), .B(nreg[280]), .Z(n21242) );
  XNOR U23291 ( .A(n21232), .B(n21243), .Z(n21234) );
  XOR U23292 ( .A(n21244), .B(n21245), .Z(n21232) );
  AND U23293 ( .A(n21246), .B(n21247), .Z(n21245) );
  XNOR U23294 ( .A(n21248), .B(n21244), .Z(n21247) );
  XOR U23295 ( .A(n21249), .B(nreg[280]), .Z(n21240) );
  IV U23296 ( .A(n21238), .Z(n21249) );
  XOR U23297 ( .A(n21250), .B(n21251), .Z(n21238) );
  AND U23298 ( .A(n21252), .B(n21253), .Z(n21251) );
  XNOR U23299 ( .A(n21250), .B(n10627), .Z(n21253) );
  XNOR U23300 ( .A(n21246), .B(n21248), .Z(n10627) );
  NAND U23301 ( .A(n21254), .B(nreg[279]), .Z(n21248) );
  NAND U23302 ( .A(n12326), .B(nreg[279]), .Z(n21254) );
  XNOR U23303 ( .A(n21244), .B(n21255), .Z(n21246) );
  XOR U23304 ( .A(n21256), .B(n21257), .Z(n21244) );
  AND U23305 ( .A(n21258), .B(n21259), .Z(n21257) );
  XNOR U23306 ( .A(n21260), .B(n21256), .Z(n21259) );
  XOR U23307 ( .A(n21261), .B(nreg[279]), .Z(n21252) );
  IV U23308 ( .A(n21250), .Z(n21261) );
  XOR U23309 ( .A(n21262), .B(n21263), .Z(n21250) );
  AND U23310 ( .A(n21264), .B(n21265), .Z(n21263) );
  XNOR U23311 ( .A(n21262), .B(n10633), .Z(n21265) );
  XNOR U23312 ( .A(n21258), .B(n21260), .Z(n10633) );
  NAND U23313 ( .A(n21266), .B(nreg[278]), .Z(n21260) );
  NAND U23314 ( .A(n12326), .B(nreg[278]), .Z(n21266) );
  XNOR U23315 ( .A(n21256), .B(n21267), .Z(n21258) );
  XOR U23316 ( .A(n21268), .B(n21269), .Z(n21256) );
  AND U23317 ( .A(n21270), .B(n21271), .Z(n21269) );
  XNOR U23318 ( .A(n21272), .B(n21268), .Z(n21271) );
  XOR U23319 ( .A(n21273), .B(nreg[278]), .Z(n21264) );
  IV U23320 ( .A(n21262), .Z(n21273) );
  XOR U23321 ( .A(n21274), .B(n21275), .Z(n21262) );
  AND U23322 ( .A(n21276), .B(n21277), .Z(n21275) );
  XNOR U23323 ( .A(n21274), .B(n10639), .Z(n21277) );
  XNOR U23324 ( .A(n21270), .B(n21272), .Z(n10639) );
  NAND U23325 ( .A(n21278), .B(nreg[277]), .Z(n21272) );
  NAND U23326 ( .A(n12326), .B(nreg[277]), .Z(n21278) );
  XNOR U23327 ( .A(n21268), .B(n21279), .Z(n21270) );
  XOR U23328 ( .A(n21280), .B(n21281), .Z(n21268) );
  AND U23329 ( .A(n21282), .B(n21283), .Z(n21281) );
  XNOR U23330 ( .A(n21284), .B(n21280), .Z(n21283) );
  XOR U23331 ( .A(n21285), .B(nreg[277]), .Z(n21276) );
  IV U23332 ( .A(n21274), .Z(n21285) );
  XOR U23333 ( .A(n21286), .B(n21287), .Z(n21274) );
  AND U23334 ( .A(n21288), .B(n21289), .Z(n21287) );
  XNOR U23335 ( .A(n21286), .B(n10645), .Z(n21289) );
  XNOR U23336 ( .A(n21282), .B(n21284), .Z(n10645) );
  NAND U23337 ( .A(n21290), .B(nreg[276]), .Z(n21284) );
  NAND U23338 ( .A(n12326), .B(nreg[276]), .Z(n21290) );
  XNOR U23339 ( .A(n21280), .B(n21291), .Z(n21282) );
  XOR U23340 ( .A(n21292), .B(n21293), .Z(n21280) );
  AND U23341 ( .A(n21294), .B(n21295), .Z(n21293) );
  XNOR U23342 ( .A(n21296), .B(n21292), .Z(n21295) );
  XOR U23343 ( .A(n21297), .B(nreg[276]), .Z(n21288) );
  IV U23344 ( .A(n21286), .Z(n21297) );
  XOR U23345 ( .A(n21298), .B(n21299), .Z(n21286) );
  AND U23346 ( .A(n21300), .B(n21301), .Z(n21299) );
  XNOR U23347 ( .A(n21298), .B(n10651), .Z(n21301) );
  XNOR U23348 ( .A(n21294), .B(n21296), .Z(n10651) );
  NAND U23349 ( .A(n21302), .B(nreg[275]), .Z(n21296) );
  NAND U23350 ( .A(n12326), .B(nreg[275]), .Z(n21302) );
  XNOR U23351 ( .A(n21292), .B(n21303), .Z(n21294) );
  XOR U23352 ( .A(n21304), .B(n21305), .Z(n21292) );
  AND U23353 ( .A(n21306), .B(n21307), .Z(n21305) );
  XNOR U23354 ( .A(n21308), .B(n21304), .Z(n21307) );
  XOR U23355 ( .A(n21309), .B(nreg[275]), .Z(n21300) );
  IV U23356 ( .A(n21298), .Z(n21309) );
  XOR U23357 ( .A(n21310), .B(n21311), .Z(n21298) );
  AND U23358 ( .A(n21312), .B(n21313), .Z(n21311) );
  XNOR U23359 ( .A(n21310), .B(n10657), .Z(n21313) );
  XNOR U23360 ( .A(n21306), .B(n21308), .Z(n10657) );
  NAND U23361 ( .A(n21314), .B(nreg[274]), .Z(n21308) );
  NAND U23362 ( .A(n12326), .B(nreg[274]), .Z(n21314) );
  XNOR U23363 ( .A(n21304), .B(n21315), .Z(n21306) );
  XOR U23364 ( .A(n21316), .B(n21317), .Z(n21304) );
  AND U23365 ( .A(n21318), .B(n21319), .Z(n21317) );
  XNOR U23366 ( .A(n21320), .B(n21316), .Z(n21319) );
  XOR U23367 ( .A(n21321), .B(nreg[274]), .Z(n21312) );
  IV U23368 ( .A(n21310), .Z(n21321) );
  XOR U23369 ( .A(n21322), .B(n21323), .Z(n21310) );
  AND U23370 ( .A(n21324), .B(n21325), .Z(n21323) );
  XNOR U23371 ( .A(n21322), .B(n10663), .Z(n21325) );
  XNOR U23372 ( .A(n21318), .B(n21320), .Z(n10663) );
  NAND U23373 ( .A(n21326), .B(nreg[273]), .Z(n21320) );
  NAND U23374 ( .A(n12326), .B(nreg[273]), .Z(n21326) );
  XNOR U23375 ( .A(n21316), .B(n21327), .Z(n21318) );
  XOR U23376 ( .A(n21328), .B(n21329), .Z(n21316) );
  AND U23377 ( .A(n21330), .B(n21331), .Z(n21329) );
  XNOR U23378 ( .A(n21332), .B(n21328), .Z(n21331) );
  XOR U23379 ( .A(n21333), .B(nreg[273]), .Z(n21324) );
  IV U23380 ( .A(n21322), .Z(n21333) );
  XOR U23381 ( .A(n21334), .B(n21335), .Z(n21322) );
  AND U23382 ( .A(n21336), .B(n21337), .Z(n21335) );
  XNOR U23383 ( .A(n21334), .B(n10669), .Z(n21337) );
  XNOR U23384 ( .A(n21330), .B(n21332), .Z(n10669) );
  NAND U23385 ( .A(n21338), .B(nreg[272]), .Z(n21332) );
  NAND U23386 ( .A(n12326), .B(nreg[272]), .Z(n21338) );
  XNOR U23387 ( .A(n21328), .B(n21339), .Z(n21330) );
  XOR U23388 ( .A(n21340), .B(n21341), .Z(n21328) );
  AND U23389 ( .A(n21342), .B(n21343), .Z(n21341) );
  XNOR U23390 ( .A(n21344), .B(n21340), .Z(n21343) );
  XOR U23391 ( .A(n21345), .B(nreg[272]), .Z(n21336) );
  IV U23392 ( .A(n21334), .Z(n21345) );
  XOR U23393 ( .A(n21346), .B(n21347), .Z(n21334) );
  AND U23394 ( .A(n21348), .B(n21349), .Z(n21347) );
  XNOR U23395 ( .A(n21346), .B(n10675), .Z(n21349) );
  XNOR U23396 ( .A(n21342), .B(n21344), .Z(n10675) );
  NAND U23397 ( .A(n21350), .B(nreg[271]), .Z(n21344) );
  NAND U23398 ( .A(n12326), .B(nreg[271]), .Z(n21350) );
  XNOR U23399 ( .A(n21340), .B(n21351), .Z(n21342) );
  XOR U23400 ( .A(n21352), .B(n21353), .Z(n21340) );
  AND U23401 ( .A(n21354), .B(n21355), .Z(n21353) );
  XNOR U23402 ( .A(n21356), .B(n21352), .Z(n21355) );
  XOR U23403 ( .A(n21357), .B(nreg[271]), .Z(n21348) );
  IV U23404 ( .A(n21346), .Z(n21357) );
  XOR U23405 ( .A(n21358), .B(n21359), .Z(n21346) );
  AND U23406 ( .A(n21360), .B(n21361), .Z(n21359) );
  XNOR U23407 ( .A(n21358), .B(n10681), .Z(n21361) );
  XNOR U23408 ( .A(n21354), .B(n21356), .Z(n10681) );
  NAND U23409 ( .A(n21362), .B(nreg[270]), .Z(n21356) );
  NAND U23410 ( .A(n12326), .B(nreg[270]), .Z(n21362) );
  XNOR U23411 ( .A(n21352), .B(n21363), .Z(n21354) );
  XOR U23412 ( .A(n21364), .B(n21365), .Z(n21352) );
  AND U23413 ( .A(n21366), .B(n21367), .Z(n21365) );
  XNOR U23414 ( .A(n21368), .B(n21364), .Z(n21367) );
  XOR U23415 ( .A(n21369), .B(nreg[270]), .Z(n21360) );
  IV U23416 ( .A(n21358), .Z(n21369) );
  XOR U23417 ( .A(n21370), .B(n21371), .Z(n21358) );
  AND U23418 ( .A(n21372), .B(n21373), .Z(n21371) );
  XNOR U23419 ( .A(n21370), .B(n10687), .Z(n21373) );
  XNOR U23420 ( .A(n21366), .B(n21368), .Z(n10687) );
  NAND U23421 ( .A(n21374), .B(nreg[269]), .Z(n21368) );
  NAND U23422 ( .A(n12326), .B(nreg[269]), .Z(n21374) );
  XNOR U23423 ( .A(n21364), .B(n21375), .Z(n21366) );
  XOR U23424 ( .A(n21376), .B(n21377), .Z(n21364) );
  AND U23425 ( .A(n21378), .B(n21379), .Z(n21377) );
  XNOR U23426 ( .A(n21380), .B(n21376), .Z(n21379) );
  XOR U23427 ( .A(n21381), .B(nreg[269]), .Z(n21372) );
  IV U23428 ( .A(n21370), .Z(n21381) );
  XOR U23429 ( .A(n21382), .B(n21383), .Z(n21370) );
  AND U23430 ( .A(n21384), .B(n21385), .Z(n21383) );
  XNOR U23431 ( .A(n21382), .B(n10693), .Z(n21385) );
  XNOR U23432 ( .A(n21378), .B(n21380), .Z(n10693) );
  NAND U23433 ( .A(n21386), .B(nreg[268]), .Z(n21380) );
  NAND U23434 ( .A(n12326), .B(nreg[268]), .Z(n21386) );
  XNOR U23435 ( .A(n21376), .B(n21387), .Z(n21378) );
  XOR U23436 ( .A(n21388), .B(n21389), .Z(n21376) );
  AND U23437 ( .A(n21390), .B(n21391), .Z(n21389) );
  XNOR U23438 ( .A(n21392), .B(n21388), .Z(n21391) );
  XOR U23439 ( .A(n21393), .B(nreg[268]), .Z(n21384) );
  IV U23440 ( .A(n21382), .Z(n21393) );
  XOR U23441 ( .A(n21394), .B(n21395), .Z(n21382) );
  AND U23442 ( .A(n21396), .B(n21397), .Z(n21395) );
  XNOR U23443 ( .A(n21394), .B(n10699), .Z(n21397) );
  XNOR U23444 ( .A(n21390), .B(n21392), .Z(n10699) );
  NAND U23445 ( .A(n21398), .B(nreg[267]), .Z(n21392) );
  NAND U23446 ( .A(n12326), .B(nreg[267]), .Z(n21398) );
  XNOR U23447 ( .A(n21388), .B(n21399), .Z(n21390) );
  XOR U23448 ( .A(n21400), .B(n21401), .Z(n21388) );
  AND U23449 ( .A(n21402), .B(n21403), .Z(n21401) );
  XNOR U23450 ( .A(n21404), .B(n21400), .Z(n21403) );
  XOR U23451 ( .A(n21405), .B(nreg[267]), .Z(n21396) );
  IV U23452 ( .A(n21394), .Z(n21405) );
  XOR U23453 ( .A(n21406), .B(n21407), .Z(n21394) );
  AND U23454 ( .A(n21408), .B(n21409), .Z(n21407) );
  XNOR U23455 ( .A(n21406), .B(n10705), .Z(n21409) );
  XNOR U23456 ( .A(n21402), .B(n21404), .Z(n10705) );
  NAND U23457 ( .A(n21410), .B(nreg[266]), .Z(n21404) );
  NAND U23458 ( .A(n12326), .B(nreg[266]), .Z(n21410) );
  XNOR U23459 ( .A(n21400), .B(n21411), .Z(n21402) );
  XOR U23460 ( .A(n21412), .B(n21413), .Z(n21400) );
  AND U23461 ( .A(n21414), .B(n21415), .Z(n21413) );
  XNOR U23462 ( .A(n21416), .B(n21412), .Z(n21415) );
  XOR U23463 ( .A(n21417), .B(nreg[266]), .Z(n21408) );
  IV U23464 ( .A(n21406), .Z(n21417) );
  XOR U23465 ( .A(n21418), .B(n21419), .Z(n21406) );
  AND U23466 ( .A(n21420), .B(n21421), .Z(n21419) );
  XNOR U23467 ( .A(n21418), .B(n10711), .Z(n21421) );
  XNOR U23468 ( .A(n21414), .B(n21416), .Z(n10711) );
  NAND U23469 ( .A(n21422), .B(nreg[265]), .Z(n21416) );
  NAND U23470 ( .A(n12326), .B(nreg[265]), .Z(n21422) );
  XNOR U23471 ( .A(n21412), .B(n21423), .Z(n21414) );
  XOR U23472 ( .A(n21424), .B(n21425), .Z(n21412) );
  AND U23473 ( .A(n21426), .B(n21427), .Z(n21425) );
  XNOR U23474 ( .A(n21428), .B(n21424), .Z(n21427) );
  XOR U23475 ( .A(n21429), .B(nreg[265]), .Z(n21420) );
  IV U23476 ( .A(n21418), .Z(n21429) );
  XOR U23477 ( .A(n21430), .B(n21431), .Z(n21418) );
  AND U23478 ( .A(n21432), .B(n21433), .Z(n21431) );
  XNOR U23479 ( .A(n21430), .B(n10717), .Z(n21433) );
  XNOR U23480 ( .A(n21426), .B(n21428), .Z(n10717) );
  NAND U23481 ( .A(n21434), .B(nreg[264]), .Z(n21428) );
  NAND U23482 ( .A(n12326), .B(nreg[264]), .Z(n21434) );
  XNOR U23483 ( .A(n21424), .B(n21435), .Z(n21426) );
  XOR U23484 ( .A(n21436), .B(n21437), .Z(n21424) );
  AND U23485 ( .A(n21438), .B(n21439), .Z(n21437) );
  XNOR U23486 ( .A(n21440), .B(n21436), .Z(n21439) );
  XOR U23487 ( .A(n21441), .B(nreg[264]), .Z(n21432) );
  IV U23488 ( .A(n21430), .Z(n21441) );
  XOR U23489 ( .A(n21442), .B(n21443), .Z(n21430) );
  AND U23490 ( .A(n21444), .B(n21445), .Z(n21443) );
  XNOR U23491 ( .A(n21442), .B(n10723), .Z(n21445) );
  XNOR U23492 ( .A(n21438), .B(n21440), .Z(n10723) );
  NAND U23493 ( .A(n21446), .B(nreg[263]), .Z(n21440) );
  NAND U23494 ( .A(n12326), .B(nreg[263]), .Z(n21446) );
  XNOR U23495 ( .A(n21436), .B(n21447), .Z(n21438) );
  XOR U23496 ( .A(n21448), .B(n21449), .Z(n21436) );
  AND U23497 ( .A(n21450), .B(n21451), .Z(n21449) );
  XNOR U23498 ( .A(n21452), .B(n21448), .Z(n21451) );
  XOR U23499 ( .A(n21453), .B(nreg[263]), .Z(n21444) );
  IV U23500 ( .A(n21442), .Z(n21453) );
  XOR U23501 ( .A(n21454), .B(n21455), .Z(n21442) );
  AND U23502 ( .A(n21456), .B(n21457), .Z(n21455) );
  XNOR U23503 ( .A(n21454), .B(n10729), .Z(n21457) );
  XNOR U23504 ( .A(n21450), .B(n21452), .Z(n10729) );
  NAND U23505 ( .A(n21458), .B(nreg[262]), .Z(n21452) );
  NAND U23506 ( .A(n12326), .B(nreg[262]), .Z(n21458) );
  XNOR U23507 ( .A(n21448), .B(n21459), .Z(n21450) );
  XOR U23508 ( .A(n21460), .B(n21461), .Z(n21448) );
  AND U23509 ( .A(n21462), .B(n21463), .Z(n21461) );
  XNOR U23510 ( .A(n21464), .B(n21460), .Z(n21463) );
  XOR U23511 ( .A(n21465), .B(nreg[262]), .Z(n21456) );
  IV U23512 ( .A(n21454), .Z(n21465) );
  XOR U23513 ( .A(n21466), .B(n21467), .Z(n21454) );
  AND U23514 ( .A(n21468), .B(n21469), .Z(n21467) );
  XNOR U23515 ( .A(n21466), .B(n10735), .Z(n21469) );
  XNOR U23516 ( .A(n21462), .B(n21464), .Z(n10735) );
  NAND U23517 ( .A(n21470), .B(nreg[261]), .Z(n21464) );
  NAND U23518 ( .A(n12326), .B(nreg[261]), .Z(n21470) );
  XNOR U23519 ( .A(n21460), .B(n21471), .Z(n21462) );
  XOR U23520 ( .A(n21472), .B(n21473), .Z(n21460) );
  AND U23521 ( .A(n21474), .B(n21475), .Z(n21473) );
  XNOR U23522 ( .A(n21476), .B(n21472), .Z(n21475) );
  XOR U23523 ( .A(n21477), .B(nreg[261]), .Z(n21468) );
  IV U23524 ( .A(n21466), .Z(n21477) );
  XOR U23525 ( .A(n21478), .B(n21479), .Z(n21466) );
  AND U23526 ( .A(n21480), .B(n21481), .Z(n21479) );
  XNOR U23527 ( .A(n21478), .B(n10741), .Z(n21481) );
  XNOR U23528 ( .A(n21474), .B(n21476), .Z(n10741) );
  NAND U23529 ( .A(n21482), .B(nreg[260]), .Z(n21476) );
  NAND U23530 ( .A(n12326), .B(nreg[260]), .Z(n21482) );
  XNOR U23531 ( .A(n21472), .B(n21483), .Z(n21474) );
  XOR U23532 ( .A(n21484), .B(n21485), .Z(n21472) );
  AND U23533 ( .A(n21486), .B(n21487), .Z(n21485) );
  XNOR U23534 ( .A(n21488), .B(n21484), .Z(n21487) );
  XOR U23535 ( .A(n21489), .B(nreg[260]), .Z(n21480) );
  IV U23536 ( .A(n21478), .Z(n21489) );
  XOR U23537 ( .A(n21490), .B(n21491), .Z(n21478) );
  AND U23538 ( .A(n21492), .B(n21493), .Z(n21491) );
  XNOR U23539 ( .A(n21490), .B(n10747), .Z(n21493) );
  XNOR U23540 ( .A(n21486), .B(n21488), .Z(n10747) );
  NAND U23541 ( .A(n21494), .B(nreg[259]), .Z(n21488) );
  NAND U23542 ( .A(n12326), .B(nreg[259]), .Z(n21494) );
  XNOR U23543 ( .A(n21484), .B(n21495), .Z(n21486) );
  XOR U23544 ( .A(n21496), .B(n21497), .Z(n21484) );
  AND U23545 ( .A(n21498), .B(n21499), .Z(n21497) );
  XNOR U23546 ( .A(n21500), .B(n21496), .Z(n21499) );
  XOR U23547 ( .A(n21501), .B(nreg[259]), .Z(n21492) );
  IV U23548 ( .A(n21490), .Z(n21501) );
  XOR U23549 ( .A(n21502), .B(n21503), .Z(n21490) );
  AND U23550 ( .A(n21504), .B(n21505), .Z(n21503) );
  XNOR U23551 ( .A(n21502), .B(n10753), .Z(n21505) );
  XNOR U23552 ( .A(n21498), .B(n21500), .Z(n10753) );
  NAND U23553 ( .A(n21506), .B(nreg[258]), .Z(n21500) );
  NAND U23554 ( .A(n12326), .B(nreg[258]), .Z(n21506) );
  XNOR U23555 ( .A(n21496), .B(n21507), .Z(n21498) );
  XOR U23556 ( .A(n21508), .B(n21509), .Z(n21496) );
  AND U23557 ( .A(n21510), .B(n21511), .Z(n21509) );
  XNOR U23558 ( .A(n21512), .B(n21508), .Z(n21511) );
  XOR U23559 ( .A(n21513), .B(nreg[258]), .Z(n21504) );
  IV U23560 ( .A(n21502), .Z(n21513) );
  XOR U23561 ( .A(n21514), .B(n21515), .Z(n21502) );
  AND U23562 ( .A(n21516), .B(n21517), .Z(n21515) );
  XNOR U23563 ( .A(n21514), .B(n10759), .Z(n21517) );
  XNOR U23564 ( .A(n21510), .B(n21512), .Z(n10759) );
  NAND U23565 ( .A(n21518), .B(nreg[257]), .Z(n21512) );
  NAND U23566 ( .A(n12326), .B(nreg[257]), .Z(n21518) );
  XNOR U23567 ( .A(n21508), .B(n21519), .Z(n21510) );
  XOR U23568 ( .A(n21520), .B(n21521), .Z(n21508) );
  AND U23569 ( .A(n21522), .B(n21523), .Z(n21521) );
  XNOR U23570 ( .A(n21524), .B(n21520), .Z(n21523) );
  XOR U23571 ( .A(n21525), .B(nreg[257]), .Z(n21516) );
  IV U23572 ( .A(n21514), .Z(n21525) );
  XOR U23573 ( .A(n21526), .B(n21527), .Z(n21514) );
  AND U23574 ( .A(n21528), .B(n21529), .Z(n21527) );
  XNOR U23575 ( .A(n21526), .B(n10765), .Z(n21529) );
  XNOR U23576 ( .A(n21522), .B(n21524), .Z(n10765) );
  NAND U23577 ( .A(n21530), .B(nreg[256]), .Z(n21524) );
  NAND U23578 ( .A(n12326), .B(nreg[256]), .Z(n21530) );
  XNOR U23579 ( .A(n21520), .B(n21531), .Z(n21522) );
  XOR U23580 ( .A(n21532), .B(n21533), .Z(n21520) );
  AND U23581 ( .A(n21534), .B(n21535), .Z(n21533) );
  XNOR U23582 ( .A(n21536), .B(n21532), .Z(n21535) );
  XOR U23583 ( .A(n21537), .B(nreg[256]), .Z(n21528) );
  IV U23584 ( .A(n21526), .Z(n21537) );
  XOR U23585 ( .A(n21538), .B(n21539), .Z(n21526) );
  AND U23586 ( .A(n21540), .B(n21541), .Z(n21539) );
  XNOR U23587 ( .A(n21538), .B(n10771), .Z(n21541) );
  XNOR U23588 ( .A(n21534), .B(n21536), .Z(n10771) );
  NAND U23589 ( .A(n21542), .B(nreg[255]), .Z(n21536) );
  NAND U23590 ( .A(n12326), .B(nreg[255]), .Z(n21542) );
  XNOR U23591 ( .A(n21532), .B(n21543), .Z(n21534) );
  XOR U23592 ( .A(n21544), .B(n21545), .Z(n21532) );
  AND U23593 ( .A(n21546), .B(n21547), .Z(n21545) );
  XNOR U23594 ( .A(n21548), .B(n21544), .Z(n21547) );
  XOR U23595 ( .A(n21549), .B(nreg[255]), .Z(n21540) );
  IV U23596 ( .A(n21538), .Z(n21549) );
  XOR U23597 ( .A(n21550), .B(n21551), .Z(n21538) );
  AND U23598 ( .A(n21552), .B(n21553), .Z(n21551) );
  XNOR U23599 ( .A(n21550), .B(n10777), .Z(n21553) );
  XNOR U23600 ( .A(n21546), .B(n21548), .Z(n10777) );
  NAND U23601 ( .A(n21554), .B(nreg[254]), .Z(n21548) );
  NAND U23602 ( .A(n12326), .B(nreg[254]), .Z(n21554) );
  XNOR U23603 ( .A(n21544), .B(n21555), .Z(n21546) );
  XOR U23604 ( .A(n21556), .B(n21557), .Z(n21544) );
  AND U23605 ( .A(n21558), .B(n21559), .Z(n21557) );
  XNOR U23606 ( .A(n21560), .B(n21556), .Z(n21559) );
  XOR U23607 ( .A(n21561), .B(nreg[254]), .Z(n21552) );
  IV U23608 ( .A(n21550), .Z(n21561) );
  XOR U23609 ( .A(n21562), .B(n21563), .Z(n21550) );
  AND U23610 ( .A(n21564), .B(n21565), .Z(n21563) );
  XNOR U23611 ( .A(n21562), .B(n10783), .Z(n21565) );
  XNOR U23612 ( .A(n21558), .B(n21560), .Z(n10783) );
  NAND U23613 ( .A(n21566), .B(nreg[253]), .Z(n21560) );
  NAND U23614 ( .A(n12326), .B(nreg[253]), .Z(n21566) );
  XNOR U23615 ( .A(n21556), .B(n21567), .Z(n21558) );
  XOR U23616 ( .A(n21568), .B(n21569), .Z(n21556) );
  AND U23617 ( .A(n21570), .B(n21571), .Z(n21569) );
  XNOR U23618 ( .A(n21572), .B(n21568), .Z(n21571) );
  XOR U23619 ( .A(n21573), .B(nreg[253]), .Z(n21564) );
  IV U23620 ( .A(n21562), .Z(n21573) );
  XOR U23621 ( .A(n21574), .B(n21575), .Z(n21562) );
  AND U23622 ( .A(n21576), .B(n21577), .Z(n21575) );
  XNOR U23623 ( .A(n21574), .B(n10789), .Z(n21577) );
  XNOR U23624 ( .A(n21570), .B(n21572), .Z(n10789) );
  NAND U23625 ( .A(n21578), .B(nreg[252]), .Z(n21572) );
  NAND U23626 ( .A(n12326), .B(nreg[252]), .Z(n21578) );
  XNOR U23627 ( .A(n21568), .B(n21579), .Z(n21570) );
  XOR U23628 ( .A(n21580), .B(n21581), .Z(n21568) );
  AND U23629 ( .A(n21582), .B(n21583), .Z(n21581) );
  XNOR U23630 ( .A(n21584), .B(n21580), .Z(n21583) );
  XOR U23631 ( .A(n21585), .B(nreg[252]), .Z(n21576) );
  IV U23632 ( .A(n21574), .Z(n21585) );
  XOR U23633 ( .A(n21586), .B(n21587), .Z(n21574) );
  AND U23634 ( .A(n21588), .B(n21589), .Z(n21587) );
  XNOR U23635 ( .A(n21586), .B(n10795), .Z(n21589) );
  XNOR U23636 ( .A(n21582), .B(n21584), .Z(n10795) );
  NAND U23637 ( .A(n21590), .B(nreg[251]), .Z(n21584) );
  NAND U23638 ( .A(n12326), .B(nreg[251]), .Z(n21590) );
  XNOR U23639 ( .A(n21580), .B(n21591), .Z(n21582) );
  XOR U23640 ( .A(n21592), .B(n21593), .Z(n21580) );
  AND U23641 ( .A(n21594), .B(n21595), .Z(n21593) );
  XNOR U23642 ( .A(n21596), .B(n21592), .Z(n21595) );
  XOR U23643 ( .A(n21597), .B(nreg[251]), .Z(n21588) );
  IV U23644 ( .A(n21586), .Z(n21597) );
  XOR U23645 ( .A(n21598), .B(n21599), .Z(n21586) );
  AND U23646 ( .A(n21600), .B(n21601), .Z(n21599) );
  XNOR U23647 ( .A(n21598), .B(n10801), .Z(n21601) );
  XNOR U23648 ( .A(n21594), .B(n21596), .Z(n10801) );
  NAND U23649 ( .A(n21602), .B(nreg[250]), .Z(n21596) );
  NAND U23650 ( .A(n12326), .B(nreg[250]), .Z(n21602) );
  XNOR U23651 ( .A(n21592), .B(n21603), .Z(n21594) );
  XOR U23652 ( .A(n21604), .B(n21605), .Z(n21592) );
  AND U23653 ( .A(n21606), .B(n21607), .Z(n21605) );
  XNOR U23654 ( .A(n21608), .B(n21604), .Z(n21607) );
  XOR U23655 ( .A(n21609), .B(nreg[250]), .Z(n21600) );
  IV U23656 ( .A(n21598), .Z(n21609) );
  XOR U23657 ( .A(n21610), .B(n21611), .Z(n21598) );
  AND U23658 ( .A(n21612), .B(n21613), .Z(n21611) );
  XNOR U23659 ( .A(n21610), .B(n10807), .Z(n21613) );
  XNOR U23660 ( .A(n21606), .B(n21608), .Z(n10807) );
  NAND U23661 ( .A(n21614), .B(nreg[249]), .Z(n21608) );
  NAND U23662 ( .A(n12326), .B(nreg[249]), .Z(n21614) );
  XNOR U23663 ( .A(n21604), .B(n21615), .Z(n21606) );
  XOR U23664 ( .A(n21616), .B(n21617), .Z(n21604) );
  AND U23665 ( .A(n21618), .B(n21619), .Z(n21617) );
  XNOR U23666 ( .A(n21620), .B(n21616), .Z(n21619) );
  XOR U23667 ( .A(n21621), .B(nreg[249]), .Z(n21612) );
  IV U23668 ( .A(n21610), .Z(n21621) );
  XOR U23669 ( .A(n21622), .B(n21623), .Z(n21610) );
  AND U23670 ( .A(n21624), .B(n21625), .Z(n21623) );
  XNOR U23671 ( .A(n21622), .B(n10813), .Z(n21625) );
  XNOR U23672 ( .A(n21618), .B(n21620), .Z(n10813) );
  NAND U23673 ( .A(n21626), .B(nreg[248]), .Z(n21620) );
  NAND U23674 ( .A(n12326), .B(nreg[248]), .Z(n21626) );
  XNOR U23675 ( .A(n21616), .B(n21627), .Z(n21618) );
  XOR U23676 ( .A(n21628), .B(n21629), .Z(n21616) );
  AND U23677 ( .A(n21630), .B(n21631), .Z(n21629) );
  XNOR U23678 ( .A(n21632), .B(n21628), .Z(n21631) );
  XOR U23679 ( .A(n21633), .B(nreg[248]), .Z(n21624) );
  IV U23680 ( .A(n21622), .Z(n21633) );
  XOR U23681 ( .A(n21634), .B(n21635), .Z(n21622) );
  AND U23682 ( .A(n21636), .B(n21637), .Z(n21635) );
  XNOR U23683 ( .A(n21634), .B(n10819), .Z(n21637) );
  XNOR U23684 ( .A(n21630), .B(n21632), .Z(n10819) );
  NAND U23685 ( .A(n21638), .B(nreg[247]), .Z(n21632) );
  NAND U23686 ( .A(n12326), .B(nreg[247]), .Z(n21638) );
  XNOR U23687 ( .A(n21628), .B(n21639), .Z(n21630) );
  XOR U23688 ( .A(n21640), .B(n21641), .Z(n21628) );
  AND U23689 ( .A(n21642), .B(n21643), .Z(n21641) );
  XNOR U23690 ( .A(n21644), .B(n21640), .Z(n21643) );
  XOR U23691 ( .A(n21645), .B(nreg[247]), .Z(n21636) );
  IV U23692 ( .A(n21634), .Z(n21645) );
  XOR U23693 ( .A(n21646), .B(n21647), .Z(n21634) );
  AND U23694 ( .A(n21648), .B(n21649), .Z(n21647) );
  XNOR U23695 ( .A(n21646), .B(n10825), .Z(n21649) );
  XNOR U23696 ( .A(n21642), .B(n21644), .Z(n10825) );
  NAND U23697 ( .A(n21650), .B(nreg[246]), .Z(n21644) );
  NAND U23698 ( .A(n12326), .B(nreg[246]), .Z(n21650) );
  XNOR U23699 ( .A(n21640), .B(n21651), .Z(n21642) );
  XOR U23700 ( .A(n21652), .B(n21653), .Z(n21640) );
  AND U23701 ( .A(n21654), .B(n21655), .Z(n21653) );
  XNOR U23702 ( .A(n21656), .B(n21652), .Z(n21655) );
  XOR U23703 ( .A(n21657), .B(nreg[246]), .Z(n21648) );
  IV U23704 ( .A(n21646), .Z(n21657) );
  XOR U23705 ( .A(n21658), .B(n21659), .Z(n21646) );
  AND U23706 ( .A(n21660), .B(n21661), .Z(n21659) );
  XNOR U23707 ( .A(n21658), .B(n10831), .Z(n21661) );
  XNOR U23708 ( .A(n21654), .B(n21656), .Z(n10831) );
  NAND U23709 ( .A(n21662), .B(nreg[245]), .Z(n21656) );
  NAND U23710 ( .A(n12326), .B(nreg[245]), .Z(n21662) );
  XNOR U23711 ( .A(n21652), .B(n21663), .Z(n21654) );
  XOR U23712 ( .A(n21664), .B(n21665), .Z(n21652) );
  AND U23713 ( .A(n21666), .B(n21667), .Z(n21665) );
  XNOR U23714 ( .A(n21668), .B(n21664), .Z(n21667) );
  XOR U23715 ( .A(n21669), .B(nreg[245]), .Z(n21660) );
  IV U23716 ( .A(n21658), .Z(n21669) );
  XOR U23717 ( .A(n21670), .B(n21671), .Z(n21658) );
  AND U23718 ( .A(n21672), .B(n21673), .Z(n21671) );
  XNOR U23719 ( .A(n21670), .B(n10837), .Z(n21673) );
  XNOR U23720 ( .A(n21666), .B(n21668), .Z(n10837) );
  NAND U23721 ( .A(n21674), .B(nreg[244]), .Z(n21668) );
  NAND U23722 ( .A(n12326), .B(nreg[244]), .Z(n21674) );
  XNOR U23723 ( .A(n21664), .B(n21675), .Z(n21666) );
  XOR U23724 ( .A(n21676), .B(n21677), .Z(n21664) );
  AND U23725 ( .A(n21678), .B(n21679), .Z(n21677) );
  XNOR U23726 ( .A(n21680), .B(n21676), .Z(n21679) );
  XOR U23727 ( .A(n21681), .B(nreg[244]), .Z(n21672) );
  IV U23728 ( .A(n21670), .Z(n21681) );
  XOR U23729 ( .A(n21682), .B(n21683), .Z(n21670) );
  AND U23730 ( .A(n21684), .B(n21685), .Z(n21683) );
  XNOR U23731 ( .A(n21682), .B(n10843), .Z(n21685) );
  XNOR U23732 ( .A(n21678), .B(n21680), .Z(n10843) );
  NAND U23733 ( .A(n21686), .B(nreg[243]), .Z(n21680) );
  NAND U23734 ( .A(n12326), .B(nreg[243]), .Z(n21686) );
  XNOR U23735 ( .A(n21676), .B(n21687), .Z(n21678) );
  XOR U23736 ( .A(n21688), .B(n21689), .Z(n21676) );
  AND U23737 ( .A(n21690), .B(n21691), .Z(n21689) );
  XNOR U23738 ( .A(n21692), .B(n21688), .Z(n21691) );
  XOR U23739 ( .A(n21693), .B(nreg[243]), .Z(n21684) );
  IV U23740 ( .A(n21682), .Z(n21693) );
  XOR U23741 ( .A(n21694), .B(n21695), .Z(n21682) );
  AND U23742 ( .A(n21696), .B(n21697), .Z(n21695) );
  XNOR U23743 ( .A(n21694), .B(n10849), .Z(n21697) );
  XNOR U23744 ( .A(n21690), .B(n21692), .Z(n10849) );
  NAND U23745 ( .A(n21698), .B(nreg[242]), .Z(n21692) );
  NAND U23746 ( .A(n12326), .B(nreg[242]), .Z(n21698) );
  XNOR U23747 ( .A(n21688), .B(n21699), .Z(n21690) );
  XOR U23748 ( .A(n21700), .B(n21701), .Z(n21688) );
  AND U23749 ( .A(n21702), .B(n21703), .Z(n21701) );
  XNOR U23750 ( .A(n21704), .B(n21700), .Z(n21703) );
  XOR U23751 ( .A(n21705), .B(nreg[242]), .Z(n21696) );
  IV U23752 ( .A(n21694), .Z(n21705) );
  XOR U23753 ( .A(n21706), .B(n21707), .Z(n21694) );
  AND U23754 ( .A(n21708), .B(n21709), .Z(n21707) );
  XNOR U23755 ( .A(n21706), .B(n10855), .Z(n21709) );
  XNOR U23756 ( .A(n21702), .B(n21704), .Z(n10855) );
  NAND U23757 ( .A(n21710), .B(nreg[241]), .Z(n21704) );
  NAND U23758 ( .A(n12326), .B(nreg[241]), .Z(n21710) );
  XNOR U23759 ( .A(n21700), .B(n21711), .Z(n21702) );
  XOR U23760 ( .A(n21712), .B(n21713), .Z(n21700) );
  AND U23761 ( .A(n21714), .B(n21715), .Z(n21713) );
  XNOR U23762 ( .A(n21716), .B(n21712), .Z(n21715) );
  XOR U23763 ( .A(n21717), .B(nreg[241]), .Z(n21708) );
  IV U23764 ( .A(n21706), .Z(n21717) );
  XOR U23765 ( .A(n21718), .B(n21719), .Z(n21706) );
  AND U23766 ( .A(n21720), .B(n21721), .Z(n21719) );
  XNOR U23767 ( .A(n21718), .B(n10861), .Z(n21721) );
  XNOR U23768 ( .A(n21714), .B(n21716), .Z(n10861) );
  NAND U23769 ( .A(n21722), .B(nreg[240]), .Z(n21716) );
  NAND U23770 ( .A(n12326), .B(nreg[240]), .Z(n21722) );
  XNOR U23771 ( .A(n21712), .B(n21723), .Z(n21714) );
  XOR U23772 ( .A(n21724), .B(n21725), .Z(n21712) );
  AND U23773 ( .A(n21726), .B(n21727), .Z(n21725) );
  XNOR U23774 ( .A(n21728), .B(n21724), .Z(n21727) );
  XOR U23775 ( .A(n21729), .B(nreg[240]), .Z(n21720) );
  IV U23776 ( .A(n21718), .Z(n21729) );
  XOR U23777 ( .A(n21730), .B(n21731), .Z(n21718) );
  AND U23778 ( .A(n21732), .B(n21733), .Z(n21731) );
  XNOR U23779 ( .A(n21730), .B(n10867), .Z(n21733) );
  XNOR U23780 ( .A(n21726), .B(n21728), .Z(n10867) );
  NAND U23781 ( .A(n21734), .B(nreg[239]), .Z(n21728) );
  NAND U23782 ( .A(n12326), .B(nreg[239]), .Z(n21734) );
  XNOR U23783 ( .A(n21724), .B(n21735), .Z(n21726) );
  XOR U23784 ( .A(n21736), .B(n21737), .Z(n21724) );
  AND U23785 ( .A(n21738), .B(n21739), .Z(n21737) );
  XNOR U23786 ( .A(n21740), .B(n21736), .Z(n21739) );
  XOR U23787 ( .A(n21741), .B(nreg[239]), .Z(n21732) );
  IV U23788 ( .A(n21730), .Z(n21741) );
  XOR U23789 ( .A(n21742), .B(n21743), .Z(n21730) );
  AND U23790 ( .A(n21744), .B(n21745), .Z(n21743) );
  XNOR U23791 ( .A(n21742), .B(n10873), .Z(n21745) );
  XNOR U23792 ( .A(n21738), .B(n21740), .Z(n10873) );
  NAND U23793 ( .A(n21746), .B(nreg[238]), .Z(n21740) );
  NAND U23794 ( .A(n12326), .B(nreg[238]), .Z(n21746) );
  XNOR U23795 ( .A(n21736), .B(n21747), .Z(n21738) );
  XOR U23796 ( .A(n21748), .B(n21749), .Z(n21736) );
  AND U23797 ( .A(n21750), .B(n21751), .Z(n21749) );
  XNOR U23798 ( .A(n21752), .B(n21748), .Z(n21751) );
  XOR U23799 ( .A(n21753), .B(nreg[238]), .Z(n21744) );
  IV U23800 ( .A(n21742), .Z(n21753) );
  XOR U23801 ( .A(n21754), .B(n21755), .Z(n21742) );
  AND U23802 ( .A(n21756), .B(n21757), .Z(n21755) );
  XNOR U23803 ( .A(n21754), .B(n10879), .Z(n21757) );
  XNOR U23804 ( .A(n21750), .B(n21752), .Z(n10879) );
  NAND U23805 ( .A(n21758), .B(nreg[237]), .Z(n21752) );
  NAND U23806 ( .A(n12326), .B(nreg[237]), .Z(n21758) );
  XNOR U23807 ( .A(n21748), .B(n21759), .Z(n21750) );
  XOR U23808 ( .A(n21760), .B(n21761), .Z(n21748) );
  AND U23809 ( .A(n21762), .B(n21763), .Z(n21761) );
  XNOR U23810 ( .A(n21764), .B(n21760), .Z(n21763) );
  XOR U23811 ( .A(n21765), .B(nreg[237]), .Z(n21756) );
  IV U23812 ( .A(n21754), .Z(n21765) );
  XOR U23813 ( .A(n21766), .B(n21767), .Z(n21754) );
  AND U23814 ( .A(n21768), .B(n21769), .Z(n21767) );
  XNOR U23815 ( .A(n21766), .B(n10885), .Z(n21769) );
  XNOR U23816 ( .A(n21762), .B(n21764), .Z(n10885) );
  NAND U23817 ( .A(n21770), .B(nreg[236]), .Z(n21764) );
  NAND U23818 ( .A(n12326), .B(nreg[236]), .Z(n21770) );
  XNOR U23819 ( .A(n21760), .B(n21771), .Z(n21762) );
  XOR U23820 ( .A(n21772), .B(n21773), .Z(n21760) );
  AND U23821 ( .A(n21774), .B(n21775), .Z(n21773) );
  XNOR U23822 ( .A(n21776), .B(n21772), .Z(n21775) );
  XOR U23823 ( .A(n21777), .B(nreg[236]), .Z(n21768) );
  IV U23824 ( .A(n21766), .Z(n21777) );
  XOR U23825 ( .A(n21778), .B(n21779), .Z(n21766) );
  AND U23826 ( .A(n21780), .B(n21781), .Z(n21779) );
  XNOR U23827 ( .A(n21778), .B(n10891), .Z(n21781) );
  XNOR U23828 ( .A(n21774), .B(n21776), .Z(n10891) );
  NAND U23829 ( .A(n21782), .B(nreg[235]), .Z(n21776) );
  NAND U23830 ( .A(n12326), .B(nreg[235]), .Z(n21782) );
  XNOR U23831 ( .A(n21772), .B(n21783), .Z(n21774) );
  XOR U23832 ( .A(n21784), .B(n21785), .Z(n21772) );
  AND U23833 ( .A(n21786), .B(n21787), .Z(n21785) );
  XNOR U23834 ( .A(n21788), .B(n21784), .Z(n21787) );
  XOR U23835 ( .A(n21789), .B(nreg[235]), .Z(n21780) );
  IV U23836 ( .A(n21778), .Z(n21789) );
  XOR U23837 ( .A(n21790), .B(n21791), .Z(n21778) );
  AND U23838 ( .A(n21792), .B(n21793), .Z(n21791) );
  XNOR U23839 ( .A(n21790), .B(n10897), .Z(n21793) );
  XNOR U23840 ( .A(n21786), .B(n21788), .Z(n10897) );
  NAND U23841 ( .A(n21794), .B(nreg[234]), .Z(n21788) );
  NAND U23842 ( .A(n12326), .B(nreg[234]), .Z(n21794) );
  XNOR U23843 ( .A(n21784), .B(n21795), .Z(n21786) );
  XOR U23844 ( .A(n21796), .B(n21797), .Z(n21784) );
  AND U23845 ( .A(n21798), .B(n21799), .Z(n21797) );
  XNOR U23846 ( .A(n21800), .B(n21796), .Z(n21799) );
  XOR U23847 ( .A(n21801), .B(nreg[234]), .Z(n21792) );
  IV U23848 ( .A(n21790), .Z(n21801) );
  XOR U23849 ( .A(n21802), .B(n21803), .Z(n21790) );
  AND U23850 ( .A(n21804), .B(n21805), .Z(n21803) );
  XNOR U23851 ( .A(n21802), .B(n10903), .Z(n21805) );
  XNOR U23852 ( .A(n21798), .B(n21800), .Z(n10903) );
  NAND U23853 ( .A(n21806), .B(nreg[233]), .Z(n21800) );
  NAND U23854 ( .A(n12326), .B(nreg[233]), .Z(n21806) );
  XNOR U23855 ( .A(n21796), .B(n21807), .Z(n21798) );
  XOR U23856 ( .A(n21808), .B(n21809), .Z(n21796) );
  AND U23857 ( .A(n21810), .B(n21811), .Z(n21809) );
  XNOR U23858 ( .A(n21812), .B(n21808), .Z(n21811) );
  XOR U23859 ( .A(n21813), .B(nreg[233]), .Z(n21804) );
  IV U23860 ( .A(n21802), .Z(n21813) );
  XOR U23861 ( .A(n21814), .B(n21815), .Z(n21802) );
  AND U23862 ( .A(n21816), .B(n21817), .Z(n21815) );
  XNOR U23863 ( .A(n21814), .B(n10909), .Z(n21817) );
  XNOR U23864 ( .A(n21810), .B(n21812), .Z(n10909) );
  NAND U23865 ( .A(n21818), .B(nreg[232]), .Z(n21812) );
  NAND U23866 ( .A(n12326), .B(nreg[232]), .Z(n21818) );
  XNOR U23867 ( .A(n21808), .B(n21819), .Z(n21810) );
  XOR U23868 ( .A(n21820), .B(n21821), .Z(n21808) );
  AND U23869 ( .A(n21822), .B(n21823), .Z(n21821) );
  XNOR U23870 ( .A(n21824), .B(n21820), .Z(n21823) );
  XOR U23871 ( .A(n21825), .B(nreg[232]), .Z(n21816) );
  IV U23872 ( .A(n21814), .Z(n21825) );
  XOR U23873 ( .A(n21826), .B(n21827), .Z(n21814) );
  AND U23874 ( .A(n21828), .B(n21829), .Z(n21827) );
  XNOR U23875 ( .A(n21826), .B(n10915), .Z(n21829) );
  XNOR U23876 ( .A(n21822), .B(n21824), .Z(n10915) );
  NAND U23877 ( .A(n21830), .B(nreg[231]), .Z(n21824) );
  NAND U23878 ( .A(n12326), .B(nreg[231]), .Z(n21830) );
  XNOR U23879 ( .A(n21820), .B(n21831), .Z(n21822) );
  XOR U23880 ( .A(n21832), .B(n21833), .Z(n21820) );
  AND U23881 ( .A(n21834), .B(n21835), .Z(n21833) );
  XNOR U23882 ( .A(n21836), .B(n21832), .Z(n21835) );
  XOR U23883 ( .A(n21837), .B(nreg[231]), .Z(n21828) );
  IV U23884 ( .A(n21826), .Z(n21837) );
  XOR U23885 ( .A(n21838), .B(n21839), .Z(n21826) );
  AND U23886 ( .A(n21840), .B(n21841), .Z(n21839) );
  XNOR U23887 ( .A(n21838), .B(n10921), .Z(n21841) );
  XNOR U23888 ( .A(n21834), .B(n21836), .Z(n10921) );
  NAND U23889 ( .A(n21842), .B(nreg[230]), .Z(n21836) );
  NAND U23890 ( .A(n12326), .B(nreg[230]), .Z(n21842) );
  XNOR U23891 ( .A(n21832), .B(n21843), .Z(n21834) );
  XOR U23892 ( .A(n21844), .B(n21845), .Z(n21832) );
  AND U23893 ( .A(n21846), .B(n21847), .Z(n21845) );
  XNOR U23894 ( .A(n21848), .B(n21844), .Z(n21847) );
  XOR U23895 ( .A(n21849), .B(nreg[230]), .Z(n21840) );
  IV U23896 ( .A(n21838), .Z(n21849) );
  XOR U23897 ( .A(n21850), .B(n21851), .Z(n21838) );
  AND U23898 ( .A(n21852), .B(n21853), .Z(n21851) );
  XNOR U23899 ( .A(n21850), .B(n10927), .Z(n21853) );
  XNOR U23900 ( .A(n21846), .B(n21848), .Z(n10927) );
  NAND U23901 ( .A(n21854), .B(nreg[229]), .Z(n21848) );
  NAND U23902 ( .A(n12326), .B(nreg[229]), .Z(n21854) );
  XNOR U23903 ( .A(n21844), .B(n21855), .Z(n21846) );
  XOR U23904 ( .A(n21856), .B(n21857), .Z(n21844) );
  AND U23905 ( .A(n21858), .B(n21859), .Z(n21857) );
  XNOR U23906 ( .A(n21860), .B(n21856), .Z(n21859) );
  XOR U23907 ( .A(n21861), .B(nreg[229]), .Z(n21852) );
  IV U23908 ( .A(n21850), .Z(n21861) );
  XOR U23909 ( .A(n21862), .B(n21863), .Z(n21850) );
  AND U23910 ( .A(n21864), .B(n21865), .Z(n21863) );
  XNOR U23911 ( .A(n21862), .B(n10933), .Z(n21865) );
  XNOR U23912 ( .A(n21858), .B(n21860), .Z(n10933) );
  NAND U23913 ( .A(n21866), .B(nreg[228]), .Z(n21860) );
  NAND U23914 ( .A(n12326), .B(nreg[228]), .Z(n21866) );
  XNOR U23915 ( .A(n21856), .B(n21867), .Z(n21858) );
  XOR U23916 ( .A(n21868), .B(n21869), .Z(n21856) );
  AND U23917 ( .A(n21870), .B(n21871), .Z(n21869) );
  XNOR U23918 ( .A(n21872), .B(n21868), .Z(n21871) );
  XOR U23919 ( .A(n21873), .B(nreg[228]), .Z(n21864) );
  IV U23920 ( .A(n21862), .Z(n21873) );
  XOR U23921 ( .A(n21874), .B(n21875), .Z(n21862) );
  AND U23922 ( .A(n21876), .B(n21877), .Z(n21875) );
  XNOR U23923 ( .A(n21874), .B(n10939), .Z(n21877) );
  XNOR U23924 ( .A(n21870), .B(n21872), .Z(n10939) );
  NAND U23925 ( .A(n21878), .B(nreg[227]), .Z(n21872) );
  NAND U23926 ( .A(n12326), .B(nreg[227]), .Z(n21878) );
  XNOR U23927 ( .A(n21868), .B(n21879), .Z(n21870) );
  XOR U23928 ( .A(n21880), .B(n21881), .Z(n21868) );
  AND U23929 ( .A(n21882), .B(n21883), .Z(n21881) );
  XNOR U23930 ( .A(n21884), .B(n21880), .Z(n21883) );
  XOR U23931 ( .A(n21885), .B(nreg[227]), .Z(n21876) );
  IV U23932 ( .A(n21874), .Z(n21885) );
  XOR U23933 ( .A(n21886), .B(n21887), .Z(n21874) );
  AND U23934 ( .A(n21888), .B(n21889), .Z(n21887) );
  XNOR U23935 ( .A(n21886), .B(n10945), .Z(n21889) );
  XNOR U23936 ( .A(n21882), .B(n21884), .Z(n10945) );
  NAND U23937 ( .A(n21890), .B(nreg[226]), .Z(n21884) );
  NAND U23938 ( .A(n12326), .B(nreg[226]), .Z(n21890) );
  XNOR U23939 ( .A(n21880), .B(n21891), .Z(n21882) );
  XOR U23940 ( .A(n21892), .B(n21893), .Z(n21880) );
  AND U23941 ( .A(n21894), .B(n21895), .Z(n21893) );
  XNOR U23942 ( .A(n21896), .B(n21892), .Z(n21895) );
  XOR U23943 ( .A(n21897), .B(nreg[226]), .Z(n21888) );
  IV U23944 ( .A(n21886), .Z(n21897) );
  XOR U23945 ( .A(n21898), .B(n21899), .Z(n21886) );
  AND U23946 ( .A(n21900), .B(n21901), .Z(n21899) );
  XNOR U23947 ( .A(n21898), .B(n10951), .Z(n21901) );
  XNOR U23948 ( .A(n21894), .B(n21896), .Z(n10951) );
  NAND U23949 ( .A(n21902), .B(nreg[225]), .Z(n21896) );
  NAND U23950 ( .A(n12326), .B(nreg[225]), .Z(n21902) );
  XNOR U23951 ( .A(n21892), .B(n21903), .Z(n21894) );
  XOR U23952 ( .A(n21904), .B(n21905), .Z(n21892) );
  AND U23953 ( .A(n21906), .B(n21907), .Z(n21905) );
  XNOR U23954 ( .A(n21908), .B(n21904), .Z(n21907) );
  XOR U23955 ( .A(n21909), .B(nreg[225]), .Z(n21900) );
  IV U23956 ( .A(n21898), .Z(n21909) );
  XOR U23957 ( .A(n21910), .B(n21911), .Z(n21898) );
  AND U23958 ( .A(n21912), .B(n21913), .Z(n21911) );
  XNOR U23959 ( .A(n21910), .B(n10957), .Z(n21913) );
  XNOR U23960 ( .A(n21906), .B(n21908), .Z(n10957) );
  NAND U23961 ( .A(n21914), .B(nreg[224]), .Z(n21908) );
  NAND U23962 ( .A(n12326), .B(nreg[224]), .Z(n21914) );
  XNOR U23963 ( .A(n21904), .B(n21915), .Z(n21906) );
  XOR U23964 ( .A(n21916), .B(n21917), .Z(n21904) );
  AND U23965 ( .A(n21918), .B(n21919), .Z(n21917) );
  XNOR U23966 ( .A(n21920), .B(n21916), .Z(n21919) );
  XOR U23967 ( .A(n21921), .B(nreg[224]), .Z(n21912) );
  IV U23968 ( .A(n21910), .Z(n21921) );
  XOR U23969 ( .A(n21922), .B(n21923), .Z(n21910) );
  AND U23970 ( .A(n21924), .B(n21925), .Z(n21923) );
  XNOR U23971 ( .A(n21922), .B(n10963), .Z(n21925) );
  XNOR U23972 ( .A(n21918), .B(n21920), .Z(n10963) );
  NAND U23973 ( .A(n21926), .B(nreg[223]), .Z(n21920) );
  NAND U23974 ( .A(n12326), .B(nreg[223]), .Z(n21926) );
  XNOR U23975 ( .A(n21916), .B(n21927), .Z(n21918) );
  XOR U23976 ( .A(n21928), .B(n21929), .Z(n21916) );
  AND U23977 ( .A(n21930), .B(n21931), .Z(n21929) );
  XNOR U23978 ( .A(n21932), .B(n21928), .Z(n21931) );
  XOR U23979 ( .A(n21933), .B(nreg[223]), .Z(n21924) );
  IV U23980 ( .A(n21922), .Z(n21933) );
  XOR U23981 ( .A(n21934), .B(n21935), .Z(n21922) );
  AND U23982 ( .A(n21936), .B(n21937), .Z(n21935) );
  XNOR U23983 ( .A(n21934), .B(n10969), .Z(n21937) );
  XNOR U23984 ( .A(n21930), .B(n21932), .Z(n10969) );
  NAND U23985 ( .A(n21938), .B(nreg[222]), .Z(n21932) );
  NAND U23986 ( .A(n12326), .B(nreg[222]), .Z(n21938) );
  XNOR U23987 ( .A(n21928), .B(n21939), .Z(n21930) );
  XOR U23988 ( .A(n21940), .B(n21941), .Z(n21928) );
  AND U23989 ( .A(n21942), .B(n21943), .Z(n21941) );
  XNOR U23990 ( .A(n21944), .B(n21940), .Z(n21943) );
  XOR U23991 ( .A(n21945), .B(nreg[222]), .Z(n21936) );
  IV U23992 ( .A(n21934), .Z(n21945) );
  XOR U23993 ( .A(n21946), .B(n21947), .Z(n21934) );
  AND U23994 ( .A(n21948), .B(n21949), .Z(n21947) );
  XNOR U23995 ( .A(n21946), .B(n10975), .Z(n21949) );
  XNOR U23996 ( .A(n21942), .B(n21944), .Z(n10975) );
  NAND U23997 ( .A(n21950), .B(nreg[221]), .Z(n21944) );
  NAND U23998 ( .A(n12326), .B(nreg[221]), .Z(n21950) );
  XNOR U23999 ( .A(n21940), .B(n21951), .Z(n21942) );
  XOR U24000 ( .A(n21952), .B(n21953), .Z(n21940) );
  AND U24001 ( .A(n21954), .B(n21955), .Z(n21953) );
  XNOR U24002 ( .A(n21956), .B(n21952), .Z(n21955) );
  XOR U24003 ( .A(n21957), .B(nreg[221]), .Z(n21948) );
  IV U24004 ( .A(n21946), .Z(n21957) );
  XOR U24005 ( .A(n21958), .B(n21959), .Z(n21946) );
  AND U24006 ( .A(n21960), .B(n21961), .Z(n21959) );
  XNOR U24007 ( .A(n21958), .B(n10981), .Z(n21961) );
  XNOR U24008 ( .A(n21954), .B(n21956), .Z(n10981) );
  NAND U24009 ( .A(n21962), .B(nreg[220]), .Z(n21956) );
  NAND U24010 ( .A(n12326), .B(nreg[220]), .Z(n21962) );
  XNOR U24011 ( .A(n21952), .B(n21963), .Z(n21954) );
  XOR U24012 ( .A(n21964), .B(n21965), .Z(n21952) );
  AND U24013 ( .A(n21966), .B(n21967), .Z(n21965) );
  XNOR U24014 ( .A(n21968), .B(n21964), .Z(n21967) );
  XOR U24015 ( .A(n21969), .B(nreg[220]), .Z(n21960) );
  IV U24016 ( .A(n21958), .Z(n21969) );
  XOR U24017 ( .A(n21970), .B(n21971), .Z(n21958) );
  AND U24018 ( .A(n21972), .B(n21973), .Z(n21971) );
  XNOR U24019 ( .A(n21970), .B(n10987), .Z(n21973) );
  XNOR U24020 ( .A(n21966), .B(n21968), .Z(n10987) );
  NAND U24021 ( .A(n21974), .B(nreg[219]), .Z(n21968) );
  NAND U24022 ( .A(n12326), .B(nreg[219]), .Z(n21974) );
  XNOR U24023 ( .A(n21964), .B(n21975), .Z(n21966) );
  XOR U24024 ( .A(n21976), .B(n21977), .Z(n21964) );
  AND U24025 ( .A(n21978), .B(n21979), .Z(n21977) );
  XNOR U24026 ( .A(n21980), .B(n21976), .Z(n21979) );
  XOR U24027 ( .A(n21981), .B(nreg[219]), .Z(n21972) );
  IV U24028 ( .A(n21970), .Z(n21981) );
  XOR U24029 ( .A(n21982), .B(n21983), .Z(n21970) );
  AND U24030 ( .A(n21984), .B(n21985), .Z(n21983) );
  XNOR U24031 ( .A(n21982), .B(n10993), .Z(n21985) );
  XNOR U24032 ( .A(n21978), .B(n21980), .Z(n10993) );
  NAND U24033 ( .A(n21986), .B(nreg[218]), .Z(n21980) );
  NAND U24034 ( .A(n12326), .B(nreg[218]), .Z(n21986) );
  XNOR U24035 ( .A(n21976), .B(n21987), .Z(n21978) );
  XOR U24036 ( .A(n21988), .B(n21989), .Z(n21976) );
  AND U24037 ( .A(n21990), .B(n21991), .Z(n21989) );
  XNOR U24038 ( .A(n21992), .B(n21988), .Z(n21991) );
  XOR U24039 ( .A(n21993), .B(nreg[218]), .Z(n21984) );
  IV U24040 ( .A(n21982), .Z(n21993) );
  XOR U24041 ( .A(n21994), .B(n21995), .Z(n21982) );
  AND U24042 ( .A(n21996), .B(n21997), .Z(n21995) );
  XNOR U24043 ( .A(n21994), .B(n10999), .Z(n21997) );
  XNOR U24044 ( .A(n21990), .B(n21992), .Z(n10999) );
  NAND U24045 ( .A(n21998), .B(nreg[217]), .Z(n21992) );
  NAND U24046 ( .A(n12326), .B(nreg[217]), .Z(n21998) );
  XNOR U24047 ( .A(n21988), .B(n21999), .Z(n21990) );
  XOR U24048 ( .A(n22000), .B(n22001), .Z(n21988) );
  AND U24049 ( .A(n22002), .B(n22003), .Z(n22001) );
  XNOR U24050 ( .A(n22004), .B(n22000), .Z(n22003) );
  XOR U24051 ( .A(n22005), .B(nreg[217]), .Z(n21996) );
  IV U24052 ( .A(n21994), .Z(n22005) );
  XOR U24053 ( .A(n22006), .B(n22007), .Z(n21994) );
  AND U24054 ( .A(n22008), .B(n22009), .Z(n22007) );
  XNOR U24055 ( .A(n22006), .B(n11005), .Z(n22009) );
  XNOR U24056 ( .A(n22002), .B(n22004), .Z(n11005) );
  NAND U24057 ( .A(n22010), .B(nreg[216]), .Z(n22004) );
  NAND U24058 ( .A(n12326), .B(nreg[216]), .Z(n22010) );
  XNOR U24059 ( .A(n22000), .B(n22011), .Z(n22002) );
  XOR U24060 ( .A(n22012), .B(n22013), .Z(n22000) );
  AND U24061 ( .A(n22014), .B(n22015), .Z(n22013) );
  XNOR U24062 ( .A(n22016), .B(n22012), .Z(n22015) );
  XOR U24063 ( .A(n22017), .B(nreg[216]), .Z(n22008) );
  IV U24064 ( .A(n22006), .Z(n22017) );
  XOR U24065 ( .A(n22018), .B(n22019), .Z(n22006) );
  AND U24066 ( .A(n22020), .B(n22021), .Z(n22019) );
  XNOR U24067 ( .A(n22018), .B(n11011), .Z(n22021) );
  XNOR U24068 ( .A(n22014), .B(n22016), .Z(n11011) );
  NAND U24069 ( .A(n22022), .B(nreg[215]), .Z(n22016) );
  NAND U24070 ( .A(n12326), .B(nreg[215]), .Z(n22022) );
  XNOR U24071 ( .A(n22012), .B(n22023), .Z(n22014) );
  XOR U24072 ( .A(n22024), .B(n22025), .Z(n22012) );
  AND U24073 ( .A(n22026), .B(n22027), .Z(n22025) );
  XNOR U24074 ( .A(n22028), .B(n22024), .Z(n22027) );
  XOR U24075 ( .A(n22029), .B(nreg[215]), .Z(n22020) );
  IV U24076 ( .A(n22018), .Z(n22029) );
  XOR U24077 ( .A(n22030), .B(n22031), .Z(n22018) );
  AND U24078 ( .A(n22032), .B(n22033), .Z(n22031) );
  XNOR U24079 ( .A(n22030), .B(n11017), .Z(n22033) );
  XNOR U24080 ( .A(n22026), .B(n22028), .Z(n11017) );
  NAND U24081 ( .A(n22034), .B(nreg[214]), .Z(n22028) );
  NAND U24082 ( .A(n12326), .B(nreg[214]), .Z(n22034) );
  XNOR U24083 ( .A(n22024), .B(n22035), .Z(n22026) );
  XOR U24084 ( .A(n22036), .B(n22037), .Z(n22024) );
  AND U24085 ( .A(n22038), .B(n22039), .Z(n22037) );
  XNOR U24086 ( .A(n22040), .B(n22036), .Z(n22039) );
  XOR U24087 ( .A(n22041), .B(nreg[214]), .Z(n22032) );
  IV U24088 ( .A(n22030), .Z(n22041) );
  XOR U24089 ( .A(n22042), .B(n22043), .Z(n22030) );
  AND U24090 ( .A(n22044), .B(n22045), .Z(n22043) );
  XNOR U24091 ( .A(n22042), .B(n11023), .Z(n22045) );
  XNOR U24092 ( .A(n22038), .B(n22040), .Z(n11023) );
  NAND U24093 ( .A(n22046), .B(nreg[213]), .Z(n22040) );
  NAND U24094 ( .A(n12326), .B(nreg[213]), .Z(n22046) );
  XNOR U24095 ( .A(n22036), .B(n22047), .Z(n22038) );
  XOR U24096 ( .A(n22048), .B(n22049), .Z(n22036) );
  AND U24097 ( .A(n22050), .B(n22051), .Z(n22049) );
  XNOR U24098 ( .A(n22052), .B(n22048), .Z(n22051) );
  XOR U24099 ( .A(n22053), .B(nreg[213]), .Z(n22044) );
  IV U24100 ( .A(n22042), .Z(n22053) );
  XOR U24101 ( .A(n22054), .B(n22055), .Z(n22042) );
  AND U24102 ( .A(n22056), .B(n22057), .Z(n22055) );
  XNOR U24103 ( .A(n22054), .B(n11029), .Z(n22057) );
  XNOR U24104 ( .A(n22050), .B(n22052), .Z(n11029) );
  NAND U24105 ( .A(n22058), .B(nreg[212]), .Z(n22052) );
  NAND U24106 ( .A(n12326), .B(nreg[212]), .Z(n22058) );
  XNOR U24107 ( .A(n22048), .B(n22059), .Z(n22050) );
  XOR U24108 ( .A(n22060), .B(n22061), .Z(n22048) );
  AND U24109 ( .A(n22062), .B(n22063), .Z(n22061) );
  XNOR U24110 ( .A(n22064), .B(n22060), .Z(n22063) );
  XOR U24111 ( .A(n22065), .B(nreg[212]), .Z(n22056) );
  IV U24112 ( .A(n22054), .Z(n22065) );
  XOR U24113 ( .A(n22066), .B(n22067), .Z(n22054) );
  AND U24114 ( .A(n22068), .B(n22069), .Z(n22067) );
  XNOR U24115 ( .A(n22066), .B(n11035), .Z(n22069) );
  XNOR U24116 ( .A(n22062), .B(n22064), .Z(n11035) );
  NAND U24117 ( .A(n22070), .B(nreg[211]), .Z(n22064) );
  NAND U24118 ( .A(n12326), .B(nreg[211]), .Z(n22070) );
  XNOR U24119 ( .A(n22060), .B(n22071), .Z(n22062) );
  XOR U24120 ( .A(n22072), .B(n22073), .Z(n22060) );
  AND U24121 ( .A(n22074), .B(n22075), .Z(n22073) );
  XNOR U24122 ( .A(n22076), .B(n22072), .Z(n22075) );
  XOR U24123 ( .A(n22077), .B(nreg[211]), .Z(n22068) );
  IV U24124 ( .A(n22066), .Z(n22077) );
  XOR U24125 ( .A(n22078), .B(n22079), .Z(n22066) );
  AND U24126 ( .A(n22080), .B(n22081), .Z(n22079) );
  XNOR U24127 ( .A(n22078), .B(n11041), .Z(n22081) );
  XNOR U24128 ( .A(n22074), .B(n22076), .Z(n11041) );
  NAND U24129 ( .A(n22082), .B(nreg[210]), .Z(n22076) );
  NAND U24130 ( .A(n12326), .B(nreg[210]), .Z(n22082) );
  XNOR U24131 ( .A(n22072), .B(n22083), .Z(n22074) );
  XOR U24132 ( .A(n22084), .B(n22085), .Z(n22072) );
  AND U24133 ( .A(n22086), .B(n22087), .Z(n22085) );
  XNOR U24134 ( .A(n22088), .B(n22084), .Z(n22087) );
  XOR U24135 ( .A(n22089), .B(nreg[210]), .Z(n22080) );
  IV U24136 ( .A(n22078), .Z(n22089) );
  XOR U24137 ( .A(n22090), .B(n22091), .Z(n22078) );
  AND U24138 ( .A(n22092), .B(n22093), .Z(n22091) );
  XNOR U24139 ( .A(n22090), .B(n11047), .Z(n22093) );
  XNOR U24140 ( .A(n22086), .B(n22088), .Z(n11047) );
  NAND U24141 ( .A(n22094), .B(nreg[209]), .Z(n22088) );
  NAND U24142 ( .A(n12326), .B(nreg[209]), .Z(n22094) );
  XNOR U24143 ( .A(n22084), .B(n22095), .Z(n22086) );
  XOR U24144 ( .A(n22096), .B(n22097), .Z(n22084) );
  AND U24145 ( .A(n22098), .B(n22099), .Z(n22097) );
  XNOR U24146 ( .A(n22100), .B(n22096), .Z(n22099) );
  XOR U24147 ( .A(n22101), .B(nreg[209]), .Z(n22092) );
  IV U24148 ( .A(n22090), .Z(n22101) );
  XOR U24149 ( .A(n22102), .B(n22103), .Z(n22090) );
  AND U24150 ( .A(n22104), .B(n22105), .Z(n22103) );
  XNOR U24151 ( .A(n22102), .B(n11053), .Z(n22105) );
  XNOR U24152 ( .A(n22098), .B(n22100), .Z(n11053) );
  NAND U24153 ( .A(n22106), .B(nreg[208]), .Z(n22100) );
  NAND U24154 ( .A(n12326), .B(nreg[208]), .Z(n22106) );
  XNOR U24155 ( .A(n22096), .B(n22107), .Z(n22098) );
  XOR U24156 ( .A(n22108), .B(n22109), .Z(n22096) );
  AND U24157 ( .A(n22110), .B(n22111), .Z(n22109) );
  XNOR U24158 ( .A(n22112), .B(n22108), .Z(n22111) );
  XOR U24159 ( .A(n22113), .B(nreg[208]), .Z(n22104) );
  IV U24160 ( .A(n22102), .Z(n22113) );
  XOR U24161 ( .A(n22114), .B(n22115), .Z(n22102) );
  AND U24162 ( .A(n22116), .B(n22117), .Z(n22115) );
  XNOR U24163 ( .A(n22114), .B(n11059), .Z(n22117) );
  XNOR U24164 ( .A(n22110), .B(n22112), .Z(n11059) );
  NAND U24165 ( .A(n22118), .B(nreg[207]), .Z(n22112) );
  NAND U24166 ( .A(n12326), .B(nreg[207]), .Z(n22118) );
  XNOR U24167 ( .A(n22108), .B(n22119), .Z(n22110) );
  XOR U24168 ( .A(n22120), .B(n22121), .Z(n22108) );
  AND U24169 ( .A(n22122), .B(n22123), .Z(n22121) );
  XNOR U24170 ( .A(n22124), .B(n22120), .Z(n22123) );
  XOR U24171 ( .A(n22125), .B(nreg[207]), .Z(n22116) );
  IV U24172 ( .A(n22114), .Z(n22125) );
  XOR U24173 ( .A(n22126), .B(n22127), .Z(n22114) );
  AND U24174 ( .A(n22128), .B(n22129), .Z(n22127) );
  XNOR U24175 ( .A(n22126), .B(n11065), .Z(n22129) );
  XNOR U24176 ( .A(n22122), .B(n22124), .Z(n11065) );
  NAND U24177 ( .A(n22130), .B(nreg[206]), .Z(n22124) );
  NAND U24178 ( .A(n12326), .B(nreg[206]), .Z(n22130) );
  XNOR U24179 ( .A(n22120), .B(n22131), .Z(n22122) );
  XOR U24180 ( .A(n22132), .B(n22133), .Z(n22120) );
  AND U24181 ( .A(n22134), .B(n22135), .Z(n22133) );
  XNOR U24182 ( .A(n22136), .B(n22132), .Z(n22135) );
  XOR U24183 ( .A(n22137), .B(nreg[206]), .Z(n22128) );
  IV U24184 ( .A(n22126), .Z(n22137) );
  XOR U24185 ( .A(n22138), .B(n22139), .Z(n22126) );
  AND U24186 ( .A(n22140), .B(n22141), .Z(n22139) );
  XNOR U24187 ( .A(n22138), .B(n11071), .Z(n22141) );
  XNOR U24188 ( .A(n22134), .B(n22136), .Z(n11071) );
  NAND U24189 ( .A(n22142), .B(nreg[205]), .Z(n22136) );
  NAND U24190 ( .A(n12326), .B(nreg[205]), .Z(n22142) );
  XNOR U24191 ( .A(n22132), .B(n22143), .Z(n22134) );
  XOR U24192 ( .A(n22144), .B(n22145), .Z(n22132) );
  AND U24193 ( .A(n22146), .B(n22147), .Z(n22145) );
  XNOR U24194 ( .A(n22148), .B(n22144), .Z(n22147) );
  XOR U24195 ( .A(n22149), .B(nreg[205]), .Z(n22140) );
  IV U24196 ( .A(n22138), .Z(n22149) );
  XOR U24197 ( .A(n22150), .B(n22151), .Z(n22138) );
  AND U24198 ( .A(n22152), .B(n22153), .Z(n22151) );
  XNOR U24199 ( .A(n22150), .B(n11077), .Z(n22153) );
  XNOR U24200 ( .A(n22146), .B(n22148), .Z(n11077) );
  NAND U24201 ( .A(n22154), .B(nreg[204]), .Z(n22148) );
  NAND U24202 ( .A(n12326), .B(nreg[204]), .Z(n22154) );
  XNOR U24203 ( .A(n22144), .B(n22155), .Z(n22146) );
  XOR U24204 ( .A(n22156), .B(n22157), .Z(n22144) );
  AND U24205 ( .A(n22158), .B(n22159), .Z(n22157) );
  XNOR U24206 ( .A(n22160), .B(n22156), .Z(n22159) );
  XOR U24207 ( .A(n22161), .B(nreg[204]), .Z(n22152) );
  IV U24208 ( .A(n22150), .Z(n22161) );
  XOR U24209 ( .A(n22162), .B(n22163), .Z(n22150) );
  AND U24210 ( .A(n22164), .B(n22165), .Z(n22163) );
  XNOR U24211 ( .A(n22162), .B(n11083), .Z(n22165) );
  XNOR U24212 ( .A(n22158), .B(n22160), .Z(n11083) );
  NAND U24213 ( .A(n22166), .B(nreg[203]), .Z(n22160) );
  NAND U24214 ( .A(n12326), .B(nreg[203]), .Z(n22166) );
  XNOR U24215 ( .A(n22156), .B(n22167), .Z(n22158) );
  XOR U24216 ( .A(n22168), .B(n22169), .Z(n22156) );
  AND U24217 ( .A(n22170), .B(n22171), .Z(n22169) );
  XNOR U24218 ( .A(n22172), .B(n22168), .Z(n22171) );
  XOR U24219 ( .A(n22173), .B(nreg[203]), .Z(n22164) );
  IV U24220 ( .A(n22162), .Z(n22173) );
  XOR U24221 ( .A(n22174), .B(n22175), .Z(n22162) );
  AND U24222 ( .A(n22176), .B(n22177), .Z(n22175) );
  XNOR U24223 ( .A(n22174), .B(n11089), .Z(n22177) );
  XNOR U24224 ( .A(n22170), .B(n22172), .Z(n11089) );
  NAND U24225 ( .A(n22178), .B(nreg[202]), .Z(n22172) );
  NAND U24226 ( .A(n12326), .B(nreg[202]), .Z(n22178) );
  XNOR U24227 ( .A(n22168), .B(n22179), .Z(n22170) );
  XOR U24228 ( .A(n22180), .B(n22181), .Z(n22168) );
  AND U24229 ( .A(n22182), .B(n22183), .Z(n22181) );
  XNOR U24230 ( .A(n22184), .B(n22180), .Z(n22183) );
  XOR U24231 ( .A(n22185), .B(nreg[202]), .Z(n22176) );
  IV U24232 ( .A(n22174), .Z(n22185) );
  XOR U24233 ( .A(n22186), .B(n22187), .Z(n22174) );
  AND U24234 ( .A(n22188), .B(n22189), .Z(n22187) );
  XNOR U24235 ( .A(n22186), .B(n11095), .Z(n22189) );
  XNOR U24236 ( .A(n22182), .B(n22184), .Z(n11095) );
  NAND U24237 ( .A(n22190), .B(nreg[201]), .Z(n22184) );
  NAND U24238 ( .A(n12326), .B(nreg[201]), .Z(n22190) );
  XNOR U24239 ( .A(n22180), .B(n22191), .Z(n22182) );
  XOR U24240 ( .A(n22192), .B(n22193), .Z(n22180) );
  AND U24241 ( .A(n22194), .B(n22195), .Z(n22193) );
  XNOR U24242 ( .A(n22196), .B(n22192), .Z(n22195) );
  XOR U24243 ( .A(n22197), .B(nreg[201]), .Z(n22188) );
  IV U24244 ( .A(n22186), .Z(n22197) );
  XOR U24245 ( .A(n22198), .B(n22199), .Z(n22186) );
  AND U24246 ( .A(n22200), .B(n22201), .Z(n22199) );
  XNOR U24247 ( .A(n22198), .B(n11101), .Z(n22201) );
  XNOR U24248 ( .A(n22194), .B(n22196), .Z(n11101) );
  NAND U24249 ( .A(n22202), .B(nreg[200]), .Z(n22196) );
  NAND U24250 ( .A(n12326), .B(nreg[200]), .Z(n22202) );
  XNOR U24251 ( .A(n22192), .B(n22203), .Z(n22194) );
  XOR U24252 ( .A(n22204), .B(n22205), .Z(n22192) );
  AND U24253 ( .A(n22206), .B(n22207), .Z(n22205) );
  XNOR U24254 ( .A(n22208), .B(n22204), .Z(n22207) );
  XOR U24255 ( .A(n22209), .B(nreg[200]), .Z(n22200) );
  IV U24256 ( .A(n22198), .Z(n22209) );
  XOR U24257 ( .A(n22210), .B(n22211), .Z(n22198) );
  AND U24258 ( .A(n22212), .B(n22213), .Z(n22211) );
  XNOR U24259 ( .A(n22210), .B(n11107), .Z(n22213) );
  XNOR U24260 ( .A(n22206), .B(n22208), .Z(n11107) );
  NAND U24261 ( .A(n22214), .B(nreg[199]), .Z(n22208) );
  NAND U24262 ( .A(n12326), .B(nreg[199]), .Z(n22214) );
  XNOR U24263 ( .A(n22204), .B(n22215), .Z(n22206) );
  XOR U24264 ( .A(n22216), .B(n22217), .Z(n22204) );
  AND U24265 ( .A(n22218), .B(n22219), .Z(n22217) );
  XNOR U24266 ( .A(n22220), .B(n22216), .Z(n22219) );
  XOR U24267 ( .A(n22221), .B(nreg[199]), .Z(n22212) );
  IV U24268 ( .A(n22210), .Z(n22221) );
  XOR U24269 ( .A(n22222), .B(n22223), .Z(n22210) );
  AND U24270 ( .A(n22224), .B(n22225), .Z(n22223) );
  XNOR U24271 ( .A(n22222), .B(n11113), .Z(n22225) );
  XNOR U24272 ( .A(n22218), .B(n22220), .Z(n11113) );
  NAND U24273 ( .A(n22226), .B(nreg[198]), .Z(n22220) );
  NAND U24274 ( .A(n12326), .B(nreg[198]), .Z(n22226) );
  XNOR U24275 ( .A(n22216), .B(n22227), .Z(n22218) );
  XOR U24276 ( .A(n22228), .B(n22229), .Z(n22216) );
  AND U24277 ( .A(n22230), .B(n22231), .Z(n22229) );
  XNOR U24278 ( .A(n22232), .B(n22228), .Z(n22231) );
  XOR U24279 ( .A(n22233), .B(nreg[198]), .Z(n22224) );
  IV U24280 ( .A(n22222), .Z(n22233) );
  XOR U24281 ( .A(n22234), .B(n22235), .Z(n22222) );
  AND U24282 ( .A(n22236), .B(n22237), .Z(n22235) );
  XNOR U24283 ( .A(n22234), .B(n11119), .Z(n22237) );
  XNOR U24284 ( .A(n22230), .B(n22232), .Z(n11119) );
  NAND U24285 ( .A(n22238), .B(nreg[197]), .Z(n22232) );
  NAND U24286 ( .A(n12326), .B(nreg[197]), .Z(n22238) );
  XNOR U24287 ( .A(n22228), .B(n22239), .Z(n22230) );
  XOR U24288 ( .A(n22240), .B(n22241), .Z(n22228) );
  AND U24289 ( .A(n22242), .B(n22243), .Z(n22241) );
  XNOR U24290 ( .A(n22244), .B(n22240), .Z(n22243) );
  XOR U24291 ( .A(n22245), .B(nreg[197]), .Z(n22236) );
  IV U24292 ( .A(n22234), .Z(n22245) );
  XOR U24293 ( .A(n22246), .B(n22247), .Z(n22234) );
  AND U24294 ( .A(n22248), .B(n22249), .Z(n22247) );
  XNOR U24295 ( .A(n22246), .B(n11125), .Z(n22249) );
  XNOR U24296 ( .A(n22242), .B(n22244), .Z(n11125) );
  NAND U24297 ( .A(n22250), .B(nreg[196]), .Z(n22244) );
  NAND U24298 ( .A(n12326), .B(nreg[196]), .Z(n22250) );
  XNOR U24299 ( .A(n22240), .B(n22251), .Z(n22242) );
  XOR U24300 ( .A(n22252), .B(n22253), .Z(n22240) );
  AND U24301 ( .A(n22254), .B(n22255), .Z(n22253) );
  XNOR U24302 ( .A(n22256), .B(n22252), .Z(n22255) );
  XOR U24303 ( .A(n22257), .B(nreg[196]), .Z(n22248) );
  IV U24304 ( .A(n22246), .Z(n22257) );
  XOR U24305 ( .A(n22258), .B(n22259), .Z(n22246) );
  AND U24306 ( .A(n22260), .B(n22261), .Z(n22259) );
  XNOR U24307 ( .A(n22258), .B(n11131), .Z(n22261) );
  XNOR U24308 ( .A(n22254), .B(n22256), .Z(n11131) );
  NAND U24309 ( .A(n22262), .B(nreg[195]), .Z(n22256) );
  NAND U24310 ( .A(n12326), .B(nreg[195]), .Z(n22262) );
  XNOR U24311 ( .A(n22252), .B(n22263), .Z(n22254) );
  XOR U24312 ( .A(n22264), .B(n22265), .Z(n22252) );
  AND U24313 ( .A(n22266), .B(n22267), .Z(n22265) );
  XNOR U24314 ( .A(n22268), .B(n22264), .Z(n22267) );
  XOR U24315 ( .A(n22269), .B(nreg[195]), .Z(n22260) );
  IV U24316 ( .A(n22258), .Z(n22269) );
  XOR U24317 ( .A(n22270), .B(n22271), .Z(n22258) );
  AND U24318 ( .A(n22272), .B(n22273), .Z(n22271) );
  XNOR U24319 ( .A(n22270), .B(n11137), .Z(n22273) );
  XNOR U24320 ( .A(n22266), .B(n22268), .Z(n11137) );
  NAND U24321 ( .A(n22274), .B(nreg[194]), .Z(n22268) );
  NAND U24322 ( .A(n12326), .B(nreg[194]), .Z(n22274) );
  XNOR U24323 ( .A(n22264), .B(n22275), .Z(n22266) );
  XOR U24324 ( .A(n22276), .B(n22277), .Z(n22264) );
  AND U24325 ( .A(n22278), .B(n22279), .Z(n22277) );
  XNOR U24326 ( .A(n22280), .B(n22276), .Z(n22279) );
  XOR U24327 ( .A(n22281), .B(nreg[194]), .Z(n22272) );
  IV U24328 ( .A(n22270), .Z(n22281) );
  XOR U24329 ( .A(n22282), .B(n22283), .Z(n22270) );
  AND U24330 ( .A(n22284), .B(n22285), .Z(n22283) );
  XNOR U24331 ( .A(n22282), .B(n11143), .Z(n22285) );
  XNOR U24332 ( .A(n22278), .B(n22280), .Z(n11143) );
  NAND U24333 ( .A(n22286), .B(nreg[193]), .Z(n22280) );
  NAND U24334 ( .A(n12326), .B(nreg[193]), .Z(n22286) );
  XNOR U24335 ( .A(n22276), .B(n22287), .Z(n22278) );
  XOR U24336 ( .A(n22288), .B(n22289), .Z(n22276) );
  AND U24337 ( .A(n22290), .B(n22291), .Z(n22289) );
  XNOR U24338 ( .A(n22292), .B(n22288), .Z(n22291) );
  XOR U24339 ( .A(n22293), .B(nreg[193]), .Z(n22284) );
  IV U24340 ( .A(n22282), .Z(n22293) );
  XOR U24341 ( .A(n22294), .B(n22295), .Z(n22282) );
  AND U24342 ( .A(n22296), .B(n22297), .Z(n22295) );
  XNOR U24343 ( .A(n22294), .B(n11149), .Z(n22297) );
  XNOR U24344 ( .A(n22290), .B(n22292), .Z(n11149) );
  NAND U24345 ( .A(n22298), .B(nreg[192]), .Z(n22292) );
  NAND U24346 ( .A(n12326), .B(nreg[192]), .Z(n22298) );
  XNOR U24347 ( .A(n22288), .B(n22299), .Z(n22290) );
  XOR U24348 ( .A(n22300), .B(n22301), .Z(n22288) );
  AND U24349 ( .A(n22302), .B(n22303), .Z(n22301) );
  XNOR U24350 ( .A(n22304), .B(n22300), .Z(n22303) );
  XOR U24351 ( .A(n22305), .B(nreg[192]), .Z(n22296) );
  IV U24352 ( .A(n22294), .Z(n22305) );
  XOR U24353 ( .A(n22306), .B(n22307), .Z(n22294) );
  AND U24354 ( .A(n22308), .B(n22309), .Z(n22307) );
  XNOR U24355 ( .A(n22306), .B(n11155), .Z(n22309) );
  XNOR U24356 ( .A(n22302), .B(n22304), .Z(n11155) );
  NAND U24357 ( .A(n22310), .B(nreg[191]), .Z(n22304) );
  NAND U24358 ( .A(n12326), .B(nreg[191]), .Z(n22310) );
  XNOR U24359 ( .A(n22300), .B(n22311), .Z(n22302) );
  XOR U24360 ( .A(n22312), .B(n22313), .Z(n22300) );
  AND U24361 ( .A(n22314), .B(n22315), .Z(n22313) );
  XNOR U24362 ( .A(n22316), .B(n22312), .Z(n22315) );
  XOR U24363 ( .A(n22317), .B(nreg[191]), .Z(n22308) );
  IV U24364 ( .A(n22306), .Z(n22317) );
  XOR U24365 ( .A(n22318), .B(n22319), .Z(n22306) );
  AND U24366 ( .A(n22320), .B(n22321), .Z(n22319) );
  XNOR U24367 ( .A(n22318), .B(n11161), .Z(n22321) );
  XNOR U24368 ( .A(n22314), .B(n22316), .Z(n11161) );
  NAND U24369 ( .A(n22322), .B(nreg[190]), .Z(n22316) );
  NAND U24370 ( .A(n12326), .B(nreg[190]), .Z(n22322) );
  XNOR U24371 ( .A(n22312), .B(n22323), .Z(n22314) );
  XOR U24372 ( .A(n22324), .B(n22325), .Z(n22312) );
  AND U24373 ( .A(n22326), .B(n22327), .Z(n22325) );
  XNOR U24374 ( .A(n22328), .B(n22324), .Z(n22327) );
  XOR U24375 ( .A(n22329), .B(nreg[190]), .Z(n22320) );
  IV U24376 ( .A(n22318), .Z(n22329) );
  XOR U24377 ( .A(n22330), .B(n22331), .Z(n22318) );
  AND U24378 ( .A(n22332), .B(n22333), .Z(n22331) );
  XNOR U24379 ( .A(n22330), .B(n11167), .Z(n22333) );
  XNOR U24380 ( .A(n22326), .B(n22328), .Z(n11167) );
  NAND U24381 ( .A(n22334), .B(nreg[189]), .Z(n22328) );
  NAND U24382 ( .A(n12326), .B(nreg[189]), .Z(n22334) );
  XNOR U24383 ( .A(n22324), .B(n22335), .Z(n22326) );
  XOR U24384 ( .A(n22336), .B(n22337), .Z(n22324) );
  AND U24385 ( .A(n22338), .B(n22339), .Z(n22337) );
  XNOR U24386 ( .A(n22340), .B(n22336), .Z(n22339) );
  XOR U24387 ( .A(n22341), .B(nreg[189]), .Z(n22332) );
  IV U24388 ( .A(n22330), .Z(n22341) );
  XOR U24389 ( .A(n22342), .B(n22343), .Z(n22330) );
  AND U24390 ( .A(n22344), .B(n22345), .Z(n22343) );
  XNOR U24391 ( .A(n22342), .B(n11173), .Z(n22345) );
  XNOR U24392 ( .A(n22338), .B(n22340), .Z(n11173) );
  NAND U24393 ( .A(n22346), .B(nreg[188]), .Z(n22340) );
  NAND U24394 ( .A(n12326), .B(nreg[188]), .Z(n22346) );
  XNOR U24395 ( .A(n22336), .B(n22347), .Z(n22338) );
  XOR U24396 ( .A(n22348), .B(n22349), .Z(n22336) );
  AND U24397 ( .A(n22350), .B(n22351), .Z(n22349) );
  XNOR U24398 ( .A(n22352), .B(n22348), .Z(n22351) );
  XOR U24399 ( .A(n22353), .B(nreg[188]), .Z(n22344) );
  IV U24400 ( .A(n22342), .Z(n22353) );
  XOR U24401 ( .A(n22354), .B(n22355), .Z(n22342) );
  AND U24402 ( .A(n22356), .B(n22357), .Z(n22355) );
  XNOR U24403 ( .A(n22354), .B(n11179), .Z(n22357) );
  XNOR U24404 ( .A(n22350), .B(n22352), .Z(n11179) );
  NAND U24405 ( .A(n22358), .B(nreg[187]), .Z(n22352) );
  NAND U24406 ( .A(n12326), .B(nreg[187]), .Z(n22358) );
  XNOR U24407 ( .A(n22348), .B(n22359), .Z(n22350) );
  XOR U24408 ( .A(n22360), .B(n22361), .Z(n22348) );
  AND U24409 ( .A(n22362), .B(n22363), .Z(n22361) );
  XNOR U24410 ( .A(n22364), .B(n22360), .Z(n22363) );
  XOR U24411 ( .A(n22365), .B(nreg[187]), .Z(n22356) );
  IV U24412 ( .A(n22354), .Z(n22365) );
  XOR U24413 ( .A(n22366), .B(n22367), .Z(n22354) );
  AND U24414 ( .A(n22368), .B(n22369), .Z(n22367) );
  XNOR U24415 ( .A(n22366), .B(n11185), .Z(n22369) );
  XNOR U24416 ( .A(n22362), .B(n22364), .Z(n11185) );
  NAND U24417 ( .A(n22370), .B(nreg[186]), .Z(n22364) );
  NAND U24418 ( .A(n12326), .B(nreg[186]), .Z(n22370) );
  XNOR U24419 ( .A(n22360), .B(n22371), .Z(n22362) );
  XOR U24420 ( .A(n22372), .B(n22373), .Z(n22360) );
  AND U24421 ( .A(n22374), .B(n22375), .Z(n22373) );
  XNOR U24422 ( .A(n22376), .B(n22372), .Z(n22375) );
  XOR U24423 ( .A(n22377), .B(nreg[186]), .Z(n22368) );
  IV U24424 ( .A(n22366), .Z(n22377) );
  XOR U24425 ( .A(n22378), .B(n22379), .Z(n22366) );
  AND U24426 ( .A(n22380), .B(n22381), .Z(n22379) );
  XNOR U24427 ( .A(n22378), .B(n11191), .Z(n22381) );
  XNOR U24428 ( .A(n22374), .B(n22376), .Z(n11191) );
  NAND U24429 ( .A(n22382), .B(nreg[185]), .Z(n22376) );
  NAND U24430 ( .A(n12326), .B(nreg[185]), .Z(n22382) );
  XNOR U24431 ( .A(n22372), .B(n22383), .Z(n22374) );
  XOR U24432 ( .A(n22384), .B(n22385), .Z(n22372) );
  AND U24433 ( .A(n22386), .B(n22387), .Z(n22385) );
  XNOR U24434 ( .A(n22388), .B(n22384), .Z(n22387) );
  XOR U24435 ( .A(n22389), .B(nreg[185]), .Z(n22380) );
  IV U24436 ( .A(n22378), .Z(n22389) );
  XOR U24437 ( .A(n22390), .B(n22391), .Z(n22378) );
  AND U24438 ( .A(n22392), .B(n22393), .Z(n22391) );
  XNOR U24439 ( .A(n22390), .B(n11197), .Z(n22393) );
  XNOR U24440 ( .A(n22386), .B(n22388), .Z(n11197) );
  NAND U24441 ( .A(n22394), .B(nreg[184]), .Z(n22388) );
  NAND U24442 ( .A(n12326), .B(nreg[184]), .Z(n22394) );
  XNOR U24443 ( .A(n22384), .B(n22395), .Z(n22386) );
  XOR U24444 ( .A(n22396), .B(n22397), .Z(n22384) );
  AND U24445 ( .A(n22398), .B(n22399), .Z(n22397) );
  XNOR U24446 ( .A(n22400), .B(n22396), .Z(n22399) );
  XOR U24447 ( .A(n22401), .B(nreg[184]), .Z(n22392) );
  IV U24448 ( .A(n22390), .Z(n22401) );
  XOR U24449 ( .A(n22402), .B(n22403), .Z(n22390) );
  AND U24450 ( .A(n22404), .B(n22405), .Z(n22403) );
  XNOR U24451 ( .A(n22402), .B(n11203), .Z(n22405) );
  XNOR U24452 ( .A(n22398), .B(n22400), .Z(n11203) );
  NAND U24453 ( .A(n22406), .B(nreg[183]), .Z(n22400) );
  NAND U24454 ( .A(n12326), .B(nreg[183]), .Z(n22406) );
  XNOR U24455 ( .A(n22396), .B(n22407), .Z(n22398) );
  XOR U24456 ( .A(n22408), .B(n22409), .Z(n22396) );
  AND U24457 ( .A(n22410), .B(n22411), .Z(n22409) );
  XNOR U24458 ( .A(n22412), .B(n22408), .Z(n22411) );
  XOR U24459 ( .A(n22413), .B(nreg[183]), .Z(n22404) );
  IV U24460 ( .A(n22402), .Z(n22413) );
  XOR U24461 ( .A(n22414), .B(n22415), .Z(n22402) );
  AND U24462 ( .A(n22416), .B(n22417), .Z(n22415) );
  XNOR U24463 ( .A(n22414), .B(n11209), .Z(n22417) );
  XNOR U24464 ( .A(n22410), .B(n22412), .Z(n11209) );
  NAND U24465 ( .A(n22418), .B(nreg[182]), .Z(n22412) );
  NAND U24466 ( .A(n12326), .B(nreg[182]), .Z(n22418) );
  XNOR U24467 ( .A(n22408), .B(n22419), .Z(n22410) );
  XOR U24468 ( .A(n22420), .B(n22421), .Z(n22408) );
  AND U24469 ( .A(n22422), .B(n22423), .Z(n22421) );
  XNOR U24470 ( .A(n22424), .B(n22420), .Z(n22423) );
  XOR U24471 ( .A(n22425), .B(nreg[182]), .Z(n22416) );
  IV U24472 ( .A(n22414), .Z(n22425) );
  XOR U24473 ( .A(n22426), .B(n22427), .Z(n22414) );
  AND U24474 ( .A(n22428), .B(n22429), .Z(n22427) );
  XNOR U24475 ( .A(n22426), .B(n11215), .Z(n22429) );
  XNOR U24476 ( .A(n22422), .B(n22424), .Z(n11215) );
  NAND U24477 ( .A(n22430), .B(nreg[181]), .Z(n22424) );
  NAND U24478 ( .A(n12326), .B(nreg[181]), .Z(n22430) );
  XNOR U24479 ( .A(n22420), .B(n22431), .Z(n22422) );
  XOR U24480 ( .A(n22432), .B(n22433), .Z(n22420) );
  AND U24481 ( .A(n22434), .B(n22435), .Z(n22433) );
  XNOR U24482 ( .A(n22436), .B(n22432), .Z(n22435) );
  XOR U24483 ( .A(n22437), .B(nreg[181]), .Z(n22428) );
  IV U24484 ( .A(n22426), .Z(n22437) );
  XOR U24485 ( .A(n22438), .B(n22439), .Z(n22426) );
  AND U24486 ( .A(n22440), .B(n22441), .Z(n22439) );
  XNOR U24487 ( .A(n22438), .B(n11221), .Z(n22441) );
  XNOR U24488 ( .A(n22434), .B(n22436), .Z(n11221) );
  NAND U24489 ( .A(n22442), .B(nreg[180]), .Z(n22436) );
  NAND U24490 ( .A(n12326), .B(nreg[180]), .Z(n22442) );
  XNOR U24491 ( .A(n22432), .B(n22443), .Z(n22434) );
  XOR U24492 ( .A(n22444), .B(n22445), .Z(n22432) );
  AND U24493 ( .A(n22446), .B(n22447), .Z(n22445) );
  XNOR U24494 ( .A(n22448), .B(n22444), .Z(n22447) );
  XOR U24495 ( .A(n22449), .B(nreg[180]), .Z(n22440) );
  IV U24496 ( .A(n22438), .Z(n22449) );
  XOR U24497 ( .A(n22450), .B(n22451), .Z(n22438) );
  AND U24498 ( .A(n22452), .B(n22453), .Z(n22451) );
  XNOR U24499 ( .A(n22450), .B(n11227), .Z(n22453) );
  XNOR U24500 ( .A(n22446), .B(n22448), .Z(n11227) );
  NAND U24501 ( .A(n22454), .B(nreg[179]), .Z(n22448) );
  NAND U24502 ( .A(n12326), .B(nreg[179]), .Z(n22454) );
  XNOR U24503 ( .A(n22444), .B(n22455), .Z(n22446) );
  XOR U24504 ( .A(n22456), .B(n22457), .Z(n22444) );
  AND U24505 ( .A(n22458), .B(n22459), .Z(n22457) );
  XNOR U24506 ( .A(n22460), .B(n22456), .Z(n22459) );
  XOR U24507 ( .A(n22461), .B(nreg[179]), .Z(n22452) );
  IV U24508 ( .A(n22450), .Z(n22461) );
  XOR U24509 ( .A(n22462), .B(n22463), .Z(n22450) );
  AND U24510 ( .A(n22464), .B(n22465), .Z(n22463) );
  XNOR U24511 ( .A(n22462), .B(n11233), .Z(n22465) );
  XNOR U24512 ( .A(n22458), .B(n22460), .Z(n11233) );
  NAND U24513 ( .A(n22466), .B(nreg[178]), .Z(n22460) );
  NAND U24514 ( .A(n12326), .B(nreg[178]), .Z(n22466) );
  XNOR U24515 ( .A(n22456), .B(n22467), .Z(n22458) );
  XOR U24516 ( .A(n22468), .B(n22469), .Z(n22456) );
  AND U24517 ( .A(n22470), .B(n22471), .Z(n22469) );
  XNOR U24518 ( .A(n22472), .B(n22468), .Z(n22471) );
  XOR U24519 ( .A(n22473), .B(nreg[178]), .Z(n22464) );
  IV U24520 ( .A(n22462), .Z(n22473) );
  XOR U24521 ( .A(n22474), .B(n22475), .Z(n22462) );
  AND U24522 ( .A(n22476), .B(n22477), .Z(n22475) );
  XNOR U24523 ( .A(n22474), .B(n11239), .Z(n22477) );
  XNOR U24524 ( .A(n22470), .B(n22472), .Z(n11239) );
  NAND U24525 ( .A(n22478), .B(nreg[177]), .Z(n22472) );
  NAND U24526 ( .A(n12326), .B(nreg[177]), .Z(n22478) );
  XNOR U24527 ( .A(n22468), .B(n22479), .Z(n22470) );
  XOR U24528 ( .A(n22480), .B(n22481), .Z(n22468) );
  AND U24529 ( .A(n22482), .B(n22483), .Z(n22481) );
  XNOR U24530 ( .A(n22484), .B(n22480), .Z(n22483) );
  XOR U24531 ( .A(n22485), .B(nreg[177]), .Z(n22476) );
  IV U24532 ( .A(n22474), .Z(n22485) );
  XOR U24533 ( .A(n22486), .B(n22487), .Z(n22474) );
  AND U24534 ( .A(n22488), .B(n22489), .Z(n22487) );
  XNOR U24535 ( .A(n22486), .B(n11245), .Z(n22489) );
  XNOR U24536 ( .A(n22482), .B(n22484), .Z(n11245) );
  NAND U24537 ( .A(n22490), .B(nreg[176]), .Z(n22484) );
  NAND U24538 ( .A(n12326), .B(nreg[176]), .Z(n22490) );
  XNOR U24539 ( .A(n22480), .B(n22491), .Z(n22482) );
  XOR U24540 ( .A(n22492), .B(n22493), .Z(n22480) );
  AND U24541 ( .A(n22494), .B(n22495), .Z(n22493) );
  XNOR U24542 ( .A(n22496), .B(n22492), .Z(n22495) );
  XOR U24543 ( .A(n22497), .B(nreg[176]), .Z(n22488) );
  IV U24544 ( .A(n22486), .Z(n22497) );
  XOR U24545 ( .A(n22498), .B(n22499), .Z(n22486) );
  AND U24546 ( .A(n22500), .B(n22501), .Z(n22499) );
  XNOR U24547 ( .A(n22498), .B(n11251), .Z(n22501) );
  XNOR U24548 ( .A(n22494), .B(n22496), .Z(n11251) );
  NAND U24549 ( .A(n22502), .B(nreg[175]), .Z(n22496) );
  NAND U24550 ( .A(n12326), .B(nreg[175]), .Z(n22502) );
  XNOR U24551 ( .A(n22492), .B(n22503), .Z(n22494) );
  XOR U24552 ( .A(n22504), .B(n22505), .Z(n22492) );
  AND U24553 ( .A(n22506), .B(n22507), .Z(n22505) );
  XNOR U24554 ( .A(n22508), .B(n22504), .Z(n22507) );
  XOR U24555 ( .A(n22509), .B(nreg[175]), .Z(n22500) );
  IV U24556 ( .A(n22498), .Z(n22509) );
  XOR U24557 ( .A(n22510), .B(n22511), .Z(n22498) );
  AND U24558 ( .A(n22512), .B(n22513), .Z(n22511) );
  XNOR U24559 ( .A(n22510), .B(n11257), .Z(n22513) );
  XNOR U24560 ( .A(n22506), .B(n22508), .Z(n11257) );
  NAND U24561 ( .A(n22514), .B(nreg[174]), .Z(n22508) );
  NAND U24562 ( .A(n12326), .B(nreg[174]), .Z(n22514) );
  XNOR U24563 ( .A(n22504), .B(n22515), .Z(n22506) );
  XOR U24564 ( .A(n22516), .B(n22517), .Z(n22504) );
  AND U24565 ( .A(n22518), .B(n22519), .Z(n22517) );
  XNOR U24566 ( .A(n22520), .B(n22516), .Z(n22519) );
  XOR U24567 ( .A(n22521), .B(nreg[174]), .Z(n22512) );
  IV U24568 ( .A(n22510), .Z(n22521) );
  XOR U24569 ( .A(n22522), .B(n22523), .Z(n22510) );
  AND U24570 ( .A(n22524), .B(n22525), .Z(n22523) );
  XNOR U24571 ( .A(n22522), .B(n11263), .Z(n22525) );
  XNOR U24572 ( .A(n22518), .B(n22520), .Z(n11263) );
  NAND U24573 ( .A(n22526), .B(nreg[173]), .Z(n22520) );
  NAND U24574 ( .A(n12326), .B(nreg[173]), .Z(n22526) );
  XNOR U24575 ( .A(n22516), .B(n22527), .Z(n22518) );
  XOR U24576 ( .A(n22528), .B(n22529), .Z(n22516) );
  AND U24577 ( .A(n22530), .B(n22531), .Z(n22529) );
  XNOR U24578 ( .A(n22532), .B(n22528), .Z(n22531) );
  XOR U24579 ( .A(n22533), .B(nreg[173]), .Z(n22524) );
  IV U24580 ( .A(n22522), .Z(n22533) );
  XOR U24581 ( .A(n22534), .B(n22535), .Z(n22522) );
  AND U24582 ( .A(n22536), .B(n22537), .Z(n22535) );
  XNOR U24583 ( .A(n22534), .B(n11269), .Z(n22537) );
  XNOR U24584 ( .A(n22530), .B(n22532), .Z(n11269) );
  NAND U24585 ( .A(n22538), .B(nreg[172]), .Z(n22532) );
  NAND U24586 ( .A(n12326), .B(nreg[172]), .Z(n22538) );
  XNOR U24587 ( .A(n22528), .B(n22539), .Z(n22530) );
  XOR U24588 ( .A(n22540), .B(n22541), .Z(n22528) );
  AND U24589 ( .A(n22542), .B(n22543), .Z(n22541) );
  XNOR U24590 ( .A(n22544), .B(n22540), .Z(n22543) );
  XOR U24591 ( .A(n22545), .B(nreg[172]), .Z(n22536) );
  IV U24592 ( .A(n22534), .Z(n22545) );
  XOR U24593 ( .A(n22546), .B(n22547), .Z(n22534) );
  AND U24594 ( .A(n22548), .B(n22549), .Z(n22547) );
  XNOR U24595 ( .A(n22546), .B(n11275), .Z(n22549) );
  XNOR U24596 ( .A(n22542), .B(n22544), .Z(n11275) );
  NAND U24597 ( .A(n22550), .B(nreg[171]), .Z(n22544) );
  NAND U24598 ( .A(n12326), .B(nreg[171]), .Z(n22550) );
  XNOR U24599 ( .A(n22540), .B(n22551), .Z(n22542) );
  XOR U24600 ( .A(n22552), .B(n22553), .Z(n22540) );
  AND U24601 ( .A(n22554), .B(n22555), .Z(n22553) );
  XNOR U24602 ( .A(n22556), .B(n22552), .Z(n22555) );
  XOR U24603 ( .A(n22557), .B(nreg[171]), .Z(n22548) );
  IV U24604 ( .A(n22546), .Z(n22557) );
  XOR U24605 ( .A(n22558), .B(n22559), .Z(n22546) );
  AND U24606 ( .A(n22560), .B(n22561), .Z(n22559) );
  XNOR U24607 ( .A(n22558), .B(n11281), .Z(n22561) );
  XNOR U24608 ( .A(n22554), .B(n22556), .Z(n11281) );
  NAND U24609 ( .A(n22562), .B(nreg[170]), .Z(n22556) );
  NAND U24610 ( .A(n12326), .B(nreg[170]), .Z(n22562) );
  XNOR U24611 ( .A(n22552), .B(n22563), .Z(n22554) );
  XOR U24612 ( .A(n22564), .B(n22565), .Z(n22552) );
  AND U24613 ( .A(n22566), .B(n22567), .Z(n22565) );
  XNOR U24614 ( .A(n22568), .B(n22564), .Z(n22567) );
  XOR U24615 ( .A(n22569), .B(nreg[170]), .Z(n22560) );
  IV U24616 ( .A(n22558), .Z(n22569) );
  XOR U24617 ( .A(n22570), .B(n22571), .Z(n22558) );
  AND U24618 ( .A(n22572), .B(n22573), .Z(n22571) );
  XNOR U24619 ( .A(n22570), .B(n11287), .Z(n22573) );
  XNOR U24620 ( .A(n22566), .B(n22568), .Z(n11287) );
  NAND U24621 ( .A(n22574), .B(nreg[169]), .Z(n22568) );
  NAND U24622 ( .A(n12326), .B(nreg[169]), .Z(n22574) );
  XNOR U24623 ( .A(n22564), .B(n22575), .Z(n22566) );
  XOR U24624 ( .A(n22576), .B(n22577), .Z(n22564) );
  AND U24625 ( .A(n22578), .B(n22579), .Z(n22577) );
  XNOR U24626 ( .A(n22580), .B(n22576), .Z(n22579) );
  XOR U24627 ( .A(n22581), .B(nreg[169]), .Z(n22572) );
  IV U24628 ( .A(n22570), .Z(n22581) );
  XOR U24629 ( .A(n22582), .B(n22583), .Z(n22570) );
  AND U24630 ( .A(n22584), .B(n22585), .Z(n22583) );
  XNOR U24631 ( .A(n22582), .B(n11293), .Z(n22585) );
  XNOR U24632 ( .A(n22578), .B(n22580), .Z(n11293) );
  NAND U24633 ( .A(n22586), .B(nreg[168]), .Z(n22580) );
  NAND U24634 ( .A(n12326), .B(nreg[168]), .Z(n22586) );
  XNOR U24635 ( .A(n22576), .B(n22587), .Z(n22578) );
  XOR U24636 ( .A(n22588), .B(n22589), .Z(n22576) );
  AND U24637 ( .A(n22590), .B(n22591), .Z(n22589) );
  XNOR U24638 ( .A(n22592), .B(n22588), .Z(n22591) );
  XOR U24639 ( .A(n22593), .B(nreg[168]), .Z(n22584) );
  IV U24640 ( .A(n22582), .Z(n22593) );
  XOR U24641 ( .A(n22594), .B(n22595), .Z(n22582) );
  AND U24642 ( .A(n22596), .B(n22597), .Z(n22595) );
  XNOR U24643 ( .A(n22594), .B(n11299), .Z(n22597) );
  XNOR U24644 ( .A(n22590), .B(n22592), .Z(n11299) );
  NAND U24645 ( .A(n22598), .B(nreg[167]), .Z(n22592) );
  NAND U24646 ( .A(n12326), .B(nreg[167]), .Z(n22598) );
  XNOR U24647 ( .A(n22588), .B(n22599), .Z(n22590) );
  XOR U24648 ( .A(n22600), .B(n22601), .Z(n22588) );
  AND U24649 ( .A(n22602), .B(n22603), .Z(n22601) );
  XNOR U24650 ( .A(n22604), .B(n22600), .Z(n22603) );
  XOR U24651 ( .A(n22605), .B(nreg[167]), .Z(n22596) );
  IV U24652 ( .A(n22594), .Z(n22605) );
  XOR U24653 ( .A(n22606), .B(n22607), .Z(n22594) );
  AND U24654 ( .A(n22608), .B(n22609), .Z(n22607) );
  XNOR U24655 ( .A(n22606), .B(n11305), .Z(n22609) );
  XNOR U24656 ( .A(n22602), .B(n22604), .Z(n11305) );
  NAND U24657 ( .A(n22610), .B(nreg[166]), .Z(n22604) );
  NAND U24658 ( .A(n12326), .B(nreg[166]), .Z(n22610) );
  XNOR U24659 ( .A(n22600), .B(n22611), .Z(n22602) );
  XOR U24660 ( .A(n22612), .B(n22613), .Z(n22600) );
  AND U24661 ( .A(n22614), .B(n22615), .Z(n22613) );
  XNOR U24662 ( .A(n22616), .B(n22612), .Z(n22615) );
  XOR U24663 ( .A(n22617), .B(nreg[166]), .Z(n22608) );
  IV U24664 ( .A(n22606), .Z(n22617) );
  XOR U24665 ( .A(n22618), .B(n22619), .Z(n22606) );
  AND U24666 ( .A(n22620), .B(n22621), .Z(n22619) );
  XNOR U24667 ( .A(n22618), .B(n11311), .Z(n22621) );
  XNOR U24668 ( .A(n22614), .B(n22616), .Z(n11311) );
  NAND U24669 ( .A(n22622), .B(nreg[165]), .Z(n22616) );
  NAND U24670 ( .A(n12326), .B(nreg[165]), .Z(n22622) );
  XNOR U24671 ( .A(n22612), .B(n22623), .Z(n22614) );
  XOR U24672 ( .A(n22624), .B(n22625), .Z(n22612) );
  AND U24673 ( .A(n22626), .B(n22627), .Z(n22625) );
  XNOR U24674 ( .A(n22628), .B(n22624), .Z(n22627) );
  XOR U24675 ( .A(n22629), .B(nreg[165]), .Z(n22620) );
  IV U24676 ( .A(n22618), .Z(n22629) );
  XOR U24677 ( .A(n22630), .B(n22631), .Z(n22618) );
  AND U24678 ( .A(n22632), .B(n22633), .Z(n22631) );
  XNOR U24679 ( .A(n22630), .B(n11317), .Z(n22633) );
  XNOR U24680 ( .A(n22626), .B(n22628), .Z(n11317) );
  NAND U24681 ( .A(n22634), .B(nreg[164]), .Z(n22628) );
  NAND U24682 ( .A(n12326), .B(nreg[164]), .Z(n22634) );
  XNOR U24683 ( .A(n22624), .B(n22635), .Z(n22626) );
  XOR U24684 ( .A(n22636), .B(n22637), .Z(n22624) );
  AND U24685 ( .A(n22638), .B(n22639), .Z(n22637) );
  XNOR U24686 ( .A(n22640), .B(n22636), .Z(n22639) );
  XOR U24687 ( .A(n22641), .B(nreg[164]), .Z(n22632) );
  IV U24688 ( .A(n22630), .Z(n22641) );
  XOR U24689 ( .A(n22642), .B(n22643), .Z(n22630) );
  AND U24690 ( .A(n22644), .B(n22645), .Z(n22643) );
  XNOR U24691 ( .A(n22642), .B(n11323), .Z(n22645) );
  XNOR U24692 ( .A(n22638), .B(n22640), .Z(n11323) );
  NAND U24693 ( .A(n22646), .B(nreg[163]), .Z(n22640) );
  NAND U24694 ( .A(n12326), .B(nreg[163]), .Z(n22646) );
  XNOR U24695 ( .A(n22636), .B(n22647), .Z(n22638) );
  XOR U24696 ( .A(n22648), .B(n22649), .Z(n22636) );
  AND U24697 ( .A(n22650), .B(n22651), .Z(n22649) );
  XNOR U24698 ( .A(n22652), .B(n22648), .Z(n22651) );
  XOR U24699 ( .A(n22653), .B(nreg[163]), .Z(n22644) );
  IV U24700 ( .A(n22642), .Z(n22653) );
  XOR U24701 ( .A(n22654), .B(n22655), .Z(n22642) );
  AND U24702 ( .A(n22656), .B(n22657), .Z(n22655) );
  XNOR U24703 ( .A(n22654), .B(n11329), .Z(n22657) );
  XNOR U24704 ( .A(n22650), .B(n22652), .Z(n11329) );
  NAND U24705 ( .A(n22658), .B(nreg[162]), .Z(n22652) );
  NAND U24706 ( .A(n12326), .B(nreg[162]), .Z(n22658) );
  XNOR U24707 ( .A(n22648), .B(n22659), .Z(n22650) );
  XOR U24708 ( .A(n22660), .B(n22661), .Z(n22648) );
  AND U24709 ( .A(n22662), .B(n22663), .Z(n22661) );
  XNOR U24710 ( .A(n22664), .B(n22660), .Z(n22663) );
  XOR U24711 ( .A(n22665), .B(nreg[162]), .Z(n22656) );
  IV U24712 ( .A(n22654), .Z(n22665) );
  XOR U24713 ( .A(n22666), .B(n22667), .Z(n22654) );
  AND U24714 ( .A(n22668), .B(n22669), .Z(n22667) );
  XNOR U24715 ( .A(n22666), .B(n11335), .Z(n22669) );
  XNOR U24716 ( .A(n22662), .B(n22664), .Z(n11335) );
  NAND U24717 ( .A(n22670), .B(nreg[161]), .Z(n22664) );
  NAND U24718 ( .A(n12326), .B(nreg[161]), .Z(n22670) );
  XNOR U24719 ( .A(n22660), .B(n22671), .Z(n22662) );
  XOR U24720 ( .A(n22672), .B(n22673), .Z(n22660) );
  AND U24721 ( .A(n22674), .B(n22675), .Z(n22673) );
  XNOR U24722 ( .A(n22676), .B(n22672), .Z(n22675) );
  XOR U24723 ( .A(n22677), .B(nreg[161]), .Z(n22668) );
  IV U24724 ( .A(n22666), .Z(n22677) );
  XOR U24725 ( .A(n22678), .B(n22679), .Z(n22666) );
  AND U24726 ( .A(n22680), .B(n22681), .Z(n22679) );
  XNOR U24727 ( .A(n22678), .B(n11341), .Z(n22681) );
  XNOR U24728 ( .A(n22674), .B(n22676), .Z(n11341) );
  NAND U24729 ( .A(n22682), .B(nreg[160]), .Z(n22676) );
  NAND U24730 ( .A(n12326), .B(nreg[160]), .Z(n22682) );
  XNOR U24731 ( .A(n22672), .B(n22683), .Z(n22674) );
  XOR U24732 ( .A(n22684), .B(n22685), .Z(n22672) );
  AND U24733 ( .A(n22686), .B(n22687), .Z(n22685) );
  XNOR U24734 ( .A(n22688), .B(n22684), .Z(n22687) );
  XOR U24735 ( .A(n22689), .B(nreg[160]), .Z(n22680) );
  IV U24736 ( .A(n22678), .Z(n22689) );
  XOR U24737 ( .A(n22690), .B(n22691), .Z(n22678) );
  AND U24738 ( .A(n22692), .B(n22693), .Z(n22691) );
  XNOR U24739 ( .A(n22690), .B(n11347), .Z(n22693) );
  XNOR U24740 ( .A(n22686), .B(n22688), .Z(n11347) );
  NAND U24741 ( .A(n22694), .B(nreg[159]), .Z(n22688) );
  NAND U24742 ( .A(n12326), .B(nreg[159]), .Z(n22694) );
  XNOR U24743 ( .A(n22684), .B(n22695), .Z(n22686) );
  XOR U24744 ( .A(n22696), .B(n22697), .Z(n22684) );
  AND U24745 ( .A(n22698), .B(n22699), .Z(n22697) );
  XNOR U24746 ( .A(n22700), .B(n22696), .Z(n22699) );
  XOR U24747 ( .A(n22701), .B(nreg[159]), .Z(n22692) );
  IV U24748 ( .A(n22690), .Z(n22701) );
  XOR U24749 ( .A(n22702), .B(n22703), .Z(n22690) );
  AND U24750 ( .A(n22704), .B(n22705), .Z(n22703) );
  XNOR U24751 ( .A(n22702), .B(n11353), .Z(n22705) );
  XNOR U24752 ( .A(n22698), .B(n22700), .Z(n11353) );
  NAND U24753 ( .A(n22706), .B(nreg[158]), .Z(n22700) );
  NAND U24754 ( .A(n12326), .B(nreg[158]), .Z(n22706) );
  XNOR U24755 ( .A(n22696), .B(n22707), .Z(n22698) );
  XOR U24756 ( .A(n22708), .B(n22709), .Z(n22696) );
  AND U24757 ( .A(n22710), .B(n22711), .Z(n22709) );
  XNOR U24758 ( .A(n22712), .B(n22708), .Z(n22711) );
  XOR U24759 ( .A(n22713), .B(nreg[158]), .Z(n22704) );
  IV U24760 ( .A(n22702), .Z(n22713) );
  XOR U24761 ( .A(n22714), .B(n22715), .Z(n22702) );
  AND U24762 ( .A(n22716), .B(n22717), .Z(n22715) );
  XNOR U24763 ( .A(n22714), .B(n11359), .Z(n22717) );
  XNOR U24764 ( .A(n22710), .B(n22712), .Z(n11359) );
  NAND U24765 ( .A(n22718), .B(nreg[157]), .Z(n22712) );
  NAND U24766 ( .A(n12326), .B(nreg[157]), .Z(n22718) );
  XNOR U24767 ( .A(n22708), .B(n22719), .Z(n22710) );
  XOR U24768 ( .A(n22720), .B(n22721), .Z(n22708) );
  AND U24769 ( .A(n22722), .B(n22723), .Z(n22721) );
  XNOR U24770 ( .A(n22724), .B(n22720), .Z(n22723) );
  XOR U24771 ( .A(n22725), .B(nreg[157]), .Z(n22716) );
  IV U24772 ( .A(n22714), .Z(n22725) );
  XOR U24773 ( .A(n22726), .B(n22727), .Z(n22714) );
  AND U24774 ( .A(n22728), .B(n22729), .Z(n22727) );
  XNOR U24775 ( .A(n22726), .B(n11365), .Z(n22729) );
  XNOR U24776 ( .A(n22722), .B(n22724), .Z(n11365) );
  NAND U24777 ( .A(n22730), .B(nreg[156]), .Z(n22724) );
  NAND U24778 ( .A(n12326), .B(nreg[156]), .Z(n22730) );
  XNOR U24779 ( .A(n22720), .B(n22731), .Z(n22722) );
  XOR U24780 ( .A(n22732), .B(n22733), .Z(n22720) );
  AND U24781 ( .A(n22734), .B(n22735), .Z(n22733) );
  XNOR U24782 ( .A(n22736), .B(n22732), .Z(n22735) );
  XOR U24783 ( .A(n22737), .B(nreg[156]), .Z(n22728) );
  IV U24784 ( .A(n22726), .Z(n22737) );
  XOR U24785 ( .A(n22738), .B(n22739), .Z(n22726) );
  AND U24786 ( .A(n22740), .B(n22741), .Z(n22739) );
  XNOR U24787 ( .A(n22738), .B(n11371), .Z(n22741) );
  XNOR U24788 ( .A(n22734), .B(n22736), .Z(n11371) );
  NAND U24789 ( .A(n22742), .B(nreg[155]), .Z(n22736) );
  NAND U24790 ( .A(n12326), .B(nreg[155]), .Z(n22742) );
  XNOR U24791 ( .A(n22732), .B(n22743), .Z(n22734) );
  XOR U24792 ( .A(n22744), .B(n22745), .Z(n22732) );
  AND U24793 ( .A(n22746), .B(n22747), .Z(n22745) );
  XNOR U24794 ( .A(n22748), .B(n22744), .Z(n22747) );
  XOR U24795 ( .A(n22749), .B(nreg[155]), .Z(n22740) );
  IV U24796 ( .A(n22738), .Z(n22749) );
  XOR U24797 ( .A(n22750), .B(n22751), .Z(n22738) );
  AND U24798 ( .A(n22752), .B(n22753), .Z(n22751) );
  XNOR U24799 ( .A(n22750), .B(n11377), .Z(n22753) );
  XNOR U24800 ( .A(n22746), .B(n22748), .Z(n11377) );
  NAND U24801 ( .A(n22754), .B(nreg[154]), .Z(n22748) );
  NAND U24802 ( .A(n12326), .B(nreg[154]), .Z(n22754) );
  XNOR U24803 ( .A(n22744), .B(n22755), .Z(n22746) );
  XOR U24804 ( .A(n22756), .B(n22757), .Z(n22744) );
  AND U24805 ( .A(n22758), .B(n22759), .Z(n22757) );
  XNOR U24806 ( .A(n22760), .B(n22756), .Z(n22759) );
  XOR U24807 ( .A(n22761), .B(nreg[154]), .Z(n22752) );
  IV U24808 ( .A(n22750), .Z(n22761) );
  XOR U24809 ( .A(n22762), .B(n22763), .Z(n22750) );
  AND U24810 ( .A(n22764), .B(n22765), .Z(n22763) );
  XNOR U24811 ( .A(n22762), .B(n11383), .Z(n22765) );
  XNOR U24812 ( .A(n22758), .B(n22760), .Z(n11383) );
  NAND U24813 ( .A(n22766), .B(nreg[153]), .Z(n22760) );
  NAND U24814 ( .A(n12326), .B(nreg[153]), .Z(n22766) );
  XNOR U24815 ( .A(n22756), .B(n22767), .Z(n22758) );
  XOR U24816 ( .A(n22768), .B(n22769), .Z(n22756) );
  AND U24817 ( .A(n22770), .B(n22771), .Z(n22769) );
  XNOR U24818 ( .A(n22772), .B(n22768), .Z(n22771) );
  XOR U24819 ( .A(n22773), .B(nreg[153]), .Z(n22764) );
  IV U24820 ( .A(n22762), .Z(n22773) );
  XOR U24821 ( .A(n22774), .B(n22775), .Z(n22762) );
  AND U24822 ( .A(n22776), .B(n22777), .Z(n22775) );
  XNOR U24823 ( .A(n22774), .B(n11389), .Z(n22777) );
  XNOR U24824 ( .A(n22770), .B(n22772), .Z(n11389) );
  NAND U24825 ( .A(n22778), .B(nreg[152]), .Z(n22772) );
  NAND U24826 ( .A(n12326), .B(nreg[152]), .Z(n22778) );
  XNOR U24827 ( .A(n22768), .B(n22779), .Z(n22770) );
  XOR U24828 ( .A(n22780), .B(n22781), .Z(n22768) );
  AND U24829 ( .A(n22782), .B(n22783), .Z(n22781) );
  XNOR U24830 ( .A(n22784), .B(n22780), .Z(n22783) );
  XOR U24831 ( .A(n22785), .B(nreg[152]), .Z(n22776) );
  IV U24832 ( .A(n22774), .Z(n22785) );
  XOR U24833 ( .A(n22786), .B(n22787), .Z(n22774) );
  AND U24834 ( .A(n22788), .B(n22789), .Z(n22787) );
  XNOR U24835 ( .A(n22786), .B(n11395), .Z(n22789) );
  XNOR U24836 ( .A(n22782), .B(n22784), .Z(n11395) );
  NAND U24837 ( .A(n22790), .B(nreg[151]), .Z(n22784) );
  NAND U24838 ( .A(n12326), .B(nreg[151]), .Z(n22790) );
  XNOR U24839 ( .A(n22780), .B(n22791), .Z(n22782) );
  XOR U24840 ( .A(n22792), .B(n22793), .Z(n22780) );
  AND U24841 ( .A(n22794), .B(n22795), .Z(n22793) );
  XNOR U24842 ( .A(n22796), .B(n22792), .Z(n22795) );
  XOR U24843 ( .A(n22797), .B(nreg[151]), .Z(n22788) );
  IV U24844 ( .A(n22786), .Z(n22797) );
  XOR U24845 ( .A(n22798), .B(n22799), .Z(n22786) );
  AND U24846 ( .A(n22800), .B(n22801), .Z(n22799) );
  XNOR U24847 ( .A(n22798), .B(n11401), .Z(n22801) );
  XNOR U24848 ( .A(n22794), .B(n22796), .Z(n11401) );
  NAND U24849 ( .A(n22802), .B(nreg[150]), .Z(n22796) );
  NAND U24850 ( .A(n12326), .B(nreg[150]), .Z(n22802) );
  XNOR U24851 ( .A(n22792), .B(n22803), .Z(n22794) );
  XOR U24852 ( .A(n22804), .B(n22805), .Z(n22792) );
  AND U24853 ( .A(n22806), .B(n22807), .Z(n22805) );
  XNOR U24854 ( .A(n22808), .B(n22804), .Z(n22807) );
  XOR U24855 ( .A(n22809), .B(nreg[150]), .Z(n22800) );
  IV U24856 ( .A(n22798), .Z(n22809) );
  XOR U24857 ( .A(n22810), .B(n22811), .Z(n22798) );
  AND U24858 ( .A(n22812), .B(n22813), .Z(n22811) );
  XNOR U24859 ( .A(n22810), .B(n11407), .Z(n22813) );
  XNOR U24860 ( .A(n22806), .B(n22808), .Z(n11407) );
  NAND U24861 ( .A(n22814), .B(nreg[149]), .Z(n22808) );
  NAND U24862 ( .A(n12326), .B(nreg[149]), .Z(n22814) );
  XNOR U24863 ( .A(n22804), .B(n22815), .Z(n22806) );
  XOR U24864 ( .A(n22816), .B(n22817), .Z(n22804) );
  AND U24865 ( .A(n22818), .B(n22819), .Z(n22817) );
  XNOR U24866 ( .A(n22820), .B(n22816), .Z(n22819) );
  XOR U24867 ( .A(n22821), .B(nreg[149]), .Z(n22812) );
  IV U24868 ( .A(n22810), .Z(n22821) );
  XOR U24869 ( .A(n22822), .B(n22823), .Z(n22810) );
  AND U24870 ( .A(n22824), .B(n22825), .Z(n22823) );
  XNOR U24871 ( .A(n22822), .B(n11413), .Z(n22825) );
  XNOR U24872 ( .A(n22818), .B(n22820), .Z(n11413) );
  NAND U24873 ( .A(n22826), .B(nreg[148]), .Z(n22820) );
  NAND U24874 ( .A(n12326), .B(nreg[148]), .Z(n22826) );
  XNOR U24875 ( .A(n22816), .B(n22827), .Z(n22818) );
  XOR U24876 ( .A(n22828), .B(n22829), .Z(n22816) );
  AND U24877 ( .A(n22830), .B(n22831), .Z(n22829) );
  XNOR U24878 ( .A(n22832), .B(n22828), .Z(n22831) );
  XOR U24879 ( .A(n22833), .B(nreg[148]), .Z(n22824) );
  IV U24880 ( .A(n22822), .Z(n22833) );
  XOR U24881 ( .A(n22834), .B(n22835), .Z(n22822) );
  AND U24882 ( .A(n22836), .B(n22837), .Z(n22835) );
  XNOR U24883 ( .A(n22834), .B(n11419), .Z(n22837) );
  XNOR U24884 ( .A(n22830), .B(n22832), .Z(n11419) );
  NAND U24885 ( .A(n22838), .B(nreg[147]), .Z(n22832) );
  NAND U24886 ( .A(n12326), .B(nreg[147]), .Z(n22838) );
  XNOR U24887 ( .A(n22828), .B(n22839), .Z(n22830) );
  XOR U24888 ( .A(n22840), .B(n22841), .Z(n22828) );
  AND U24889 ( .A(n22842), .B(n22843), .Z(n22841) );
  XNOR U24890 ( .A(n22844), .B(n22840), .Z(n22843) );
  XOR U24891 ( .A(n22845), .B(nreg[147]), .Z(n22836) );
  IV U24892 ( .A(n22834), .Z(n22845) );
  XOR U24893 ( .A(n22846), .B(n22847), .Z(n22834) );
  AND U24894 ( .A(n22848), .B(n22849), .Z(n22847) );
  XNOR U24895 ( .A(n22846), .B(n11425), .Z(n22849) );
  XNOR U24896 ( .A(n22842), .B(n22844), .Z(n11425) );
  NAND U24897 ( .A(n22850), .B(nreg[146]), .Z(n22844) );
  NAND U24898 ( .A(n12326), .B(nreg[146]), .Z(n22850) );
  XNOR U24899 ( .A(n22840), .B(n22851), .Z(n22842) );
  XOR U24900 ( .A(n22852), .B(n22853), .Z(n22840) );
  AND U24901 ( .A(n22854), .B(n22855), .Z(n22853) );
  XNOR U24902 ( .A(n22856), .B(n22852), .Z(n22855) );
  XOR U24903 ( .A(n22857), .B(nreg[146]), .Z(n22848) );
  IV U24904 ( .A(n22846), .Z(n22857) );
  XOR U24905 ( .A(n22858), .B(n22859), .Z(n22846) );
  AND U24906 ( .A(n22860), .B(n22861), .Z(n22859) );
  XNOR U24907 ( .A(n22858), .B(n11431), .Z(n22861) );
  XNOR U24908 ( .A(n22854), .B(n22856), .Z(n11431) );
  NAND U24909 ( .A(n22862), .B(nreg[145]), .Z(n22856) );
  NAND U24910 ( .A(n12326), .B(nreg[145]), .Z(n22862) );
  XNOR U24911 ( .A(n22852), .B(n22863), .Z(n22854) );
  XOR U24912 ( .A(n22864), .B(n22865), .Z(n22852) );
  AND U24913 ( .A(n22866), .B(n22867), .Z(n22865) );
  XNOR U24914 ( .A(n22868), .B(n22864), .Z(n22867) );
  XOR U24915 ( .A(n22869), .B(nreg[145]), .Z(n22860) );
  IV U24916 ( .A(n22858), .Z(n22869) );
  XOR U24917 ( .A(n22870), .B(n22871), .Z(n22858) );
  AND U24918 ( .A(n22872), .B(n22873), .Z(n22871) );
  XNOR U24919 ( .A(n22870), .B(n11437), .Z(n22873) );
  XNOR U24920 ( .A(n22866), .B(n22868), .Z(n11437) );
  NAND U24921 ( .A(n22874), .B(nreg[144]), .Z(n22868) );
  NAND U24922 ( .A(n12326), .B(nreg[144]), .Z(n22874) );
  XNOR U24923 ( .A(n22864), .B(n22875), .Z(n22866) );
  XOR U24924 ( .A(n22876), .B(n22877), .Z(n22864) );
  AND U24925 ( .A(n22878), .B(n22879), .Z(n22877) );
  XNOR U24926 ( .A(n22880), .B(n22876), .Z(n22879) );
  XOR U24927 ( .A(n22881), .B(nreg[144]), .Z(n22872) );
  IV U24928 ( .A(n22870), .Z(n22881) );
  XOR U24929 ( .A(n22882), .B(n22883), .Z(n22870) );
  AND U24930 ( .A(n22884), .B(n22885), .Z(n22883) );
  XNOR U24931 ( .A(n22882), .B(n11443), .Z(n22885) );
  XNOR U24932 ( .A(n22878), .B(n22880), .Z(n11443) );
  NAND U24933 ( .A(n22886), .B(nreg[143]), .Z(n22880) );
  NAND U24934 ( .A(n12326), .B(nreg[143]), .Z(n22886) );
  XNOR U24935 ( .A(n22876), .B(n22887), .Z(n22878) );
  XOR U24936 ( .A(n22888), .B(n22889), .Z(n22876) );
  AND U24937 ( .A(n22890), .B(n22891), .Z(n22889) );
  XNOR U24938 ( .A(n22892), .B(n22888), .Z(n22891) );
  XOR U24939 ( .A(n22893), .B(nreg[143]), .Z(n22884) );
  IV U24940 ( .A(n22882), .Z(n22893) );
  XOR U24941 ( .A(n22894), .B(n22895), .Z(n22882) );
  AND U24942 ( .A(n22896), .B(n22897), .Z(n22895) );
  XNOR U24943 ( .A(n22894), .B(n11449), .Z(n22897) );
  XNOR U24944 ( .A(n22890), .B(n22892), .Z(n11449) );
  NAND U24945 ( .A(n22898), .B(nreg[142]), .Z(n22892) );
  NAND U24946 ( .A(n12326), .B(nreg[142]), .Z(n22898) );
  XNOR U24947 ( .A(n22888), .B(n22899), .Z(n22890) );
  XOR U24948 ( .A(n22900), .B(n22901), .Z(n22888) );
  AND U24949 ( .A(n22902), .B(n22903), .Z(n22901) );
  XNOR U24950 ( .A(n22904), .B(n22900), .Z(n22903) );
  XOR U24951 ( .A(n22905), .B(nreg[142]), .Z(n22896) );
  IV U24952 ( .A(n22894), .Z(n22905) );
  XOR U24953 ( .A(n22906), .B(n22907), .Z(n22894) );
  AND U24954 ( .A(n22908), .B(n22909), .Z(n22907) );
  XNOR U24955 ( .A(n22906), .B(n11455), .Z(n22909) );
  XNOR U24956 ( .A(n22902), .B(n22904), .Z(n11455) );
  NAND U24957 ( .A(n22910), .B(nreg[141]), .Z(n22904) );
  NAND U24958 ( .A(n12326), .B(nreg[141]), .Z(n22910) );
  XNOR U24959 ( .A(n22900), .B(n22911), .Z(n22902) );
  XOR U24960 ( .A(n22912), .B(n22913), .Z(n22900) );
  AND U24961 ( .A(n22914), .B(n22915), .Z(n22913) );
  XNOR U24962 ( .A(n22916), .B(n22912), .Z(n22915) );
  XOR U24963 ( .A(n22917), .B(nreg[141]), .Z(n22908) );
  IV U24964 ( .A(n22906), .Z(n22917) );
  XOR U24965 ( .A(n22918), .B(n22919), .Z(n22906) );
  AND U24966 ( .A(n22920), .B(n22921), .Z(n22919) );
  XNOR U24967 ( .A(n22918), .B(n11461), .Z(n22921) );
  XNOR U24968 ( .A(n22914), .B(n22916), .Z(n11461) );
  NAND U24969 ( .A(n22922), .B(nreg[140]), .Z(n22916) );
  NAND U24970 ( .A(n12326), .B(nreg[140]), .Z(n22922) );
  XNOR U24971 ( .A(n22912), .B(n22923), .Z(n22914) );
  XOR U24972 ( .A(n22924), .B(n22925), .Z(n22912) );
  AND U24973 ( .A(n22926), .B(n22927), .Z(n22925) );
  XNOR U24974 ( .A(n22928), .B(n22924), .Z(n22927) );
  XOR U24975 ( .A(n22929), .B(nreg[140]), .Z(n22920) );
  IV U24976 ( .A(n22918), .Z(n22929) );
  XOR U24977 ( .A(n22930), .B(n22931), .Z(n22918) );
  AND U24978 ( .A(n22932), .B(n22933), .Z(n22931) );
  XNOR U24979 ( .A(n22930), .B(n11467), .Z(n22933) );
  XNOR U24980 ( .A(n22926), .B(n22928), .Z(n11467) );
  NAND U24981 ( .A(n22934), .B(nreg[139]), .Z(n22928) );
  NAND U24982 ( .A(n12326), .B(nreg[139]), .Z(n22934) );
  XNOR U24983 ( .A(n22924), .B(n22935), .Z(n22926) );
  XOR U24984 ( .A(n22936), .B(n22937), .Z(n22924) );
  AND U24985 ( .A(n22938), .B(n22939), .Z(n22937) );
  XNOR U24986 ( .A(n22940), .B(n22936), .Z(n22939) );
  XOR U24987 ( .A(n22941), .B(nreg[139]), .Z(n22932) );
  IV U24988 ( .A(n22930), .Z(n22941) );
  XOR U24989 ( .A(n22942), .B(n22943), .Z(n22930) );
  AND U24990 ( .A(n22944), .B(n22945), .Z(n22943) );
  XNOR U24991 ( .A(n22942), .B(n11473), .Z(n22945) );
  XNOR U24992 ( .A(n22938), .B(n22940), .Z(n11473) );
  NAND U24993 ( .A(n22946), .B(nreg[138]), .Z(n22940) );
  NAND U24994 ( .A(n12326), .B(nreg[138]), .Z(n22946) );
  XNOR U24995 ( .A(n22936), .B(n22947), .Z(n22938) );
  XOR U24996 ( .A(n22948), .B(n22949), .Z(n22936) );
  AND U24997 ( .A(n22950), .B(n22951), .Z(n22949) );
  XNOR U24998 ( .A(n22952), .B(n22948), .Z(n22951) );
  XOR U24999 ( .A(n22953), .B(nreg[138]), .Z(n22944) );
  IV U25000 ( .A(n22942), .Z(n22953) );
  XOR U25001 ( .A(n22954), .B(n22955), .Z(n22942) );
  AND U25002 ( .A(n22956), .B(n22957), .Z(n22955) );
  XNOR U25003 ( .A(n22954), .B(n11479), .Z(n22957) );
  XNOR U25004 ( .A(n22950), .B(n22952), .Z(n11479) );
  NAND U25005 ( .A(n22958), .B(nreg[137]), .Z(n22952) );
  NAND U25006 ( .A(n12326), .B(nreg[137]), .Z(n22958) );
  XNOR U25007 ( .A(n22948), .B(n22959), .Z(n22950) );
  XOR U25008 ( .A(n22960), .B(n22961), .Z(n22948) );
  AND U25009 ( .A(n22962), .B(n22963), .Z(n22961) );
  XNOR U25010 ( .A(n22964), .B(n22960), .Z(n22963) );
  XOR U25011 ( .A(n22965), .B(nreg[137]), .Z(n22956) );
  IV U25012 ( .A(n22954), .Z(n22965) );
  XOR U25013 ( .A(n22966), .B(n22967), .Z(n22954) );
  AND U25014 ( .A(n22968), .B(n22969), .Z(n22967) );
  XNOR U25015 ( .A(n22966), .B(n11485), .Z(n22969) );
  XNOR U25016 ( .A(n22962), .B(n22964), .Z(n11485) );
  NAND U25017 ( .A(n22970), .B(nreg[136]), .Z(n22964) );
  NAND U25018 ( .A(n12326), .B(nreg[136]), .Z(n22970) );
  XNOR U25019 ( .A(n22960), .B(n22971), .Z(n22962) );
  XOR U25020 ( .A(n22972), .B(n22973), .Z(n22960) );
  AND U25021 ( .A(n22974), .B(n22975), .Z(n22973) );
  XNOR U25022 ( .A(n22976), .B(n22972), .Z(n22975) );
  XOR U25023 ( .A(n22977), .B(nreg[136]), .Z(n22968) );
  IV U25024 ( .A(n22966), .Z(n22977) );
  XOR U25025 ( .A(n22978), .B(n22979), .Z(n22966) );
  AND U25026 ( .A(n22980), .B(n22981), .Z(n22979) );
  XNOR U25027 ( .A(n22978), .B(n11491), .Z(n22981) );
  XNOR U25028 ( .A(n22974), .B(n22976), .Z(n11491) );
  NAND U25029 ( .A(n22982), .B(nreg[135]), .Z(n22976) );
  NAND U25030 ( .A(n12326), .B(nreg[135]), .Z(n22982) );
  XNOR U25031 ( .A(n22972), .B(n22983), .Z(n22974) );
  XOR U25032 ( .A(n22984), .B(n22985), .Z(n22972) );
  AND U25033 ( .A(n22986), .B(n22987), .Z(n22985) );
  XNOR U25034 ( .A(n22988), .B(n22984), .Z(n22987) );
  XOR U25035 ( .A(n22989), .B(nreg[135]), .Z(n22980) );
  IV U25036 ( .A(n22978), .Z(n22989) );
  XOR U25037 ( .A(n22990), .B(n22991), .Z(n22978) );
  AND U25038 ( .A(n22992), .B(n22993), .Z(n22991) );
  XNOR U25039 ( .A(n22990), .B(n11497), .Z(n22993) );
  XNOR U25040 ( .A(n22986), .B(n22988), .Z(n11497) );
  NAND U25041 ( .A(n22994), .B(nreg[134]), .Z(n22988) );
  NAND U25042 ( .A(n12326), .B(nreg[134]), .Z(n22994) );
  XNOR U25043 ( .A(n22984), .B(n22995), .Z(n22986) );
  XOR U25044 ( .A(n22996), .B(n22997), .Z(n22984) );
  AND U25045 ( .A(n22998), .B(n22999), .Z(n22997) );
  XNOR U25046 ( .A(n23000), .B(n22996), .Z(n22999) );
  XOR U25047 ( .A(n23001), .B(nreg[134]), .Z(n22992) );
  IV U25048 ( .A(n22990), .Z(n23001) );
  XOR U25049 ( .A(n23002), .B(n23003), .Z(n22990) );
  AND U25050 ( .A(n23004), .B(n23005), .Z(n23003) );
  XNOR U25051 ( .A(n23002), .B(n11503), .Z(n23005) );
  XNOR U25052 ( .A(n22998), .B(n23000), .Z(n11503) );
  NAND U25053 ( .A(n23006), .B(nreg[133]), .Z(n23000) );
  NAND U25054 ( .A(n12326), .B(nreg[133]), .Z(n23006) );
  XNOR U25055 ( .A(n22996), .B(n23007), .Z(n22998) );
  XOR U25056 ( .A(n23008), .B(n23009), .Z(n22996) );
  AND U25057 ( .A(n23010), .B(n23011), .Z(n23009) );
  XNOR U25058 ( .A(n23012), .B(n23008), .Z(n23011) );
  XOR U25059 ( .A(n23013), .B(nreg[133]), .Z(n23004) );
  IV U25060 ( .A(n23002), .Z(n23013) );
  XOR U25061 ( .A(n23014), .B(n23015), .Z(n23002) );
  AND U25062 ( .A(n23016), .B(n23017), .Z(n23015) );
  XNOR U25063 ( .A(n23014), .B(n11509), .Z(n23017) );
  XNOR U25064 ( .A(n23010), .B(n23012), .Z(n11509) );
  NAND U25065 ( .A(n23018), .B(nreg[132]), .Z(n23012) );
  NAND U25066 ( .A(n12326), .B(nreg[132]), .Z(n23018) );
  XNOR U25067 ( .A(n23008), .B(n23019), .Z(n23010) );
  XOR U25068 ( .A(n23020), .B(n23021), .Z(n23008) );
  AND U25069 ( .A(n23022), .B(n23023), .Z(n23021) );
  XNOR U25070 ( .A(n23024), .B(n23020), .Z(n23023) );
  XOR U25071 ( .A(n23025), .B(nreg[132]), .Z(n23016) );
  IV U25072 ( .A(n23014), .Z(n23025) );
  XOR U25073 ( .A(n23026), .B(n23027), .Z(n23014) );
  AND U25074 ( .A(n23028), .B(n23029), .Z(n23027) );
  XNOR U25075 ( .A(n23026), .B(n11515), .Z(n23029) );
  XNOR U25076 ( .A(n23022), .B(n23024), .Z(n11515) );
  NAND U25077 ( .A(n23030), .B(nreg[131]), .Z(n23024) );
  NAND U25078 ( .A(n12326), .B(nreg[131]), .Z(n23030) );
  XNOR U25079 ( .A(n23020), .B(n23031), .Z(n23022) );
  XOR U25080 ( .A(n23032), .B(n23033), .Z(n23020) );
  AND U25081 ( .A(n23034), .B(n23035), .Z(n23033) );
  XNOR U25082 ( .A(n23036), .B(n23032), .Z(n23035) );
  XOR U25083 ( .A(n23037), .B(nreg[131]), .Z(n23028) );
  IV U25084 ( .A(n23026), .Z(n23037) );
  XOR U25085 ( .A(n23038), .B(n23039), .Z(n23026) );
  AND U25086 ( .A(n23040), .B(n23041), .Z(n23039) );
  XNOR U25087 ( .A(n23038), .B(n11521), .Z(n23041) );
  XNOR U25088 ( .A(n23034), .B(n23036), .Z(n11521) );
  NAND U25089 ( .A(n23042), .B(nreg[130]), .Z(n23036) );
  NAND U25090 ( .A(n12326), .B(nreg[130]), .Z(n23042) );
  XNOR U25091 ( .A(n23032), .B(n23043), .Z(n23034) );
  XOR U25092 ( .A(n23044), .B(n23045), .Z(n23032) );
  AND U25093 ( .A(n23046), .B(n23047), .Z(n23045) );
  XNOR U25094 ( .A(n23048), .B(n23044), .Z(n23047) );
  XOR U25095 ( .A(n23049), .B(nreg[130]), .Z(n23040) );
  IV U25096 ( .A(n23038), .Z(n23049) );
  XOR U25097 ( .A(n23050), .B(n23051), .Z(n23038) );
  AND U25098 ( .A(n23052), .B(n23053), .Z(n23051) );
  XNOR U25099 ( .A(n23050), .B(n11527), .Z(n23053) );
  XNOR U25100 ( .A(n23046), .B(n23048), .Z(n11527) );
  NAND U25101 ( .A(n23054), .B(nreg[129]), .Z(n23048) );
  NAND U25102 ( .A(n12326), .B(nreg[129]), .Z(n23054) );
  XNOR U25103 ( .A(n23044), .B(n23055), .Z(n23046) );
  XOR U25104 ( .A(n23056), .B(n23057), .Z(n23044) );
  AND U25105 ( .A(n23058), .B(n23059), .Z(n23057) );
  XNOR U25106 ( .A(n23060), .B(n23056), .Z(n23059) );
  XOR U25107 ( .A(n23061), .B(nreg[129]), .Z(n23052) );
  IV U25108 ( .A(n23050), .Z(n23061) );
  XOR U25109 ( .A(n23062), .B(n23063), .Z(n23050) );
  AND U25110 ( .A(n23064), .B(n23065), .Z(n23063) );
  XNOR U25111 ( .A(n23062), .B(n11533), .Z(n23065) );
  XNOR U25112 ( .A(n23058), .B(n23060), .Z(n11533) );
  NAND U25113 ( .A(n23066), .B(nreg[128]), .Z(n23060) );
  NAND U25114 ( .A(n12326), .B(nreg[128]), .Z(n23066) );
  XNOR U25115 ( .A(n23056), .B(n23067), .Z(n23058) );
  XOR U25116 ( .A(n23068), .B(n23069), .Z(n23056) );
  AND U25117 ( .A(n23070), .B(n23071), .Z(n23069) );
  XNOR U25118 ( .A(n23072), .B(n23068), .Z(n23071) );
  XOR U25119 ( .A(n23073), .B(nreg[128]), .Z(n23064) );
  IV U25120 ( .A(n23062), .Z(n23073) );
  XOR U25121 ( .A(n23074), .B(n23075), .Z(n23062) );
  AND U25122 ( .A(n23076), .B(n23077), .Z(n23075) );
  XNOR U25123 ( .A(n23074), .B(n11539), .Z(n23077) );
  XNOR U25124 ( .A(n23070), .B(n23072), .Z(n11539) );
  NAND U25125 ( .A(n23078), .B(nreg[127]), .Z(n23072) );
  NAND U25126 ( .A(n12326), .B(nreg[127]), .Z(n23078) );
  XNOR U25127 ( .A(n23068), .B(n23079), .Z(n23070) );
  XOR U25128 ( .A(n23080), .B(n23081), .Z(n23068) );
  AND U25129 ( .A(n23082), .B(n23083), .Z(n23081) );
  XNOR U25130 ( .A(n23084), .B(n23080), .Z(n23083) );
  XOR U25131 ( .A(n23085), .B(nreg[127]), .Z(n23076) );
  IV U25132 ( .A(n23074), .Z(n23085) );
  XOR U25133 ( .A(n23086), .B(n23087), .Z(n23074) );
  AND U25134 ( .A(n23088), .B(n23089), .Z(n23087) );
  XNOR U25135 ( .A(n23086), .B(n11545), .Z(n23089) );
  XNOR U25136 ( .A(n23082), .B(n23084), .Z(n11545) );
  NAND U25137 ( .A(n23090), .B(nreg[126]), .Z(n23084) );
  NAND U25138 ( .A(n12326), .B(nreg[126]), .Z(n23090) );
  XNOR U25139 ( .A(n23080), .B(n23091), .Z(n23082) );
  XOR U25140 ( .A(n23092), .B(n23093), .Z(n23080) );
  AND U25141 ( .A(n23094), .B(n23095), .Z(n23093) );
  XNOR U25142 ( .A(n23096), .B(n23092), .Z(n23095) );
  XOR U25143 ( .A(n23097), .B(nreg[126]), .Z(n23088) );
  IV U25144 ( .A(n23086), .Z(n23097) );
  XOR U25145 ( .A(n23098), .B(n23099), .Z(n23086) );
  AND U25146 ( .A(n23100), .B(n23101), .Z(n23099) );
  XNOR U25147 ( .A(n23098), .B(n11551), .Z(n23101) );
  XNOR U25148 ( .A(n23094), .B(n23096), .Z(n11551) );
  NAND U25149 ( .A(n23102), .B(nreg[125]), .Z(n23096) );
  NAND U25150 ( .A(n12326), .B(nreg[125]), .Z(n23102) );
  XNOR U25151 ( .A(n23092), .B(n23103), .Z(n23094) );
  XOR U25152 ( .A(n23104), .B(n23105), .Z(n23092) );
  AND U25153 ( .A(n23106), .B(n23107), .Z(n23105) );
  XNOR U25154 ( .A(n23108), .B(n23104), .Z(n23107) );
  XOR U25155 ( .A(n23109), .B(nreg[125]), .Z(n23100) );
  IV U25156 ( .A(n23098), .Z(n23109) );
  XOR U25157 ( .A(n23110), .B(n23111), .Z(n23098) );
  AND U25158 ( .A(n23112), .B(n23113), .Z(n23111) );
  XNOR U25159 ( .A(n23110), .B(n11557), .Z(n23113) );
  XNOR U25160 ( .A(n23106), .B(n23108), .Z(n11557) );
  NAND U25161 ( .A(n23114), .B(nreg[124]), .Z(n23108) );
  NAND U25162 ( .A(n12326), .B(nreg[124]), .Z(n23114) );
  XNOR U25163 ( .A(n23104), .B(n23115), .Z(n23106) );
  XOR U25164 ( .A(n23116), .B(n23117), .Z(n23104) );
  AND U25165 ( .A(n23118), .B(n23119), .Z(n23117) );
  XNOR U25166 ( .A(n23120), .B(n23116), .Z(n23119) );
  XOR U25167 ( .A(n23121), .B(nreg[124]), .Z(n23112) );
  IV U25168 ( .A(n23110), .Z(n23121) );
  XOR U25169 ( .A(n23122), .B(n23123), .Z(n23110) );
  AND U25170 ( .A(n23124), .B(n23125), .Z(n23123) );
  XNOR U25171 ( .A(n23122), .B(n11563), .Z(n23125) );
  XNOR U25172 ( .A(n23118), .B(n23120), .Z(n11563) );
  NAND U25173 ( .A(n23126), .B(nreg[123]), .Z(n23120) );
  NAND U25174 ( .A(n12326), .B(nreg[123]), .Z(n23126) );
  XNOR U25175 ( .A(n23116), .B(n23127), .Z(n23118) );
  XOR U25176 ( .A(n23128), .B(n23129), .Z(n23116) );
  AND U25177 ( .A(n23130), .B(n23131), .Z(n23129) );
  XNOR U25178 ( .A(n23132), .B(n23128), .Z(n23131) );
  XOR U25179 ( .A(n23133), .B(nreg[123]), .Z(n23124) );
  IV U25180 ( .A(n23122), .Z(n23133) );
  XOR U25181 ( .A(n23134), .B(n23135), .Z(n23122) );
  AND U25182 ( .A(n23136), .B(n23137), .Z(n23135) );
  XNOR U25183 ( .A(n23134), .B(n11569), .Z(n23137) );
  XNOR U25184 ( .A(n23130), .B(n23132), .Z(n11569) );
  NAND U25185 ( .A(n23138), .B(nreg[122]), .Z(n23132) );
  NAND U25186 ( .A(n12326), .B(nreg[122]), .Z(n23138) );
  XNOR U25187 ( .A(n23128), .B(n23139), .Z(n23130) );
  XOR U25188 ( .A(n23140), .B(n23141), .Z(n23128) );
  AND U25189 ( .A(n23142), .B(n23143), .Z(n23141) );
  XNOR U25190 ( .A(n23144), .B(n23140), .Z(n23143) );
  XOR U25191 ( .A(n23145), .B(nreg[122]), .Z(n23136) );
  IV U25192 ( .A(n23134), .Z(n23145) );
  XOR U25193 ( .A(n23146), .B(n23147), .Z(n23134) );
  AND U25194 ( .A(n23148), .B(n23149), .Z(n23147) );
  XNOR U25195 ( .A(n23146), .B(n11575), .Z(n23149) );
  XNOR U25196 ( .A(n23142), .B(n23144), .Z(n11575) );
  NAND U25197 ( .A(n23150), .B(nreg[121]), .Z(n23144) );
  NAND U25198 ( .A(n12326), .B(nreg[121]), .Z(n23150) );
  XNOR U25199 ( .A(n23140), .B(n23151), .Z(n23142) );
  XOR U25200 ( .A(n23152), .B(n23153), .Z(n23140) );
  AND U25201 ( .A(n23154), .B(n23155), .Z(n23153) );
  XNOR U25202 ( .A(n23156), .B(n23152), .Z(n23155) );
  XOR U25203 ( .A(n23157), .B(nreg[121]), .Z(n23148) );
  IV U25204 ( .A(n23146), .Z(n23157) );
  XOR U25205 ( .A(n23158), .B(n23159), .Z(n23146) );
  AND U25206 ( .A(n23160), .B(n23161), .Z(n23159) );
  XNOR U25207 ( .A(n23158), .B(n11581), .Z(n23161) );
  XNOR U25208 ( .A(n23154), .B(n23156), .Z(n11581) );
  NAND U25209 ( .A(n23162), .B(nreg[120]), .Z(n23156) );
  NAND U25210 ( .A(n12326), .B(nreg[120]), .Z(n23162) );
  XNOR U25211 ( .A(n23152), .B(n23163), .Z(n23154) );
  XOR U25212 ( .A(n23164), .B(n23165), .Z(n23152) );
  AND U25213 ( .A(n23166), .B(n23167), .Z(n23165) );
  XNOR U25214 ( .A(n23168), .B(n23164), .Z(n23167) );
  XOR U25215 ( .A(n23169), .B(nreg[120]), .Z(n23160) );
  IV U25216 ( .A(n23158), .Z(n23169) );
  XOR U25217 ( .A(n23170), .B(n23171), .Z(n23158) );
  AND U25218 ( .A(n23172), .B(n23173), .Z(n23171) );
  XNOR U25219 ( .A(n23170), .B(n11587), .Z(n23173) );
  XNOR U25220 ( .A(n23166), .B(n23168), .Z(n11587) );
  NAND U25221 ( .A(n23174), .B(nreg[119]), .Z(n23168) );
  NAND U25222 ( .A(n12326), .B(nreg[119]), .Z(n23174) );
  XNOR U25223 ( .A(n23164), .B(n23175), .Z(n23166) );
  XOR U25224 ( .A(n23176), .B(n23177), .Z(n23164) );
  AND U25225 ( .A(n23178), .B(n23179), .Z(n23177) );
  XNOR U25226 ( .A(n23180), .B(n23176), .Z(n23179) );
  XOR U25227 ( .A(n23181), .B(nreg[119]), .Z(n23172) );
  IV U25228 ( .A(n23170), .Z(n23181) );
  XOR U25229 ( .A(n23182), .B(n23183), .Z(n23170) );
  AND U25230 ( .A(n23184), .B(n23185), .Z(n23183) );
  XNOR U25231 ( .A(n23182), .B(n11593), .Z(n23185) );
  XNOR U25232 ( .A(n23178), .B(n23180), .Z(n11593) );
  NAND U25233 ( .A(n23186), .B(nreg[118]), .Z(n23180) );
  NAND U25234 ( .A(n12326), .B(nreg[118]), .Z(n23186) );
  XNOR U25235 ( .A(n23176), .B(n23187), .Z(n23178) );
  XOR U25236 ( .A(n23188), .B(n23189), .Z(n23176) );
  AND U25237 ( .A(n23190), .B(n23191), .Z(n23189) );
  XNOR U25238 ( .A(n23192), .B(n23188), .Z(n23191) );
  XOR U25239 ( .A(n23193), .B(nreg[118]), .Z(n23184) );
  IV U25240 ( .A(n23182), .Z(n23193) );
  XOR U25241 ( .A(n23194), .B(n23195), .Z(n23182) );
  AND U25242 ( .A(n23196), .B(n23197), .Z(n23195) );
  XNOR U25243 ( .A(n23194), .B(n11599), .Z(n23197) );
  XNOR U25244 ( .A(n23190), .B(n23192), .Z(n11599) );
  NAND U25245 ( .A(n23198), .B(nreg[117]), .Z(n23192) );
  NAND U25246 ( .A(n12326), .B(nreg[117]), .Z(n23198) );
  XNOR U25247 ( .A(n23188), .B(n23199), .Z(n23190) );
  XOR U25248 ( .A(n23200), .B(n23201), .Z(n23188) );
  AND U25249 ( .A(n23202), .B(n23203), .Z(n23201) );
  XNOR U25250 ( .A(n23204), .B(n23200), .Z(n23203) );
  XOR U25251 ( .A(n23205), .B(nreg[117]), .Z(n23196) );
  IV U25252 ( .A(n23194), .Z(n23205) );
  XOR U25253 ( .A(n23206), .B(n23207), .Z(n23194) );
  AND U25254 ( .A(n23208), .B(n23209), .Z(n23207) );
  XNOR U25255 ( .A(n23206), .B(n11605), .Z(n23209) );
  XNOR U25256 ( .A(n23202), .B(n23204), .Z(n11605) );
  NAND U25257 ( .A(n23210), .B(nreg[116]), .Z(n23204) );
  NAND U25258 ( .A(n12326), .B(nreg[116]), .Z(n23210) );
  XNOR U25259 ( .A(n23200), .B(n23211), .Z(n23202) );
  XOR U25260 ( .A(n23212), .B(n23213), .Z(n23200) );
  AND U25261 ( .A(n23214), .B(n23215), .Z(n23213) );
  XNOR U25262 ( .A(n23216), .B(n23212), .Z(n23215) );
  XOR U25263 ( .A(n23217), .B(nreg[116]), .Z(n23208) );
  IV U25264 ( .A(n23206), .Z(n23217) );
  XOR U25265 ( .A(n23218), .B(n23219), .Z(n23206) );
  AND U25266 ( .A(n23220), .B(n23221), .Z(n23219) );
  XNOR U25267 ( .A(n23218), .B(n11611), .Z(n23221) );
  XNOR U25268 ( .A(n23214), .B(n23216), .Z(n11611) );
  NAND U25269 ( .A(n23222), .B(nreg[115]), .Z(n23216) );
  NAND U25270 ( .A(n12326), .B(nreg[115]), .Z(n23222) );
  XNOR U25271 ( .A(n23212), .B(n23223), .Z(n23214) );
  XOR U25272 ( .A(n23224), .B(n23225), .Z(n23212) );
  AND U25273 ( .A(n23226), .B(n23227), .Z(n23225) );
  XNOR U25274 ( .A(n23228), .B(n23224), .Z(n23227) );
  XOR U25275 ( .A(n23229), .B(nreg[115]), .Z(n23220) );
  IV U25276 ( .A(n23218), .Z(n23229) );
  XOR U25277 ( .A(n23230), .B(n23231), .Z(n23218) );
  AND U25278 ( .A(n23232), .B(n23233), .Z(n23231) );
  XNOR U25279 ( .A(n23230), .B(n11617), .Z(n23233) );
  XNOR U25280 ( .A(n23226), .B(n23228), .Z(n11617) );
  NAND U25281 ( .A(n23234), .B(nreg[114]), .Z(n23228) );
  NAND U25282 ( .A(n12326), .B(nreg[114]), .Z(n23234) );
  XNOR U25283 ( .A(n23224), .B(n23235), .Z(n23226) );
  XOR U25284 ( .A(n23236), .B(n23237), .Z(n23224) );
  AND U25285 ( .A(n23238), .B(n23239), .Z(n23237) );
  XNOR U25286 ( .A(n23240), .B(n23236), .Z(n23239) );
  XOR U25287 ( .A(n23241), .B(nreg[114]), .Z(n23232) );
  IV U25288 ( .A(n23230), .Z(n23241) );
  XOR U25289 ( .A(n23242), .B(n23243), .Z(n23230) );
  AND U25290 ( .A(n23244), .B(n23245), .Z(n23243) );
  XNOR U25291 ( .A(n23242), .B(n11623), .Z(n23245) );
  XNOR U25292 ( .A(n23238), .B(n23240), .Z(n11623) );
  NAND U25293 ( .A(n23246), .B(nreg[113]), .Z(n23240) );
  NAND U25294 ( .A(n12326), .B(nreg[113]), .Z(n23246) );
  XNOR U25295 ( .A(n23236), .B(n23247), .Z(n23238) );
  XOR U25296 ( .A(n23248), .B(n23249), .Z(n23236) );
  AND U25297 ( .A(n23250), .B(n23251), .Z(n23249) );
  XNOR U25298 ( .A(n23252), .B(n23248), .Z(n23251) );
  XOR U25299 ( .A(n23253), .B(nreg[113]), .Z(n23244) );
  IV U25300 ( .A(n23242), .Z(n23253) );
  XOR U25301 ( .A(n23254), .B(n23255), .Z(n23242) );
  AND U25302 ( .A(n23256), .B(n23257), .Z(n23255) );
  XNOR U25303 ( .A(n23254), .B(n11629), .Z(n23257) );
  XNOR U25304 ( .A(n23250), .B(n23252), .Z(n11629) );
  NAND U25305 ( .A(n23258), .B(nreg[112]), .Z(n23252) );
  NAND U25306 ( .A(n12326), .B(nreg[112]), .Z(n23258) );
  XNOR U25307 ( .A(n23248), .B(n23259), .Z(n23250) );
  XOR U25308 ( .A(n23260), .B(n23261), .Z(n23248) );
  AND U25309 ( .A(n23262), .B(n23263), .Z(n23261) );
  XNOR U25310 ( .A(n23264), .B(n23260), .Z(n23263) );
  XOR U25311 ( .A(n23265), .B(nreg[112]), .Z(n23256) );
  IV U25312 ( .A(n23254), .Z(n23265) );
  XOR U25313 ( .A(n23266), .B(n23267), .Z(n23254) );
  AND U25314 ( .A(n23268), .B(n23269), .Z(n23267) );
  XNOR U25315 ( .A(n23266), .B(n11635), .Z(n23269) );
  XNOR U25316 ( .A(n23262), .B(n23264), .Z(n11635) );
  NAND U25317 ( .A(n23270), .B(nreg[111]), .Z(n23264) );
  NAND U25318 ( .A(n12326), .B(nreg[111]), .Z(n23270) );
  XNOR U25319 ( .A(n23260), .B(n23271), .Z(n23262) );
  XOR U25320 ( .A(n23272), .B(n23273), .Z(n23260) );
  AND U25321 ( .A(n23274), .B(n23275), .Z(n23273) );
  XNOR U25322 ( .A(n23276), .B(n23272), .Z(n23275) );
  XOR U25323 ( .A(n23277), .B(nreg[111]), .Z(n23268) );
  IV U25324 ( .A(n23266), .Z(n23277) );
  XOR U25325 ( .A(n23278), .B(n23279), .Z(n23266) );
  AND U25326 ( .A(n23280), .B(n23281), .Z(n23279) );
  XNOR U25327 ( .A(n23278), .B(n11641), .Z(n23281) );
  XNOR U25328 ( .A(n23274), .B(n23276), .Z(n11641) );
  NAND U25329 ( .A(n23282), .B(nreg[110]), .Z(n23276) );
  NAND U25330 ( .A(n12326), .B(nreg[110]), .Z(n23282) );
  XNOR U25331 ( .A(n23272), .B(n23283), .Z(n23274) );
  XOR U25332 ( .A(n23284), .B(n23285), .Z(n23272) );
  AND U25333 ( .A(n23286), .B(n23287), .Z(n23285) );
  XNOR U25334 ( .A(n23288), .B(n23284), .Z(n23287) );
  XOR U25335 ( .A(n23289), .B(nreg[110]), .Z(n23280) );
  IV U25336 ( .A(n23278), .Z(n23289) );
  XOR U25337 ( .A(n23290), .B(n23291), .Z(n23278) );
  AND U25338 ( .A(n23292), .B(n23293), .Z(n23291) );
  XNOR U25339 ( .A(n23290), .B(n11647), .Z(n23293) );
  XNOR U25340 ( .A(n23286), .B(n23288), .Z(n11647) );
  NAND U25341 ( .A(n23294), .B(nreg[109]), .Z(n23288) );
  NAND U25342 ( .A(n12326), .B(nreg[109]), .Z(n23294) );
  XNOR U25343 ( .A(n23284), .B(n23295), .Z(n23286) );
  XOR U25344 ( .A(n23296), .B(n23297), .Z(n23284) );
  AND U25345 ( .A(n23298), .B(n23299), .Z(n23297) );
  XNOR U25346 ( .A(n23300), .B(n23296), .Z(n23299) );
  XOR U25347 ( .A(n23301), .B(nreg[109]), .Z(n23292) );
  IV U25348 ( .A(n23290), .Z(n23301) );
  XOR U25349 ( .A(n23302), .B(n23303), .Z(n23290) );
  AND U25350 ( .A(n23304), .B(n23305), .Z(n23303) );
  XNOR U25351 ( .A(n23302), .B(n11653), .Z(n23305) );
  XNOR U25352 ( .A(n23298), .B(n23300), .Z(n11653) );
  NAND U25353 ( .A(n23306), .B(nreg[108]), .Z(n23300) );
  NAND U25354 ( .A(n12326), .B(nreg[108]), .Z(n23306) );
  XNOR U25355 ( .A(n23296), .B(n23307), .Z(n23298) );
  XOR U25356 ( .A(n23308), .B(n23309), .Z(n23296) );
  AND U25357 ( .A(n23310), .B(n23311), .Z(n23309) );
  XNOR U25358 ( .A(n23312), .B(n23308), .Z(n23311) );
  XOR U25359 ( .A(n23313), .B(nreg[108]), .Z(n23304) );
  IV U25360 ( .A(n23302), .Z(n23313) );
  XOR U25361 ( .A(n23314), .B(n23315), .Z(n23302) );
  AND U25362 ( .A(n23316), .B(n23317), .Z(n23315) );
  XNOR U25363 ( .A(n23314), .B(n11659), .Z(n23317) );
  XNOR U25364 ( .A(n23310), .B(n23312), .Z(n11659) );
  NAND U25365 ( .A(n23318), .B(nreg[107]), .Z(n23312) );
  NAND U25366 ( .A(n12326), .B(nreg[107]), .Z(n23318) );
  XNOR U25367 ( .A(n23308), .B(n23319), .Z(n23310) );
  XOR U25368 ( .A(n23320), .B(n23321), .Z(n23308) );
  AND U25369 ( .A(n23322), .B(n23323), .Z(n23321) );
  XNOR U25370 ( .A(n23324), .B(n23320), .Z(n23323) );
  XOR U25371 ( .A(n23325), .B(nreg[107]), .Z(n23316) );
  IV U25372 ( .A(n23314), .Z(n23325) );
  XOR U25373 ( .A(n23326), .B(n23327), .Z(n23314) );
  AND U25374 ( .A(n23328), .B(n23329), .Z(n23327) );
  XNOR U25375 ( .A(n23326), .B(n11665), .Z(n23329) );
  XNOR U25376 ( .A(n23322), .B(n23324), .Z(n11665) );
  NAND U25377 ( .A(n23330), .B(nreg[106]), .Z(n23324) );
  NAND U25378 ( .A(n12326), .B(nreg[106]), .Z(n23330) );
  XNOR U25379 ( .A(n23320), .B(n23331), .Z(n23322) );
  XOR U25380 ( .A(n23332), .B(n23333), .Z(n23320) );
  AND U25381 ( .A(n23334), .B(n23335), .Z(n23333) );
  XNOR U25382 ( .A(n23336), .B(n23332), .Z(n23335) );
  XOR U25383 ( .A(n23337), .B(nreg[106]), .Z(n23328) );
  IV U25384 ( .A(n23326), .Z(n23337) );
  XOR U25385 ( .A(n23338), .B(n23339), .Z(n23326) );
  AND U25386 ( .A(n23340), .B(n23341), .Z(n23339) );
  XNOR U25387 ( .A(n23338), .B(n11671), .Z(n23341) );
  XNOR U25388 ( .A(n23334), .B(n23336), .Z(n11671) );
  NAND U25389 ( .A(n23342), .B(nreg[105]), .Z(n23336) );
  NAND U25390 ( .A(n12326), .B(nreg[105]), .Z(n23342) );
  XNOR U25391 ( .A(n23332), .B(n23343), .Z(n23334) );
  XOR U25392 ( .A(n23344), .B(n23345), .Z(n23332) );
  AND U25393 ( .A(n23346), .B(n23347), .Z(n23345) );
  XNOR U25394 ( .A(n23348), .B(n23344), .Z(n23347) );
  XOR U25395 ( .A(n23349), .B(nreg[105]), .Z(n23340) );
  IV U25396 ( .A(n23338), .Z(n23349) );
  XOR U25397 ( .A(n23350), .B(n23351), .Z(n23338) );
  AND U25398 ( .A(n23352), .B(n23353), .Z(n23351) );
  XNOR U25399 ( .A(n23350), .B(n11677), .Z(n23353) );
  XNOR U25400 ( .A(n23346), .B(n23348), .Z(n11677) );
  NAND U25401 ( .A(n23354), .B(nreg[104]), .Z(n23348) );
  NAND U25402 ( .A(n12326), .B(nreg[104]), .Z(n23354) );
  XNOR U25403 ( .A(n23344), .B(n23355), .Z(n23346) );
  XOR U25404 ( .A(n23356), .B(n23357), .Z(n23344) );
  AND U25405 ( .A(n23358), .B(n23359), .Z(n23357) );
  XNOR U25406 ( .A(n23360), .B(n23356), .Z(n23359) );
  XOR U25407 ( .A(n23361), .B(nreg[104]), .Z(n23352) );
  IV U25408 ( .A(n23350), .Z(n23361) );
  XOR U25409 ( .A(n23362), .B(n23363), .Z(n23350) );
  AND U25410 ( .A(n23364), .B(n23365), .Z(n23363) );
  XNOR U25411 ( .A(n23362), .B(n11683), .Z(n23365) );
  XNOR U25412 ( .A(n23358), .B(n23360), .Z(n11683) );
  NAND U25413 ( .A(n23366), .B(nreg[103]), .Z(n23360) );
  NAND U25414 ( .A(n12326), .B(nreg[103]), .Z(n23366) );
  XNOR U25415 ( .A(n23356), .B(n23367), .Z(n23358) );
  XOR U25416 ( .A(n23368), .B(n23369), .Z(n23356) );
  AND U25417 ( .A(n23370), .B(n23371), .Z(n23369) );
  XNOR U25418 ( .A(n23372), .B(n23368), .Z(n23371) );
  XOR U25419 ( .A(n23373), .B(nreg[103]), .Z(n23364) );
  IV U25420 ( .A(n23362), .Z(n23373) );
  XOR U25421 ( .A(n23374), .B(n23375), .Z(n23362) );
  AND U25422 ( .A(n23376), .B(n23377), .Z(n23375) );
  XNOR U25423 ( .A(n23374), .B(n11689), .Z(n23377) );
  XNOR U25424 ( .A(n23370), .B(n23372), .Z(n11689) );
  NAND U25425 ( .A(n23378), .B(nreg[102]), .Z(n23372) );
  NAND U25426 ( .A(n12326), .B(nreg[102]), .Z(n23378) );
  XNOR U25427 ( .A(n23368), .B(n23379), .Z(n23370) );
  XOR U25428 ( .A(n23380), .B(n23381), .Z(n23368) );
  AND U25429 ( .A(n23382), .B(n23383), .Z(n23381) );
  XNOR U25430 ( .A(n23384), .B(n23380), .Z(n23383) );
  XOR U25431 ( .A(n23385), .B(nreg[102]), .Z(n23376) );
  IV U25432 ( .A(n23374), .Z(n23385) );
  XOR U25433 ( .A(n23386), .B(n23387), .Z(n23374) );
  AND U25434 ( .A(n23388), .B(n23389), .Z(n23387) );
  XNOR U25435 ( .A(n23386), .B(n11695), .Z(n23389) );
  XNOR U25436 ( .A(n23382), .B(n23384), .Z(n11695) );
  NAND U25437 ( .A(n23390), .B(nreg[101]), .Z(n23384) );
  NAND U25438 ( .A(n12326), .B(nreg[101]), .Z(n23390) );
  XNOR U25439 ( .A(n23380), .B(n23391), .Z(n23382) );
  XOR U25440 ( .A(n23392), .B(n23393), .Z(n23380) );
  AND U25441 ( .A(n23394), .B(n23395), .Z(n23393) );
  XNOR U25442 ( .A(n23396), .B(n23392), .Z(n23395) );
  XOR U25443 ( .A(n23397), .B(nreg[101]), .Z(n23388) );
  IV U25444 ( .A(n23386), .Z(n23397) );
  XOR U25445 ( .A(n23398), .B(n23399), .Z(n23386) );
  AND U25446 ( .A(n23400), .B(n23401), .Z(n23399) );
  XNOR U25447 ( .A(n23398), .B(n11701), .Z(n23401) );
  XNOR U25448 ( .A(n23394), .B(n23396), .Z(n11701) );
  NAND U25449 ( .A(n23402), .B(nreg[100]), .Z(n23396) );
  NAND U25450 ( .A(n12326), .B(nreg[100]), .Z(n23402) );
  XNOR U25451 ( .A(n23392), .B(n23403), .Z(n23394) );
  XOR U25452 ( .A(n23404), .B(n23405), .Z(n23392) );
  AND U25453 ( .A(n23406), .B(n23407), .Z(n23405) );
  XNOR U25454 ( .A(n23408), .B(n23404), .Z(n23407) );
  XOR U25455 ( .A(n23409), .B(nreg[100]), .Z(n23400) );
  IV U25456 ( .A(n23398), .Z(n23409) );
  XOR U25457 ( .A(n23410), .B(n23411), .Z(n23398) );
  AND U25458 ( .A(n23412), .B(n23413), .Z(n23411) );
  XNOR U25459 ( .A(n23410), .B(n11707), .Z(n23413) );
  XNOR U25460 ( .A(n23406), .B(n23408), .Z(n11707) );
  NAND U25461 ( .A(n23414), .B(nreg[99]), .Z(n23408) );
  NAND U25462 ( .A(n12326), .B(nreg[99]), .Z(n23414) );
  XNOR U25463 ( .A(n23404), .B(n23415), .Z(n23406) );
  XOR U25464 ( .A(n23416), .B(n23417), .Z(n23404) );
  AND U25465 ( .A(n23418), .B(n23419), .Z(n23417) );
  XNOR U25466 ( .A(n23420), .B(n23416), .Z(n23419) );
  XOR U25467 ( .A(n23421), .B(nreg[99]), .Z(n23412) );
  IV U25468 ( .A(n23410), .Z(n23421) );
  XOR U25469 ( .A(n23422), .B(n23423), .Z(n23410) );
  AND U25470 ( .A(n23424), .B(n23425), .Z(n23423) );
  XNOR U25471 ( .A(n23422), .B(n11713), .Z(n23425) );
  XNOR U25472 ( .A(n23418), .B(n23420), .Z(n11713) );
  NAND U25473 ( .A(n23426), .B(nreg[98]), .Z(n23420) );
  NAND U25474 ( .A(n12326), .B(nreg[98]), .Z(n23426) );
  XNOR U25475 ( .A(n23416), .B(n23427), .Z(n23418) );
  XOR U25476 ( .A(n23428), .B(n23429), .Z(n23416) );
  AND U25477 ( .A(n23430), .B(n23431), .Z(n23429) );
  XNOR U25478 ( .A(n23432), .B(n23428), .Z(n23431) );
  XOR U25479 ( .A(n23433), .B(nreg[98]), .Z(n23424) );
  IV U25480 ( .A(n23422), .Z(n23433) );
  XOR U25481 ( .A(n23434), .B(n23435), .Z(n23422) );
  AND U25482 ( .A(n23436), .B(n23437), .Z(n23435) );
  XNOR U25483 ( .A(n23434), .B(n11722), .Z(n23437) );
  XNOR U25484 ( .A(n23430), .B(n23432), .Z(n11722) );
  NAND U25485 ( .A(n23438), .B(nreg[97]), .Z(n23432) );
  NAND U25486 ( .A(n12326), .B(nreg[97]), .Z(n23438) );
  XNOR U25487 ( .A(n23428), .B(n23439), .Z(n23430) );
  XOR U25488 ( .A(n23440), .B(n23441), .Z(n23428) );
  AND U25489 ( .A(n23442), .B(n23443), .Z(n23441) );
  XNOR U25490 ( .A(n23444), .B(n23440), .Z(n23443) );
  XOR U25491 ( .A(n23445), .B(nreg[97]), .Z(n23436) );
  IV U25492 ( .A(n23434), .Z(n23445) );
  XOR U25493 ( .A(n23446), .B(n23447), .Z(n23434) );
  AND U25494 ( .A(n23448), .B(n23449), .Z(n23447) );
  XNOR U25495 ( .A(n23446), .B(n11727), .Z(n23449) );
  XNOR U25496 ( .A(n23442), .B(n23444), .Z(n11727) );
  NAND U25497 ( .A(n23450), .B(nreg[96]), .Z(n23444) );
  NAND U25498 ( .A(n12326), .B(nreg[96]), .Z(n23450) );
  XNOR U25499 ( .A(n23440), .B(n23451), .Z(n23442) );
  XOR U25500 ( .A(n23452), .B(n23453), .Z(n23440) );
  AND U25501 ( .A(n23454), .B(n23455), .Z(n23453) );
  XNOR U25502 ( .A(n23456), .B(n23452), .Z(n23455) );
  XOR U25503 ( .A(n23457), .B(nreg[96]), .Z(n23448) );
  IV U25504 ( .A(n23446), .Z(n23457) );
  XOR U25505 ( .A(n23458), .B(n23459), .Z(n23446) );
  AND U25506 ( .A(n23460), .B(n23461), .Z(n23459) );
  XNOR U25507 ( .A(n23458), .B(n11733), .Z(n23461) );
  XNOR U25508 ( .A(n23454), .B(n23456), .Z(n11733) );
  NAND U25509 ( .A(n23462), .B(nreg[95]), .Z(n23456) );
  NAND U25510 ( .A(n12326), .B(nreg[95]), .Z(n23462) );
  XNOR U25511 ( .A(n23452), .B(n23463), .Z(n23454) );
  XOR U25512 ( .A(n23464), .B(n23465), .Z(n23452) );
  AND U25513 ( .A(n23466), .B(n23467), .Z(n23465) );
  XNOR U25514 ( .A(n23468), .B(n23464), .Z(n23467) );
  XOR U25515 ( .A(n23469), .B(nreg[95]), .Z(n23460) );
  IV U25516 ( .A(n23458), .Z(n23469) );
  XOR U25517 ( .A(n23470), .B(n23471), .Z(n23458) );
  AND U25518 ( .A(n23472), .B(n23473), .Z(n23471) );
  XNOR U25519 ( .A(n23470), .B(n11739), .Z(n23473) );
  XNOR U25520 ( .A(n23466), .B(n23468), .Z(n11739) );
  NAND U25521 ( .A(n23474), .B(nreg[94]), .Z(n23468) );
  NAND U25522 ( .A(n12326), .B(nreg[94]), .Z(n23474) );
  XNOR U25523 ( .A(n23464), .B(n23475), .Z(n23466) );
  XOR U25524 ( .A(n23476), .B(n23477), .Z(n23464) );
  AND U25525 ( .A(n23478), .B(n23479), .Z(n23477) );
  XNOR U25526 ( .A(n23480), .B(n23476), .Z(n23479) );
  XOR U25527 ( .A(n23481), .B(nreg[94]), .Z(n23472) );
  IV U25528 ( .A(n23470), .Z(n23481) );
  XOR U25529 ( .A(n23482), .B(n23483), .Z(n23470) );
  AND U25530 ( .A(n23484), .B(n23485), .Z(n23483) );
  XNOR U25531 ( .A(n23482), .B(n11745), .Z(n23485) );
  XNOR U25532 ( .A(n23478), .B(n23480), .Z(n11745) );
  NAND U25533 ( .A(n23486), .B(nreg[93]), .Z(n23480) );
  NAND U25534 ( .A(n12326), .B(nreg[93]), .Z(n23486) );
  XNOR U25535 ( .A(n23476), .B(n23487), .Z(n23478) );
  XOR U25536 ( .A(n23488), .B(n23489), .Z(n23476) );
  AND U25537 ( .A(n23490), .B(n23491), .Z(n23489) );
  XNOR U25538 ( .A(n23492), .B(n23488), .Z(n23491) );
  XOR U25539 ( .A(n23493), .B(nreg[93]), .Z(n23484) );
  IV U25540 ( .A(n23482), .Z(n23493) );
  XOR U25541 ( .A(n23494), .B(n23495), .Z(n23482) );
  AND U25542 ( .A(n23496), .B(n23497), .Z(n23495) );
  XNOR U25543 ( .A(n23494), .B(n11751), .Z(n23497) );
  XNOR U25544 ( .A(n23490), .B(n23492), .Z(n11751) );
  NAND U25545 ( .A(n23498), .B(nreg[92]), .Z(n23492) );
  NAND U25546 ( .A(n12326), .B(nreg[92]), .Z(n23498) );
  XNOR U25547 ( .A(n23488), .B(n23499), .Z(n23490) );
  XOR U25548 ( .A(n23500), .B(n23501), .Z(n23488) );
  AND U25549 ( .A(n23502), .B(n23503), .Z(n23501) );
  XNOR U25550 ( .A(n23504), .B(n23500), .Z(n23503) );
  XOR U25551 ( .A(n23505), .B(nreg[92]), .Z(n23496) );
  IV U25552 ( .A(n23494), .Z(n23505) );
  XOR U25553 ( .A(n23506), .B(n23507), .Z(n23494) );
  AND U25554 ( .A(n23508), .B(n23509), .Z(n23507) );
  XNOR U25555 ( .A(n23506), .B(n11757), .Z(n23509) );
  XNOR U25556 ( .A(n23502), .B(n23504), .Z(n11757) );
  NAND U25557 ( .A(n23510), .B(nreg[91]), .Z(n23504) );
  NAND U25558 ( .A(n12326), .B(nreg[91]), .Z(n23510) );
  XNOR U25559 ( .A(n23500), .B(n23511), .Z(n23502) );
  XOR U25560 ( .A(n23512), .B(n23513), .Z(n23500) );
  AND U25561 ( .A(n23514), .B(n23515), .Z(n23513) );
  XNOR U25562 ( .A(n23516), .B(n23512), .Z(n23515) );
  XOR U25563 ( .A(n23517), .B(nreg[91]), .Z(n23508) );
  IV U25564 ( .A(n23506), .Z(n23517) );
  XOR U25565 ( .A(n23518), .B(n23519), .Z(n23506) );
  AND U25566 ( .A(n23520), .B(n23521), .Z(n23519) );
  XNOR U25567 ( .A(n23518), .B(n11763), .Z(n23521) );
  XNOR U25568 ( .A(n23514), .B(n23516), .Z(n11763) );
  NAND U25569 ( .A(n23522), .B(nreg[90]), .Z(n23516) );
  NAND U25570 ( .A(n12326), .B(nreg[90]), .Z(n23522) );
  XNOR U25571 ( .A(n23512), .B(n23523), .Z(n23514) );
  XOR U25572 ( .A(n23524), .B(n23525), .Z(n23512) );
  AND U25573 ( .A(n23526), .B(n23527), .Z(n23525) );
  XNOR U25574 ( .A(n23528), .B(n23524), .Z(n23527) );
  XOR U25575 ( .A(n23529), .B(nreg[90]), .Z(n23520) );
  IV U25576 ( .A(n23518), .Z(n23529) );
  XOR U25577 ( .A(n23530), .B(n23531), .Z(n23518) );
  AND U25578 ( .A(n23532), .B(n23533), .Z(n23531) );
  XNOR U25579 ( .A(n23530), .B(n11769), .Z(n23533) );
  XNOR U25580 ( .A(n23526), .B(n23528), .Z(n11769) );
  NAND U25581 ( .A(n23534), .B(nreg[89]), .Z(n23528) );
  NAND U25582 ( .A(n12326), .B(nreg[89]), .Z(n23534) );
  XNOR U25583 ( .A(n23524), .B(n23535), .Z(n23526) );
  XOR U25584 ( .A(n23536), .B(n23537), .Z(n23524) );
  AND U25585 ( .A(n23538), .B(n23539), .Z(n23537) );
  XNOR U25586 ( .A(n23540), .B(n23536), .Z(n23539) );
  XOR U25587 ( .A(n23541), .B(nreg[89]), .Z(n23532) );
  IV U25588 ( .A(n23530), .Z(n23541) );
  XOR U25589 ( .A(n23542), .B(n23543), .Z(n23530) );
  AND U25590 ( .A(n23544), .B(n23545), .Z(n23543) );
  XNOR U25591 ( .A(n23542), .B(n11775), .Z(n23545) );
  XNOR U25592 ( .A(n23538), .B(n23540), .Z(n11775) );
  NAND U25593 ( .A(n23546), .B(nreg[88]), .Z(n23540) );
  NAND U25594 ( .A(n12326), .B(nreg[88]), .Z(n23546) );
  XNOR U25595 ( .A(n23536), .B(n23547), .Z(n23538) );
  XOR U25596 ( .A(n23548), .B(n23549), .Z(n23536) );
  AND U25597 ( .A(n23550), .B(n23551), .Z(n23549) );
  XNOR U25598 ( .A(n23552), .B(n23548), .Z(n23551) );
  XOR U25599 ( .A(n23553), .B(nreg[88]), .Z(n23544) );
  IV U25600 ( .A(n23542), .Z(n23553) );
  XOR U25601 ( .A(n23554), .B(n23555), .Z(n23542) );
  AND U25602 ( .A(n23556), .B(n23557), .Z(n23555) );
  XNOR U25603 ( .A(n23554), .B(n11781), .Z(n23557) );
  XNOR U25604 ( .A(n23550), .B(n23552), .Z(n11781) );
  NAND U25605 ( .A(n23558), .B(nreg[87]), .Z(n23552) );
  NAND U25606 ( .A(n12326), .B(nreg[87]), .Z(n23558) );
  XNOR U25607 ( .A(n23548), .B(n23559), .Z(n23550) );
  XOR U25608 ( .A(n23560), .B(n23561), .Z(n23548) );
  AND U25609 ( .A(n23562), .B(n23563), .Z(n23561) );
  XNOR U25610 ( .A(n23564), .B(n23560), .Z(n23563) );
  XOR U25611 ( .A(n23565), .B(nreg[87]), .Z(n23556) );
  IV U25612 ( .A(n23554), .Z(n23565) );
  XOR U25613 ( .A(n23566), .B(n23567), .Z(n23554) );
  AND U25614 ( .A(n23568), .B(n23569), .Z(n23567) );
  XNOR U25615 ( .A(n23566), .B(n11787), .Z(n23569) );
  XNOR U25616 ( .A(n23562), .B(n23564), .Z(n11787) );
  NAND U25617 ( .A(n23570), .B(nreg[86]), .Z(n23564) );
  NAND U25618 ( .A(n12326), .B(nreg[86]), .Z(n23570) );
  XNOR U25619 ( .A(n23560), .B(n23571), .Z(n23562) );
  XOR U25620 ( .A(n23572), .B(n23573), .Z(n23560) );
  AND U25621 ( .A(n23574), .B(n23575), .Z(n23573) );
  XNOR U25622 ( .A(n23576), .B(n23572), .Z(n23575) );
  XOR U25623 ( .A(n23577), .B(nreg[86]), .Z(n23568) );
  IV U25624 ( .A(n23566), .Z(n23577) );
  XOR U25625 ( .A(n23578), .B(n23579), .Z(n23566) );
  AND U25626 ( .A(n23580), .B(n23581), .Z(n23579) );
  XNOR U25627 ( .A(n23578), .B(n11793), .Z(n23581) );
  XNOR U25628 ( .A(n23574), .B(n23576), .Z(n11793) );
  NAND U25629 ( .A(n23582), .B(nreg[85]), .Z(n23576) );
  NAND U25630 ( .A(n12326), .B(nreg[85]), .Z(n23582) );
  XNOR U25631 ( .A(n23572), .B(n23583), .Z(n23574) );
  XOR U25632 ( .A(n23584), .B(n23585), .Z(n23572) );
  AND U25633 ( .A(n23586), .B(n23587), .Z(n23585) );
  XNOR U25634 ( .A(n23588), .B(n23584), .Z(n23587) );
  XOR U25635 ( .A(n23589), .B(nreg[85]), .Z(n23580) );
  IV U25636 ( .A(n23578), .Z(n23589) );
  XOR U25637 ( .A(n23590), .B(n23591), .Z(n23578) );
  AND U25638 ( .A(n23592), .B(n23593), .Z(n23591) );
  XNOR U25639 ( .A(n23590), .B(n11799), .Z(n23593) );
  XNOR U25640 ( .A(n23586), .B(n23588), .Z(n11799) );
  NAND U25641 ( .A(n23594), .B(nreg[84]), .Z(n23588) );
  NAND U25642 ( .A(n12326), .B(nreg[84]), .Z(n23594) );
  XNOR U25643 ( .A(n23584), .B(n23595), .Z(n23586) );
  XOR U25644 ( .A(n23596), .B(n23597), .Z(n23584) );
  AND U25645 ( .A(n23598), .B(n23599), .Z(n23597) );
  XNOR U25646 ( .A(n23600), .B(n23596), .Z(n23599) );
  XOR U25647 ( .A(n23601), .B(nreg[84]), .Z(n23592) );
  IV U25648 ( .A(n23590), .Z(n23601) );
  XOR U25649 ( .A(n23602), .B(n23603), .Z(n23590) );
  AND U25650 ( .A(n23604), .B(n23605), .Z(n23603) );
  XNOR U25651 ( .A(n23602), .B(n11805), .Z(n23605) );
  XNOR U25652 ( .A(n23598), .B(n23600), .Z(n11805) );
  NAND U25653 ( .A(n23606), .B(nreg[83]), .Z(n23600) );
  NAND U25654 ( .A(n12326), .B(nreg[83]), .Z(n23606) );
  XNOR U25655 ( .A(n23596), .B(n23607), .Z(n23598) );
  XOR U25656 ( .A(n23608), .B(n23609), .Z(n23596) );
  AND U25657 ( .A(n23610), .B(n23611), .Z(n23609) );
  XNOR U25658 ( .A(n23612), .B(n23608), .Z(n23611) );
  XOR U25659 ( .A(n23613), .B(nreg[83]), .Z(n23604) );
  IV U25660 ( .A(n23602), .Z(n23613) );
  XOR U25661 ( .A(n23614), .B(n23615), .Z(n23602) );
  AND U25662 ( .A(n23616), .B(n23617), .Z(n23615) );
  XNOR U25663 ( .A(n23614), .B(n11811), .Z(n23617) );
  XNOR U25664 ( .A(n23610), .B(n23612), .Z(n11811) );
  NAND U25665 ( .A(n23618), .B(nreg[82]), .Z(n23612) );
  NAND U25666 ( .A(n12326), .B(nreg[82]), .Z(n23618) );
  XNOR U25667 ( .A(n23608), .B(n23619), .Z(n23610) );
  XOR U25668 ( .A(n23620), .B(n23621), .Z(n23608) );
  AND U25669 ( .A(n23622), .B(n23623), .Z(n23621) );
  XNOR U25670 ( .A(n23624), .B(n23620), .Z(n23623) );
  XOR U25671 ( .A(n23625), .B(nreg[82]), .Z(n23616) );
  IV U25672 ( .A(n23614), .Z(n23625) );
  XOR U25673 ( .A(n23626), .B(n23627), .Z(n23614) );
  AND U25674 ( .A(n23628), .B(n23629), .Z(n23627) );
  XNOR U25675 ( .A(n23626), .B(n11817), .Z(n23629) );
  XNOR U25676 ( .A(n23622), .B(n23624), .Z(n11817) );
  NAND U25677 ( .A(n23630), .B(nreg[81]), .Z(n23624) );
  NAND U25678 ( .A(n12326), .B(nreg[81]), .Z(n23630) );
  XNOR U25679 ( .A(n23620), .B(n23631), .Z(n23622) );
  XOR U25680 ( .A(n23632), .B(n23633), .Z(n23620) );
  AND U25681 ( .A(n23634), .B(n23635), .Z(n23633) );
  XNOR U25682 ( .A(n23636), .B(n23632), .Z(n23635) );
  XOR U25683 ( .A(n23637), .B(nreg[81]), .Z(n23628) );
  IV U25684 ( .A(n23626), .Z(n23637) );
  XOR U25685 ( .A(n23638), .B(n23639), .Z(n23626) );
  AND U25686 ( .A(n23640), .B(n23641), .Z(n23639) );
  XNOR U25687 ( .A(n23638), .B(n11823), .Z(n23641) );
  XNOR U25688 ( .A(n23634), .B(n23636), .Z(n11823) );
  NAND U25689 ( .A(n23642), .B(nreg[80]), .Z(n23636) );
  NAND U25690 ( .A(n12326), .B(nreg[80]), .Z(n23642) );
  XNOR U25691 ( .A(n23632), .B(n23643), .Z(n23634) );
  XOR U25692 ( .A(n23644), .B(n23645), .Z(n23632) );
  AND U25693 ( .A(n23646), .B(n23647), .Z(n23645) );
  XNOR U25694 ( .A(n23648), .B(n23644), .Z(n23647) );
  XOR U25695 ( .A(n23649), .B(nreg[80]), .Z(n23640) );
  IV U25696 ( .A(n23638), .Z(n23649) );
  XOR U25697 ( .A(n23650), .B(n23651), .Z(n23638) );
  AND U25698 ( .A(n23652), .B(n23653), .Z(n23651) );
  XNOR U25699 ( .A(n23650), .B(n11829), .Z(n23653) );
  XNOR U25700 ( .A(n23646), .B(n23648), .Z(n11829) );
  NAND U25701 ( .A(n23654), .B(nreg[79]), .Z(n23648) );
  NAND U25702 ( .A(n12326), .B(nreg[79]), .Z(n23654) );
  XNOR U25703 ( .A(n23644), .B(n23655), .Z(n23646) );
  XOR U25704 ( .A(n23656), .B(n23657), .Z(n23644) );
  AND U25705 ( .A(n23658), .B(n23659), .Z(n23657) );
  XNOR U25706 ( .A(n23660), .B(n23656), .Z(n23659) );
  XOR U25707 ( .A(n23661), .B(nreg[79]), .Z(n23652) );
  IV U25708 ( .A(n23650), .Z(n23661) );
  XOR U25709 ( .A(n23662), .B(n23663), .Z(n23650) );
  AND U25710 ( .A(n23664), .B(n23665), .Z(n23663) );
  XNOR U25711 ( .A(n23662), .B(n11835), .Z(n23665) );
  XNOR U25712 ( .A(n23658), .B(n23660), .Z(n11835) );
  NAND U25713 ( .A(n23666), .B(nreg[78]), .Z(n23660) );
  NAND U25714 ( .A(n12326), .B(nreg[78]), .Z(n23666) );
  XNOR U25715 ( .A(n23656), .B(n23667), .Z(n23658) );
  XOR U25716 ( .A(n23668), .B(n23669), .Z(n23656) );
  AND U25717 ( .A(n23670), .B(n23671), .Z(n23669) );
  XNOR U25718 ( .A(n23672), .B(n23668), .Z(n23671) );
  XOR U25719 ( .A(n23673), .B(nreg[78]), .Z(n23664) );
  IV U25720 ( .A(n23662), .Z(n23673) );
  XOR U25721 ( .A(n23674), .B(n23675), .Z(n23662) );
  AND U25722 ( .A(n23676), .B(n23677), .Z(n23675) );
  XNOR U25723 ( .A(n23674), .B(n11841), .Z(n23677) );
  XNOR U25724 ( .A(n23670), .B(n23672), .Z(n11841) );
  NAND U25725 ( .A(n23678), .B(nreg[77]), .Z(n23672) );
  NAND U25726 ( .A(n12326), .B(nreg[77]), .Z(n23678) );
  XNOR U25727 ( .A(n23668), .B(n23679), .Z(n23670) );
  XOR U25728 ( .A(n23680), .B(n23681), .Z(n23668) );
  AND U25729 ( .A(n23682), .B(n23683), .Z(n23681) );
  XNOR U25730 ( .A(n23684), .B(n23680), .Z(n23683) );
  XOR U25731 ( .A(n23685), .B(nreg[77]), .Z(n23676) );
  IV U25732 ( .A(n23674), .Z(n23685) );
  XOR U25733 ( .A(n23686), .B(n23687), .Z(n23674) );
  AND U25734 ( .A(n23688), .B(n23689), .Z(n23687) );
  XNOR U25735 ( .A(n23686), .B(n11847), .Z(n23689) );
  XNOR U25736 ( .A(n23682), .B(n23684), .Z(n11847) );
  NAND U25737 ( .A(n23690), .B(nreg[76]), .Z(n23684) );
  NAND U25738 ( .A(n12326), .B(nreg[76]), .Z(n23690) );
  XNOR U25739 ( .A(n23680), .B(n23691), .Z(n23682) );
  XOR U25740 ( .A(n23692), .B(n23693), .Z(n23680) );
  AND U25741 ( .A(n23694), .B(n23695), .Z(n23693) );
  XNOR U25742 ( .A(n23696), .B(n23692), .Z(n23695) );
  XOR U25743 ( .A(n23697), .B(nreg[76]), .Z(n23688) );
  IV U25744 ( .A(n23686), .Z(n23697) );
  XOR U25745 ( .A(n23698), .B(n23699), .Z(n23686) );
  AND U25746 ( .A(n23700), .B(n23701), .Z(n23699) );
  XNOR U25747 ( .A(n23698), .B(n11853), .Z(n23701) );
  XNOR U25748 ( .A(n23694), .B(n23696), .Z(n11853) );
  NAND U25749 ( .A(n23702), .B(nreg[75]), .Z(n23696) );
  NAND U25750 ( .A(n12326), .B(nreg[75]), .Z(n23702) );
  XNOR U25751 ( .A(n23692), .B(n23703), .Z(n23694) );
  XOR U25752 ( .A(n23704), .B(n23705), .Z(n23692) );
  AND U25753 ( .A(n23706), .B(n23707), .Z(n23705) );
  XNOR U25754 ( .A(n23708), .B(n23704), .Z(n23707) );
  XOR U25755 ( .A(n23709), .B(nreg[75]), .Z(n23700) );
  IV U25756 ( .A(n23698), .Z(n23709) );
  XOR U25757 ( .A(n23710), .B(n23711), .Z(n23698) );
  AND U25758 ( .A(n23712), .B(n23713), .Z(n23711) );
  XNOR U25759 ( .A(n23710), .B(n11859), .Z(n23713) );
  XNOR U25760 ( .A(n23706), .B(n23708), .Z(n11859) );
  NAND U25761 ( .A(n23714), .B(nreg[74]), .Z(n23708) );
  NAND U25762 ( .A(n12326), .B(nreg[74]), .Z(n23714) );
  XNOR U25763 ( .A(n23704), .B(n23715), .Z(n23706) );
  XOR U25764 ( .A(n23716), .B(n23717), .Z(n23704) );
  AND U25765 ( .A(n23718), .B(n23719), .Z(n23717) );
  XNOR U25766 ( .A(n23720), .B(n23716), .Z(n23719) );
  XOR U25767 ( .A(n23721), .B(nreg[74]), .Z(n23712) );
  IV U25768 ( .A(n23710), .Z(n23721) );
  XOR U25769 ( .A(n23722), .B(n23723), .Z(n23710) );
  AND U25770 ( .A(n23724), .B(n23725), .Z(n23723) );
  XNOR U25771 ( .A(n23722), .B(n11865), .Z(n23725) );
  XNOR U25772 ( .A(n23718), .B(n23720), .Z(n11865) );
  NAND U25773 ( .A(n23726), .B(nreg[73]), .Z(n23720) );
  NAND U25774 ( .A(n12326), .B(nreg[73]), .Z(n23726) );
  XNOR U25775 ( .A(n23716), .B(n23727), .Z(n23718) );
  XOR U25776 ( .A(n23728), .B(n23729), .Z(n23716) );
  AND U25777 ( .A(n23730), .B(n23731), .Z(n23729) );
  XNOR U25778 ( .A(n23732), .B(n23728), .Z(n23731) );
  XOR U25779 ( .A(n23733), .B(nreg[73]), .Z(n23724) );
  IV U25780 ( .A(n23722), .Z(n23733) );
  XOR U25781 ( .A(n23734), .B(n23735), .Z(n23722) );
  AND U25782 ( .A(n23736), .B(n23737), .Z(n23735) );
  XNOR U25783 ( .A(n23734), .B(n11871), .Z(n23737) );
  XNOR U25784 ( .A(n23730), .B(n23732), .Z(n11871) );
  NAND U25785 ( .A(n23738), .B(nreg[72]), .Z(n23732) );
  NAND U25786 ( .A(n12326), .B(nreg[72]), .Z(n23738) );
  XNOR U25787 ( .A(n23728), .B(n23739), .Z(n23730) );
  XOR U25788 ( .A(n23740), .B(n23741), .Z(n23728) );
  AND U25789 ( .A(n23742), .B(n23743), .Z(n23741) );
  XNOR U25790 ( .A(n23744), .B(n23740), .Z(n23743) );
  XOR U25791 ( .A(n23745), .B(nreg[72]), .Z(n23736) );
  IV U25792 ( .A(n23734), .Z(n23745) );
  XOR U25793 ( .A(n23746), .B(n23747), .Z(n23734) );
  AND U25794 ( .A(n23748), .B(n23749), .Z(n23747) );
  XNOR U25795 ( .A(n23746), .B(n11877), .Z(n23749) );
  XNOR U25796 ( .A(n23742), .B(n23744), .Z(n11877) );
  NAND U25797 ( .A(n23750), .B(nreg[71]), .Z(n23744) );
  NAND U25798 ( .A(n12326), .B(nreg[71]), .Z(n23750) );
  XNOR U25799 ( .A(n23740), .B(n23751), .Z(n23742) );
  XOR U25800 ( .A(n23752), .B(n23753), .Z(n23740) );
  AND U25801 ( .A(n23754), .B(n23755), .Z(n23753) );
  XNOR U25802 ( .A(n23756), .B(n23752), .Z(n23755) );
  XOR U25803 ( .A(n23757), .B(nreg[71]), .Z(n23748) );
  IV U25804 ( .A(n23746), .Z(n23757) );
  XOR U25805 ( .A(n23758), .B(n23759), .Z(n23746) );
  AND U25806 ( .A(n23760), .B(n23761), .Z(n23759) );
  XNOR U25807 ( .A(n23758), .B(n11883), .Z(n23761) );
  XNOR U25808 ( .A(n23754), .B(n23756), .Z(n11883) );
  NAND U25809 ( .A(n23762), .B(nreg[70]), .Z(n23756) );
  NAND U25810 ( .A(n12326), .B(nreg[70]), .Z(n23762) );
  XNOR U25811 ( .A(n23752), .B(n23763), .Z(n23754) );
  XOR U25812 ( .A(n23764), .B(n23765), .Z(n23752) );
  AND U25813 ( .A(n23766), .B(n23767), .Z(n23765) );
  XNOR U25814 ( .A(n23768), .B(n23764), .Z(n23767) );
  XOR U25815 ( .A(n23769), .B(nreg[70]), .Z(n23760) );
  IV U25816 ( .A(n23758), .Z(n23769) );
  XOR U25817 ( .A(n23770), .B(n23771), .Z(n23758) );
  AND U25818 ( .A(n23772), .B(n23773), .Z(n23771) );
  XNOR U25819 ( .A(n23770), .B(n11889), .Z(n23773) );
  XNOR U25820 ( .A(n23766), .B(n23768), .Z(n11889) );
  NAND U25821 ( .A(n23774), .B(nreg[69]), .Z(n23768) );
  NAND U25822 ( .A(n12326), .B(nreg[69]), .Z(n23774) );
  XNOR U25823 ( .A(n23764), .B(n23775), .Z(n23766) );
  XOR U25824 ( .A(n23776), .B(n23777), .Z(n23764) );
  AND U25825 ( .A(n23778), .B(n23779), .Z(n23777) );
  XNOR U25826 ( .A(n23780), .B(n23776), .Z(n23779) );
  XOR U25827 ( .A(n23781), .B(nreg[69]), .Z(n23772) );
  IV U25828 ( .A(n23770), .Z(n23781) );
  XOR U25829 ( .A(n23782), .B(n23783), .Z(n23770) );
  AND U25830 ( .A(n23784), .B(n23785), .Z(n23783) );
  XNOR U25831 ( .A(n23782), .B(n11895), .Z(n23785) );
  XNOR U25832 ( .A(n23778), .B(n23780), .Z(n11895) );
  NAND U25833 ( .A(n23786), .B(nreg[68]), .Z(n23780) );
  NAND U25834 ( .A(n12326), .B(nreg[68]), .Z(n23786) );
  XNOR U25835 ( .A(n23776), .B(n23787), .Z(n23778) );
  XOR U25836 ( .A(n23788), .B(n23789), .Z(n23776) );
  AND U25837 ( .A(n23790), .B(n23791), .Z(n23789) );
  XNOR U25838 ( .A(n23792), .B(n23788), .Z(n23791) );
  XOR U25839 ( .A(n23793), .B(nreg[68]), .Z(n23784) );
  IV U25840 ( .A(n23782), .Z(n23793) );
  XOR U25841 ( .A(n23794), .B(n23795), .Z(n23782) );
  AND U25842 ( .A(n23796), .B(n23797), .Z(n23795) );
  XNOR U25843 ( .A(n23794), .B(n11901), .Z(n23797) );
  XNOR U25844 ( .A(n23790), .B(n23792), .Z(n11901) );
  NAND U25845 ( .A(n23798), .B(nreg[67]), .Z(n23792) );
  NAND U25846 ( .A(n12326), .B(nreg[67]), .Z(n23798) );
  XNOR U25847 ( .A(n23788), .B(n23799), .Z(n23790) );
  XOR U25848 ( .A(n23800), .B(n23801), .Z(n23788) );
  AND U25849 ( .A(n23802), .B(n23803), .Z(n23801) );
  XNOR U25850 ( .A(n23804), .B(n23800), .Z(n23803) );
  XOR U25851 ( .A(n23805), .B(nreg[67]), .Z(n23796) );
  IV U25852 ( .A(n23794), .Z(n23805) );
  XOR U25853 ( .A(n23806), .B(n23807), .Z(n23794) );
  AND U25854 ( .A(n23808), .B(n23809), .Z(n23807) );
  XNOR U25855 ( .A(n23806), .B(n11907), .Z(n23809) );
  XNOR U25856 ( .A(n23802), .B(n23804), .Z(n11907) );
  NAND U25857 ( .A(n23810), .B(nreg[66]), .Z(n23804) );
  NAND U25858 ( .A(n12326), .B(nreg[66]), .Z(n23810) );
  XNOR U25859 ( .A(n23800), .B(n23811), .Z(n23802) );
  XOR U25860 ( .A(n23812), .B(n23813), .Z(n23800) );
  AND U25861 ( .A(n23814), .B(n23815), .Z(n23813) );
  XNOR U25862 ( .A(n23816), .B(n23812), .Z(n23815) );
  XOR U25863 ( .A(n23817), .B(nreg[66]), .Z(n23808) );
  IV U25864 ( .A(n23806), .Z(n23817) );
  XOR U25865 ( .A(n23818), .B(n23819), .Z(n23806) );
  AND U25866 ( .A(n23820), .B(n23821), .Z(n23819) );
  XNOR U25867 ( .A(n23818), .B(n11913), .Z(n23821) );
  XNOR U25868 ( .A(n23814), .B(n23816), .Z(n11913) );
  NAND U25869 ( .A(n23822), .B(nreg[65]), .Z(n23816) );
  NAND U25870 ( .A(n12326), .B(nreg[65]), .Z(n23822) );
  XNOR U25871 ( .A(n23812), .B(n23823), .Z(n23814) );
  XOR U25872 ( .A(n23824), .B(n23825), .Z(n23812) );
  AND U25873 ( .A(n23826), .B(n23827), .Z(n23825) );
  XNOR U25874 ( .A(n23828), .B(n23824), .Z(n23827) );
  XOR U25875 ( .A(n23829), .B(nreg[65]), .Z(n23820) );
  IV U25876 ( .A(n23818), .Z(n23829) );
  XOR U25877 ( .A(n23830), .B(n23831), .Z(n23818) );
  AND U25878 ( .A(n23832), .B(n23833), .Z(n23831) );
  XNOR U25879 ( .A(n23830), .B(n11919), .Z(n23833) );
  XNOR U25880 ( .A(n23826), .B(n23828), .Z(n11919) );
  NAND U25881 ( .A(n23834), .B(nreg[64]), .Z(n23828) );
  NAND U25882 ( .A(n12326), .B(nreg[64]), .Z(n23834) );
  XNOR U25883 ( .A(n23824), .B(n23835), .Z(n23826) );
  XOR U25884 ( .A(n23836), .B(n23837), .Z(n23824) );
  AND U25885 ( .A(n23838), .B(n23839), .Z(n23837) );
  XNOR U25886 ( .A(n23840), .B(n23836), .Z(n23839) );
  XOR U25887 ( .A(n23841), .B(nreg[64]), .Z(n23832) );
  IV U25888 ( .A(n23830), .Z(n23841) );
  XOR U25889 ( .A(n23842), .B(n23843), .Z(n23830) );
  AND U25890 ( .A(n23844), .B(n23845), .Z(n23843) );
  XNOR U25891 ( .A(n23842), .B(n11925), .Z(n23845) );
  XNOR U25892 ( .A(n23838), .B(n23840), .Z(n11925) );
  NAND U25893 ( .A(n23846), .B(nreg[63]), .Z(n23840) );
  NAND U25894 ( .A(n12326), .B(nreg[63]), .Z(n23846) );
  XNOR U25895 ( .A(n23836), .B(n23847), .Z(n23838) );
  XOR U25896 ( .A(n23848), .B(n23849), .Z(n23836) );
  AND U25897 ( .A(n23850), .B(n23851), .Z(n23849) );
  XNOR U25898 ( .A(n23852), .B(n23848), .Z(n23851) );
  XOR U25899 ( .A(n23853), .B(nreg[63]), .Z(n23844) );
  IV U25900 ( .A(n23842), .Z(n23853) );
  XOR U25901 ( .A(n23854), .B(n23855), .Z(n23842) );
  AND U25902 ( .A(n23856), .B(n23857), .Z(n23855) );
  XNOR U25903 ( .A(n23854), .B(n11931), .Z(n23857) );
  XNOR U25904 ( .A(n23850), .B(n23852), .Z(n11931) );
  NAND U25905 ( .A(n23858), .B(nreg[62]), .Z(n23852) );
  NAND U25906 ( .A(n12326), .B(nreg[62]), .Z(n23858) );
  XNOR U25907 ( .A(n23848), .B(n23859), .Z(n23850) );
  XOR U25908 ( .A(n23860), .B(n23861), .Z(n23848) );
  AND U25909 ( .A(n23862), .B(n23863), .Z(n23861) );
  XNOR U25910 ( .A(n23864), .B(n23860), .Z(n23863) );
  XOR U25911 ( .A(n23865), .B(nreg[62]), .Z(n23856) );
  IV U25912 ( .A(n23854), .Z(n23865) );
  XOR U25913 ( .A(n23866), .B(n23867), .Z(n23854) );
  AND U25914 ( .A(n23868), .B(n23869), .Z(n23867) );
  XNOR U25915 ( .A(n23866), .B(n11937), .Z(n23869) );
  XNOR U25916 ( .A(n23862), .B(n23864), .Z(n11937) );
  NAND U25917 ( .A(n23870), .B(nreg[61]), .Z(n23864) );
  NAND U25918 ( .A(n12326), .B(nreg[61]), .Z(n23870) );
  XNOR U25919 ( .A(n23860), .B(n23871), .Z(n23862) );
  XOR U25920 ( .A(n23872), .B(n23873), .Z(n23860) );
  AND U25921 ( .A(n23874), .B(n23875), .Z(n23873) );
  XNOR U25922 ( .A(n23876), .B(n23872), .Z(n23875) );
  XOR U25923 ( .A(n23877), .B(nreg[61]), .Z(n23868) );
  IV U25924 ( .A(n23866), .Z(n23877) );
  XOR U25925 ( .A(n23878), .B(n23879), .Z(n23866) );
  AND U25926 ( .A(n23880), .B(n23881), .Z(n23879) );
  XNOR U25927 ( .A(n23878), .B(n11943), .Z(n23881) );
  XNOR U25928 ( .A(n23874), .B(n23876), .Z(n11943) );
  NAND U25929 ( .A(n23882), .B(nreg[60]), .Z(n23876) );
  NAND U25930 ( .A(n12326), .B(nreg[60]), .Z(n23882) );
  XNOR U25931 ( .A(n23872), .B(n23883), .Z(n23874) );
  XOR U25932 ( .A(n23884), .B(n23885), .Z(n23872) );
  AND U25933 ( .A(n23886), .B(n23887), .Z(n23885) );
  XNOR U25934 ( .A(n23888), .B(n23884), .Z(n23887) );
  XOR U25935 ( .A(n23889), .B(nreg[60]), .Z(n23880) );
  IV U25936 ( .A(n23878), .Z(n23889) );
  XOR U25937 ( .A(n23890), .B(n23891), .Z(n23878) );
  AND U25938 ( .A(n23892), .B(n23893), .Z(n23891) );
  XNOR U25939 ( .A(n23890), .B(n11949), .Z(n23893) );
  XNOR U25940 ( .A(n23886), .B(n23888), .Z(n11949) );
  NAND U25941 ( .A(n23894), .B(nreg[59]), .Z(n23888) );
  NAND U25942 ( .A(n12326), .B(nreg[59]), .Z(n23894) );
  XNOR U25943 ( .A(n23884), .B(n23895), .Z(n23886) );
  XOR U25944 ( .A(n23896), .B(n23897), .Z(n23884) );
  AND U25945 ( .A(n23898), .B(n23899), .Z(n23897) );
  XNOR U25946 ( .A(n23900), .B(n23896), .Z(n23899) );
  XOR U25947 ( .A(n23901), .B(nreg[59]), .Z(n23892) );
  IV U25948 ( .A(n23890), .Z(n23901) );
  XOR U25949 ( .A(n23902), .B(n23903), .Z(n23890) );
  AND U25950 ( .A(n23904), .B(n23905), .Z(n23903) );
  XNOR U25951 ( .A(n23902), .B(n11955), .Z(n23905) );
  XNOR U25952 ( .A(n23898), .B(n23900), .Z(n11955) );
  NAND U25953 ( .A(n23906), .B(nreg[58]), .Z(n23900) );
  NAND U25954 ( .A(n12326), .B(nreg[58]), .Z(n23906) );
  XNOR U25955 ( .A(n23896), .B(n23907), .Z(n23898) );
  XOR U25956 ( .A(n23908), .B(n23909), .Z(n23896) );
  AND U25957 ( .A(n23910), .B(n23911), .Z(n23909) );
  XNOR U25958 ( .A(n23912), .B(n23908), .Z(n23911) );
  XOR U25959 ( .A(n23913), .B(nreg[58]), .Z(n23904) );
  IV U25960 ( .A(n23902), .Z(n23913) );
  XOR U25961 ( .A(n23914), .B(n23915), .Z(n23902) );
  AND U25962 ( .A(n23916), .B(n23917), .Z(n23915) );
  XNOR U25963 ( .A(n23914), .B(n11961), .Z(n23917) );
  XNOR U25964 ( .A(n23910), .B(n23912), .Z(n11961) );
  NAND U25965 ( .A(n23918), .B(nreg[57]), .Z(n23912) );
  NAND U25966 ( .A(n12326), .B(nreg[57]), .Z(n23918) );
  XNOR U25967 ( .A(n23908), .B(n23919), .Z(n23910) );
  XOR U25968 ( .A(n23920), .B(n23921), .Z(n23908) );
  AND U25969 ( .A(n23922), .B(n23923), .Z(n23921) );
  XNOR U25970 ( .A(n23924), .B(n23920), .Z(n23923) );
  XOR U25971 ( .A(n23925), .B(nreg[57]), .Z(n23916) );
  IV U25972 ( .A(n23914), .Z(n23925) );
  XOR U25973 ( .A(n23926), .B(n23927), .Z(n23914) );
  AND U25974 ( .A(n23928), .B(n23929), .Z(n23927) );
  XNOR U25975 ( .A(n23926), .B(n11967), .Z(n23929) );
  XNOR U25976 ( .A(n23922), .B(n23924), .Z(n11967) );
  NAND U25977 ( .A(n23930), .B(nreg[56]), .Z(n23924) );
  NAND U25978 ( .A(n12326), .B(nreg[56]), .Z(n23930) );
  XNOR U25979 ( .A(n23920), .B(n23931), .Z(n23922) );
  XOR U25980 ( .A(n23932), .B(n23933), .Z(n23920) );
  AND U25981 ( .A(n23934), .B(n23935), .Z(n23933) );
  XNOR U25982 ( .A(n23936), .B(n23932), .Z(n23935) );
  XOR U25983 ( .A(n23937), .B(nreg[56]), .Z(n23928) );
  IV U25984 ( .A(n23926), .Z(n23937) );
  XOR U25985 ( .A(n23938), .B(n23939), .Z(n23926) );
  AND U25986 ( .A(n23940), .B(n23941), .Z(n23939) );
  XNOR U25987 ( .A(n23938), .B(n11973), .Z(n23941) );
  XNOR U25988 ( .A(n23934), .B(n23936), .Z(n11973) );
  NAND U25989 ( .A(n23942), .B(nreg[55]), .Z(n23936) );
  NAND U25990 ( .A(n12326), .B(nreg[55]), .Z(n23942) );
  XNOR U25991 ( .A(n23932), .B(n23943), .Z(n23934) );
  XOR U25992 ( .A(n23944), .B(n23945), .Z(n23932) );
  AND U25993 ( .A(n23946), .B(n23947), .Z(n23945) );
  XNOR U25994 ( .A(n23948), .B(n23944), .Z(n23947) );
  XOR U25995 ( .A(n23949), .B(nreg[55]), .Z(n23940) );
  IV U25996 ( .A(n23938), .Z(n23949) );
  XOR U25997 ( .A(n23950), .B(n23951), .Z(n23938) );
  AND U25998 ( .A(n23952), .B(n23953), .Z(n23951) );
  XNOR U25999 ( .A(n23950), .B(n11979), .Z(n23953) );
  XNOR U26000 ( .A(n23946), .B(n23948), .Z(n11979) );
  NAND U26001 ( .A(n23954), .B(nreg[54]), .Z(n23948) );
  NAND U26002 ( .A(n12326), .B(nreg[54]), .Z(n23954) );
  XNOR U26003 ( .A(n23944), .B(n23955), .Z(n23946) );
  XOR U26004 ( .A(n23956), .B(n23957), .Z(n23944) );
  AND U26005 ( .A(n23958), .B(n23959), .Z(n23957) );
  XNOR U26006 ( .A(n23960), .B(n23956), .Z(n23959) );
  XOR U26007 ( .A(n23961), .B(nreg[54]), .Z(n23952) );
  IV U26008 ( .A(n23950), .Z(n23961) );
  XOR U26009 ( .A(n23962), .B(n23963), .Z(n23950) );
  AND U26010 ( .A(n23964), .B(n23965), .Z(n23963) );
  XNOR U26011 ( .A(n23962), .B(n11985), .Z(n23965) );
  XNOR U26012 ( .A(n23958), .B(n23960), .Z(n11985) );
  NAND U26013 ( .A(n23966), .B(nreg[53]), .Z(n23960) );
  NAND U26014 ( .A(n12326), .B(nreg[53]), .Z(n23966) );
  XNOR U26015 ( .A(n23956), .B(n23967), .Z(n23958) );
  XOR U26016 ( .A(n23968), .B(n23969), .Z(n23956) );
  AND U26017 ( .A(n23970), .B(n23971), .Z(n23969) );
  XNOR U26018 ( .A(n23972), .B(n23968), .Z(n23971) );
  XOR U26019 ( .A(n23973), .B(nreg[53]), .Z(n23964) );
  IV U26020 ( .A(n23962), .Z(n23973) );
  XOR U26021 ( .A(n23974), .B(n23975), .Z(n23962) );
  AND U26022 ( .A(n23976), .B(n23977), .Z(n23975) );
  XNOR U26023 ( .A(n23974), .B(n11991), .Z(n23977) );
  XNOR U26024 ( .A(n23970), .B(n23972), .Z(n11991) );
  NAND U26025 ( .A(n23978), .B(nreg[52]), .Z(n23972) );
  NAND U26026 ( .A(n12326), .B(nreg[52]), .Z(n23978) );
  XNOR U26027 ( .A(n23968), .B(n23979), .Z(n23970) );
  XOR U26028 ( .A(n23980), .B(n23981), .Z(n23968) );
  AND U26029 ( .A(n23982), .B(n23983), .Z(n23981) );
  XNOR U26030 ( .A(n23984), .B(n23980), .Z(n23983) );
  XOR U26031 ( .A(n23985), .B(nreg[52]), .Z(n23976) );
  IV U26032 ( .A(n23974), .Z(n23985) );
  XOR U26033 ( .A(n23986), .B(n23987), .Z(n23974) );
  AND U26034 ( .A(n23988), .B(n23989), .Z(n23987) );
  XNOR U26035 ( .A(n23986), .B(n11997), .Z(n23989) );
  XNOR U26036 ( .A(n23982), .B(n23984), .Z(n11997) );
  NAND U26037 ( .A(n23990), .B(nreg[51]), .Z(n23984) );
  NAND U26038 ( .A(n12326), .B(nreg[51]), .Z(n23990) );
  XNOR U26039 ( .A(n23980), .B(n23991), .Z(n23982) );
  XOR U26040 ( .A(n23992), .B(n23993), .Z(n23980) );
  AND U26041 ( .A(n23994), .B(n23995), .Z(n23993) );
  XNOR U26042 ( .A(n23996), .B(n23992), .Z(n23995) );
  XOR U26043 ( .A(n23997), .B(nreg[51]), .Z(n23988) );
  IV U26044 ( .A(n23986), .Z(n23997) );
  XOR U26045 ( .A(n23998), .B(n23999), .Z(n23986) );
  AND U26046 ( .A(n24000), .B(n24001), .Z(n23999) );
  XNOR U26047 ( .A(n23998), .B(n12003), .Z(n24001) );
  XNOR U26048 ( .A(n23994), .B(n23996), .Z(n12003) );
  NAND U26049 ( .A(n24002), .B(nreg[50]), .Z(n23996) );
  NAND U26050 ( .A(n12326), .B(nreg[50]), .Z(n24002) );
  XNOR U26051 ( .A(n23992), .B(n24003), .Z(n23994) );
  XOR U26052 ( .A(n24004), .B(n24005), .Z(n23992) );
  AND U26053 ( .A(n24006), .B(n24007), .Z(n24005) );
  XNOR U26054 ( .A(n24008), .B(n24004), .Z(n24007) );
  XOR U26055 ( .A(n24009), .B(nreg[50]), .Z(n24000) );
  IV U26056 ( .A(n23998), .Z(n24009) );
  XOR U26057 ( .A(n24010), .B(n24011), .Z(n23998) );
  AND U26058 ( .A(n24012), .B(n24013), .Z(n24011) );
  XNOR U26059 ( .A(n24010), .B(n12009), .Z(n24013) );
  XNOR U26060 ( .A(n24006), .B(n24008), .Z(n12009) );
  NAND U26061 ( .A(n24014), .B(nreg[49]), .Z(n24008) );
  NAND U26062 ( .A(n12326), .B(nreg[49]), .Z(n24014) );
  XNOR U26063 ( .A(n24004), .B(n24015), .Z(n24006) );
  XOR U26064 ( .A(n24016), .B(n24017), .Z(n24004) );
  AND U26065 ( .A(n24018), .B(n24019), .Z(n24017) );
  XNOR U26066 ( .A(n24020), .B(n24016), .Z(n24019) );
  XOR U26067 ( .A(n24021), .B(nreg[49]), .Z(n24012) );
  IV U26068 ( .A(n24010), .Z(n24021) );
  XOR U26069 ( .A(n24022), .B(n24023), .Z(n24010) );
  AND U26070 ( .A(n24024), .B(n24025), .Z(n24023) );
  XNOR U26071 ( .A(n24022), .B(n12015), .Z(n24025) );
  XNOR U26072 ( .A(n24018), .B(n24020), .Z(n12015) );
  NAND U26073 ( .A(n24026), .B(nreg[48]), .Z(n24020) );
  NAND U26074 ( .A(n12326), .B(nreg[48]), .Z(n24026) );
  XNOR U26075 ( .A(n24016), .B(n24027), .Z(n24018) );
  XOR U26076 ( .A(n24028), .B(n24029), .Z(n24016) );
  AND U26077 ( .A(n24030), .B(n24031), .Z(n24029) );
  XNOR U26078 ( .A(n24032), .B(n24028), .Z(n24031) );
  XOR U26079 ( .A(n24033), .B(nreg[48]), .Z(n24024) );
  IV U26080 ( .A(n24022), .Z(n24033) );
  XOR U26081 ( .A(n24034), .B(n24035), .Z(n24022) );
  AND U26082 ( .A(n24036), .B(n24037), .Z(n24035) );
  XNOR U26083 ( .A(n24034), .B(n12021), .Z(n24037) );
  XNOR U26084 ( .A(n24030), .B(n24032), .Z(n12021) );
  NAND U26085 ( .A(n24038), .B(nreg[47]), .Z(n24032) );
  NAND U26086 ( .A(n12326), .B(nreg[47]), .Z(n24038) );
  XNOR U26087 ( .A(n24028), .B(n24039), .Z(n24030) );
  XOR U26088 ( .A(n24040), .B(n24041), .Z(n24028) );
  AND U26089 ( .A(n24042), .B(n24043), .Z(n24041) );
  XNOR U26090 ( .A(n24044), .B(n24040), .Z(n24043) );
  XOR U26091 ( .A(n24045), .B(nreg[47]), .Z(n24036) );
  IV U26092 ( .A(n24034), .Z(n24045) );
  XOR U26093 ( .A(n24046), .B(n24047), .Z(n24034) );
  AND U26094 ( .A(n24048), .B(n24049), .Z(n24047) );
  XNOR U26095 ( .A(n24046), .B(n12027), .Z(n24049) );
  XNOR U26096 ( .A(n24042), .B(n24044), .Z(n12027) );
  NAND U26097 ( .A(n24050), .B(nreg[46]), .Z(n24044) );
  NAND U26098 ( .A(n12326), .B(nreg[46]), .Z(n24050) );
  XNOR U26099 ( .A(n24040), .B(n24051), .Z(n24042) );
  XOR U26100 ( .A(n24052), .B(n24053), .Z(n24040) );
  AND U26101 ( .A(n24054), .B(n24055), .Z(n24053) );
  XNOR U26102 ( .A(n24056), .B(n24052), .Z(n24055) );
  XOR U26103 ( .A(n24057), .B(nreg[46]), .Z(n24048) );
  IV U26104 ( .A(n24046), .Z(n24057) );
  XOR U26105 ( .A(n24058), .B(n24059), .Z(n24046) );
  AND U26106 ( .A(n24060), .B(n24061), .Z(n24059) );
  XNOR U26107 ( .A(n24058), .B(n12033), .Z(n24061) );
  XNOR U26108 ( .A(n24054), .B(n24056), .Z(n12033) );
  NAND U26109 ( .A(n24062), .B(nreg[45]), .Z(n24056) );
  NAND U26110 ( .A(n12326), .B(nreg[45]), .Z(n24062) );
  XNOR U26111 ( .A(n24052), .B(n24063), .Z(n24054) );
  XOR U26112 ( .A(n24064), .B(n24065), .Z(n24052) );
  AND U26113 ( .A(n24066), .B(n24067), .Z(n24065) );
  XNOR U26114 ( .A(n24068), .B(n24064), .Z(n24067) );
  XOR U26115 ( .A(n24069), .B(nreg[45]), .Z(n24060) );
  IV U26116 ( .A(n24058), .Z(n24069) );
  XOR U26117 ( .A(n24070), .B(n24071), .Z(n24058) );
  AND U26118 ( .A(n24072), .B(n24073), .Z(n24071) );
  XNOR U26119 ( .A(n24070), .B(n12039), .Z(n24073) );
  XNOR U26120 ( .A(n24066), .B(n24068), .Z(n12039) );
  NAND U26121 ( .A(n24074), .B(nreg[44]), .Z(n24068) );
  NAND U26122 ( .A(n12326), .B(nreg[44]), .Z(n24074) );
  XNOR U26123 ( .A(n24064), .B(n24075), .Z(n24066) );
  XOR U26124 ( .A(n24076), .B(n24077), .Z(n24064) );
  AND U26125 ( .A(n24078), .B(n24079), .Z(n24077) );
  XNOR U26126 ( .A(n24080), .B(n24076), .Z(n24079) );
  XOR U26127 ( .A(n24081), .B(nreg[44]), .Z(n24072) );
  IV U26128 ( .A(n24070), .Z(n24081) );
  XOR U26129 ( .A(n24082), .B(n24083), .Z(n24070) );
  AND U26130 ( .A(n24084), .B(n24085), .Z(n24083) );
  XNOR U26131 ( .A(n24082), .B(n12045), .Z(n24085) );
  XNOR U26132 ( .A(n24078), .B(n24080), .Z(n12045) );
  NAND U26133 ( .A(n24086), .B(nreg[43]), .Z(n24080) );
  NAND U26134 ( .A(n12326), .B(nreg[43]), .Z(n24086) );
  XNOR U26135 ( .A(n24076), .B(n24087), .Z(n24078) );
  XOR U26136 ( .A(n24088), .B(n24089), .Z(n24076) );
  AND U26137 ( .A(n24090), .B(n24091), .Z(n24089) );
  XNOR U26138 ( .A(n24092), .B(n24088), .Z(n24091) );
  XOR U26139 ( .A(n24093), .B(nreg[43]), .Z(n24084) );
  IV U26140 ( .A(n24082), .Z(n24093) );
  XOR U26141 ( .A(n24094), .B(n24095), .Z(n24082) );
  AND U26142 ( .A(n24096), .B(n24097), .Z(n24095) );
  XNOR U26143 ( .A(n24094), .B(n12051), .Z(n24097) );
  XNOR U26144 ( .A(n24090), .B(n24092), .Z(n12051) );
  NAND U26145 ( .A(n24098), .B(nreg[42]), .Z(n24092) );
  NAND U26146 ( .A(n12326), .B(nreg[42]), .Z(n24098) );
  XNOR U26147 ( .A(n24088), .B(n24099), .Z(n24090) );
  XOR U26148 ( .A(n24100), .B(n24101), .Z(n24088) );
  AND U26149 ( .A(n24102), .B(n24103), .Z(n24101) );
  XNOR U26150 ( .A(n24104), .B(n24100), .Z(n24103) );
  XOR U26151 ( .A(n24105), .B(nreg[42]), .Z(n24096) );
  IV U26152 ( .A(n24094), .Z(n24105) );
  XOR U26153 ( .A(n24106), .B(n24107), .Z(n24094) );
  AND U26154 ( .A(n24108), .B(n24109), .Z(n24107) );
  XNOR U26155 ( .A(n24106), .B(n12057), .Z(n24109) );
  XNOR U26156 ( .A(n24102), .B(n24104), .Z(n12057) );
  NAND U26157 ( .A(n24110), .B(nreg[41]), .Z(n24104) );
  NAND U26158 ( .A(n12326), .B(nreg[41]), .Z(n24110) );
  XNOR U26159 ( .A(n24100), .B(n24111), .Z(n24102) );
  XOR U26160 ( .A(n24112), .B(n24113), .Z(n24100) );
  AND U26161 ( .A(n24114), .B(n24115), .Z(n24113) );
  XNOR U26162 ( .A(n24116), .B(n24112), .Z(n24115) );
  XOR U26163 ( .A(n24117), .B(nreg[41]), .Z(n24108) );
  IV U26164 ( .A(n24106), .Z(n24117) );
  XOR U26165 ( .A(n24118), .B(n24119), .Z(n24106) );
  AND U26166 ( .A(n24120), .B(n24121), .Z(n24119) );
  XNOR U26167 ( .A(n24118), .B(n12063), .Z(n24121) );
  XNOR U26168 ( .A(n24114), .B(n24116), .Z(n12063) );
  NAND U26169 ( .A(n24122), .B(nreg[40]), .Z(n24116) );
  NAND U26170 ( .A(n12326), .B(nreg[40]), .Z(n24122) );
  XNOR U26171 ( .A(n24112), .B(n24123), .Z(n24114) );
  XOR U26172 ( .A(n24124), .B(n24125), .Z(n24112) );
  AND U26173 ( .A(n24126), .B(n24127), .Z(n24125) );
  XNOR U26174 ( .A(n24128), .B(n24124), .Z(n24127) );
  XOR U26175 ( .A(n24129), .B(nreg[40]), .Z(n24120) );
  IV U26176 ( .A(n24118), .Z(n24129) );
  XOR U26177 ( .A(n24130), .B(n24131), .Z(n24118) );
  AND U26178 ( .A(n24132), .B(n24133), .Z(n24131) );
  XNOR U26179 ( .A(n24130), .B(n12069), .Z(n24133) );
  XNOR U26180 ( .A(n24126), .B(n24128), .Z(n12069) );
  NAND U26181 ( .A(n24134), .B(nreg[39]), .Z(n24128) );
  NAND U26182 ( .A(n12326), .B(nreg[39]), .Z(n24134) );
  XNOR U26183 ( .A(n24124), .B(n24135), .Z(n24126) );
  XOR U26184 ( .A(n24136), .B(n24137), .Z(n24124) );
  AND U26185 ( .A(n24138), .B(n24139), .Z(n24137) );
  XNOR U26186 ( .A(n24140), .B(n24136), .Z(n24139) );
  XOR U26187 ( .A(n24141), .B(nreg[39]), .Z(n24132) );
  IV U26188 ( .A(n24130), .Z(n24141) );
  XOR U26189 ( .A(n24142), .B(n24143), .Z(n24130) );
  AND U26190 ( .A(n24144), .B(n24145), .Z(n24143) );
  XNOR U26191 ( .A(n24142), .B(n12075), .Z(n24145) );
  XNOR U26192 ( .A(n24138), .B(n24140), .Z(n12075) );
  NAND U26193 ( .A(n24146), .B(nreg[38]), .Z(n24140) );
  NAND U26194 ( .A(n12326), .B(nreg[38]), .Z(n24146) );
  XNOR U26195 ( .A(n24136), .B(n24147), .Z(n24138) );
  XOR U26196 ( .A(n24148), .B(n24149), .Z(n24136) );
  AND U26197 ( .A(n24150), .B(n24151), .Z(n24149) );
  XNOR U26198 ( .A(n24152), .B(n24148), .Z(n24151) );
  XOR U26199 ( .A(n24153), .B(nreg[38]), .Z(n24144) );
  IV U26200 ( .A(n24142), .Z(n24153) );
  XOR U26201 ( .A(n24154), .B(n24155), .Z(n24142) );
  AND U26202 ( .A(n24156), .B(n24157), .Z(n24155) );
  XNOR U26203 ( .A(n24154), .B(n12081), .Z(n24157) );
  XNOR U26204 ( .A(n24150), .B(n24152), .Z(n12081) );
  NAND U26205 ( .A(n24158), .B(nreg[37]), .Z(n24152) );
  NAND U26206 ( .A(n12326), .B(nreg[37]), .Z(n24158) );
  XNOR U26207 ( .A(n24148), .B(n24159), .Z(n24150) );
  XOR U26208 ( .A(n24160), .B(n24161), .Z(n24148) );
  AND U26209 ( .A(n24162), .B(n24163), .Z(n24161) );
  XNOR U26210 ( .A(n24164), .B(n24160), .Z(n24163) );
  XOR U26211 ( .A(n24165), .B(nreg[37]), .Z(n24156) );
  IV U26212 ( .A(n24154), .Z(n24165) );
  XOR U26213 ( .A(n24166), .B(n24167), .Z(n24154) );
  AND U26214 ( .A(n24168), .B(n24169), .Z(n24167) );
  XNOR U26215 ( .A(n24166), .B(n12087), .Z(n24169) );
  XNOR U26216 ( .A(n24162), .B(n24164), .Z(n12087) );
  NAND U26217 ( .A(n24170), .B(nreg[36]), .Z(n24164) );
  NAND U26218 ( .A(n12326), .B(nreg[36]), .Z(n24170) );
  XNOR U26219 ( .A(n24160), .B(n24171), .Z(n24162) );
  XOR U26220 ( .A(n24172), .B(n24173), .Z(n24160) );
  AND U26221 ( .A(n24174), .B(n24175), .Z(n24173) );
  XNOR U26222 ( .A(n24176), .B(n24172), .Z(n24175) );
  XOR U26223 ( .A(n24177), .B(nreg[36]), .Z(n24168) );
  IV U26224 ( .A(n24166), .Z(n24177) );
  XOR U26225 ( .A(n24178), .B(n24179), .Z(n24166) );
  AND U26226 ( .A(n24180), .B(n24181), .Z(n24179) );
  XNOR U26227 ( .A(n24178), .B(n12093), .Z(n24181) );
  XNOR U26228 ( .A(n24174), .B(n24176), .Z(n12093) );
  NAND U26229 ( .A(n24182), .B(nreg[35]), .Z(n24176) );
  NAND U26230 ( .A(n12326), .B(nreg[35]), .Z(n24182) );
  XNOR U26231 ( .A(n24172), .B(n24183), .Z(n24174) );
  XOR U26232 ( .A(n24184), .B(n24185), .Z(n24172) );
  AND U26233 ( .A(n24186), .B(n24187), .Z(n24185) );
  XNOR U26234 ( .A(n24188), .B(n24184), .Z(n24187) );
  XOR U26235 ( .A(n24189), .B(nreg[35]), .Z(n24180) );
  IV U26236 ( .A(n24178), .Z(n24189) );
  XOR U26237 ( .A(n24190), .B(n24191), .Z(n24178) );
  AND U26238 ( .A(n24192), .B(n24193), .Z(n24191) );
  XNOR U26239 ( .A(n24190), .B(n12099), .Z(n24193) );
  XNOR U26240 ( .A(n24186), .B(n24188), .Z(n12099) );
  NAND U26241 ( .A(n24194), .B(nreg[34]), .Z(n24188) );
  NAND U26242 ( .A(n12326), .B(nreg[34]), .Z(n24194) );
  XNOR U26243 ( .A(n24184), .B(n24195), .Z(n24186) );
  XOR U26244 ( .A(n24196), .B(n24197), .Z(n24184) );
  AND U26245 ( .A(n24198), .B(n24199), .Z(n24197) );
  XNOR U26246 ( .A(n24200), .B(n24196), .Z(n24199) );
  XOR U26247 ( .A(n24201), .B(nreg[34]), .Z(n24192) );
  IV U26248 ( .A(n24190), .Z(n24201) );
  XOR U26249 ( .A(n24202), .B(n24203), .Z(n24190) );
  AND U26250 ( .A(n24204), .B(n24205), .Z(n24203) );
  XNOR U26251 ( .A(n24202), .B(n12105), .Z(n24205) );
  XNOR U26252 ( .A(n24198), .B(n24200), .Z(n12105) );
  NAND U26253 ( .A(n24206), .B(nreg[33]), .Z(n24200) );
  NAND U26254 ( .A(n12326), .B(nreg[33]), .Z(n24206) );
  XNOR U26255 ( .A(n24196), .B(n24207), .Z(n24198) );
  XOR U26256 ( .A(n24208), .B(n24209), .Z(n24196) );
  AND U26257 ( .A(n24210), .B(n24211), .Z(n24209) );
  XNOR U26258 ( .A(n24212), .B(n24208), .Z(n24211) );
  XOR U26259 ( .A(n24213), .B(nreg[33]), .Z(n24204) );
  IV U26260 ( .A(n24202), .Z(n24213) );
  XOR U26261 ( .A(n24214), .B(n24215), .Z(n24202) );
  AND U26262 ( .A(n24216), .B(n24217), .Z(n24215) );
  XNOR U26263 ( .A(n24214), .B(n12111), .Z(n24217) );
  XNOR U26264 ( .A(n24210), .B(n24212), .Z(n12111) );
  NAND U26265 ( .A(n24218), .B(nreg[32]), .Z(n24212) );
  NAND U26266 ( .A(n12326), .B(nreg[32]), .Z(n24218) );
  XNOR U26267 ( .A(n24208), .B(n24219), .Z(n24210) );
  XOR U26268 ( .A(n24220), .B(n24221), .Z(n24208) );
  AND U26269 ( .A(n24222), .B(n24223), .Z(n24221) );
  XNOR U26270 ( .A(n24224), .B(n24220), .Z(n24223) );
  XOR U26271 ( .A(n24225), .B(nreg[32]), .Z(n24216) );
  IV U26272 ( .A(n24214), .Z(n24225) );
  XOR U26273 ( .A(n24226), .B(n24227), .Z(n24214) );
  AND U26274 ( .A(n24228), .B(n24229), .Z(n24227) );
  XNOR U26275 ( .A(n24226), .B(n12117), .Z(n24229) );
  XNOR U26276 ( .A(n24222), .B(n24224), .Z(n12117) );
  NAND U26277 ( .A(n24230), .B(nreg[31]), .Z(n24224) );
  NAND U26278 ( .A(n12326), .B(nreg[31]), .Z(n24230) );
  XNOR U26279 ( .A(n24220), .B(n24231), .Z(n24222) );
  XOR U26280 ( .A(n24232), .B(n24233), .Z(n24220) );
  AND U26281 ( .A(n24234), .B(n24235), .Z(n24233) );
  XNOR U26282 ( .A(n24236), .B(n24232), .Z(n24235) );
  XOR U26283 ( .A(n24237), .B(nreg[31]), .Z(n24228) );
  IV U26284 ( .A(n24226), .Z(n24237) );
  XOR U26285 ( .A(n24238), .B(n24239), .Z(n24226) );
  AND U26286 ( .A(n24240), .B(n24241), .Z(n24239) );
  XNOR U26287 ( .A(n24238), .B(n12123), .Z(n24241) );
  XNOR U26288 ( .A(n24234), .B(n24236), .Z(n12123) );
  NAND U26289 ( .A(n24242), .B(nreg[30]), .Z(n24236) );
  NAND U26290 ( .A(n12326), .B(nreg[30]), .Z(n24242) );
  XNOR U26291 ( .A(n24232), .B(n24243), .Z(n24234) );
  XOR U26292 ( .A(n24244), .B(n24245), .Z(n24232) );
  AND U26293 ( .A(n24246), .B(n24247), .Z(n24245) );
  XNOR U26294 ( .A(n24248), .B(n24244), .Z(n24247) );
  XOR U26295 ( .A(n24249), .B(nreg[30]), .Z(n24240) );
  IV U26296 ( .A(n24238), .Z(n24249) );
  XOR U26297 ( .A(n24250), .B(n24251), .Z(n24238) );
  AND U26298 ( .A(n24252), .B(n24253), .Z(n24251) );
  XNOR U26299 ( .A(n24250), .B(n12129), .Z(n24253) );
  XNOR U26300 ( .A(n24246), .B(n24248), .Z(n12129) );
  NAND U26301 ( .A(n24254), .B(nreg[29]), .Z(n24248) );
  NAND U26302 ( .A(n12326), .B(nreg[29]), .Z(n24254) );
  XNOR U26303 ( .A(n24244), .B(n24255), .Z(n24246) );
  XOR U26304 ( .A(n24256), .B(n24257), .Z(n24244) );
  AND U26305 ( .A(n24258), .B(n24259), .Z(n24257) );
  XNOR U26306 ( .A(n24260), .B(n24256), .Z(n24259) );
  XOR U26307 ( .A(n24261), .B(nreg[29]), .Z(n24252) );
  IV U26308 ( .A(n24250), .Z(n24261) );
  XOR U26309 ( .A(n24262), .B(n24263), .Z(n24250) );
  AND U26310 ( .A(n24264), .B(n24265), .Z(n24263) );
  XNOR U26311 ( .A(n24262), .B(n12135), .Z(n24265) );
  XNOR U26312 ( .A(n24258), .B(n24260), .Z(n12135) );
  NAND U26313 ( .A(n24266), .B(nreg[28]), .Z(n24260) );
  NAND U26314 ( .A(n12326), .B(nreg[28]), .Z(n24266) );
  XNOR U26315 ( .A(n24256), .B(n24267), .Z(n24258) );
  XOR U26316 ( .A(n24268), .B(n24269), .Z(n24256) );
  AND U26317 ( .A(n24270), .B(n24271), .Z(n24269) );
  XNOR U26318 ( .A(n24272), .B(n24268), .Z(n24271) );
  XOR U26319 ( .A(n24273), .B(nreg[28]), .Z(n24264) );
  IV U26320 ( .A(n24262), .Z(n24273) );
  XOR U26321 ( .A(n24274), .B(n24275), .Z(n24262) );
  AND U26322 ( .A(n24276), .B(n24277), .Z(n24275) );
  XNOR U26323 ( .A(n24274), .B(n12141), .Z(n24277) );
  XNOR U26324 ( .A(n24270), .B(n24272), .Z(n12141) );
  NAND U26325 ( .A(n24278), .B(nreg[27]), .Z(n24272) );
  NAND U26326 ( .A(n12326), .B(nreg[27]), .Z(n24278) );
  XNOR U26327 ( .A(n24268), .B(n24279), .Z(n24270) );
  XOR U26328 ( .A(n24280), .B(n24281), .Z(n24268) );
  AND U26329 ( .A(n24282), .B(n24283), .Z(n24281) );
  XNOR U26330 ( .A(n24284), .B(n24280), .Z(n24283) );
  XOR U26331 ( .A(n24285), .B(nreg[27]), .Z(n24276) );
  IV U26332 ( .A(n24274), .Z(n24285) );
  XOR U26333 ( .A(n24286), .B(n24287), .Z(n24274) );
  AND U26334 ( .A(n24288), .B(n24289), .Z(n24287) );
  XNOR U26335 ( .A(n24286), .B(n12147), .Z(n24289) );
  XNOR U26336 ( .A(n24282), .B(n24284), .Z(n12147) );
  NAND U26337 ( .A(n24290), .B(nreg[26]), .Z(n24284) );
  NAND U26338 ( .A(n12326), .B(nreg[26]), .Z(n24290) );
  XNOR U26339 ( .A(n24280), .B(n24291), .Z(n24282) );
  XOR U26340 ( .A(n24292), .B(n24293), .Z(n24280) );
  AND U26341 ( .A(n24294), .B(n24295), .Z(n24293) );
  XNOR U26342 ( .A(n24296), .B(n24292), .Z(n24295) );
  XOR U26343 ( .A(n24297), .B(nreg[26]), .Z(n24288) );
  IV U26344 ( .A(n24286), .Z(n24297) );
  XOR U26345 ( .A(n24298), .B(n24299), .Z(n24286) );
  AND U26346 ( .A(n24300), .B(n24301), .Z(n24299) );
  XNOR U26347 ( .A(n24298), .B(n12153), .Z(n24301) );
  XNOR U26348 ( .A(n24294), .B(n24296), .Z(n12153) );
  NAND U26349 ( .A(n24302), .B(nreg[25]), .Z(n24296) );
  NAND U26350 ( .A(n12326), .B(nreg[25]), .Z(n24302) );
  XNOR U26351 ( .A(n24292), .B(n24303), .Z(n24294) );
  XOR U26352 ( .A(n24304), .B(n24305), .Z(n24292) );
  AND U26353 ( .A(n24306), .B(n24307), .Z(n24305) );
  XNOR U26354 ( .A(n24308), .B(n24304), .Z(n24307) );
  XOR U26355 ( .A(n24309), .B(nreg[25]), .Z(n24300) );
  IV U26356 ( .A(n24298), .Z(n24309) );
  XOR U26357 ( .A(n24310), .B(n24311), .Z(n24298) );
  AND U26358 ( .A(n24312), .B(n24313), .Z(n24311) );
  XNOR U26359 ( .A(n24310), .B(n12159), .Z(n24313) );
  XNOR U26360 ( .A(n24306), .B(n24308), .Z(n12159) );
  NAND U26361 ( .A(n24314), .B(nreg[24]), .Z(n24308) );
  NAND U26362 ( .A(n12326), .B(nreg[24]), .Z(n24314) );
  XNOR U26363 ( .A(n24304), .B(n24315), .Z(n24306) );
  XOR U26364 ( .A(n24316), .B(n24317), .Z(n24304) );
  AND U26365 ( .A(n24318), .B(n24319), .Z(n24317) );
  XNOR U26366 ( .A(n24320), .B(n24316), .Z(n24319) );
  XOR U26367 ( .A(n24321), .B(nreg[24]), .Z(n24312) );
  IV U26368 ( .A(n24310), .Z(n24321) );
  XOR U26369 ( .A(n24322), .B(n24323), .Z(n24310) );
  AND U26370 ( .A(n24324), .B(n24325), .Z(n24323) );
  XNOR U26371 ( .A(n24322), .B(n12165), .Z(n24325) );
  XNOR U26372 ( .A(n24318), .B(n24320), .Z(n12165) );
  NAND U26373 ( .A(n24326), .B(nreg[23]), .Z(n24320) );
  NAND U26374 ( .A(n12326), .B(nreg[23]), .Z(n24326) );
  XNOR U26375 ( .A(n24316), .B(n24327), .Z(n24318) );
  XOR U26376 ( .A(n24328), .B(n24329), .Z(n24316) );
  AND U26377 ( .A(n24330), .B(n24331), .Z(n24329) );
  XNOR U26378 ( .A(n24332), .B(n24328), .Z(n24331) );
  XOR U26379 ( .A(n24333), .B(nreg[23]), .Z(n24324) );
  IV U26380 ( .A(n24322), .Z(n24333) );
  XOR U26381 ( .A(n24334), .B(n24335), .Z(n24322) );
  AND U26382 ( .A(n24336), .B(n24337), .Z(n24335) );
  XNOR U26383 ( .A(n24334), .B(n12171), .Z(n24337) );
  XNOR U26384 ( .A(n24330), .B(n24332), .Z(n12171) );
  NAND U26385 ( .A(n24338), .B(nreg[22]), .Z(n24332) );
  NAND U26386 ( .A(n12326), .B(nreg[22]), .Z(n24338) );
  XNOR U26387 ( .A(n24328), .B(n24339), .Z(n24330) );
  XOR U26388 ( .A(n24340), .B(n24341), .Z(n24328) );
  AND U26389 ( .A(n24342), .B(n24343), .Z(n24341) );
  XNOR U26390 ( .A(n24344), .B(n24340), .Z(n24343) );
  XOR U26391 ( .A(n24345), .B(nreg[22]), .Z(n24336) );
  IV U26392 ( .A(n24334), .Z(n24345) );
  XOR U26393 ( .A(n24346), .B(n24347), .Z(n24334) );
  AND U26394 ( .A(n24348), .B(n24349), .Z(n24347) );
  XNOR U26395 ( .A(n24346), .B(n12177), .Z(n24349) );
  XNOR U26396 ( .A(n24342), .B(n24344), .Z(n12177) );
  NAND U26397 ( .A(n24350), .B(nreg[21]), .Z(n24344) );
  NAND U26398 ( .A(n12326), .B(nreg[21]), .Z(n24350) );
  XNOR U26399 ( .A(n24340), .B(n24351), .Z(n24342) );
  XOR U26400 ( .A(n24352), .B(n24353), .Z(n24340) );
  AND U26401 ( .A(n24354), .B(n24355), .Z(n24353) );
  XNOR U26402 ( .A(n24356), .B(n24352), .Z(n24355) );
  XOR U26403 ( .A(n24357), .B(nreg[21]), .Z(n24348) );
  IV U26404 ( .A(n24346), .Z(n24357) );
  XOR U26405 ( .A(n24358), .B(n24359), .Z(n24346) );
  AND U26406 ( .A(n24360), .B(n24361), .Z(n24359) );
  XNOR U26407 ( .A(n24358), .B(n12183), .Z(n24361) );
  XNOR U26408 ( .A(n24354), .B(n24356), .Z(n12183) );
  NAND U26409 ( .A(n24362), .B(nreg[20]), .Z(n24356) );
  NAND U26410 ( .A(n12326), .B(nreg[20]), .Z(n24362) );
  XNOR U26411 ( .A(n24352), .B(n24363), .Z(n24354) );
  XOR U26412 ( .A(n24364), .B(n24365), .Z(n24352) );
  AND U26413 ( .A(n24366), .B(n24367), .Z(n24365) );
  XNOR U26414 ( .A(n24368), .B(n24364), .Z(n24367) );
  XOR U26415 ( .A(n24369), .B(nreg[20]), .Z(n24360) );
  IV U26416 ( .A(n24358), .Z(n24369) );
  XOR U26417 ( .A(n24370), .B(n24371), .Z(n24358) );
  AND U26418 ( .A(n24372), .B(n24373), .Z(n24371) );
  XNOR U26419 ( .A(n24370), .B(n12189), .Z(n24373) );
  XNOR U26420 ( .A(n24366), .B(n24368), .Z(n12189) );
  NAND U26421 ( .A(n24374), .B(nreg[19]), .Z(n24368) );
  NAND U26422 ( .A(n12326), .B(nreg[19]), .Z(n24374) );
  XNOR U26423 ( .A(n24364), .B(n24375), .Z(n24366) );
  XOR U26424 ( .A(n24376), .B(n24377), .Z(n24364) );
  AND U26425 ( .A(n24378), .B(n24379), .Z(n24377) );
  XNOR U26426 ( .A(n24380), .B(n24376), .Z(n24379) );
  XOR U26427 ( .A(n24381), .B(nreg[19]), .Z(n24372) );
  IV U26428 ( .A(n24370), .Z(n24381) );
  XOR U26429 ( .A(n24382), .B(n24383), .Z(n24370) );
  AND U26430 ( .A(n24384), .B(n24385), .Z(n24383) );
  XNOR U26431 ( .A(n24382), .B(n12195), .Z(n24385) );
  XNOR U26432 ( .A(n24378), .B(n24380), .Z(n12195) );
  NAND U26433 ( .A(n24386), .B(nreg[18]), .Z(n24380) );
  NAND U26434 ( .A(n12326), .B(nreg[18]), .Z(n24386) );
  XNOR U26435 ( .A(n24376), .B(n24387), .Z(n24378) );
  XOR U26436 ( .A(n24388), .B(n24389), .Z(n24376) );
  AND U26437 ( .A(n24390), .B(n24391), .Z(n24389) );
  XNOR U26438 ( .A(n24392), .B(n24388), .Z(n24391) );
  XOR U26439 ( .A(n24393), .B(nreg[18]), .Z(n24384) );
  IV U26440 ( .A(n24382), .Z(n24393) );
  XOR U26441 ( .A(n24394), .B(n24395), .Z(n24382) );
  AND U26442 ( .A(n24396), .B(n24397), .Z(n24395) );
  XNOR U26443 ( .A(n24394), .B(n12201), .Z(n24397) );
  XNOR U26444 ( .A(n24390), .B(n24392), .Z(n12201) );
  NAND U26445 ( .A(n24398), .B(nreg[17]), .Z(n24392) );
  NAND U26446 ( .A(n12326), .B(nreg[17]), .Z(n24398) );
  XNOR U26447 ( .A(n24388), .B(n24399), .Z(n24390) );
  XOR U26448 ( .A(n24400), .B(n24401), .Z(n24388) );
  AND U26449 ( .A(n24402), .B(n24403), .Z(n24401) );
  XNOR U26450 ( .A(n24404), .B(n24400), .Z(n24403) );
  XOR U26451 ( .A(n24405), .B(nreg[17]), .Z(n24396) );
  IV U26452 ( .A(n24394), .Z(n24405) );
  XOR U26453 ( .A(n24406), .B(n24407), .Z(n24394) );
  AND U26454 ( .A(n24408), .B(n24409), .Z(n24407) );
  XNOR U26455 ( .A(n24406), .B(n12207), .Z(n24409) );
  XNOR U26456 ( .A(n24402), .B(n24404), .Z(n12207) );
  NAND U26457 ( .A(n24410), .B(nreg[16]), .Z(n24404) );
  NAND U26458 ( .A(n12326), .B(nreg[16]), .Z(n24410) );
  XNOR U26459 ( .A(n24400), .B(n24411), .Z(n24402) );
  XOR U26460 ( .A(n24412), .B(n24413), .Z(n24400) );
  AND U26461 ( .A(n24414), .B(n24415), .Z(n24413) );
  XNOR U26462 ( .A(n24416), .B(n24412), .Z(n24415) );
  XOR U26463 ( .A(n24417), .B(nreg[16]), .Z(n24408) );
  IV U26464 ( .A(n24406), .Z(n24417) );
  XOR U26465 ( .A(n24418), .B(n24419), .Z(n24406) );
  AND U26466 ( .A(n24420), .B(n24421), .Z(n24419) );
  XNOR U26467 ( .A(n24418), .B(n12213), .Z(n24421) );
  XNOR U26468 ( .A(n24414), .B(n24416), .Z(n12213) );
  NAND U26469 ( .A(n24422), .B(nreg[15]), .Z(n24416) );
  NAND U26470 ( .A(n12326), .B(nreg[15]), .Z(n24422) );
  XNOR U26471 ( .A(n24412), .B(n24423), .Z(n24414) );
  XOR U26472 ( .A(n24424), .B(n24425), .Z(n24412) );
  AND U26473 ( .A(n24426), .B(n24427), .Z(n24425) );
  XNOR U26474 ( .A(n24428), .B(n24424), .Z(n24427) );
  XOR U26475 ( .A(n24429), .B(nreg[15]), .Z(n24420) );
  IV U26476 ( .A(n24418), .Z(n24429) );
  XOR U26477 ( .A(n24430), .B(n24431), .Z(n24418) );
  AND U26478 ( .A(n24432), .B(n24433), .Z(n24431) );
  XNOR U26479 ( .A(n24430), .B(n12219), .Z(n24433) );
  XNOR U26480 ( .A(n24426), .B(n24428), .Z(n12219) );
  NAND U26481 ( .A(n24434), .B(nreg[14]), .Z(n24428) );
  NAND U26482 ( .A(n12326), .B(nreg[14]), .Z(n24434) );
  XNOR U26483 ( .A(n24424), .B(n24435), .Z(n24426) );
  XOR U26484 ( .A(n24436), .B(n24437), .Z(n24424) );
  AND U26485 ( .A(n24438), .B(n24439), .Z(n24437) );
  XNOR U26486 ( .A(n24440), .B(n24436), .Z(n24439) );
  XOR U26487 ( .A(n24441), .B(nreg[14]), .Z(n24432) );
  IV U26488 ( .A(n24430), .Z(n24441) );
  XOR U26489 ( .A(n24442), .B(n24443), .Z(n24430) );
  AND U26490 ( .A(n24444), .B(n24445), .Z(n24443) );
  XNOR U26491 ( .A(n24442), .B(n12225), .Z(n24445) );
  XNOR U26492 ( .A(n24438), .B(n24440), .Z(n12225) );
  NAND U26493 ( .A(n24446), .B(nreg[13]), .Z(n24440) );
  NAND U26494 ( .A(n12326), .B(nreg[13]), .Z(n24446) );
  XNOR U26495 ( .A(n24436), .B(n24447), .Z(n24438) );
  XOR U26496 ( .A(n24448), .B(n24449), .Z(n24436) );
  AND U26497 ( .A(n24450), .B(n24451), .Z(n24449) );
  XNOR U26498 ( .A(n24452), .B(n24448), .Z(n24451) );
  XOR U26499 ( .A(n24453), .B(nreg[13]), .Z(n24444) );
  IV U26500 ( .A(n24442), .Z(n24453) );
  XOR U26501 ( .A(n24454), .B(n24455), .Z(n24442) );
  AND U26502 ( .A(n24456), .B(n24457), .Z(n24455) );
  XNOR U26503 ( .A(n24454), .B(n12231), .Z(n24457) );
  XNOR U26504 ( .A(n24450), .B(n24452), .Z(n12231) );
  NAND U26505 ( .A(n24458), .B(nreg[12]), .Z(n24452) );
  NAND U26506 ( .A(n12326), .B(nreg[12]), .Z(n24458) );
  XNOR U26507 ( .A(n24448), .B(n24459), .Z(n24450) );
  XOR U26508 ( .A(n24460), .B(n24461), .Z(n24448) );
  AND U26509 ( .A(n24462), .B(n24463), .Z(n24461) );
  XNOR U26510 ( .A(n24464), .B(n24460), .Z(n24463) );
  XOR U26511 ( .A(n24465), .B(nreg[12]), .Z(n24456) );
  IV U26512 ( .A(n24454), .Z(n24465) );
  XOR U26513 ( .A(n24466), .B(n24467), .Z(n24454) );
  AND U26514 ( .A(n24468), .B(n24469), .Z(n24467) );
  XNOR U26515 ( .A(n24466), .B(n12237), .Z(n24469) );
  XNOR U26516 ( .A(n24462), .B(n24464), .Z(n12237) );
  NAND U26517 ( .A(n24470), .B(nreg[11]), .Z(n24464) );
  NAND U26518 ( .A(n12326), .B(nreg[11]), .Z(n24470) );
  XNOR U26519 ( .A(n24460), .B(n24471), .Z(n24462) );
  XOR U26520 ( .A(n24472), .B(n24473), .Z(n24460) );
  AND U26521 ( .A(n24474), .B(n24475), .Z(n24473) );
  XNOR U26522 ( .A(n24476), .B(n24472), .Z(n24475) );
  XOR U26523 ( .A(n24477), .B(nreg[11]), .Z(n24468) );
  IV U26524 ( .A(n24466), .Z(n24477) );
  XOR U26525 ( .A(n24478), .B(n24479), .Z(n24466) );
  AND U26526 ( .A(n24480), .B(n24481), .Z(n24479) );
  XNOR U26527 ( .A(n24478), .B(n12243), .Z(n24481) );
  XNOR U26528 ( .A(n24474), .B(n24476), .Z(n12243) );
  NAND U26529 ( .A(n24482), .B(nreg[10]), .Z(n24476) );
  NAND U26530 ( .A(n12326), .B(nreg[10]), .Z(n24482) );
  XNOR U26531 ( .A(n24472), .B(n24483), .Z(n24474) );
  XOR U26532 ( .A(n24484), .B(n24485), .Z(n24472) );
  AND U26533 ( .A(n24486), .B(n24487), .Z(n24485) );
  XNOR U26534 ( .A(n24488), .B(n24484), .Z(n24487) );
  XOR U26535 ( .A(n24489), .B(nreg[10]), .Z(n24480) );
  IV U26536 ( .A(n24478), .Z(n24489) );
  XOR U26537 ( .A(n24490), .B(n24491), .Z(n24478) );
  AND U26538 ( .A(n24492), .B(n24493), .Z(n24491) );
  XNOR U26539 ( .A(n12249), .B(n24490), .Z(n24493) );
  XNOR U26540 ( .A(n24486), .B(n24488), .Z(n12249) );
  NAND U26541 ( .A(n24494), .B(nreg[9]), .Z(n24488) );
  NAND U26542 ( .A(n12326), .B(nreg[9]), .Z(n24494) );
  XNOR U26543 ( .A(n24484), .B(n24495), .Z(n24486) );
  XOR U26544 ( .A(n24496), .B(n24497), .Z(n24484) );
  AND U26545 ( .A(n24498), .B(n24499), .Z(n24497) );
  XNOR U26546 ( .A(n24500), .B(n24496), .Z(n24499) );
  XOR U26547 ( .A(n24501), .B(nreg[9]), .Z(n24492) );
  IV U26548 ( .A(n24490), .Z(n24501) );
  XOR U26549 ( .A(n24502), .B(n24503), .Z(n24490) );
  AND U26550 ( .A(n24504), .B(n24505), .Z(n24503) );
  XNOR U26551 ( .A(n24502), .B(n12255), .Z(n24505) );
  XNOR U26552 ( .A(n24498), .B(n24500), .Z(n12255) );
  NAND U26553 ( .A(n24506), .B(nreg[8]), .Z(n24500) );
  NAND U26554 ( .A(n12326), .B(nreg[8]), .Z(n24506) );
  XNOR U26555 ( .A(n24496), .B(n24507), .Z(n24498) );
  XOR U26556 ( .A(n24508), .B(n24509), .Z(n24496) );
  AND U26557 ( .A(n24510), .B(n24511), .Z(n24509) );
  XNOR U26558 ( .A(n24512), .B(n24508), .Z(n24511) );
  XOR U26559 ( .A(n24513), .B(nreg[8]), .Z(n24504) );
  IV U26560 ( .A(n24502), .Z(n24513) );
  XOR U26561 ( .A(n24514), .B(n24515), .Z(n24502) );
  AND U26562 ( .A(n24516), .B(n24517), .Z(n24515) );
  XNOR U26563 ( .A(n24514), .B(n12264), .Z(n24517) );
  XNOR U26564 ( .A(n24510), .B(n24512), .Z(n12264) );
  NAND U26565 ( .A(n24518), .B(nreg[7]), .Z(n24512) );
  NAND U26566 ( .A(n12326), .B(nreg[7]), .Z(n24518) );
  XNOR U26567 ( .A(n24508), .B(n24519), .Z(n24510) );
  XOR U26568 ( .A(n24520), .B(n24521), .Z(n24508) );
  AND U26569 ( .A(n24522), .B(n24523), .Z(n24521) );
  XNOR U26570 ( .A(n24524), .B(n24520), .Z(n24523) );
  XOR U26571 ( .A(n24525), .B(nreg[7]), .Z(n24516) );
  IV U26572 ( .A(n24514), .Z(n24525) );
  XOR U26573 ( .A(n24526), .B(n24527), .Z(n24514) );
  AND U26574 ( .A(n24528), .B(n24529), .Z(n24527) );
  XNOR U26575 ( .A(n24526), .B(n12269), .Z(n24529) );
  XNOR U26576 ( .A(n24522), .B(n24524), .Z(n12269) );
  NAND U26577 ( .A(n24530), .B(nreg[6]), .Z(n24524) );
  NAND U26578 ( .A(n12326), .B(nreg[6]), .Z(n24530) );
  XNOR U26579 ( .A(n24520), .B(n24531), .Z(n24522) );
  XOR U26580 ( .A(n24532), .B(n24533), .Z(n24520) );
  AND U26581 ( .A(n24534), .B(n24535), .Z(n24533) );
  XNOR U26582 ( .A(n24536), .B(n24532), .Z(n24535) );
  XOR U26583 ( .A(n24537), .B(nreg[6]), .Z(n24528) );
  IV U26584 ( .A(n24526), .Z(n24537) );
  XOR U26585 ( .A(n24538), .B(n24539), .Z(n24526) );
  AND U26586 ( .A(n24540), .B(n24541), .Z(n24539) );
  XNOR U26587 ( .A(n24538), .B(n12275), .Z(n24541) );
  XNOR U26588 ( .A(n24534), .B(n24536), .Z(n12275) );
  NAND U26589 ( .A(n24542), .B(nreg[5]), .Z(n24536) );
  NAND U26590 ( .A(n12326), .B(nreg[5]), .Z(n24542) );
  XNOR U26591 ( .A(n24532), .B(n24543), .Z(n24534) );
  XOR U26592 ( .A(n24544), .B(n24545), .Z(n24532) );
  AND U26593 ( .A(n24546), .B(n24547), .Z(n24545) );
  XNOR U26594 ( .A(n24548), .B(n24544), .Z(n24547) );
  XOR U26595 ( .A(n24549), .B(nreg[5]), .Z(n24540) );
  IV U26596 ( .A(n24538), .Z(n24549) );
  XOR U26597 ( .A(n24550), .B(n24551), .Z(n24538) );
  AND U26598 ( .A(n24552), .B(n24553), .Z(n24551) );
  XNOR U26599 ( .A(n24550), .B(n12281), .Z(n24553) );
  XNOR U26600 ( .A(n24546), .B(n24548), .Z(n12281) );
  NAND U26601 ( .A(n24554), .B(nreg[4]), .Z(n24548) );
  NAND U26602 ( .A(n12326), .B(nreg[4]), .Z(n24554) );
  XNOR U26603 ( .A(n24544), .B(n24555), .Z(n24546) );
  XOR U26604 ( .A(n24556), .B(n24557), .Z(n24544) );
  AND U26605 ( .A(n24558), .B(n24559), .Z(n24557) );
  XNOR U26606 ( .A(n24560), .B(n24556), .Z(n24559) );
  XOR U26607 ( .A(n24561), .B(nreg[4]), .Z(n24552) );
  IV U26608 ( .A(n24550), .Z(n24561) );
  XOR U26609 ( .A(n24562), .B(n24563), .Z(n24550) );
  AND U26610 ( .A(n24564), .B(n24565), .Z(n24563) );
  XNOR U26611 ( .A(n24562), .B(n12287), .Z(n24565) );
  XNOR U26612 ( .A(n24558), .B(n24560), .Z(n12287) );
  NAND U26613 ( .A(n24566), .B(nreg[3]), .Z(n24560) );
  NAND U26614 ( .A(n12326), .B(nreg[3]), .Z(n24566) );
  XNOR U26615 ( .A(n24556), .B(n24567), .Z(n24558) );
  XOR U26616 ( .A(n24568), .B(n24569), .Z(n24556) );
  AND U26617 ( .A(n24570), .B(n24571), .Z(n24569) );
  XNOR U26618 ( .A(n24572), .B(n24568), .Z(n24571) );
  XOR U26619 ( .A(n24573), .B(nreg[3]), .Z(n24564) );
  IV U26620 ( .A(n24562), .Z(n24573) );
  XNOR U26621 ( .A(n24574), .B(n24575), .Z(n24562) );
  AND U26622 ( .A(n24576), .B(n24577), .Z(n24575) );
  XOR U26623 ( .A(n24574), .B(n12292), .Z(n24577) );
  XNOR U26624 ( .A(n24570), .B(n24572), .Z(n12292) );
  NAND U26625 ( .A(n24578), .B(nreg[2]), .Z(n24572) );
  NAND U26626 ( .A(n12326), .B(nreg[2]), .Z(n24578) );
  XOR U26627 ( .A(n24568), .B(n24579), .Z(n24570) );
  XOR U26628 ( .A(n24580), .B(n24581), .Z(n24568) );
  NANDN U26629 ( .B(n24582), .A(n24583), .Z(n24580) );
  XOR U26630 ( .A(n24581), .B(n24584), .Z(n24583) );
  XOR U26631 ( .A(n24574), .B(nreg[2]), .Z(n24576) );
  XOR U26632 ( .A(n24585), .B(n24586), .Z(n24574) );
  NAND U26633 ( .A(n24587), .B(n24588), .Z(n24585) );
  XOR U26634 ( .A(n24586), .B(n12299), .Z(n24588) );
  XNOR U26635 ( .A(n24586), .B(nreg[1]), .Z(n24587) );
  NOR U26636 ( .A(nreg[0]), .B(n5663), .Z(n24586) );
  XOR U26637 ( .A(n24589), .B(n24590), .Z(n5663) );
  XNOR U26638 ( .A(n24582), .B(n24584), .Z(n12299) );
  NAND U26639 ( .A(n24591), .B(nreg[1]), .Z(n24584) );
  NAND U26640 ( .A(n12326), .B(nreg[1]), .Z(n24591) );
  XNOR U26641 ( .A(n24592), .B(n24581), .Z(n24582) );
  OR U26642 ( .A(n24589), .B(n24590), .Z(n24581) );
  NAND U26643 ( .A(n24593), .B(nreg[0]), .Z(n24590) );
  NAND U26644 ( .A(n12326), .B(nreg[0]), .Z(n24593) );
  NAND U26645 ( .A(n24594), .B(n24595), .Z(n12326) );
  NAND U26646 ( .A(n24596), .B(n24595), .Z(n24594) );
  XOR U26647 ( .A(n12309), .B(n24595), .Z(n24596) );
  AND U26648 ( .A(n24597), .B(n24598), .Z(n24595) );
  NAND U26649 ( .A(n24599), .B(n24598), .Z(n24597) );
  XNOR U26650 ( .A(n12315), .B(n24598), .Z(n24599) );
  XOR U26651 ( .A(n24600), .B(n24601), .Z(n24598) );
  AND U26652 ( .A(n24602), .B(n24603), .Z(n24601) );
  XOR U26653 ( .A(nreg[1023]), .B(n24600), .Z(n24603) );
  XNOR U26654 ( .A(n12327), .B(n24600), .Z(n24602) );
  XOR U26655 ( .A(n24604), .B(n24605), .Z(n12327) );
  XOR U26656 ( .A(n24606), .B(n24607), .Z(n24600) );
  AND U26657 ( .A(n24608), .B(n24609), .Z(n24607) );
  XOR U26658 ( .A(nreg[1022]), .B(n24606), .Z(n24609) );
  XNOR U26659 ( .A(n12339), .B(n24606), .Z(n24608) );
  XOR U26660 ( .A(n24610), .B(n24611), .Z(n12339) );
  XOR U26661 ( .A(n24612), .B(n24613), .Z(n24606) );
  AND U26662 ( .A(n24614), .B(n24615), .Z(n24613) );
  XOR U26663 ( .A(nreg[1021]), .B(n24612), .Z(n24615) );
  XNOR U26664 ( .A(n12351), .B(n24612), .Z(n24614) );
  XOR U26665 ( .A(n24616), .B(n24617), .Z(n12351) );
  XOR U26666 ( .A(n24618), .B(n24619), .Z(n24612) );
  AND U26667 ( .A(n24620), .B(n24621), .Z(n24619) );
  XOR U26668 ( .A(nreg[1020]), .B(n24618), .Z(n24621) );
  XNOR U26669 ( .A(n12363), .B(n24618), .Z(n24620) );
  XOR U26670 ( .A(n24622), .B(n24623), .Z(n12363) );
  XOR U26671 ( .A(n24624), .B(n24625), .Z(n24618) );
  AND U26672 ( .A(n24626), .B(n24627), .Z(n24625) );
  XOR U26673 ( .A(nreg[1019]), .B(n24624), .Z(n24627) );
  XNOR U26674 ( .A(n12375), .B(n24624), .Z(n24626) );
  XOR U26675 ( .A(n24628), .B(n24629), .Z(n12375) );
  XOR U26676 ( .A(n24630), .B(n24631), .Z(n24624) );
  AND U26677 ( .A(n24632), .B(n24633), .Z(n24631) );
  XOR U26678 ( .A(nreg[1018]), .B(n24630), .Z(n24633) );
  XNOR U26679 ( .A(n12387), .B(n24630), .Z(n24632) );
  XOR U26680 ( .A(n24634), .B(n24635), .Z(n12387) );
  XOR U26681 ( .A(n24636), .B(n24637), .Z(n24630) );
  AND U26682 ( .A(n24638), .B(n24639), .Z(n24637) );
  XOR U26683 ( .A(nreg[1017]), .B(n24636), .Z(n24639) );
  XNOR U26684 ( .A(n12399), .B(n24636), .Z(n24638) );
  XOR U26685 ( .A(n24640), .B(n24641), .Z(n12399) );
  XOR U26686 ( .A(n24642), .B(n24643), .Z(n24636) );
  AND U26687 ( .A(n24644), .B(n24645), .Z(n24643) );
  XOR U26688 ( .A(nreg[1016]), .B(n24642), .Z(n24645) );
  XNOR U26689 ( .A(n12411), .B(n24642), .Z(n24644) );
  XOR U26690 ( .A(n24646), .B(n24647), .Z(n12411) );
  XOR U26691 ( .A(n24648), .B(n24649), .Z(n24642) );
  AND U26692 ( .A(n24650), .B(n24651), .Z(n24649) );
  XOR U26693 ( .A(nreg[1015]), .B(n24648), .Z(n24651) );
  XNOR U26694 ( .A(n12423), .B(n24648), .Z(n24650) );
  XOR U26695 ( .A(n24652), .B(n24653), .Z(n12423) );
  XOR U26696 ( .A(n24654), .B(n24655), .Z(n24648) );
  AND U26697 ( .A(n24656), .B(n24657), .Z(n24655) );
  XOR U26698 ( .A(nreg[1014]), .B(n24654), .Z(n24657) );
  XNOR U26699 ( .A(n12435), .B(n24654), .Z(n24656) );
  XOR U26700 ( .A(n24658), .B(n24659), .Z(n12435) );
  XOR U26701 ( .A(n24660), .B(n24661), .Z(n24654) );
  AND U26702 ( .A(n24662), .B(n24663), .Z(n24661) );
  XOR U26703 ( .A(nreg[1013]), .B(n24660), .Z(n24663) );
  XNOR U26704 ( .A(n12447), .B(n24660), .Z(n24662) );
  XOR U26705 ( .A(n24664), .B(n24665), .Z(n12447) );
  XOR U26706 ( .A(n24666), .B(n24667), .Z(n24660) );
  AND U26707 ( .A(n24668), .B(n24669), .Z(n24667) );
  XOR U26708 ( .A(nreg[1012]), .B(n24666), .Z(n24669) );
  XNOR U26709 ( .A(n12459), .B(n24666), .Z(n24668) );
  XOR U26710 ( .A(n24670), .B(n24671), .Z(n12459) );
  XOR U26711 ( .A(n24672), .B(n24673), .Z(n24666) );
  AND U26712 ( .A(n24674), .B(n24675), .Z(n24673) );
  XOR U26713 ( .A(nreg[1011]), .B(n24672), .Z(n24675) );
  XNOR U26714 ( .A(n12471), .B(n24672), .Z(n24674) );
  XOR U26715 ( .A(n24676), .B(n24677), .Z(n12471) );
  XOR U26716 ( .A(n24678), .B(n24679), .Z(n24672) );
  AND U26717 ( .A(n24680), .B(n24681), .Z(n24679) );
  XOR U26718 ( .A(nreg[1010]), .B(n24678), .Z(n24681) );
  XNOR U26719 ( .A(n12483), .B(n24678), .Z(n24680) );
  XOR U26720 ( .A(n24682), .B(n24683), .Z(n12483) );
  XOR U26721 ( .A(n24684), .B(n24685), .Z(n24678) );
  AND U26722 ( .A(n24686), .B(n24687), .Z(n24685) );
  XOR U26723 ( .A(nreg[1009]), .B(n24684), .Z(n24687) );
  XNOR U26724 ( .A(n12495), .B(n24684), .Z(n24686) );
  XOR U26725 ( .A(n24688), .B(n24689), .Z(n12495) );
  XOR U26726 ( .A(n24690), .B(n24691), .Z(n24684) );
  AND U26727 ( .A(n24692), .B(n24693), .Z(n24691) );
  XOR U26728 ( .A(nreg[1008]), .B(n24690), .Z(n24693) );
  XNOR U26729 ( .A(n12507), .B(n24690), .Z(n24692) );
  XOR U26730 ( .A(n24694), .B(n24695), .Z(n12507) );
  XOR U26731 ( .A(n24696), .B(n24697), .Z(n24690) );
  AND U26732 ( .A(n24698), .B(n24699), .Z(n24697) );
  XOR U26733 ( .A(nreg[1007]), .B(n24696), .Z(n24699) );
  XNOR U26734 ( .A(n12519), .B(n24696), .Z(n24698) );
  XOR U26735 ( .A(n24700), .B(n24701), .Z(n12519) );
  XOR U26736 ( .A(n24702), .B(n24703), .Z(n24696) );
  AND U26737 ( .A(n24704), .B(n24705), .Z(n24703) );
  XOR U26738 ( .A(nreg[1006]), .B(n24702), .Z(n24705) );
  XNOR U26739 ( .A(n12531), .B(n24702), .Z(n24704) );
  XOR U26740 ( .A(n24706), .B(n24707), .Z(n12531) );
  XOR U26741 ( .A(n24708), .B(n24709), .Z(n24702) );
  AND U26742 ( .A(n24710), .B(n24711), .Z(n24709) );
  XOR U26743 ( .A(nreg[1005]), .B(n24708), .Z(n24711) );
  XNOR U26744 ( .A(n12543), .B(n24708), .Z(n24710) );
  XOR U26745 ( .A(n24712), .B(n24713), .Z(n12543) );
  XOR U26746 ( .A(n24714), .B(n24715), .Z(n24708) );
  AND U26747 ( .A(n24716), .B(n24717), .Z(n24715) );
  XOR U26748 ( .A(nreg[1004]), .B(n24714), .Z(n24717) );
  XNOR U26749 ( .A(n12555), .B(n24714), .Z(n24716) );
  XOR U26750 ( .A(n24718), .B(n24719), .Z(n12555) );
  XOR U26751 ( .A(n24720), .B(n24721), .Z(n24714) );
  AND U26752 ( .A(n24722), .B(n24723), .Z(n24721) );
  XOR U26753 ( .A(nreg[1003]), .B(n24720), .Z(n24723) );
  XNOR U26754 ( .A(n12567), .B(n24720), .Z(n24722) );
  XOR U26755 ( .A(n24724), .B(n24725), .Z(n12567) );
  XOR U26756 ( .A(n24726), .B(n24727), .Z(n24720) );
  AND U26757 ( .A(n24728), .B(n24729), .Z(n24727) );
  XOR U26758 ( .A(nreg[1002]), .B(n24726), .Z(n24729) );
  XNOR U26759 ( .A(n12579), .B(n24726), .Z(n24728) );
  XOR U26760 ( .A(n24730), .B(n24731), .Z(n12579) );
  XOR U26761 ( .A(n24732), .B(n24733), .Z(n24726) );
  AND U26762 ( .A(n24734), .B(n24735), .Z(n24733) );
  XOR U26763 ( .A(nreg[1001]), .B(n24732), .Z(n24735) );
  XNOR U26764 ( .A(n12591), .B(n24732), .Z(n24734) );
  XOR U26765 ( .A(n24736), .B(n24737), .Z(n12591) );
  XOR U26766 ( .A(n24738), .B(n24739), .Z(n24732) );
  AND U26767 ( .A(n24740), .B(n24741), .Z(n24739) );
  XOR U26768 ( .A(nreg[1000]), .B(n24738), .Z(n24741) );
  XNOR U26769 ( .A(n12603), .B(n24738), .Z(n24740) );
  XOR U26770 ( .A(n24742), .B(n24743), .Z(n12603) );
  XOR U26771 ( .A(n24744), .B(n24745), .Z(n24738) );
  AND U26772 ( .A(n24746), .B(n24747), .Z(n24745) );
  XOR U26773 ( .A(nreg[999]), .B(n24744), .Z(n24747) );
  XNOR U26774 ( .A(n12615), .B(n24744), .Z(n24746) );
  XOR U26775 ( .A(n24748), .B(n24749), .Z(n12615) );
  XOR U26776 ( .A(n24750), .B(n24751), .Z(n24744) );
  AND U26777 ( .A(n24752), .B(n24753), .Z(n24751) );
  XOR U26778 ( .A(nreg[998]), .B(n24750), .Z(n24753) );
  XNOR U26779 ( .A(n12627), .B(n24750), .Z(n24752) );
  XOR U26780 ( .A(n24754), .B(n24755), .Z(n12627) );
  XOR U26781 ( .A(n24756), .B(n24757), .Z(n24750) );
  AND U26782 ( .A(n24758), .B(n24759), .Z(n24757) );
  XOR U26783 ( .A(nreg[997]), .B(n24756), .Z(n24759) );
  XNOR U26784 ( .A(n12639), .B(n24756), .Z(n24758) );
  XOR U26785 ( .A(n24760), .B(n24761), .Z(n12639) );
  XOR U26786 ( .A(n24762), .B(n24763), .Z(n24756) );
  AND U26787 ( .A(n24764), .B(n24765), .Z(n24763) );
  XOR U26788 ( .A(nreg[996]), .B(n24762), .Z(n24765) );
  XNOR U26789 ( .A(n12651), .B(n24762), .Z(n24764) );
  XOR U26790 ( .A(n24766), .B(n24767), .Z(n12651) );
  XOR U26791 ( .A(n24768), .B(n24769), .Z(n24762) );
  AND U26792 ( .A(n24770), .B(n24771), .Z(n24769) );
  XOR U26793 ( .A(nreg[995]), .B(n24768), .Z(n24771) );
  XNOR U26794 ( .A(n12663), .B(n24768), .Z(n24770) );
  XOR U26795 ( .A(n24772), .B(n24773), .Z(n12663) );
  XOR U26796 ( .A(n24774), .B(n24775), .Z(n24768) );
  AND U26797 ( .A(n24776), .B(n24777), .Z(n24775) );
  XOR U26798 ( .A(nreg[994]), .B(n24774), .Z(n24777) );
  XNOR U26799 ( .A(n12675), .B(n24774), .Z(n24776) );
  XOR U26800 ( .A(n24778), .B(n24779), .Z(n12675) );
  XOR U26801 ( .A(n24780), .B(n24781), .Z(n24774) );
  AND U26802 ( .A(n24782), .B(n24783), .Z(n24781) );
  XOR U26803 ( .A(nreg[993]), .B(n24780), .Z(n24783) );
  XNOR U26804 ( .A(n12687), .B(n24780), .Z(n24782) );
  XOR U26805 ( .A(n24784), .B(n24785), .Z(n12687) );
  XOR U26806 ( .A(n24786), .B(n24787), .Z(n24780) );
  AND U26807 ( .A(n24788), .B(n24789), .Z(n24787) );
  XOR U26808 ( .A(nreg[992]), .B(n24786), .Z(n24789) );
  XNOR U26809 ( .A(n12699), .B(n24786), .Z(n24788) );
  XOR U26810 ( .A(n24790), .B(n24791), .Z(n12699) );
  XOR U26811 ( .A(n24792), .B(n24793), .Z(n24786) );
  AND U26812 ( .A(n24794), .B(n24795), .Z(n24793) );
  XOR U26813 ( .A(nreg[991]), .B(n24792), .Z(n24795) );
  XNOR U26814 ( .A(n12711), .B(n24792), .Z(n24794) );
  XOR U26815 ( .A(n24796), .B(n24797), .Z(n12711) );
  XOR U26816 ( .A(n24798), .B(n24799), .Z(n24792) );
  AND U26817 ( .A(n24800), .B(n24801), .Z(n24799) );
  XOR U26818 ( .A(nreg[990]), .B(n24798), .Z(n24801) );
  XNOR U26819 ( .A(n12723), .B(n24798), .Z(n24800) );
  XOR U26820 ( .A(n24802), .B(n24803), .Z(n12723) );
  XOR U26821 ( .A(n24804), .B(n24805), .Z(n24798) );
  AND U26822 ( .A(n24806), .B(n24807), .Z(n24805) );
  XOR U26823 ( .A(nreg[989]), .B(n24804), .Z(n24807) );
  XNOR U26824 ( .A(n12735), .B(n24804), .Z(n24806) );
  XOR U26825 ( .A(n24808), .B(n24809), .Z(n12735) );
  XOR U26826 ( .A(n24810), .B(n24811), .Z(n24804) );
  AND U26827 ( .A(n24812), .B(n24813), .Z(n24811) );
  XOR U26828 ( .A(nreg[988]), .B(n24810), .Z(n24813) );
  XNOR U26829 ( .A(n12747), .B(n24810), .Z(n24812) );
  XOR U26830 ( .A(n24814), .B(n24815), .Z(n12747) );
  XOR U26831 ( .A(n24816), .B(n24817), .Z(n24810) );
  AND U26832 ( .A(n24818), .B(n24819), .Z(n24817) );
  XOR U26833 ( .A(nreg[987]), .B(n24816), .Z(n24819) );
  XNOR U26834 ( .A(n12759), .B(n24816), .Z(n24818) );
  XOR U26835 ( .A(n24820), .B(n24821), .Z(n12759) );
  XOR U26836 ( .A(n24822), .B(n24823), .Z(n24816) );
  AND U26837 ( .A(n24824), .B(n24825), .Z(n24823) );
  XOR U26838 ( .A(nreg[986]), .B(n24822), .Z(n24825) );
  XNOR U26839 ( .A(n12771), .B(n24822), .Z(n24824) );
  XOR U26840 ( .A(n24826), .B(n24827), .Z(n12771) );
  XOR U26841 ( .A(n24828), .B(n24829), .Z(n24822) );
  AND U26842 ( .A(n24830), .B(n24831), .Z(n24829) );
  XOR U26843 ( .A(nreg[985]), .B(n24828), .Z(n24831) );
  XNOR U26844 ( .A(n12783), .B(n24828), .Z(n24830) );
  XOR U26845 ( .A(n24832), .B(n24833), .Z(n12783) );
  XOR U26846 ( .A(n24834), .B(n24835), .Z(n24828) );
  AND U26847 ( .A(n24836), .B(n24837), .Z(n24835) );
  XOR U26848 ( .A(nreg[984]), .B(n24834), .Z(n24837) );
  XNOR U26849 ( .A(n12795), .B(n24834), .Z(n24836) );
  XOR U26850 ( .A(n24838), .B(n24839), .Z(n12795) );
  XOR U26851 ( .A(n24840), .B(n24841), .Z(n24834) );
  AND U26852 ( .A(n24842), .B(n24843), .Z(n24841) );
  XOR U26853 ( .A(nreg[983]), .B(n24840), .Z(n24843) );
  XNOR U26854 ( .A(n12807), .B(n24840), .Z(n24842) );
  XOR U26855 ( .A(n24844), .B(n24845), .Z(n12807) );
  XOR U26856 ( .A(n24846), .B(n24847), .Z(n24840) );
  AND U26857 ( .A(n24848), .B(n24849), .Z(n24847) );
  XOR U26858 ( .A(nreg[982]), .B(n24846), .Z(n24849) );
  XNOR U26859 ( .A(n12819), .B(n24846), .Z(n24848) );
  XOR U26860 ( .A(n24850), .B(n24851), .Z(n12819) );
  XOR U26861 ( .A(n24852), .B(n24853), .Z(n24846) );
  AND U26862 ( .A(n24854), .B(n24855), .Z(n24853) );
  XOR U26863 ( .A(nreg[981]), .B(n24852), .Z(n24855) );
  XNOR U26864 ( .A(n12831), .B(n24852), .Z(n24854) );
  XOR U26865 ( .A(n24856), .B(n24857), .Z(n12831) );
  XOR U26866 ( .A(n24858), .B(n24859), .Z(n24852) );
  AND U26867 ( .A(n24860), .B(n24861), .Z(n24859) );
  XOR U26868 ( .A(nreg[980]), .B(n24858), .Z(n24861) );
  XNOR U26869 ( .A(n12843), .B(n24858), .Z(n24860) );
  XOR U26870 ( .A(n24862), .B(n24863), .Z(n12843) );
  XOR U26871 ( .A(n24864), .B(n24865), .Z(n24858) );
  AND U26872 ( .A(n24866), .B(n24867), .Z(n24865) );
  XOR U26873 ( .A(nreg[979]), .B(n24864), .Z(n24867) );
  XNOR U26874 ( .A(n12855), .B(n24864), .Z(n24866) );
  XOR U26875 ( .A(n24868), .B(n24869), .Z(n12855) );
  XOR U26876 ( .A(n24870), .B(n24871), .Z(n24864) );
  AND U26877 ( .A(n24872), .B(n24873), .Z(n24871) );
  XOR U26878 ( .A(nreg[978]), .B(n24870), .Z(n24873) );
  XNOR U26879 ( .A(n12867), .B(n24870), .Z(n24872) );
  XOR U26880 ( .A(n24874), .B(n24875), .Z(n12867) );
  XOR U26881 ( .A(n24876), .B(n24877), .Z(n24870) );
  AND U26882 ( .A(n24878), .B(n24879), .Z(n24877) );
  XOR U26883 ( .A(nreg[977]), .B(n24876), .Z(n24879) );
  XNOR U26884 ( .A(n12879), .B(n24876), .Z(n24878) );
  XOR U26885 ( .A(n24880), .B(n24881), .Z(n12879) );
  XOR U26886 ( .A(n24882), .B(n24883), .Z(n24876) );
  AND U26887 ( .A(n24884), .B(n24885), .Z(n24883) );
  XOR U26888 ( .A(nreg[976]), .B(n24882), .Z(n24885) );
  XNOR U26889 ( .A(n12891), .B(n24882), .Z(n24884) );
  XOR U26890 ( .A(n24886), .B(n24887), .Z(n12891) );
  XOR U26891 ( .A(n24888), .B(n24889), .Z(n24882) );
  AND U26892 ( .A(n24890), .B(n24891), .Z(n24889) );
  XOR U26893 ( .A(nreg[975]), .B(n24888), .Z(n24891) );
  XNOR U26894 ( .A(n12903), .B(n24888), .Z(n24890) );
  XOR U26895 ( .A(n24892), .B(n24893), .Z(n12903) );
  XOR U26896 ( .A(n24894), .B(n24895), .Z(n24888) );
  AND U26897 ( .A(n24896), .B(n24897), .Z(n24895) );
  XOR U26898 ( .A(nreg[974]), .B(n24894), .Z(n24897) );
  XNOR U26899 ( .A(n12915), .B(n24894), .Z(n24896) );
  XOR U26900 ( .A(n24898), .B(n24899), .Z(n12915) );
  XOR U26901 ( .A(n24900), .B(n24901), .Z(n24894) );
  AND U26902 ( .A(n24902), .B(n24903), .Z(n24901) );
  XOR U26903 ( .A(nreg[973]), .B(n24900), .Z(n24903) );
  XNOR U26904 ( .A(n12927), .B(n24900), .Z(n24902) );
  XOR U26905 ( .A(n24904), .B(n24905), .Z(n12927) );
  XOR U26906 ( .A(n24906), .B(n24907), .Z(n24900) );
  AND U26907 ( .A(n24908), .B(n24909), .Z(n24907) );
  XOR U26908 ( .A(nreg[972]), .B(n24906), .Z(n24909) );
  XNOR U26909 ( .A(n12939), .B(n24906), .Z(n24908) );
  XOR U26910 ( .A(n24910), .B(n24911), .Z(n12939) );
  XOR U26911 ( .A(n24912), .B(n24913), .Z(n24906) );
  AND U26912 ( .A(n24914), .B(n24915), .Z(n24913) );
  XOR U26913 ( .A(nreg[971]), .B(n24912), .Z(n24915) );
  XNOR U26914 ( .A(n12951), .B(n24912), .Z(n24914) );
  XOR U26915 ( .A(n24916), .B(n24917), .Z(n12951) );
  XOR U26916 ( .A(n24918), .B(n24919), .Z(n24912) );
  AND U26917 ( .A(n24920), .B(n24921), .Z(n24919) );
  XOR U26918 ( .A(nreg[970]), .B(n24918), .Z(n24921) );
  XNOR U26919 ( .A(n12963), .B(n24918), .Z(n24920) );
  XOR U26920 ( .A(n24922), .B(n24923), .Z(n12963) );
  XOR U26921 ( .A(n24924), .B(n24925), .Z(n24918) );
  AND U26922 ( .A(n24926), .B(n24927), .Z(n24925) );
  XOR U26923 ( .A(nreg[969]), .B(n24924), .Z(n24927) );
  XNOR U26924 ( .A(n12975), .B(n24924), .Z(n24926) );
  XOR U26925 ( .A(n24928), .B(n24929), .Z(n12975) );
  XOR U26926 ( .A(n24930), .B(n24931), .Z(n24924) );
  AND U26927 ( .A(n24932), .B(n24933), .Z(n24931) );
  XOR U26928 ( .A(nreg[968]), .B(n24930), .Z(n24933) );
  XNOR U26929 ( .A(n12987), .B(n24930), .Z(n24932) );
  XOR U26930 ( .A(n24934), .B(n24935), .Z(n12987) );
  XOR U26931 ( .A(n24936), .B(n24937), .Z(n24930) );
  AND U26932 ( .A(n24938), .B(n24939), .Z(n24937) );
  XOR U26933 ( .A(nreg[967]), .B(n24936), .Z(n24939) );
  XNOR U26934 ( .A(n12999), .B(n24936), .Z(n24938) );
  XOR U26935 ( .A(n24940), .B(n24941), .Z(n12999) );
  XOR U26936 ( .A(n24942), .B(n24943), .Z(n24936) );
  AND U26937 ( .A(n24944), .B(n24945), .Z(n24943) );
  XOR U26938 ( .A(nreg[966]), .B(n24942), .Z(n24945) );
  XNOR U26939 ( .A(n13011), .B(n24942), .Z(n24944) );
  XOR U26940 ( .A(n24946), .B(n24947), .Z(n13011) );
  XOR U26941 ( .A(n24948), .B(n24949), .Z(n24942) );
  AND U26942 ( .A(n24950), .B(n24951), .Z(n24949) );
  XOR U26943 ( .A(nreg[965]), .B(n24948), .Z(n24951) );
  XNOR U26944 ( .A(n13023), .B(n24948), .Z(n24950) );
  XOR U26945 ( .A(n24952), .B(n24953), .Z(n13023) );
  XOR U26946 ( .A(n24954), .B(n24955), .Z(n24948) );
  AND U26947 ( .A(n24956), .B(n24957), .Z(n24955) );
  XOR U26948 ( .A(nreg[964]), .B(n24954), .Z(n24957) );
  XNOR U26949 ( .A(n13035), .B(n24954), .Z(n24956) );
  XOR U26950 ( .A(n24958), .B(n24959), .Z(n13035) );
  XOR U26951 ( .A(n24960), .B(n24961), .Z(n24954) );
  AND U26952 ( .A(n24962), .B(n24963), .Z(n24961) );
  XOR U26953 ( .A(nreg[963]), .B(n24960), .Z(n24963) );
  XNOR U26954 ( .A(n13047), .B(n24960), .Z(n24962) );
  XOR U26955 ( .A(n24964), .B(n24965), .Z(n13047) );
  XOR U26956 ( .A(n24966), .B(n24967), .Z(n24960) );
  AND U26957 ( .A(n24968), .B(n24969), .Z(n24967) );
  XOR U26958 ( .A(nreg[962]), .B(n24966), .Z(n24969) );
  XNOR U26959 ( .A(n13059), .B(n24966), .Z(n24968) );
  XOR U26960 ( .A(n24970), .B(n24971), .Z(n13059) );
  XOR U26961 ( .A(n24972), .B(n24973), .Z(n24966) );
  AND U26962 ( .A(n24974), .B(n24975), .Z(n24973) );
  XOR U26963 ( .A(nreg[961]), .B(n24972), .Z(n24975) );
  XNOR U26964 ( .A(n13071), .B(n24972), .Z(n24974) );
  XOR U26965 ( .A(n24976), .B(n24977), .Z(n13071) );
  XOR U26966 ( .A(n24978), .B(n24979), .Z(n24972) );
  AND U26967 ( .A(n24980), .B(n24981), .Z(n24979) );
  XOR U26968 ( .A(nreg[960]), .B(n24978), .Z(n24981) );
  XNOR U26969 ( .A(n13083), .B(n24978), .Z(n24980) );
  XOR U26970 ( .A(n24982), .B(n24983), .Z(n13083) );
  XOR U26971 ( .A(n24984), .B(n24985), .Z(n24978) );
  AND U26972 ( .A(n24986), .B(n24987), .Z(n24985) );
  XOR U26973 ( .A(nreg[959]), .B(n24984), .Z(n24987) );
  XNOR U26974 ( .A(n13095), .B(n24984), .Z(n24986) );
  XOR U26975 ( .A(n24988), .B(n24989), .Z(n13095) );
  XOR U26976 ( .A(n24990), .B(n24991), .Z(n24984) );
  AND U26977 ( .A(n24992), .B(n24993), .Z(n24991) );
  XOR U26978 ( .A(nreg[958]), .B(n24990), .Z(n24993) );
  XNOR U26979 ( .A(n13107), .B(n24990), .Z(n24992) );
  XOR U26980 ( .A(n24994), .B(n24995), .Z(n13107) );
  XOR U26981 ( .A(n24996), .B(n24997), .Z(n24990) );
  AND U26982 ( .A(n24998), .B(n24999), .Z(n24997) );
  XOR U26983 ( .A(nreg[957]), .B(n24996), .Z(n24999) );
  XNOR U26984 ( .A(n13119), .B(n24996), .Z(n24998) );
  XOR U26985 ( .A(n25000), .B(n25001), .Z(n13119) );
  XOR U26986 ( .A(n25002), .B(n25003), .Z(n24996) );
  AND U26987 ( .A(n25004), .B(n25005), .Z(n25003) );
  XOR U26988 ( .A(nreg[956]), .B(n25002), .Z(n25005) );
  XNOR U26989 ( .A(n13131), .B(n25002), .Z(n25004) );
  XOR U26990 ( .A(n25006), .B(n25007), .Z(n13131) );
  XOR U26991 ( .A(n25008), .B(n25009), .Z(n25002) );
  AND U26992 ( .A(n25010), .B(n25011), .Z(n25009) );
  XOR U26993 ( .A(nreg[955]), .B(n25008), .Z(n25011) );
  XNOR U26994 ( .A(n13143), .B(n25008), .Z(n25010) );
  XOR U26995 ( .A(n25012), .B(n25013), .Z(n13143) );
  XOR U26996 ( .A(n25014), .B(n25015), .Z(n25008) );
  AND U26997 ( .A(n25016), .B(n25017), .Z(n25015) );
  XOR U26998 ( .A(nreg[954]), .B(n25014), .Z(n25017) );
  XNOR U26999 ( .A(n13155), .B(n25014), .Z(n25016) );
  XOR U27000 ( .A(n25018), .B(n25019), .Z(n13155) );
  XOR U27001 ( .A(n25020), .B(n25021), .Z(n25014) );
  AND U27002 ( .A(n25022), .B(n25023), .Z(n25021) );
  XOR U27003 ( .A(nreg[953]), .B(n25020), .Z(n25023) );
  XNOR U27004 ( .A(n13167), .B(n25020), .Z(n25022) );
  XOR U27005 ( .A(n25024), .B(n25025), .Z(n13167) );
  XOR U27006 ( .A(n25026), .B(n25027), .Z(n25020) );
  AND U27007 ( .A(n25028), .B(n25029), .Z(n25027) );
  XOR U27008 ( .A(nreg[952]), .B(n25026), .Z(n25029) );
  XNOR U27009 ( .A(n13179), .B(n25026), .Z(n25028) );
  XOR U27010 ( .A(n25030), .B(n25031), .Z(n13179) );
  XOR U27011 ( .A(n25032), .B(n25033), .Z(n25026) );
  AND U27012 ( .A(n25034), .B(n25035), .Z(n25033) );
  XOR U27013 ( .A(nreg[951]), .B(n25032), .Z(n25035) );
  XNOR U27014 ( .A(n13191), .B(n25032), .Z(n25034) );
  XOR U27015 ( .A(n25036), .B(n25037), .Z(n13191) );
  XOR U27016 ( .A(n25038), .B(n25039), .Z(n25032) );
  AND U27017 ( .A(n25040), .B(n25041), .Z(n25039) );
  XOR U27018 ( .A(nreg[950]), .B(n25038), .Z(n25041) );
  XNOR U27019 ( .A(n13203), .B(n25038), .Z(n25040) );
  XOR U27020 ( .A(n25042), .B(n25043), .Z(n13203) );
  XOR U27021 ( .A(n25044), .B(n25045), .Z(n25038) );
  AND U27022 ( .A(n25046), .B(n25047), .Z(n25045) );
  XOR U27023 ( .A(nreg[949]), .B(n25044), .Z(n25047) );
  XNOR U27024 ( .A(n13215), .B(n25044), .Z(n25046) );
  XOR U27025 ( .A(n25048), .B(n25049), .Z(n13215) );
  XOR U27026 ( .A(n25050), .B(n25051), .Z(n25044) );
  AND U27027 ( .A(n25052), .B(n25053), .Z(n25051) );
  XOR U27028 ( .A(nreg[948]), .B(n25050), .Z(n25053) );
  XNOR U27029 ( .A(n13227), .B(n25050), .Z(n25052) );
  XOR U27030 ( .A(n25054), .B(n25055), .Z(n13227) );
  XOR U27031 ( .A(n25056), .B(n25057), .Z(n25050) );
  AND U27032 ( .A(n25058), .B(n25059), .Z(n25057) );
  XOR U27033 ( .A(nreg[947]), .B(n25056), .Z(n25059) );
  XNOR U27034 ( .A(n13239), .B(n25056), .Z(n25058) );
  XOR U27035 ( .A(n25060), .B(n25061), .Z(n13239) );
  XOR U27036 ( .A(n25062), .B(n25063), .Z(n25056) );
  AND U27037 ( .A(n25064), .B(n25065), .Z(n25063) );
  XOR U27038 ( .A(nreg[946]), .B(n25062), .Z(n25065) );
  XNOR U27039 ( .A(n13251), .B(n25062), .Z(n25064) );
  XOR U27040 ( .A(n25066), .B(n25067), .Z(n13251) );
  XOR U27041 ( .A(n25068), .B(n25069), .Z(n25062) );
  AND U27042 ( .A(n25070), .B(n25071), .Z(n25069) );
  XOR U27043 ( .A(nreg[945]), .B(n25068), .Z(n25071) );
  XNOR U27044 ( .A(n13263), .B(n25068), .Z(n25070) );
  XOR U27045 ( .A(n25072), .B(n25073), .Z(n13263) );
  XOR U27046 ( .A(n25074), .B(n25075), .Z(n25068) );
  AND U27047 ( .A(n25076), .B(n25077), .Z(n25075) );
  XOR U27048 ( .A(nreg[944]), .B(n25074), .Z(n25077) );
  XNOR U27049 ( .A(n13275), .B(n25074), .Z(n25076) );
  XOR U27050 ( .A(n25078), .B(n25079), .Z(n13275) );
  XOR U27051 ( .A(n25080), .B(n25081), .Z(n25074) );
  AND U27052 ( .A(n25082), .B(n25083), .Z(n25081) );
  XOR U27053 ( .A(nreg[943]), .B(n25080), .Z(n25083) );
  XNOR U27054 ( .A(n13287), .B(n25080), .Z(n25082) );
  XOR U27055 ( .A(n25084), .B(n25085), .Z(n13287) );
  XOR U27056 ( .A(n25086), .B(n25087), .Z(n25080) );
  AND U27057 ( .A(n25088), .B(n25089), .Z(n25087) );
  XOR U27058 ( .A(nreg[942]), .B(n25086), .Z(n25089) );
  XNOR U27059 ( .A(n13299), .B(n25086), .Z(n25088) );
  XOR U27060 ( .A(n25090), .B(n25091), .Z(n13299) );
  XOR U27061 ( .A(n25092), .B(n25093), .Z(n25086) );
  AND U27062 ( .A(n25094), .B(n25095), .Z(n25093) );
  XOR U27063 ( .A(nreg[941]), .B(n25092), .Z(n25095) );
  XNOR U27064 ( .A(n13311), .B(n25092), .Z(n25094) );
  XOR U27065 ( .A(n25096), .B(n25097), .Z(n13311) );
  XOR U27066 ( .A(n25098), .B(n25099), .Z(n25092) );
  AND U27067 ( .A(n25100), .B(n25101), .Z(n25099) );
  XOR U27068 ( .A(nreg[940]), .B(n25098), .Z(n25101) );
  XNOR U27069 ( .A(n13323), .B(n25098), .Z(n25100) );
  XOR U27070 ( .A(n25102), .B(n25103), .Z(n13323) );
  XOR U27071 ( .A(n25104), .B(n25105), .Z(n25098) );
  AND U27072 ( .A(n25106), .B(n25107), .Z(n25105) );
  XOR U27073 ( .A(nreg[939]), .B(n25104), .Z(n25107) );
  XNOR U27074 ( .A(n13335), .B(n25104), .Z(n25106) );
  XOR U27075 ( .A(n25108), .B(n25109), .Z(n13335) );
  XOR U27076 ( .A(n25110), .B(n25111), .Z(n25104) );
  AND U27077 ( .A(n25112), .B(n25113), .Z(n25111) );
  XOR U27078 ( .A(nreg[938]), .B(n25110), .Z(n25113) );
  XNOR U27079 ( .A(n13347), .B(n25110), .Z(n25112) );
  XOR U27080 ( .A(n25114), .B(n25115), .Z(n13347) );
  XOR U27081 ( .A(n25116), .B(n25117), .Z(n25110) );
  AND U27082 ( .A(n25118), .B(n25119), .Z(n25117) );
  XOR U27083 ( .A(nreg[937]), .B(n25116), .Z(n25119) );
  XNOR U27084 ( .A(n13359), .B(n25116), .Z(n25118) );
  XOR U27085 ( .A(n25120), .B(n25121), .Z(n13359) );
  XOR U27086 ( .A(n25122), .B(n25123), .Z(n25116) );
  AND U27087 ( .A(n25124), .B(n25125), .Z(n25123) );
  XOR U27088 ( .A(nreg[936]), .B(n25122), .Z(n25125) );
  XNOR U27089 ( .A(n13371), .B(n25122), .Z(n25124) );
  XOR U27090 ( .A(n25126), .B(n25127), .Z(n13371) );
  XOR U27091 ( .A(n25128), .B(n25129), .Z(n25122) );
  AND U27092 ( .A(n25130), .B(n25131), .Z(n25129) );
  XOR U27093 ( .A(nreg[935]), .B(n25128), .Z(n25131) );
  XNOR U27094 ( .A(n13383), .B(n25128), .Z(n25130) );
  XOR U27095 ( .A(n25132), .B(n25133), .Z(n13383) );
  XOR U27096 ( .A(n25134), .B(n25135), .Z(n25128) );
  AND U27097 ( .A(n25136), .B(n25137), .Z(n25135) );
  XOR U27098 ( .A(nreg[934]), .B(n25134), .Z(n25137) );
  XNOR U27099 ( .A(n13395), .B(n25134), .Z(n25136) );
  XOR U27100 ( .A(n25138), .B(n25139), .Z(n13395) );
  XOR U27101 ( .A(n25140), .B(n25141), .Z(n25134) );
  AND U27102 ( .A(n25142), .B(n25143), .Z(n25141) );
  XOR U27103 ( .A(nreg[933]), .B(n25140), .Z(n25143) );
  XNOR U27104 ( .A(n13407), .B(n25140), .Z(n25142) );
  XOR U27105 ( .A(n25144), .B(n25145), .Z(n13407) );
  XOR U27106 ( .A(n25146), .B(n25147), .Z(n25140) );
  AND U27107 ( .A(n25148), .B(n25149), .Z(n25147) );
  XOR U27108 ( .A(nreg[932]), .B(n25146), .Z(n25149) );
  XNOR U27109 ( .A(n13419), .B(n25146), .Z(n25148) );
  XOR U27110 ( .A(n25150), .B(n25151), .Z(n13419) );
  XOR U27111 ( .A(n25152), .B(n25153), .Z(n25146) );
  AND U27112 ( .A(n25154), .B(n25155), .Z(n25153) );
  XOR U27113 ( .A(nreg[931]), .B(n25152), .Z(n25155) );
  XNOR U27114 ( .A(n13431), .B(n25152), .Z(n25154) );
  XOR U27115 ( .A(n25156), .B(n25157), .Z(n13431) );
  XOR U27116 ( .A(n25158), .B(n25159), .Z(n25152) );
  AND U27117 ( .A(n25160), .B(n25161), .Z(n25159) );
  XOR U27118 ( .A(nreg[930]), .B(n25158), .Z(n25161) );
  XNOR U27119 ( .A(n13443), .B(n25158), .Z(n25160) );
  XOR U27120 ( .A(n25162), .B(n25163), .Z(n13443) );
  XOR U27121 ( .A(n25164), .B(n25165), .Z(n25158) );
  AND U27122 ( .A(n25166), .B(n25167), .Z(n25165) );
  XOR U27123 ( .A(nreg[929]), .B(n25164), .Z(n25167) );
  XNOR U27124 ( .A(n13455), .B(n25164), .Z(n25166) );
  XOR U27125 ( .A(n25168), .B(n25169), .Z(n13455) );
  XOR U27126 ( .A(n25170), .B(n25171), .Z(n25164) );
  AND U27127 ( .A(n25172), .B(n25173), .Z(n25171) );
  XOR U27128 ( .A(nreg[928]), .B(n25170), .Z(n25173) );
  XNOR U27129 ( .A(n13467), .B(n25170), .Z(n25172) );
  XOR U27130 ( .A(n25174), .B(n25175), .Z(n13467) );
  XOR U27131 ( .A(n25176), .B(n25177), .Z(n25170) );
  AND U27132 ( .A(n25178), .B(n25179), .Z(n25177) );
  XOR U27133 ( .A(nreg[927]), .B(n25176), .Z(n25179) );
  XNOR U27134 ( .A(n13479), .B(n25176), .Z(n25178) );
  XOR U27135 ( .A(n25180), .B(n25181), .Z(n13479) );
  XOR U27136 ( .A(n25182), .B(n25183), .Z(n25176) );
  AND U27137 ( .A(n25184), .B(n25185), .Z(n25183) );
  XOR U27138 ( .A(nreg[926]), .B(n25182), .Z(n25185) );
  XNOR U27139 ( .A(n13491), .B(n25182), .Z(n25184) );
  XOR U27140 ( .A(n25186), .B(n25187), .Z(n13491) );
  XOR U27141 ( .A(n25188), .B(n25189), .Z(n25182) );
  AND U27142 ( .A(n25190), .B(n25191), .Z(n25189) );
  XOR U27143 ( .A(nreg[925]), .B(n25188), .Z(n25191) );
  XNOR U27144 ( .A(n13503), .B(n25188), .Z(n25190) );
  XOR U27145 ( .A(n25192), .B(n25193), .Z(n13503) );
  XOR U27146 ( .A(n25194), .B(n25195), .Z(n25188) );
  AND U27147 ( .A(n25196), .B(n25197), .Z(n25195) );
  XOR U27148 ( .A(nreg[924]), .B(n25194), .Z(n25197) );
  XNOR U27149 ( .A(n13515), .B(n25194), .Z(n25196) );
  XOR U27150 ( .A(n25198), .B(n25199), .Z(n13515) );
  XOR U27151 ( .A(n25200), .B(n25201), .Z(n25194) );
  AND U27152 ( .A(n25202), .B(n25203), .Z(n25201) );
  XOR U27153 ( .A(nreg[923]), .B(n25200), .Z(n25203) );
  XNOR U27154 ( .A(n13527), .B(n25200), .Z(n25202) );
  XOR U27155 ( .A(n25204), .B(n25205), .Z(n13527) );
  XOR U27156 ( .A(n25206), .B(n25207), .Z(n25200) );
  AND U27157 ( .A(n25208), .B(n25209), .Z(n25207) );
  XOR U27158 ( .A(nreg[922]), .B(n25206), .Z(n25209) );
  XNOR U27159 ( .A(n13539), .B(n25206), .Z(n25208) );
  XOR U27160 ( .A(n25210), .B(n25211), .Z(n13539) );
  XOR U27161 ( .A(n25212), .B(n25213), .Z(n25206) );
  AND U27162 ( .A(n25214), .B(n25215), .Z(n25213) );
  XOR U27163 ( .A(nreg[921]), .B(n25212), .Z(n25215) );
  XNOR U27164 ( .A(n13551), .B(n25212), .Z(n25214) );
  XOR U27165 ( .A(n25216), .B(n25217), .Z(n13551) );
  XOR U27166 ( .A(n25218), .B(n25219), .Z(n25212) );
  AND U27167 ( .A(n25220), .B(n25221), .Z(n25219) );
  XOR U27168 ( .A(nreg[920]), .B(n25218), .Z(n25221) );
  XNOR U27169 ( .A(n13563), .B(n25218), .Z(n25220) );
  XOR U27170 ( .A(n25222), .B(n25223), .Z(n13563) );
  XOR U27171 ( .A(n25224), .B(n25225), .Z(n25218) );
  AND U27172 ( .A(n25226), .B(n25227), .Z(n25225) );
  XOR U27173 ( .A(nreg[919]), .B(n25224), .Z(n25227) );
  XNOR U27174 ( .A(n13575), .B(n25224), .Z(n25226) );
  XOR U27175 ( .A(n25228), .B(n25229), .Z(n13575) );
  XOR U27176 ( .A(n25230), .B(n25231), .Z(n25224) );
  AND U27177 ( .A(n25232), .B(n25233), .Z(n25231) );
  XOR U27178 ( .A(nreg[918]), .B(n25230), .Z(n25233) );
  XNOR U27179 ( .A(n13587), .B(n25230), .Z(n25232) );
  XOR U27180 ( .A(n25234), .B(n25235), .Z(n13587) );
  XOR U27181 ( .A(n25236), .B(n25237), .Z(n25230) );
  AND U27182 ( .A(n25238), .B(n25239), .Z(n25237) );
  XOR U27183 ( .A(nreg[917]), .B(n25236), .Z(n25239) );
  XNOR U27184 ( .A(n13599), .B(n25236), .Z(n25238) );
  XOR U27185 ( .A(n25240), .B(n25241), .Z(n13599) );
  XOR U27186 ( .A(n25242), .B(n25243), .Z(n25236) );
  AND U27187 ( .A(n25244), .B(n25245), .Z(n25243) );
  XOR U27188 ( .A(nreg[916]), .B(n25242), .Z(n25245) );
  XNOR U27189 ( .A(n13611), .B(n25242), .Z(n25244) );
  XOR U27190 ( .A(n25246), .B(n25247), .Z(n13611) );
  XOR U27191 ( .A(n25248), .B(n25249), .Z(n25242) );
  AND U27192 ( .A(n25250), .B(n25251), .Z(n25249) );
  XOR U27193 ( .A(nreg[915]), .B(n25248), .Z(n25251) );
  XNOR U27194 ( .A(n13623), .B(n25248), .Z(n25250) );
  XOR U27195 ( .A(n25252), .B(n25253), .Z(n13623) );
  XOR U27196 ( .A(n25254), .B(n25255), .Z(n25248) );
  AND U27197 ( .A(n25256), .B(n25257), .Z(n25255) );
  XOR U27198 ( .A(nreg[914]), .B(n25254), .Z(n25257) );
  XNOR U27199 ( .A(n13635), .B(n25254), .Z(n25256) );
  XOR U27200 ( .A(n25258), .B(n25259), .Z(n13635) );
  XOR U27201 ( .A(n25260), .B(n25261), .Z(n25254) );
  AND U27202 ( .A(n25262), .B(n25263), .Z(n25261) );
  XOR U27203 ( .A(nreg[913]), .B(n25260), .Z(n25263) );
  XNOR U27204 ( .A(n13647), .B(n25260), .Z(n25262) );
  XOR U27205 ( .A(n25264), .B(n25265), .Z(n13647) );
  XOR U27206 ( .A(n25266), .B(n25267), .Z(n25260) );
  AND U27207 ( .A(n25268), .B(n25269), .Z(n25267) );
  XOR U27208 ( .A(nreg[912]), .B(n25266), .Z(n25269) );
  XNOR U27209 ( .A(n13659), .B(n25266), .Z(n25268) );
  XOR U27210 ( .A(n25270), .B(n25271), .Z(n13659) );
  XOR U27211 ( .A(n25272), .B(n25273), .Z(n25266) );
  AND U27212 ( .A(n25274), .B(n25275), .Z(n25273) );
  XOR U27213 ( .A(nreg[911]), .B(n25272), .Z(n25275) );
  XNOR U27214 ( .A(n13671), .B(n25272), .Z(n25274) );
  XOR U27215 ( .A(n25276), .B(n25277), .Z(n13671) );
  XOR U27216 ( .A(n25278), .B(n25279), .Z(n25272) );
  AND U27217 ( .A(n25280), .B(n25281), .Z(n25279) );
  XOR U27218 ( .A(nreg[910]), .B(n25278), .Z(n25281) );
  XNOR U27219 ( .A(n13683), .B(n25278), .Z(n25280) );
  XOR U27220 ( .A(n25282), .B(n25283), .Z(n13683) );
  XOR U27221 ( .A(n25284), .B(n25285), .Z(n25278) );
  AND U27222 ( .A(n25286), .B(n25287), .Z(n25285) );
  XOR U27223 ( .A(nreg[909]), .B(n25284), .Z(n25287) );
  XNOR U27224 ( .A(n13695), .B(n25284), .Z(n25286) );
  XOR U27225 ( .A(n25288), .B(n25289), .Z(n13695) );
  XOR U27226 ( .A(n25290), .B(n25291), .Z(n25284) );
  AND U27227 ( .A(n25292), .B(n25293), .Z(n25291) );
  XOR U27228 ( .A(nreg[908]), .B(n25290), .Z(n25293) );
  XNOR U27229 ( .A(n13707), .B(n25290), .Z(n25292) );
  XOR U27230 ( .A(n25294), .B(n25295), .Z(n13707) );
  XOR U27231 ( .A(n25296), .B(n25297), .Z(n25290) );
  AND U27232 ( .A(n25298), .B(n25299), .Z(n25297) );
  XOR U27233 ( .A(nreg[907]), .B(n25296), .Z(n25299) );
  XNOR U27234 ( .A(n13719), .B(n25296), .Z(n25298) );
  XOR U27235 ( .A(n25300), .B(n25301), .Z(n13719) );
  XOR U27236 ( .A(n25302), .B(n25303), .Z(n25296) );
  AND U27237 ( .A(n25304), .B(n25305), .Z(n25303) );
  XOR U27238 ( .A(nreg[906]), .B(n25302), .Z(n25305) );
  XNOR U27239 ( .A(n13731), .B(n25302), .Z(n25304) );
  XOR U27240 ( .A(n25306), .B(n25307), .Z(n13731) );
  XOR U27241 ( .A(n25308), .B(n25309), .Z(n25302) );
  AND U27242 ( .A(n25310), .B(n25311), .Z(n25309) );
  XOR U27243 ( .A(nreg[905]), .B(n25308), .Z(n25311) );
  XNOR U27244 ( .A(n13743), .B(n25308), .Z(n25310) );
  XOR U27245 ( .A(n25312), .B(n25313), .Z(n13743) );
  XOR U27246 ( .A(n25314), .B(n25315), .Z(n25308) );
  AND U27247 ( .A(n25316), .B(n25317), .Z(n25315) );
  XOR U27248 ( .A(nreg[904]), .B(n25314), .Z(n25317) );
  XNOR U27249 ( .A(n13755), .B(n25314), .Z(n25316) );
  XOR U27250 ( .A(n25318), .B(n25319), .Z(n13755) );
  XOR U27251 ( .A(n25320), .B(n25321), .Z(n25314) );
  AND U27252 ( .A(n25322), .B(n25323), .Z(n25321) );
  XOR U27253 ( .A(nreg[903]), .B(n25320), .Z(n25323) );
  XNOR U27254 ( .A(n13767), .B(n25320), .Z(n25322) );
  XOR U27255 ( .A(n25324), .B(n25325), .Z(n13767) );
  XOR U27256 ( .A(n25326), .B(n25327), .Z(n25320) );
  AND U27257 ( .A(n25328), .B(n25329), .Z(n25327) );
  XOR U27258 ( .A(nreg[902]), .B(n25326), .Z(n25329) );
  XNOR U27259 ( .A(n13779), .B(n25326), .Z(n25328) );
  XOR U27260 ( .A(n25330), .B(n25331), .Z(n13779) );
  XOR U27261 ( .A(n25332), .B(n25333), .Z(n25326) );
  AND U27262 ( .A(n25334), .B(n25335), .Z(n25333) );
  XOR U27263 ( .A(nreg[901]), .B(n25332), .Z(n25335) );
  XNOR U27264 ( .A(n13791), .B(n25332), .Z(n25334) );
  XOR U27265 ( .A(n25336), .B(n25337), .Z(n13791) );
  XOR U27266 ( .A(n25338), .B(n25339), .Z(n25332) );
  AND U27267 ( .A(n25340), .B(n25341), .Z(n25339) );
  XOR U27268 ( .A(nreg[900]), .B(n25338), .Z(n25341) );
  XNOR U27269 ( .A(n13803), .B(n25338), .Z(n25340) );
  XOR U27270 ( .A(n25342), .B(n25343), .Z(n13803) );
  XOR U27271 ( .A(n25344), .B(n25345), .Z(n25338) );
  AND U27272 ( .A(n25346), .B(n25347), .Z(n25345) );
  XOR U27273 ( .A(nreg[899]), .B(n25344), .Z(n25347) );
  XNOR U27274 ( .A(n13815), .B(n25344), .Z(n25346) );
  XOR U27275 ( .A(n25348), .B(n25349), .Z(n13815) );
  XOR U27276 ( .A(n25350), .B(n25351), .Z(n25344) );
  AND U27277 ( .A(n25352), .B(n25353), .Z(n25351) );
  XOR U27278 ( .A(nreg[898]), .B(n25350), .Z(n25353) );
  XNOR U27279 ( .A(n13827), .B(n25350), .Z(n25352) );
  XOR U27280 ( .A(n25354), .B(n25355), .Z(n13827) );
  XOR U27281 ( .A(n25356), .B(n25357), .Z(n25350) );
  AND U27282 ( .A(n25358), .B(n25359), .Z(n25357) );
  XOR U27283 ( .A(nreg[897]), .B(n25356), .Z(n25359) );
  XNOR U27284 ( .A(n13839), .B(n25356), .Z(n25358) );
  XOR U27285 ( .A(n25360), .B(n25361), .Z(n13839) );
  XOR U27286 ( .A(n25362), .B(n25363), .Z(n25356) );
  AND U27287 ( .A(n25364), .B(n25365), .Z(n25363) );
  XOR U27288 ( .A(nreg[896]), .B(n25362), .Z(n25365) );
  XNOR U27289 ( .A(n13851), .B(n25362), .Z(n25364) );
  XOR U27290 ( .A(n25366), .B(n25367), .Z(n13851) );
  XOR U27291 ( .A(n25368), .B(n25369), .Z(n25362) );
  AND U27292 ( .A(n25370), .B(n25371), .Z(n25369) );
  XOR U27293 ( .A(nreg[895]), .B(n25368), .Z(n25371) );
  XNOR U27294 ( .A(n13863), .B(n25368), .Z(n25370) );
  XOR U27295 ( .A(n25372), .B(n25373), .Z(n13863) );
  XOR U27296 ( .A(n25374), .B(n25375), .Z(n25368) );
  AND U27297 ( .A(n25376), .B(n25377), .Z(n25375) );
  XOR U27298 ( .A(nreg[894]), .B(n25374), .Z(n25377) );
  XNOR U27299 ( .A(n13875), .B(n25374), .Z(n25376) );
  XOR U27300 ( .A(n25378), .B(n25379), .Z(n13875) );
  XOR U27301 ( .A(n25380), .B(n25381), .Z(n25374) );
  AND U27302 ( .A(n25382), .B(n25383), .Z(n25381) );
  XOR U27303 ( .A(nreg[893]), .B(n25380), .Z(n25383) );
  XNOR U27304 ( .A(n13887), .B(n25380), .Z(n25382) );
  XOR U27305 ( .A(n25384), .B(n25385), .Z(n13887) );
  XOR U27306 ( .A(n25386), .B(n25387), .Z(n25380) );
  AND U27307 ( .A(n25388), .B(n25389), .Z(n25387) );
  XOR U27308 ( .A(nreg[892]), .B(n25386), .Z(n25389) );
  XNOR U27309 ( .A(n13899), .B(n25386), .Z(n25388) );
  XOR U27310 ( .A(n25390), .B(n25391), .Z(n13899) );
  XOR U27311 ( .A(n25392), .B(n25393), .Z(n25386) );
  AND U27312 ( .A(n25394), .B(n25395), .Z(n25393) );
  XOR U27313 ( .A(nreg[891]), .B(n25392), .Z(n25395) );
  XNOR U27314 ( .A(n13911), .B(n25392), .Z(n25394) );
  XOR U27315 ( .A(n25396), .B(n25397), .Z(n13911) );
  XOR U27316 ( .A(n25398), .B(n25399), .Z(n25392) );
  AND U27317 ( .A(n25400), .B(n25401), .Z(n25399) );
  XOR U27318 ( .A(nreg[890]), .B(n25398), .Z(n25401) );
  XNOR U27319 ( .A(n13923), .B(n25398), .Z(n25400) );
  XOR U27320 ( .A(n25402), .B(n25403), .Z(n13923) );
  XOR U27321 ( .A(n25404), .B(n25405), .Z(n25398) );
  AND U27322 ( .A(n25406), .B(n25407), .Z(n25405) );
  XOR U27323 ( .A(nreg[889]), .B(n25404), .Z(n25407) );
  XNOR U27324 ( .A(n13935), .B(n25404), .Z(n25406) );
  XOR U27325 ( .A(n25408), .B(n25409), .Z(n13935) );
  XOR U27326 ( .A(n25410), .B(n25411), .Z(n25404) );
  AND U27327 ( .A(n25412), .B(n25413), .Z(n25411) );
  XOR U27328 ( .A(nreg[888]), .B(n25410), .Z(n25413) );
  XNOR U27329 ( .A(n13947), .B(n25410), .Z(n25412) );
  XOR U27330 ( .A(n25414), .B(n25415), .Z(n13947) );
  XOR U27331 ( .A(n25416), .B(n25417), .Z(n25410) );
  AND U27332 ( .A(n25418), .B(n25419), .Z(n25417) );
  XOR U27333 ( .A(nreg[887]), .B(n25416), .Z(n25419) );
  XNOR U27334 ( .A(n13959), .B(n25416), .Z(n25418) );
  XOR U27335 ( .A(n25420), .B(n25421), .Z(n13959) );
  XOR U27336 ( .A(n25422), .B(n25423), .Z(n25416) );
  AND U27337 ( .A(n25424), .B(n25425), .Z(n25423) );
  XOR U27338 ( .A(nreg[886]), .B(n25422), .Z(n25425) );
  XNOR U27339 ( .A(n13971), .B(n25422), .Z(n25424) );
  XOR U27340 ( .A(n25426), .B(n25427), .Z(n13971) );
  XOR U27341 ( .A(n25428), .B(n25429), .Z(n25422) );
  AND U27342 ( .A(n25430), .B(n25431), .Z(n25429) );
  XOR U27343 ( .A(nreg[885]), .B(n25428), .Z(n25431) );
  XNOR U27344 ( .A(n13983), .B(n25428), .Z(n25430) );
  XOR U27345 ( .A(n25432), .B(n25433), .Z(n13983) );
  XOR U27346 ( .A(n25434), .B(n25435), .Z(n25428) );
  AND U27347 ( .A(n25436), .B(n25437), .Z(n25435) );
  XOR U27348 ( .A(nreg[884]), .B(n25434), .Z(n25437) );
  XNOR U27349 ( .A(n13995), .B(n25434), .Z(n25436) );
  XOR U27350 ( .A(n25438), .B(n25439), .Z(n13995) );
  XOR U27351 ( .A(n25440), .B(n25441), .Z(n25434) );
  AND U27352 ( .A(n25442), .B(n25443), .Z(n25441) );
  XOR U27353 ( .A(nreg[883]), .B(n25440), .Z(n25443) );
  XNOR U27354 ( .A(n14007), .B(n25440), .Z(n25442) );
  XOR U27355 ( .A(n25444), .B(n25445), .Z(n14007) );
  XOR U27356 ( .A(n25446), .B(n25447), .Z(n25440) );
  AND U27357 ( .A(n25448), .B(n25449), .Z(n25447) );
  XOR U27358 ( .A(nreg[882]), .B(n25446), .Z(n25449) );
  XNOR U27359 ( .A(n14019), .B(n25446), .Z(n25448) );
  XOR U27360 ( .A(n25450), .B(n25451), .Z(n14019) );
  XOR U27361 ( .A(n25452), .B(n25453), .Z(n25446) );
  AND U27362 ( .A(n25454), .B(n25455), .Z(n25453) );
  XOR U27363 ( .A(nreg[881]), .B(n25452), .Z(n25455) );
  XNOR U27364 ( .A(n14031), .B(n25452), .Z(n25454) );
  XOR U27365 ( .A(n25456), .B(n25457), .Z(n14031) );
  XOR U27366 ( .A(n25458), .B(n25459), .Z(n25452) );
  AND U27367 ( .A(n25460), .B(n25461), .Z(n25459) );
  XOR U27368 ( .A(nreg[880]), .B(n25458), .Z(n25461) );
  XNOR U27369 ( .A(n14043), .B(n25458), .Z(n25460) );
  XOR U27370 ( .A(n25462), .B(n25463), .Z(n14043) );
  XOR U27371 ( .A(n25464), .B(n25465), .Z(n25458) );
  AND U27372 ( .A(n25466), .B(n25467), .Z(n25465) );
  XOR U27373 ( .A(nreg[879]), .B(n25464), .Z(n25467) );
  XNOR U27374 ( .A(n14055), .B(n25464), .Z(n25466) );
  XOR U27375 ( .A(n25468), .B(n25469), .Z(n14055) );
  XOR U27376 ( .A(n25470), .B(n25471), .Z(n25464) );
  AND U27377 ( .A(n25472), .B(n25473), .Z(n25471) );
  XOR U27378 ( .A(nreg[878]), .B(n25470), .Z(n25473) );
  XNOR U27379 ( .A(n14067), .B(n25470), .Z(n25472) );
  XOR U27380 ( .A(n25474), .B(n25475), .Z(n14067) );
  XOR U27381 ( .A(n25476), .B(n25477), .Z(n25470) );
  AND U27382 ( .A(n25478), .B(n25479), .Z(n25477) );
  XOR U27383 ( .A(nreg[877]), .B(n25476), .Z(n25479) );
  XNOR U27384 ( .A(n14079), .B(n25476), .Z(n25478) );
  XOR U27385 ( .A(n25480), .B(n25481), .Z(n14079) );
  XOR U27386 ( .A(n25482), .B(n25483), .Z(n25476) );
  AND U27387 ( .A(n25484), .B(n25485), .Z(n25483) );
  XOR U27388 ( .A(nreg[876]), .B(n25482), .Z(n25485) );
  XNOR U27389 ( .A(n14091), .B(n25482), .Z(n25484) );
  XOR U27390 ( .A(n25486), .B(n25487), .Z(n14091) );
  XOR U27391 ( .A(n25488), .B(n25489), .Z(n25482) );
  AND U27392 ( .A(n25490), .B(n25491), .Z(n25489) );
  XOR U27393 ( .A(nreg[875]), .B(n25488), .Z(n25491) );
  XNOR U27394 ( .A(n14103), .B(n25488), .Z(n25490) );
  XOR U27395 ( .A(n25492), .B(n25493), .Z(n14103) );
  XOR U27396 ( .A(n25494), .B(n25495), .Z(n25488) );
  AND U27397 ( .A(n25496), .B(n25497), .Z(n25495) );
  XOR U27398 ( .A(nreg[874]), .B(n25494), .Z(n25497) );
  XNOR U27399 ( .A(n14115), .B(n25494), .Z(n25496) );
  XOR U27400 ( .A(n25498), .B(n25499), .Z(n14115) );
  XOR U27401 ( .A(n25500), .B(n25501), .Z(n25494) );
  AND U27402 ( .A(n25502), .B(n25503), .Z(n25501) );
  XOR U27403 ( .A(nreg[873]), .B(n25500), .Z(n25503) );
  XNOR U27404 ( .A(n14127), .B(n25500), .Z(n25502) );
  XOR U27405 ( .A(n25504), .B(n25505), .Z(n14127) );
  XOR U27406 ( .A(n25506), .B(n25507), .Z(n25500) );
  AND U27407 ( .A(n25508), .B(n25509), .Z(n25507) );
  XOR U27408 ( .A(nreg[872]), .B(n25506), .Z(n25509) );
  XNOR U27409 ( .A(n14139), .B(n25506), .Z(n25508) );
  XOR U27410 ( .A(n25510), .B(n25511), .Z(n14139) );
  XOR U27411 ( .A(n25512), .B(n25513), .Z(n25506) );
  AND U27412 ( .A(n25514), .B(n25515), .Z(n25513) );
  XOR U27413 ( .A(nreg[871]), .B(n25512), .Z(n25515) );
  XNOR U27414 ( .A(n14151), .B(n25512), .Z(n25514) );
  XOR U27415 ( .A(n25516), .B(n25517), .Z(n14151) );
  XOR U27416 ( .A(n25518), .B(n25519), .Z(n25512) );
  AND U27417 ( .A(n25520), .B(n25521), .Z(n25519) );
  XOR U27418 ( .A(nreg[870]), .B(n25518), .Z(n25521) );
  XNOR U27419 ( .A(n14163), .B(n25518), .Z(n25520) );
  XOR U27420 ( .A(n25522), .B(n25523), .Z(n14163) );
  XOR U27421 ( .A(n25524), .B(n25525), .Z(n25518) );
  AND U27422 ( .A(n25526), .B(n25527), .Z(n25525) );
  XOR U27423 ( .A(nreg[869]), .B(n25524), .Z(n25527) );
  XNOR U27424 ( .A(n14175), .B(n25524), .Z(n25526) );
  XOR U27425 ( .A(n25528), .B(n25529), .Z(n14175) );
  XOR U27426 ( .A(n25530), .B(n25531), .Z(n25524) );
  AND U27427 ( .A(n25532), .B(n25533), .Z(n25531) );
  XOR U27428 ( .A(nreg[868]), .B(n25530), .Z(n25533) );
  XNOR U27429 ( .A(n14187), .B(n25530), .Z(n25532) );
  XOR U27430 ( .A(n25534), .B(n25535), .Z(n14187) );
  XOR U27431 ( .A(n25536), .B(n25537), .Z(n25530) );
  AND U27432 ( .A(n25538), .B(n25539), .Z(n25537) );
  XOR U27433 ( .A(nreg[867]), .B(n25536), .Z(n25539) );
  XNOR U27434 ( .A(n14199), .B(n25536), .Z(n25538) );
  XOR U27435 ( .A(n25540), .B(n25541), .Z(n14199) );
  XOR U27436 ( .A(n25542), .B(n25543), .Z(n25536) );
  AND U27437 ( .A(n25544), .B(n25545), .Z(n25543) );
  XOR U27438 ( .A(nreg[866]), .B(n25542), .Z(n25545) );
  XNOR U27439 ( .A(n14211), .B(n25542), .Z(n25544) );
  XOR U27440 ( .A(n25546), .B(n25547), .Z(n14211) );
  XOR U27441 ( .A(n25548), .B(n25549), .Z(n25542) );
  AND U27442 ( .A(n25550), .B(n25551), .Z(n25549) );
  XOR U27443 ( .A(nreg[865]), .B(n25548), .Z(n25551) );
  XNOR U27444 ( .A(n14223), .B(n25548), .Z(n25550) );
  XOR U27445 ( .A(n25552), .B(n25553), .Z(n14223) );
  XOR U27446 ( .A(n25554), .B(n25555), .Z(n25548) );
  AND U27447 ( .A(n25556), .B(n25557), .Z(n25555) );
  XOR U27448 ( .A(nreg[864]), .B(n25554), .Z(n25557) );
  XNOR U27449 ( .A(n14235), .B(n25554), .Z(n25556) );
  XOR U27450 ( .A(n25558), .B(n25559), .Z(n14235) );
  XOR U27451 ( .A(n25560), .B(n25561), .Z(n25554) );
  AND U27452 ( .A(n25562), .B(n25563), .Z(n25561) );
  XOR U27453 ( .A(nreg[863]), .B(n25560), .Z(n25563) );
  XNOR U27454 ( .A(n14247), .B(n25560), .Z(n25562) );
  XOR U27455 ( .A(n25564), .B(n25565), .Z(n14247) );
  XOR U27456 ( .A(n25566), .B(n25567), .Z(n25560) );
  AND U27457 ( .A(n25568), .B(n25569), .Z(n25567) );
  XOR U27458 ( .A(nreg[862]), .B(n25566), .Z(n25569) );
  XNOR U27459 ( .A(n14259), .B(n25566), .Z(n25568) );
  XOR U27460 ( .A(n25570), .B(n25571), .Z(n14259) );
  XOR U27461 ( .A(n25572), .B(n25573), .Z(n25566) );
  AND U27462 ( .A(n25574), .B(n25575), .Z(n25573) );
  XOR U27463 ( .A(nreg[861]), .B(n25572), .Z(n25575) );
  XNOR U27464 ( .A(n14271), .B(n25572), .Z(n25574) );
  XOR U27465 ( .A(n25576), .B(n25577), .Z(n14271) );
  XOR U27466 ( .A(n25578), .B(n25579), .Z(n25572) );
  AND U27467 ( .A(n25580), .B(n25581), .Z(n25579) );
  XOR U27468 ( .A(nreg[860]), .B(n25578), .Z(n25581) );
  XNOR U27469 ( .A(n14283), .B(n25578), .Z(n25580) );
  XOR U27470 ( .A(n25582), .B(n25583), .Z(n14283) );
  XOR U27471 ( .A(n25584), .B(n25585), .Z(n25578) );
  AND U27472 ( .A(n25586), .B(n25587), .Z(n25585) );
  XOR U27473 ( .A(nreg[859]), .B(n25584), .Z(n25587) );
  XNOR U27474 ( .A(n14295), .B(n25584), .Z(n25586) );
  XOR U27475 ( .A(n25588), .B(n25589), .Z(n14295) );
  XOR U27476 ( .A(n25590), .B(n25591), .Z(n25584) );
  AND U27477 ( .A(n25592), .B(n25593), .Z(n25591) );
  XOR U27478 ( .A(nreg[858]), .B(n25590), .Z(n25593) );
  XNOR U27479 ( .A(n14307), .B(n25590), .Z(n25592) );
  XOR U27480 ( .A(n25594), .B(n25595), .Z(n14307) );
  XOR U27481 ( .A(n25596), .B(n25597), .Z(n25590) );
  AND U27482 ( .A(n25598), .B(n25599), .Z(n25597) );
  XOR U27483 ( .A(nreg[857]), .B(n25596), .Z(n25599) );
  XNOR U27484 ( .A(n14319), .B(n25596), .Z(n25598) );
  XOR U27485 ( .A(n25600), .B(n25601), .Z(n14319) );
  XOR U27486 ( .A(n25602), .B(n25603), .Z(n25596) );
  AND U27487 ( .A(n25604), .B(n25605), .Z(n25603) );
  XOR U27488 ( .A(nreg[856]), .B(n25602), .Z(n25605) );
  XNOR U27489 ( .A(n14331), .B(n25602), .Z(n25604) );
  XOR U27490 ( .A(n25606), .B(n25607), .Z(n14331) );
  XOR U27491 ( .A(n25608), .B(n25609), .Z(n25602) );
  AND U27492 ( .A(n25610), .B(n25611), .Z(n25609) );
  XOR U27493 ( .A(nreg[855]), .B(n25608), .Z(n25611) );
  XNOR U27494 ( .A(n14343), .B(n25608), .Z(n25610) );
  XOR U27495 ( .A(n25612), .B(n25613), .Z(n14343) );
  XOR U27496 ( .A(n25614), .B(n25615), .Z(n25608) );
  AND U27497 ( .A(n25616), .B(n25617), .Z(n25615) );
  XOR U27498 ( .A(nreg[854]), .B(n25614), .Z(n25617) );
  XNOR U27499 ( .A(n14355), .B(n25614), .Z(n25616) );
  XOR U27500 ( .A(n25618), .B(n25619), .Z(n14355) );
  XOR U27501 ( .A(n25620), .B(n25621), .Z(n25614) );
  AND U27502 ( .A(n25622), .B(n25623), .Z(n25621) );
  XOR U27503 ( .A(nreg[853]), .B(n25620), .Z(n25623) );
  XNOR U27504 ( .A(n14367), .B(n25620), .Z(n25622) );
  XOR U27505 ( .A(n25624), .B(n25625), .Z(n14367) );
  XOR U27506 ( .A(n25626), .B(n25627), .Z(n25620) );
  AND U27507 ( .A(n25628), .B(n25629), .Z(n25627) );
  XOR U27508 ( .A(nreg[852]), .B(n25626), .Z(n25629) );
  XNOR U27509 ( .A(n14379), .B(n25626), .Z(n25628) );
  XOR U27510 ( .A(n25630), .B(n25631), .Z(n14379) );
  XOR U27511 ( .A(n25632), .B(n25633), .Z(n25626) );
  AND U27512 ( .A(n25634), .B(n25635), .Z(n25633) );
  XOR U27513 ( .A(nreg[851]), .B(n25632), .Z(n25635) );
  XNOR U27514 ( .A(n14391), .B(n25632), .Z(n25634) );
  XOR U27515 ( .A(n25636), .B(n25637), .Z(n14391) );
  XOR U27516 ( .A(n25638), .B(n25639), .Z(n25632) );
  AND U27517 ( .A(n25640), .B(n25641), .Z(n25639) );
  XOR U27518 ( .A(nreg[850]), .B(n25638), .Z(n25641) );
  XNOR U27519 ( .A(n14403), .B(n25638), .Z(n25640) );
  XOR U27520 ( .A(n25642), .B(n25643), .Z(n14403) );
  XOR U27521 ( .A(n25644), .B(n25645), .Z(n25638) );
  AND U27522 ( .A(n25646), .B(n25647), .Z(n25645) );
  XOR U27523 ( .A(nreg[849]), .B(n25644), .Z(n25647) );
  XNOR U27524 ( .A(n14415), .B(n25644), .Z(n25646) );
  XOR U27525 ( .A(n25648), .B(n25649), .Z(n14415) );
  XOR U27526 ( .A(n25650), .B(n25651), .Z(n25644) );
  AND U27527 ( .A(n25652), .B(n25653), .Z(n25651) );
  XOR U27528 ( .A(nreg[848]), .B(n25650), .Z(n25653) );
  XNOR U27529 ( .A(n14427), .B(n25650), .Z(n25652) );
  XOR U27530 ( .A(n25654), .B(n25655), .Z(n14427) );
  XOR U27531 ( .A(n25656), .B(n25657), .Z(n25650) );
  AND U27532 ( .A(n25658), .B(n25659), .Z(n25657) );
  XOR U27533 ( .A(nreg[847]), .B(n25656), .Z(n25659) );
  XNOR U27534 ( .A(n14439), .B(n25656), .Z(n25658) );
  XOR U27535 ( .A(n25660), .B(n25661), .Z(n14439) );
  XOR U27536 ( .A(n25662), .B(n25663), .Z(n25656) );
  AND U27537 ( .A(n25664), .B(n25665), .Z(n25663) );
  XOR U27538 ( .A(nreg[846]), .B(n25662), .Z(n25665) );
  XNOR U27539 ( .A(n14451), .B(n25662), .Z(n25664) );
  XOR U27540 ( .A(n25666), .B(n25667), .Z(n14451) );
  XOR U27541 ( .A(n25668), .B(n25669), .Z(n25662) );
  AND U27542 ( .A(n25670), .B(n25671), .Z(n25669) );
  XOR U27543 ( .A(nreg[845]), .B(n25668), .Z(n25671) );
  XNOR U27544 ( .A(n14463), .B(n25668), .Z(n25670) );
  XOR U27545 ( .A(n25672), .B(n25673), .Z(n14463) );
  XOR U27546 ( .A(n25674), .B(n25675), .Z(n25668) );
  AND U27547 ( .A(n25676), .B(n25677), .Z(n25675) );
  XOR U27548 ( .A(nreg[844]), .B(n25674), .Z(n25677) );
  XNOR U27549 ( .A(n14475), .B(n25674), .Z(n25676) );
  XOR U27550 ( .A(n25678), .B(n25679), .Z(n14475) );
  XOR U27551 ( .A(n25680), .B(n25681), .Z(n25674) );
  AND U27552 ( .A(n25682), .B(n25683), .Z(n25681) );
  XOR U27553 ( .A(nreg[843]), .B(n25680), .Z(n25683) );
  XNOR U27554 ( .A(n14487), .B(n25680), .Z(n25682) );
  XOR U27555 ( .A(n25684), .B(n25685), .Z(n14487) );
  XOR U27556 ( .A(n25686), .B(n25687), .Z(n25680) );
  AND U27557 ( .A(n25688), .B(n25689), .Z(n25687) );
  XOR U27558 ( .A(nreg[842]), .B(n25686), .Z(n25689) );
  XNOR U27559 ( .A(n14499), .B(n25686), .Z(n25688) );
  XOR U27560 ( .A(n25690), .B(n25691), .Z(n14499) );
  XOR U27561 ( .A(n25692), .B(n25693), .Z(n25686) );
  AND U27562 ( .A(n25694), .B(n25695), .Z(n25693) );
  XOR U27563 ( .A(nreg[841]), .B(n25692), .Z(n25695) );
  XNOR U27564 ( .A(n14511), .B(n25692), .Z(n25694) );
  XOR U27565 ( .A(n25696), .B(n25697), .Z(n14511) );
  XOR U27566 ( .A(n25698), .B(n25699), .Z(n25692) );
  AND U27567 ( .A(n25700), .B(n25701), .Z(n25699) );
  XOR U27568 ( .A(nreg[840]), .B(n25698), .Z(n25701) );
  XNOR U27569 ( .A(n14523), .B(n25698), .Z(n25700) );
  XOR U27570 ( .A(n25702), .B(n25703), .Z(n14523) );
  XOR U27571 ( .A(n25704), .B(n25705), .Z(n25698) );
  AND U27572 ( .A(n25706), .B(n25707), .Z(n25705) );
  XOR U27573 ( .A(nreg[839]), .B(n25704), .Z(n25707) );
  XNOR U27574 ( .A(n14535), .B(n25704), .Z(n25706) );
  XOR U27575 ( .A(n25708), .B(n25709), .Z(n14535) );
  XOR U27576 ( .A(n25710), .B(n25711), .Z(n25704) );
  AND U27577 ( .A(n25712), .B(n25713), .Z(n25711) );
  XOR U27578 ( .A(nreg[838]), .B(n25710), .Z(n25713) );
  XNOR U27579 ( .A(n14547), .B(n25710), .Z(n25712) );
  XOR U27580 ( .A(n25714), .B(n25715), .Z(n14547) );
  XOR U27581 ( .A(n25716), .B(n25717), .Z(n25710) );
  AND U27582 ( .A(n25718), .B(n25719), .Z(n25717) );
  XOR U27583 ( .A(nreg[837]), .B(n25716), .Z(n25719) );
  XNOR U27584 ( .A(n14559), .B(n25716), .Z(n25718) );
  XOR U27585 ( .A(n25720), .B(n25721), .Z(n14559) );
  XOR U27586 ( .A(n25722), .B(n25723), .Z(n25716) );
  AND U27587 ( .A(n25724), .B(n25725), .Z(n25723) );
  XOR U27588 ( .A(nreg[836]), .B(n25722), .Z(n25725) );
  XNOR U27589 ( .A(n14571), .B(n25722), .Z(n25724) );
  XOR U27590 ( .A(n25726), .B(n25727), .Z(n14571) );
  XOR U27591 ( .A(n25728), .B(n25729), .Z(n25722) );
  AND U27592 ( .A(n25730), .B(n25731), .Z(n25729) );
  XOR U27593 ( .A(nreg[835]), .B(n25728), .Z(n25731) );
  XNOR U27594 ( .A(n14583), .B(n25728), .Z(n25730) );
  XOR U27595 ( .A(n25732), .B(n25733), .Z(n14583) );
  XOR U27596 ( .A(n25734), .B(n25735), .Z(n25728) );
  AND U27597 ( .A(n25736), .B(n25737), .Z(n25735) );
  XOR U27598 ( .A(nreg[834]), .B(n25734), .Z(n25737) );
  XNOR U27599 ( .A(n14595), .B(n25734), .Z(n25736) );
  XOR U27600 ( .A(n25738), .B(n25739), .Z(n14595) );
  XOR U27601 ( .A(n25740), .B(n25741), .Z(n25734) );
  AND U27602 ( .A(n25742), .B(n25743), .Z(n25741) );
  XOR U27603 ( .A(nreg[833]), .B(n25740), .Z(n25743) );
  XNOR U27604 ( .A(n14607), .B(n25740), .Z(n25742) );
  XOR U27605 ( .A(n25744), .B(n25745), .Z(n14607) );
  XOR U27606 ( .A(n25746), .B(n25747), .Z(n25740) );
  AND U27607 ( .A(n25748), .B(n25749), .Z(n25747) );
  XOR U27608 ( .A(nreg[832]), .B(n25746), .Z(n25749) );
  XNOR U27609 ( .A(n14619), .B(n25746), .Z(n25748) );
  XOR U27610 ( .A(n25750), .B(n25751), .Z(n14619) );
  XOR U27611 ( .A(n25752), .B(n25753), .Z(n25746) );
  AND U27612 ( .A(n25754), .B(n25755), .Z(n25753) );
  XOR U27613 ( .A(nreg[831]), .B(n25752), .Z(n25755) );
  XNOR U27614 ( .A(n14631), .B(n25752), .Z(n25754) );
  XOR U27615 ( .A(n25756), .B(n25757), .Z(n14631) );
  XOR U27616 ( .A(n25758), .B(n25759), .Z(n25752) );
  AND U27617 ( .A(n25760), .B(n25761), .Z(n25759) );
  XOR U27618 ( .A(nreg[830]), .B(n25758), .Z(n25761) );
  XNOR U27619 ( .A(n14643), .B(n25758), .Z(n25760) );
  XOR U27620 ( .A(n25762), .B(n25763), .Z(n14643) );
  XOR U27621 ( .A(n25764), .B(n25765), .Z(n25758) );
  AND U27622 ( .A(n25766), .B(n25767), .Z(n25765) );
  XOR U27623 ( .A(nreg[829]), .B(n25764), .Z(n25767) );
  XNOR U27624 ( .A(n14655), .B(n25764), .Z(n25766) );
  XOR U27625 ( .A(n25768), .B(n25769), .Z(n14655) );
  XOR U27626 ( .A(n25770), .B(n25771), .Z(n25764) );
  AND U27627 ( .A(n25772), .B(n25773), .Z(n25771) );
  XOR U27628 ( .A(nreg[828]), .B(n25770), .Z(n25773) );
  XNOR U27629 ( .A(n14667), .B(n25770), .Z(n25772) );
  XOR U27630 ( .A(n25774), .B(n25775), .Z(n14667) );
  XOR U27631 ( .A(n25776), .B(n25777), .Z(n25770) );
  AND U27632 ( .A(n25778), .B(n25779), .Z(n25777) );
  XOR U27633 ( .A(nreg[827]), .B(n25776), .Z(n25779) );
  XNOR U27634 ( .A(n14679), .B(n25776), .Z(n25778) );
  XOR U27635 ( .A(n25780), .B(n25781), .Z(n14679) );
  XOR U27636 ( .A(n25782), .B(n25783), .Z(n25776) );
  AND U27637 ( .A(n25784), .B(n25785), .Z(n25783) );
  XOR U27638 ( .A(nreg[826]), .B(n25782), .Z(n25785) );
  XNOR U27639 ( .A(n14691), .B(n25782), .Z(n25784) );
  XOR U27640 ( .A(n25786), .B(n25787), .Z(n14691) );
  XOR U27641 ( .A(n25788), .B(n25789), .Z(n25782) );
  AND U27642 ( .A(n25790), .B(n25791), .Z(n25789) );
  XOR U27643 ( .A(nreg[825]), .B(n25788), .Z(n25791) );
  XNOR U27644 ( .A(n14703), .B(n25788), .Z(n25790) );
  XOR U27645 ( .A(n25792), .B(n25793), .Z(n14703) );
  XOR U27646 ( .A(n25794), .B(n25795), .Z(n25788) );
  AND U27647 ( .A(n25796), .B(n25797), .Z(n25795) );
  XOR U27648 ( .A(nreg[824]), .B(n25794), .Z(n25797) );
  XNOR U27649 ( .A(n14715), .B(n25794), .Z(n25796) );
  XOR U27650 ( .A(n25798), .B(n25799), .Z(n14715) );
  XOR U27651 ( .A(n25800), .B(n25801), .Z(n25794) );
  AND U27652 ( .A(n25802), .B(n25803), .Z(n25801) );
  XOR U27653 ( .A(nreg[823]), .B(n25800), .Z(n25803) );
  XNOR U27654 ( .A(n14727), .B(n25800), .Z(n25802) );
  XOR U27655 ( .A(n25804), .B(n25805), .Z(n14727) );
  XOR U27656 ( .A(n25806), .B(n25807), .Z(n25800) );
  AND U27657 ( .A(n25808), .B(n25809), .Z(n25807) );
  XOR U27658 ( .A(nreg[822]), .B(n25806), .Z(n25809) );
  XNOR U27659 ( .A(n14739), .B(n25806), .Z(n25808) );
  XOR U27660 ( .A(n25810), .B(n25811), .Z(n14739) );
  XOR U27661 ( .A(n25812), .B(n25813), .Z(n25806) );
  AND U27662 ( .A(n25814), .B(n25815), .Z(n25813) );
  XOR U27663 ( .A(nreg[821]), .B(n25812), .Z(n25815) );
  XNOR U27664 ( .A(n14751), .B(n25812), .Z(n25814) );
  XOR U27665 ( .A(n25816), .B(n25817), .Z(n14751) );
  XOR U27666 ( .A(n25818), .B(n25819), .Z(n25812) );
  AND U27667 ( .A(n25820), .B(n25821), .Z(n25819) );
  XOR U27668 ( .A(nreg[820]), .B(n25818), .Z(n25821) );
  XNOR U27669 ( .A(n14763), .B(n25818), .Z(n25820) );
  XOR U27670 ( .A(n25822), .B(n25823), .Z(n14763) );
  XOR U27671 ( .A(n25824), .B(n25825), .Z(n25818) );
  AND U27672 ( .A(n25826), .B(n25827), .Z(n25825) );
  XOR U27673 ( .A(nreg[819]), .B(n25824), .Z(n25827) );
  XNOR U27674 ( .A(n14775), .B(n25824), .Z(n25826) );
  XOR U27675 ( .A(n25828), .B(n25829), .Z(n14775) );
  XOR U27676 ( .A(n25830), .B(n25831), .Z(n25824) );
  AND U27677 ( .A(n25832), .B(n25833), .Z(n25831) );
  XOR U27678 ( .A(nreg[818]), .B(n25830), .Z(n25833) );
  XNOR U27679 ( .A(n14787), .B(n25830), .Z(n25832) );
  XOR U27680 ( .A(n25834), .B(n25835), .Z(n14787) );
  XOR U27681 ( .A(n25836), .B(n25837), .Z(n25830) );
  AND U27682 ( .A(n25838), .B(n25839), .Z(n25837) );
  XOR U27683 ( .A(nreg[817]), .B(n25836), .Z(n25839) );
  XNOR U27684 ( .A(n14799), .B(n25836), .Z(n25838) );
  XOR U27685 ( .A(n25840), .B(n25841), .Z(n14799) );
  XOR U27686 ( .A(n25842), .B(n25843), .Z(n25836) );
  AND U27687 ( .A(n25844), .B(n25845), .Z(n25843) );
  XOR U27688 ( .A(nreg[816]), .B(n25842), .Z(n25845) );
  XNOR U27689 ( .A(n14811), .B(n25842), .Z(n25844) );
  XOR U27690 ( .A(n25846), .B(n25847), .Z(n14811) );
  XOR U27691 ( .A(n25848), .B(n25849), .Z(n25842) );
  AND U27692 ( .A(n25850), .B(n25851), .Z(n25849) );
  XOR U27693 ( .A(nreg[815]), .B(n25848), .Z(n25851) );
  XNOR U27694 ( .A(n14823), .B(n25848), .Z(n25850) );
  XOR U27695 ( .A(n25852), .B(n25853), .Z(n14823) );
  XOR U27696 ( .A(n25854), .B(n25855), .Z(n25848) );
  AND U27697 ( .A(n25856), .B(n25857), .Z(n25855) );
  XOR U27698 ( .A(nreg[814]), .B(n25854), .Z(n25857) );
  XNOR U27699 ( .A(n14835), .B(n25854), .Z(n25856) );
  XOR U27700 ( .A(n25858), .B(n25859), .Z(n14835) );
  XOR U27701 ( .A(n25860), .B(n25861), .Z(n25854) );
  AND U27702 ( .A(n25862), .B(n25863), .Z(n25861) );
  XOR U27703 ( .A(nreg[813]), .B(n25860), .Z(n25863) );
  XNOR U27704 ( .A(n14847), .B(n25860), .Z(n25862) );
  XOR U27705 ( .A(n25864), .B(n25865), .Z(n14847) );
  XOR U27706 ( .A(n25866), .B(n25867), .Z(n25860) );
  AND U27707 ( .A(n25868), .B(n25869), .Z(n25867) );
  XOR U27708 ( .A(nreg[812]), .B(n25866), .Z(n25869) );
  XNOR U27709 ( .A(n14859), .B(n25866), .Z(n25868) );
  XOR U27710 ( .A(n25870), .B(n25871), .Z(n14859) );
  XOR U27711 ( .A(n25872), .B(n25873), .Z(n25866) );
  AND U27712 ( .A(n25874), .B(n25875), .Z(n25873) );
  XOR U27713 ( .A(nreg[811]), .B(n25872), .Z(n25875) );
  XNOR U27714 ( .A(n14871), .B(n25872), .Z(n25874) );
  XOR U27715 ( .A(n25876), .B(n25877), .Z(n14871) );
  XOR U27716 ( .A(n25878), .B(n25879), .Z(n25872) );
  AND U27717 ( .A(n25880), .B(n25881), .Z(n25879) );
  XOR U27718 ( .A(nreg[810]), .B(n25878), .Z(n25881) );
  XNOR U27719 ( .A(n14883), .B(n25878), .Z(n25880) );
  XOR U27720 ( .A(n25882), .B(n25883), .Z(n14883) );
  XOR U27721 ( .A(n25884), .B(n25885), .Z(n25878) );
  AND U27722 ( .A(n25886), .B(n25887), .Z(n25885) );
  XOR U27723 ( .A(nreg[809]), .B(n25884), .Z(n25887) );
  XNOR U27724 ( .A(n14895), .B(n25884), .Z(n25886) );
  XOR U27725 ( .A(n25888), .B(n25889), .Z(n14895) );
  XOR U27726 ( .A(n25890), .B(n25891), .Z(n25884) );
  AND U27727 ( .A(n25892), .B(n25893), .Z(n25891) );
  XOR U27728 ( .A(nreg[808]), .B(n25890), .Z(n25893) );
  XNOR U27729 ( .A(n14907), .B(n25890), .Z(n25892) );
  XOR U27730 ( .A(n25894), .B(n25895), .Z(n14907) );
  XOR U27731 ( .A(n25896), .B(n25897), .Z(n25890) );
  AND U27732 ( .A(n25898), .B(n25899), .Z(n25897) );
  XOR U27733 ( .A(nreg[807]), .B(n25896), .Z(n25899) );
  XNOR U27734 ( .A(n14919), .B(n25896), .Z(n25898) );
  XOR U27735 ( .A(n25900), .B(n25901), .Z(n14919) );
  XOR U27736 ( .A(n25902), .B(n25903), .Z(n25896) );
  AND U27737 ( .A(n25904), .B(n25905), .Z(n25903) );
  XOR U27738 ( .A(nreg[806]), .B(n25902), .Z(n25905) );
  XNOR U27739 ( .A(n14931), .B(n25902), .Z(n25904) );
  XOR U27740 ( .A(n25906), .B(n25907), .Z(n14931) );
  XOR U27741 ( .A(n25908), .B(n25909), .Z(n25902) );
  AND U27742 ( .A(n25910), .B(n25911), .Z(n25909) );
  XOR U27743 ( .A(nreg[805]), .B(n25908), .Z(n25911) );
  XNOR U27744 ( .A(n14943), .B(n25908), .Z(n25910) );
  XOR U27745 ( .A(n25912), .B(n25913), .Z(n14943) );
  XOR U27746 ( .A(n25914), .B(n25915), .Z(n25908) );
  AND U27747 ( .A(n25916), .B(n25917), .Z(n25915) );
  XOR U27748 ( .A(nreg[804]), .B(n25914), .Z(n25917) );
  XNOR U27749 ( .A(n14955), .B(n25914), .Z(n25916) );
  XOR U27750 ( .A(n25918), .B(n25919), .Z(n14955) );
  XOR U27751 ( .A(n25920), .B(n25921), .Z(n25914) );
  AND U27752 ( .A(n25922), .B(n25923), .Z(n25921) );
  XOR U27753 ( .A(nreg[803]), .B(n25920), .Z(n25923) );
  XNOR U27754 ( .A(n14967), .B(n25920), .Z(n25922) );
  XOR U27755 ( .A(n25924), .B(n25925), .Z(n14967) );
  XOR U27756 ( .A(n25926), .B(n25927), .Z(n25920) );
  AND U27757 ( .A(n25928), .B(n25929), .Z(n25927) );
  XOR U27758 ( .A(nreg[802]), .B(n25926), .Z(n25929) );
  XNOR U27759 ( .A(n14979), .B(n25926), .Z(n25928) );
  XOR U27760 ( .A(n25930), .B(n25931), .Z(n14979) );
  XOR U27761 ( .A(n25932), .B(n25933), .Z(n25926) );
  AND U27762 ( .A(n25934), .B(n25935), .Z(n25933) );
  XOR U27763 ( .A(nreg[801]), .B(n25932), .Z(n25935) );
  XNOR U27764 ( .A(n14991), .B(n25932), .Z(n25934) );
  XOR U27765 ( .A(n25936), .B(n25937), .Z(n14991) );
  XOR U27766 ( .A(n25938), .B(n25939), .Z(n25932) );
  AND U27767 ( .A(n25940), .B(n25941), .Z(n25939) );
  XOR U27768 ( .A(nreg[800]), .B(n25938), .Z(n25941) );
  XNOR U27769 ( .A(n15003), .B(n25938), .Z(n25940) );
  XOR U27770 ( .A(n25942), .B(n25943), .Z(n15003) );
  XOR U27771 ( .A(n25944), .B(n25945), .Z(n25938) );
  AND U27772 ( .A(n25946), .B(n25947), .Z(n25945) );
  XOR U27773 ( .A(nreg[799]), .B(n25944), .Z(n25947) );
  XNOR U27774 ( .A(n15015), .B(n25944), .Z(n25946) );
  XOR U27775 ( .A(n25948), .B(n25949), .Z(n15015) );
  XOR U27776 ( .A(n25950), .B(n25951), .Z(n25944) );
  AND U27777 ( .A(n25952), .B(n25953), .Z(n25951) );
  XOR U27778 ( .A(nreg[798]), .B(n25950), .Z(n25953) );
  XNOR U27779 ( .A(n15027), .B(n25950), .Z(n25952) );
  XOR U27780 ( .A(n25954), .B(n25955), .Z(n15027) );
  XOR U27781 ( .A(n25956), .B(n25957), .Z(n25950) );
  AND U27782 ( .A(n25958), .B(n25959), .Z(n25957) );
  XOR U27783 ( .A(nreg[797]), .B(n25956), .Z(n25959) );
  XNOR U27784 ( .A(n15039), .B(n25956), .Z(n25958) );
  XOR U27785 ( .A(n25960), .B(n25961), .Z(n15039) );
  XOR U27786 ( .A(n25962), .B(n25963), .Z(n25956) );
  AND U27787 ( .A(n25964), .B(n25965), .Z(n25963) );
  XOR U27788 ( .A(nreg[796]), .B(n25962), .Z(n25965) );
  XNOR U27789 ( .A(n15051), .B(n25962), .Z(n25964) );
  XOR U27790 ( .A(n25966), .B(n25967), .Z(n15051) );
  XOR U27791 ( .A(n25968), .B(n25969), .Z(n25962) );
  AND U27792 ( .A(n25970), .B(n25971), .Z(n25969) );
  XOR U27793 ( .A(nreg[795]), .B(n25968), .Z(n25971) );
  XNOR U27794 ( .A(n15063), .B(n25968), .Z(n25970) );
  XOR U27795 ( .A(n25972), .B(n25973), .Z(n15063) );
  XOR U27796 ( .A(n25974), .B(n25975), .Z(n25968) );
  AND U27797 ( .A(n25976), .B(n25977), .Z(n25975) );
  XOR U27798 ( .A(nreg[794]), .B(n25974), .Z(n25977) );
  XNOR U27799 ( .A(n15075), .B(n25974), .Z(n25976) );
  XOR U27800 ( .A(n25978), .B(n25979), .Z(n15075) );
  XOR U27801 ( .A(n25980), .B(n25981), .Z(n25974) );
  AND U27802 ( .A(n25982), .B(n25983), .Z(n25981) );
  XOR U27803 ( .A(nreg[793]), .B(n25980), .Z(n25983) );
  XNOR U27804 ( .A(n15087), .B(n25980), .Z(n25982) );
  XOR U27805 ( .A(n25984), .B(n25985), .Z(n15087) );
  XOR U27806 ( .A(n25986), .B(n25987), .Z(n25980) );
  AND U27807 ( .A(n25988), .B(n25989), .Z(n25987) );
  XOR U27808 ( .A(nreg[792]), .B(n25986), .Z(n25989) );
  XNOR U27809 ( .A(n15099), .B(n25986), .Z(n25988) );
  XOR U27810 ( .A(n25990), .B(n25991), .Z(n15099) );
  XOR U27811 ( .A(n25992), .B(n25993), .Z(n25986) );
  AND U27812 ( .A(n25994), .B(n25995), .Z(n25993) );
  XOR U27813 ( .A(nreg[791]), .B(n25992), .Z(n25995) );
  XNOR U27814 ( .A(n15111), .B(n25992), .Z(n25994) );
  XOR U27815 ( .A(n25996), .B(n25997), .Z(n15111) );
  XOR U27816 ( .A(n25998), .B(n25999), .Z(n25992) );
  AND U27817 ( .A(n26000), .B(n26001), .Z(n25999) );
  XOR U27818 ( .A(nreg[790]), .B(n25998), .Z(n26001) );
  XNOR U27819 ( .A(n15123), .B(n25998), .Z(n26000) );
  XOR U27820 ( .A(n26002), .B(n26003), .Z(n15123) );
  XOR U27821 ( .A(n26004), .B(n26005), .Z(n25998) );
  AND U27822 ( .A(n26006), .B(n26007), .Z(n26005) );
  XOR U27823 ( .A(nreg[789]), .B(n26004), .Z(n26007) );
  XNOR U27824 ( .A(n15135), .B(n26004), .Z(n26006) );
  XOR U27825 ( .A(n26008), .B(n26009), .Z(n15135) );
  XOR U27826 ( .A(n26010), .B(n26011), .Z(n26004) );
  AND U27827 ( .A(n26012), .B(n26013), .Z(n26011) );
  XOR U27828 ( .A(nreg[788]), .B(n26010), .Z(n26013) );
  XNOR U27829 ( .A(n15147), .B(n26010), .Z(n26012) );
  XOR U27830 ( .A(n26014), .B(n26015), .Z(n15147) );
  XOR U27831 ( .A(n26016), .B(n26017), .Z(n26010) );
  AND U27832 ( .A(n26018), .B(n26019), .Z(n26017) );
  XOR U27833 ( .A(nreg[787]), .B(n26016), .Z(n26019) );
  XNOR U27834 ( .A(n15159), .B(n26016), .Z(n26018) );
  XOR U27835 ( .A(n26020), .B(n26021), .Z(n15159) );
  XOR U27836 ( .A(n26022), .B(n26023), .Z(n26016) );
  AND U27837 ( .A(n26024), .B(n26025), .Z(n26023) );
  XOR U27838 ( .A(nreg[786]), .B(n26022), .Z(n26025) );
  XNOR U27839 ( .A(n15171), .B(n26022), .Z(n26024) );
  XOR U27840 ( .A(n26026), .B(n26027), .Z(n15171) );
  XOR U27841 ( .A(n26028), .B(n26029), .Z(n26022) );
  AND U27842 ( .A(n26030), .B(n26031), .Z(n26029) );
  XOR U27843 ( .A(nreg[785]), .B(n26028), .Z(n26031) );
  XNOR U27844 ( .A(n15183), .B(n26028), .Z(n26030) );
  XOR U27845 ( .A(n26032), .B(n26033), .Z(n15183) );
  XOR U27846 ( .A(n26034), .B(n26035), .Z(n26028) );
  AND U27847 ( .A(n26036), .B(n26037), .Z(n26035) );
  XOR U27848 ( .A(nreg[784]), .B(n26034), .Z(n26037) );
  XNOR U27849 ( .A(n15195), .B(n26034), .Z(n26036) );
  XOR U27850 ( .A(n26038), .B(n26039), .Z(n15195) );
  XOR U27851 ( .A(n26040), .B(n26041), .Z(n26034) );
  AND U27852 ( .A(n26042), .B(n26043), .Z(n26041) );
  XOR U27853 ( .A(nreg[783]), .B(n26040), .Z(n26043) );
  XNOR U27854 ( .A(n15207), .B(n26040), .Z(n26042) );
  XOR U27855 ( .A(n26044), .B(n26045), .Z(n15207) );
  XOR U27856 ( .A(n26046), .B(n26047), .Z(n26040) );
  AND U27857 ( .A(n26048), .B(n26049), .Z(n26047) );
  XOR U27858 ( .A(nreg[782]), .B(n26046), .Z(n26049) );
  XNOR U27859 ( .A(n15219), .B(n26046), .Z(n26048) );
  XOR U27860 ( .A(n26050), .B(n26051), .Z(n15219) );
  XOR U27861 ( .A(n26052), .B(n26053), .Z(n26046) );
  AND U27862 ( .A(n26054), .B(n26055), .Z(n26053) );
  XOR U27863 ( .A(nreg[781]), .B(n26052), .Z(n26055) );
  XNOR U27864 ( .A(n15231), .B(n26052), .Z(n26054) );
  XOR U27865 ( .A(n26056), .B(n26057), .Z(n15231) );
  XOR U27866 ( .A(n26058), .B(n26059), .Z(n26052) );
  AND U27867 ( .A(n26060), .B(n26061), .Z(n26059) );
  XOR U27868 ( .A(nreg[780]), .B(n26058), .Z(n26061) );
  XNOR U27869 ( .A(n15243), .B(n26058), .Z(n26060) );
  XOR U27870 ( .A(n26062), .B(n26063), .Z(n15243) );
  XOR U27871 ( .A(n26064), .B(n26065), .Z(n26058) );
  AND U27872 ( .A(n26066), .B(n26067), .Z(n26065) );
  XOR U27873 ( .A(nreg[779]), .B(n26064), .Z(n26067) );
  XNOR U27874 ( .A(n15255), .B(n26064), .Z(n26066) );
  XOR U27875 ( .A(n26068), .B(n26069), .Z(n15255) );
  XOR U27876 ( .A(n26070), .B(n26071), .Z(n26064) );
  AND U27877 ( .A(n26072), .B(n26073), .Z(n26071) );
  XOR U27878 ( .A(nreg[778]), .B(n26070), .Z(n26073) );
  XNOR U27879 ( .A(n15267), .B(n26070), .Z(n26072) );
  XOR U27880 ( .A(n26074), .B(n26075), .Z(n15267) );
  XOR U27881 ( .A(n26076), .B(n26077), .Z(n26070) );
  AND U27882 ( .A(n26078), .B(n26079), .Z(n26077) );
  XOR U27883 ( .A(nreg[777]), .B(n26076), .Z(n26079) );
  XNOR U27884 ( .A(n15279), .B(n26076), .Z(n26078) );
  XOR U27885 ( .A(n26080), .B(n26081), .Z(n15279) );
  XOR U27886 ( .A(n26082), .B(n26083), .Z(n26076) );
  AND U27887 ( .A(n26084), .B(n26085), .Z(n26083) );
  XOR U27888 ( .A(nreg[776]), .B(n26082), .Z(n26085) );
  XNOR U27889 ( .A(n15291), .B(n26082), .Z(n26084) );
  XOR U27890 ( .A(n26086), .B(n26087), .Z(n15291) );
  XOR U27891 ( .A(n26088), .B(n26089), .Z(n26082) );
  AND U27892 ( .A(n26090), .B(n26091), .Z(n26089) );
  XOR U27893 ( .A(nreg[775]), .B(n26088), .Z(n26091) );
  XNOR U27894 ( .A(n15303), .B(n26088), .Z(n26090) );
  XOR U27895 ( .A(n26092), .B(n26093), .Z(n15303) );
  XOR U27896 ( .A(n26094), .B(n26095), .Z(n26088) );
  AND U27897 ( .A(n26096), .B(n26097), .Z(n26095) );
  XOR U27898 ( .A(nreg[774]), .B(n26094), .Z(n26097) );
  XNOR U27899 ( .A(n15315), .B(n26094), .Z(n26096) );
  XOR U27900 ( .A(n26098), .B(n26099), .Z(n15315) );
  XOR U27901 ( .A(n26100), .B(n26101), .Z(n26094) );
  AND U27902 ( .A(n26102), .B(n26103), .Z(n26101) );
  XOR U27903 ( .A(nreg[773]), .B(n26100), .Z(n26103) );
  XNOR U27904 ( .A(n15327), .B(n26100), .Z(n26102) );
  XOR U27905 ( .A(n26104), .B(n26105), .Z(n15327) );
  XOR U27906 ( .A(n26106), .B(n26107), .Z(n26100) );
  AND U27907 ( .A(n26108), .B(n26109), .Z(n26107) );
  XOR U27908 ( .A(nreg[772]), .B(n26106), .Z(n26109) );
  XNOR U27909 ( .A(n15339), .B(n26106), .Z(n26108) );
  XOR U27910 ( .A(n26110), .B(n26111), .Z(n15339) );
  XOR U27911 ( .A(n26112), .B(n26113), .Z(n26106) );
  AND U27912 ( .A(n26114), .B(n26115), .Z(n26113) );
  XOR U27913 ( .A(nreg[771]), .B(n26112), .Z(n26115) );
  XNOR U27914 ( .A(n15351), .B(n26112), .Z(n26114) );
  XOR U27915 ( .A(n26116), .B(n26117), .Z(n15351) );
  XOR U27916 ( .A(n26118), .B(n26119), .Z(n26112) );
  AND U27917 ( .A(n26120), .B(n26121), .Z(n26119) );
  XOR U27918 ( .A(nreg[770]), .B(n26118), .Z(n26121) );
  XNOR U27919 ( .A(n15363), .B(n26118), .Z(n26120) );
  XOR U27920 ( .A(n26122), .B(n26123), .Z(n15363) );
  XOR U27921 ( .A(n26124), .B(n26125), .Z(n26118) );
  AND U27922 ( .A(n26126), .B(n26127), .Z(n26125) );
  XOR U27923 ( .A(nreg[769]), .B(n26124), .Z(n26127) );
  XNOR U27924 ( .A(n15375), .B(n26124), .Z(n26126) );
  XOR U27925 ( .A(n26128), .B(n26129), .Z(n15375) );
  XOR U27926 ( .A(n26130), .B(n26131), .Z(n26124) );
  AND U27927 ( .A(n26132), .B(n26133), .Z(n26131) );
  XOR U27928 ( .A(nreg[768]), .B(n26130), .Z(n26133) );
  XNOR U27929 ( .A(n15387), .B(n26130), .Z(n26132) );
  XOR U27930 ( .A(n26134), .B(n26135), .Z(n15387) );
  XOR U27931 ( .A(n26136), .B(n26137), .Z(n26130) );
  AND U27932 ( .A(n26138), .B(n26139), .Z(n26137) );
  XOR U27933 ( .A(nreg[767]), .B(n26136), .Z(n26139) );
  XNOR U27934 ( .A(n15399), .B(n26136), .Z(n26138) );
  XOR U27935 ( .A(n26140), .B(n26141), .Z(n15399) );
  XOR U27936 ( .A(n26142), .B(n26143), .Z(n26136) );
  AND U27937 ( .A(n26144), .B(n26145), .Z(n26143) );
  XOR U27938 ( .A(nreg[766]), .B(n26142), .Z(n26145) );
  XNOR U27939 ( .A(n15411), .B(n26142), .Z(n26144) );
  XOR U27940 ( .A(n26146), .B(n26147), .Z(n15411) );
  XOR U27941 ( .A(n26148), .B(n26149), .Z(n26142) );
  AND U27942 ( .A(n26150), .B(n26151), .Z(n26149) );
  XOR U27943 ( .A(nreg[765]), .B(n26148), .Z(n26151) );
  XNOR U27944 ( .A(n15423), .B(n26148), .Z(n26150) );
  XOR U27945 ( .A(n26152), .B(n26153), .Z(n15423) );
  XOR U27946 ( .A(n26154), .B(n26155), .Z(n26148) );
  AND U27947 ( .A(n26156), .B(n26157), .Z(n26155) );
  XOR U27948 ( .A(nreg[764]), .B(n26154), .Z(n26157) );
  XNOR U27949 ( .A(n15435), .B(n26154), .Z(n26156) );
  XOR U27950 ( .A(n26158), .B(n26159), .Z(n15435) );
  XOR U27951 ( .A(n26160), .B(n26161), .Z(n26154) );
  AND U27952 ( .A(n26162), .B(n26163), .Z(n26161) );
  XOR U27953 ( .A(nreg[763]), .B(n26160), .Z(n26163) );
  XNOR U27954 ( .A(n15447), .B(n26160), .Z(n26162) );
  XOR U27955 ( .A(n26164), .B(n26165), .Z(n15447) );
  XOR U27956 ( .A(n26166), .B(n26167), .Z(n26160) );
  AND U27957 ( .A(n26168), .B(n26169), .Z(n26167) );
  XOR U27958 ( .A(nreg[762]), .B(n26166), .Z(n26169) );
  XNOR U27959 ( .A(n15459), .B(n26166), .Z(n26168) );
  XOR U27960 ( .A(n26170), .B(n26171), .Z(n15459) );
  XOR U27961 ( .A(n26172), .B(n26173), .Z(n26166) );
  AND U27962 ( .A(n26174), .B(n26175), .Z(n26173) );
  XOR U27963 ( .A(nreg[761]), .B(n26172), .Z(n26175) );
  XNOR U27964 ( .A(n15471), .B(n26172), .Z(n26174) );
  XOR U27965 ( .A(n26176), .B(n26177), .Z(n15471) );
  XOR U27966 ( .A(n26178), .B(n26179), .Z(n26172) );
  AND U27967 ( .A(n26180), .B(n26181), .Z(n26179) );
  XOR U27968 ( .A(nreg[760]), .B(n26178), .Z(n26181) );
  XNOR U27969 ( .A(n15483), .B(n26178), .Z(n26180) );
  XOR U27970 ( .A(n26182), .B(n26183), .Z(n15483) );
  XOR U27971 ( .A(n26184), .B(n26185), .Z(n26178) );
  AND U27972 ( .A(n26186), .B(n26187), .Z(n26185) );
  XOR U27973 ( .A(nreg[759]), .B(n26184), .Z(n26187) );
  XNOR U27974 ( .A(n15495), .B(n26184), .Z(n26186) );
  XOR U27975 ( .A(n26188), .B(n26189), .Z(n15495) );
  XOR U27976 ( .A(n26190), .B(n26191), .Z(n26184) );
  AND U27977 ( .A(n26192), .B(n26193), .Z(n26191) );
  XOR U27978 ( .A(nreg[758]), .B(n26190), .Z(n26193) );
  XNOR U27979 ( .A(n15507), .B(n26190), .Z(n26192) );
  XOR U27980 ( .A(n26194), .B(n26195), .Z(n15507) );
  XOR U27981 ( .A(n26196), .B(n26197), .Z(n26190) );
  AND U27982 ( .A(n26198), .B(n26199), .Z(n26197) );
  XOR U27983 ( .A(nreg[757]), .B(n26196), .Z(n26199) );
  XNOR U27984 ( .A(n15519), .B(n26196), .Z(n26198) );
  XOR U27985 ( .A(n26200), .B(n26201), .Z(n15519) );
  XOR U27986 ( .A(n26202), .B(n26203), .Z(n26196) );
  AND U27987 ( .A(n26204), .B(n26205), .Z(n26203) );
  XOR U27988 ( .A(nreg[756]), .B(n26202), .Z(n26205) );
  XNOR U27989 ( .A(n15531), .B(n26202), .Z(n26204) );
  XOR U27990 ( .A(n26206), .B(n26207), .Z(n15531) );
  XOR U27991 ( .A(n26208), .B(n26209), .Z(n26202) );
  AND U27992 ( .A(n26210), .B(n26211), .Z(n26209) );
  XOR U27993 ( .A(nreg[755]), .B(n26208), .Z(n26211) );
  XNOR U27994 ( .A(n15543), .B(n26208), .Z(n26210) );
  XOR U27995 ( .A(n26212), .B(n26213), .Z(n15543) );
  XOR U27996 ( .A(n26214), .B(n26215), .Z(n26208) );
  AND U27997 ( .A(n26216), .B(n26217), .Z(n26215) );
  XOR U27998 ( .A(nreg[754]), .B(n26214), .Z(n26217) );
  XNOR U27999 ( .A(n15555), .B(n26214), .Z(n26216) );
  XOR U28000 ( .A(n26218), .B(n26219), .Z(n15555) );
  XOR U28001 ( .A(n26220), .B(n26221), .Z(n26214) );
  AND U28002 ( .A(n26222), .B(n26223), .Z(n26221) );
  XOR U28003 ( .A(nreg[753]), .B(n26220), .Z(n26223) );
  XNOR U28004 ( .A(n15567), .B(n26220), .Z(n26222) );
  XOR U28005 ( .A(n26224), .B(n26225), .Z(n15567) );
  XOR U28006 ( .A(n26226), .B(n26227), .Z(n26220) );
  AND U28007 ( .A(n26228), .B(n26229), .Z(n26227) );
  XOR U28008 ( .A(nreg[752]), .B(n26226), .Z(n26229) );
  XNOR U28009 ( .A(n15579), .B(n26226), .Z(n26228) );
  XOR U28010 ( .A(n26230), .B(n26231), .Z(n15579) );
  XOR U28011 ( .A(n26232), .B(n26233), .Z(n26226) );
  AND U28012 ( .A(n26234), .B(n26235), .Z(n26233) );
  XOR U28013 ( .A(nreg[751]), .B(n26232), .Z(n26235) );
  XNOR U28014 ( .A(n15591), .B(n26232), .Z(n26234) );
  XOR U28015 ( .A(n26236), .B(n26237), .Z(n15591) );
  XOR U28016 ( .A(n26238), .B(n26239), .Z(n26232) );
  AND U28017 ( .A(n26240), .B(n26241), .Z(n26239) );
  XOR U28018 ( .A(nreg[750]), .B(n26238), .Z(n26241) );
  XNOR U28019 ( .A(n15603), .B(n26238), .Z(n26240) );
  XOR U28020 ( .A(n26242), .B(n26243), .Z(n15603) );
  XOR U28021 ( .A(n26244), .B(n26245), .Z(n26238) );
  AND U28022 ( .A(n26246), .B(n26247), .Z(n26245) );
  XOR U28023 ( .A(nreg[749]), .B(n26244), .Z(n26247) );
  XNOR U28024 ( .A(n15615), .B(n26244), .Z(n26246) );
  XOR U28025 ( .A(n26248), .B(n26249), .Z(n15615) );
  XOR U28026 ( .A(n26250), .B(n26251), .Z(n26244) );
  AND U28027 ( .A(n26252), .B(n26253), .Z(n26251) );
  XOR U28028 ( .A(nreg[748]), .B(n26250), .Z(n26253) );
  XNOR U28029 ( .A(n15627), .B(n26250), .Z(n26252) );
  XOR U28030 ( .A(n26254), .B(n26255), .Z(n15627) );
  XOR U28031 ( .A(n26256), .B(n26257), .Z(n26250) );
  AND U28032 ( .A(n26258), .B(n26259), .Z(n26257) );
  XOR U28033 ( .A(nreg[747]), .B(n26256), .Z(n26259) );
  XNOR U28034 ( .A(n15639), .B(n26256), .Z(n26258) );
  XOR U28035 ( .A(n26260), .B(n26261), .Z(n15639) );
  XOR U28036 ( .A(n26262), .B(n26263), .Z(n26256) );
  AND U28037 ( .A(n26264), .B(n26265), .Z(n26263) );
  XOR U28038 ( .A(nreg[746]), .B(n26262), .Z(n26265) );
  XNOR U28039 ( .A(n15651), .B(n26262), .Z(n26264) );
  XOR U28040 ( .A(n26266), .B(n26267), .Z(n15651) );
  XOR U28041 ( .A(n26268), .B(n26269), .Z(n26262) );
  AND U28042 ( .A(n26270), .B(n26271), .Z(n26269) );
  XOR U28043 ( .A(nreg[745]), .B(n26268), .Z(n26271) );
  XNOR U28044 ( .A(n15663), .B(n26268), .Z(n26270) );
  XOR U28045 ( .A(n26272), .B(n26273), .Z(n15663) );
  XOR U28046 ( .A(n26274), .B(n26275), .Z(n26268) );
  AND U28047 ( .A(n26276), .B(n26277), .Z(n26275) );
  XOR U28048 ( .A(nreg[744]), .B(n26274), .Z(n26277) );
  XNOR U28049 ( .A(n15675), .B(n26274), .Z(n26276) );
  XOR U28050 ( .A(n26278), .B(n26279), .Z(n15675) );
  XOR U28051 ( .A(n26280), .B(n26281), .Z(n26274) );
  AND U28052 ( .A(n26282), .B(n26283), .Z(n26281) );
  XOR U28053 ( .A(nreg[743]), .B(n26280), .Z(n26283) );
  XNOR U28054 ( .A(n15687), .B(n26280), .Z(n26282) );
  XOR U28055 ( .A(n26284), .B(n26285), .Z(n15687) );
  XOR U28056 ( .A(n26286), .B(n26287), .Z(n26280) );
  AND U28057 ( .A(n26288), .B(n26289), .Z(n26287) );
  XOR U28058 ( .A(nreg[742]), .B(n26286), .Z(n26289) );
  XNOR U28059 ( .A(n15699), .B(n26286), .Z(n26288) );
  XOR U28060 ( .A(n26290), .B(n26291), .Z(n15699) );
  XOR U28061 ( .A(n26292), .B(n26293), .Z(n26286) );
  AND U28062 ( .A(n26294), .B(n26295), .Z(n26293) );
  XOR U28063 ( .A(nreg[741]), .B(n26292), .Z(n26295) );
  XNOR U28064 ( .A(n15711), .B(n26292), .Z(n26294) );
  XOR U28065 ( .A(n26296), .B(n26297), .Z(n15711) );
  XOR U28066 ( .A(n26298), .B(n26299), .Z(n26292) );
  AND U28067 ( .A(n26300), .B(n26301), .Z(n26299) );
  XOR U28068 ( .A(nreg[740]), .B(n26298), .Z(n26301) );
  XNOR U28069 ( .A(n15723), .B(n26298), .Z(n26300) );
  XOR U28070 ( .A(n26302), .B(n26303), .Z(n15723) );
  XOR U28071 ( .A(n26304), .B(n26305), .Z(n26298) );
  AND U28072 ( .A(n26306), .B(n26307), .Z(n26305) );
  XOR U28073 ( .A(nreg[739]), .B(n26304), .Z(n26307) );
  XNOR U28074 ( .A(n15735), .B(n26304), .Z(n26306) );
  XOR U28075 ( .A(n26308), .B(n26309), .Z(n15735) );
  XOR U28076 ( .A(n26310), .B(n26311), .Z(n26304) );
  AND U28077 ( .A(n26312), .B(n26313), .Z(n26311) );
  XOR U28078 ( .A(nreg[738]), .B(n26310), .Z(n26313) );
  XNOR U28079 ( .A(n15747), .B(n26310), .Z(n26312) );
  XOR U28080 ( .A(n26314), .B(n26315), .Z(n15747) );
  XOR U28081 ( .A(n26316), .B(n26317), .Z(n26310) );
  AND U28082 ( .A(n26318), .B(n26319), .Z(n26317) );
  XOR U28083 ( .A(nreg[737]), .B(n26316), .Z(n26319) );
  XNOR U28084 ( .A(n15759), .B(n26316), .Z(n26318) );
  XOR U28085 ( .A(n26320), .B(n26321), .Z(n15759) );
  XOR U28086 ( .A(n26322), .B(n26323), .Z(n26316) );
  AND U28087 ( .A(n26324), .B(n26325), .Z(n26323) );
  XOR U28088 ( .A(nreg[736]), .B(n26322), .Z(n26325) );
  XNOR U28089 ( .A(n15771), .B(n26322), .Z(n26324) );
  XOR U28090 ( .A(n26326), .B(n26327), .Z(n15771) );
  XOR U28091 ( .A(n26328), .B(n26329), .Z(n26322) );
  AND U28092 ( .A(n26330), .B(n26331), .Z(n26329) );
  XOR U28093 ( .A(nreg[735]), .B(n26328), .Z(n26331) );
  XNOR U28094 ( .A(n15783), .B(n26328), .Z(n26330) );
  XOR U28095 ( .A(n26332), .B(n26333), .Z(n15783) );
  XOR U28096 ( .A(n26334), .B(n26335), .Z(n26328) );
  AND U28097 ( .A(n26336), .B(n26337), .Z(n26335) );
  XOR U28098 ( .A(nreg[734]), .B(n26334), .Z(n26337) );
  XNOR U28099 ( .A(n15795), .B(n26334), .Z(n26336) );
  XOR U28100 ( .A(n26338), .B(n26339), .Z(n15795) );
  XOR U28101 ( .A(n26340), .B(n26341), .Z(n26334) );
  AND U28102 ( .A(n26342), .B(n26343), .Z(n26341) );
  XOR U28103 ( .A(nreg[733]), .B(n26340), .Z(n26343) );
  XNOR U28104 ( .A(n15807), .B(n26340), .Z(n26342) );
  XOR U28105 ( .A(n26344), .B(n26345), .Z(n15807) );
  XOR U28106 ( .A(n26346), .B(n26347), .Z(n26340) );
  AND U28107 ( .A(n26348), .B(n26349), .Z(n26347) );
  XOR U28108 ( .A(nreg[732]), .B(n26346), .Z(n26349) );
  XNOR U28109 ( .A(n15819), .B(n26346), .Z(n26348) );
  XOR U28110 ( .A(n26350), .B(n26351), .Z(n15819) );
  XOR U28111 ( .A(n26352), .B(n26353), .Z(n26346) );
  AND U28112 ( .A(n26354), .B(n26355), .Z(n26353) );
  XOR U28113 ( .A(nreg[731]), .B(n26352), .Z(n26355) );
  XNOR U28114 ( .A(n15831), .B(n26352), .Z(n26354) );
  XOR U28115 ( .A(n26356), .B(n26357), .Z(n15831) );
  XOR U28116 ( .A(n26358), .B(n26359), .Z(n26352) );
  AND U28117 ( .A(n26360), .B(n26361), .Z(n26359) );
  XOR U28118 ( .A(nreg[730]), .B(n26358), .Z(n26361) );
  XNOR U28119 ( .A(n15843), .B(n26358), .Z(n26360) );
  XOR U28120 ( .A(n26362), .B(n26363), .Z(n15843) );
  XOR U28121 ( .A(n26364), .B(n26365), .Z(n26358) );
  AND U28122 ( .A(n26366), .B(n26367), .Z(n26365) );
  XOR U28123 ( .A(nreg[729]), .B(n26364), .Z(n26367) );
  XNOR U28124 ( .A(n15855), .B(n26364), .Z(n26366) );
  XOR U28125 ( .A(n26368), .B(n26369), .Z(n15855) );
  XOR U28126 ( .A(n26370), .B(n26371), .Z(n26364) );
  AND U28127 ( .A(n26372), .B(n26373), .Z(n26371) );
  XOR U28128 ( .A(nreg[728]), .B(n26370), .Z(n26373) );
  XNOR U28129 ( .A(n15867), .B(n26370), .Z(n26372) );
  XOR U28130 ( .A(n26374), .B(n26375), .Z(n15867) );
  XOR U28131 ( .A(n26376), .B(n26377), .Z(n26370) );
  AND U28132 ( .A(n26378), .B(n26379), .Z(n26377) );
  XOR U28133 ( .A(nreg[727]), .B(n26376), .Z(n26379) );
  XNOR U28134 ( .A(n15879), .B(n26376), .Z(n26378) );
  XOR U28135 ( .A(n26380), .B(n26381), .Z(n15879) );
  XOR U28136 ( .A(n26382), .B(n26383), .Z(n26376) );
  AND U28137 ( .A(n26384), .B(n26385), .Z(n26383) );
  XOR U28138 ( .A(nreg[726]), .B(n26382), .Z(n26385) );
  XNOR U28139 ( .A(n15891), .B(n26382), .Z(n26384) );
  XOR U28140 ( .A(n26386), .B(n26387), .Z(n15891) );
  XOR U28141 ( .A(n26388), .B(n26389), .Z(n26382) );
  AND U28142 ( .A(n26390), .B(n26391), .Z(n26389) );
  XOR U28143 ( .A(nreg[725]), .B(n26388), .Z(n26391) );
  XNOR U28144 ( .A(n15903), .B(n26388), .Z(n26390) );
  XOR U28145 ( .A(n26392), .B(n26393), .Z(n15903) );
  XOR U28146 ( .A(n26394), .B(n26395), .Z(n26388) );
  AND U28147 ( .A(n26396), .B(n26397), .Z(n26395) );
  XOR U28148 ( .A(nreg[724]), .B(n26394), .Z(n26397) );
  XNOR U28149 ( .A(n15915), .B(n26394), .Z(n26396) );
  XOR U28150 ( .A(n26398), .B(n26399), .Z(n15915) );
  XOR U28151 ( .A(n26400), .B(n26401), .Z(n26394) );
  AND U28152 ( .A(n26402), .B(n26403), .Z(n26401) );
  XOR U28153 ( .A(nreg[723]), .B(n26400), .Z(n26403) );
  XNOR U28154 ( .A(n15927), .B(n26400), .Z(n26402) );
  XOR U28155 ( .A(n26404), .B(n26405), .Z(n15927) );
  XOR U28156 ( .A(n26406), .B(n26407), .Z(n26400) );
  AND U28157 ( .A(n26408), .B(n26409), .Z(n26407) );
  XOR U28158 ( .A(nreg[722]), .B(n26406), .Z(n26409) );
  XNOR U28159 ( .A(n15939), .B(n26406), .Z(n26408) );
  XOR U28160 ( .A(n26410), .B(n26411), .Z(n15939) );
  XOR U28161 ( .A(n26412), .B(n26413), .Z(n26406) );
  AND U28162 ( .A(n26414), .B(n26415), .Z(n26413) );
  XOR U28163 ( .A(nreg[721]), .B(n26412), .Z(n26415) );
  XNOR U28164 ( .A(n15951), .B(n26412), .Z(n26414) );
  XOR U28165 ( .A(n26416), .B(n26417), .Z(n15951) );
  XOR U28166 ( .A(n26418), .B(n26419), .Z(n26412) );
  AND U28167 ( .A(n26420), .B(n26421), .Z(n26419) );
  XOR U28168 ( .A(nreg[720]), .B(n26418), .Z(n26421) );
  XNOR U28169 ( .A(n15963), .B(n26418), .Z(n26420) );
  XOR U28170 ( .A(n26422), .B(n26423), .Z(n15963) );
  XOR U28171 ( .A(n26424), .B(n26425), .Z(n26418) );
  AND U28172 ( .A(n26426), .B(n26427), .Z(n26425) );
  XOR U28173 ( .A(nreg[719]), .B(n26424), .Z(n26427) );
  XNOR U28174 ( .A(n15975), .B(n26424), .Z(n26426) );
  XOR U28175 ( .A(n26428), .B(n26429), .Z(n15975) );
  XOR U28176 ( .A(n26430), .B(n26431), .Z(n26424) );
  AND U28177 ( .A(n26432), .B(n26433), .Z(n26431) );
  XOR U28178 ( .A(nreg[718]), .B(n26430), .Z(n26433) );
  XNOR U28179 ( .A(n15987), .B(n26430), .Z(n26432) );
  XOR U28180 ( .A(n26434), .B(n26435), .Z(n15987) );
  XOR U28181 ( .A(n26436), .B(n26437), .Z(n26430) );
  AND U28182 ( .A(n26438), .B(n26439), .Z(n26437) );
  XOR U28183 ( .A(nreg[717]), .B(n26436), .Z(n26439) );
  XNOR U28184 ( .A(n15999), .B(n26436), .Z(n26438) );
  XOR U28185 ( .A(n26440), .B(n26441), .Z(n15999) );
  XOR U28186 ( .A(n26442), .B(n26443), .Z(n26436) );
  AND U28187 ( .A(n26444), .B(n26445), .Z(n26443) );
  XOR U28188 ( .A(nreg[716]), .B(n26442), .Z(n26445) );
  XNOR U28189 ( .A(n16011), .B(n26442), .Z(n26444) );
  XOR U28190 ( .A(n26446), .B(n26447), .Z(n16011) );
  XOR U28191 ( .A(n26448), .B(n26449), .Z(n26442) );
  AND U28192 ( .A(n26450), .B(n26451), .Z(n26449) );
  XOR U28193 ( .A(nreg[715]), .B(n26448), .Z(n26451) );
  XNOR U28194 ( .A(n16023), .B(n26448), .Z(n26450) );
  XOR U28195 ( .A(n26452), .B(n26453), .Z(n16023) );
  XOR U28196 ( .A(n26454), .B(n26455), .Z(n26448) );
  AND U28197 ( .A(n26456), .B(n26457), .Z(n26455) );
  XOR U28198 ( .A(nreg[714]), .B(n26454), .Z(n26457) );
  XNOR U28199 ( .A(n16035), .B(n26454), .Z(n26456) );
  XOR U28200 ( .A(n26458), .B(n26459), .Z(n16035) );
  XOR U28201 ( .A(n26460), .B(n26461), .Z(n26454) );
  AND U28202 ( .A(n26462), .B(n26463), .Z(n26461) );
  XOR U28203 ( .A(nreg[713]), .B(n26460), .Z(n26463) );
  XNOR U28204 ( .A(n16047), .B(n26460), .Z(n26462) );
  XOR U28205 ( .A(n26464), .B(n26465), .Z(n16047) );
  XOR U28206 ( .A(n26466), .B(n26467), .Z(n26460) );
  AND U28207 ( .A(n26468), .B(n26469), .Z(n26467) );
  XOR U28208 ( .A(nreg[712]), .B(n26466), .Z(n26469) );
  XNOR U28209 ( .A(n16059), .B(n26466), .Z(n26468) );
  XOR U28210 ( .A(n26470), .B(n26471), .Z(n16059) );
  XOR U28211 ( .A(n26472), .B(n26473), .Z(n26466) );
  AND U28212 ( .A(n26474), .B(n26475), .Z(n26473) );
  XOR U28213 ( .A(nreg[711]), .B(n26472), .Z(n26475) );
  XNOR U28214 ( .A(n16071), .B(n26472), .Z(n26474) );
  XOR U28215 ( .A(n26476), .B(n26477), .Z(n16071) );
  XOR U28216 ( .A(n26478), .B(n26479), .Z(n26472) );
  AND U28217 ( .A(n26480), .B(n26481), .Z(n26479) );
  XOR U28218 ( .A(nreg[710]), .B(n26478), .Z(n26481) );
  XNOR U28219 ( .A(n16083), .B(n26478), .Z(n26480) );
  XOR U28220 ( .A(n26482), .B(n26483), .Z(n16083) );
  XOR U28221 ( .A(n26484), .B(n26485), .Z(n26478) );
  AND U28222 ( .A(n26486), .B(n26487), .Z(n26485) );
  XOR U28223 ( .A(nreg[709]), .B(n26484), .Z(n26487) );
  XNOR U28224 ( .A(n16095), .B(n26484), .Z(n26486) );
  XOR U28225 ( .A(n26488), .B(n26489), .Z(n16095) );
  XOR U28226 ( .A(n26490), .B(n26491), .Z(n26484) );
  AND U28227 ( .A(n26492), .B(n26493), .Z(n26491) );
  XOR U28228 ( .A(nreg[708]), .B(n26490), .Z(n26493) );
  XNOR U28229 ( .A(n16107), .B(n26490), .Z(n26492) );
  XOR U28230 ( .A(n26494), .B(n26495), .Z(n16107) );
  XOR U28231 ( .A(n26496), .B(n26497), .Z(n26490) );
  AND U28232 ( .A(n26498), .B(n26499), .Z(n26497) );
  XOR U28233 ( .A(nreg[707]), .B(n26496), .Z(n26499) );
  XNOR U28234 ( .A(n16119), .B(n26496), .Z(n26498) );
  XOR U28235 ( .A(n26500), .B(n26501), .Z(n16119) );
  XOR U28236 ( .A(n26502), .B(n26503), .Z(n26496) );
  AND U28237 ( .A(n26504), .B(n26505), .Z(n26503) );
  XOR U28238 ( .A(nreg[706]), .B(n26502), .Z(n26505) );
  XNOR U28239 ( .A(n16131), .B(n26502), .Z(n26504) );
  XOR U28240 ( .A(n26506), .B(n26507), .Z(n16131) );
  XOR U28241 ( .A(n26508), .B(n26509), .Z(n26502) );
  AND U28242 ( .A(n26510), .B(n26511), .Z(n26509) );
  XOR U28243 ( .A(nreg[705]), .B(n26508), .Z(n26511) );
  XNOR U28244 ( .A(n16143), .B(n26508), .Z(n26510) );
  XOR U28245 ( .A(n26512), .B(n26513), .Z(n16143) );
  XOR U28246 ( .A(n26514), .B(n26515), .Z(n26508) );
  AND U28247 ( .A(n26516), .B(n26517), .Z(n26515) );
  XOR U28248 ( .A(nreg[704]), .B(n26514), .Z(n26517) );
  XNOR U28249 ( .A(n16155), .B(n26514), .Z(n26516) );
  XOR U28250 ( .A(n26518), .B(n26519), .Z(n16155) );
  XOR U28251 ( .A(n26520), .B(n26521), .Z(n26514) );
  AND U28252 ( .A(n26522), .B(n26523), .Z(n26521) );
  XOR U28253 ( .A(nreg[703]), .B(n26520), .Z(n26523) );
  XNOR U28254 ( .A(n16167), .B(n26520), .Z(n26522) );
  XOR U28255 ( .A(n26524), .B(n26525), .Z(n16167) );
  XOR U28256 ( .A(n26526), .B(n26527), .Z(n26520) );
  AND U28257 ( .A(n26528), .B(n26529), .Z(n26527) );
  XOR U28258 ( .A(nreg[702]), .B(n26526), .Z(n26529) );
  XNOR U28259 ( .A(n16179), .B(n26526), .Z(n26528) );
  XOR U28260 ( .A(n26530), .B(n26531), .Z(n16179) );
  XOR U28261 ( .A(n26532), .B(n26533), .Z(n26526) );
  AND U28262 ( .A(n26534), .B(n26535), .Z(n26533) );
  XOR U28263 ( .A(nreg[701]), .B(n26532), .Z(n26535) );
  XNOR U28264 ( .A(n16191), .B(n26532), .Z(n26534) );
  XOR U28265 ( .A(n26536), .B(n26537), .Z(n16191) );
  XOR U28266 ( .A(n26538), .B(n26539), .Z(n26532) );
  AND U28267 ( .A(n26540), .B(n26541), .Z(n26539) );
  XOR U28268 ( .A(nreg[700]), .B(n26538), .Z(n26541) );
  XNOR U28269 ( .A(n16203), .B(n26538), .Z(n26540) );
  XOR U28270 ( .A(n26542), .B(n26543), .Z(n16203) );
  XOR U28271 ( .A(n26544), .B(n26545), .Z(n26538) );
  AND U28272 ( .A(n26546), .B(n26547), .Z(n26545) );
  XOR U28273 ( .A(nreg[699]), .B(n26544), .Z(n26547) );
  XNOR U28274 ( .A(n16215), .B(n26544), .Z(n26546) );
  XOR U28275 ( .A(n26548), .B(n26549), .Z(n16215) );
  XOR U28276 ( .A(n26550), .B(n26551), .Z(n26544) );
  AND U28277 ( .A(n26552), .B(n26553), .Z(n26551) );
  XOR U28278 ( .A(nreg[698]), .B(n26550), .Z(n26553) );
  XNOR U28279 ( .A(n16227), .B(n26550), .Z(n26552) );
  XOR U28280 ( .A(n26554), .B(n26555), .Z(n16227) );
  XOR U28281 ( .A(n26556), .B(n26557), .Z(n26550) );
  AND U28282 ( .A(n26558), .B(n26559), .Z(n26557) );
  XOR U28283 ( .A(nreg[697]), .B(n26556), .Z(n26559) );
  XNOR U28284 ( .A(n16239), .B(n26556), .Z(n26558) );
  XOR U28285 ( .A(n26560), .B(n26561), .Z(n16239) );
  XOR U28286 ( .A(n26562), .B(n26563), .Z(n26556) );
  AND U28287 ( .A(n26564), .B(n26565), .Z(n26563) );
  XOR U28288 ( .A(nreg[696]), .B(n26562), .Z(n26565) );
  XNOR U28289 ( .A(n16251), .B(n26562), .Z(n26564) );
  XOR U28290 ( .A(n26566), .B(n26567), .Z(n16251) );
  XOR U28291 ( .A(n26568), .B(n26569), .Z(n26562) );
  AND U28292 ( .A(n26570), .B(n26571), .Z(n26569) );
  XOR U28293 ( .A(nreg[695]), .B(n26568), .Z(n26571) );
  XNOR U28294 ( .A(n16263), .B(n26568), .Z(n26570) );
  XOR U28295 ( .A(n26572), .B(n26573), .Z(n16263) );
  XOR U28296 ( .A(n26574), .B(n26575), .Z(n26568) );
  AND U28297 ( .A(n26576), .B(n26577), .Z(n26575) );
  XOR U28298 ( .A(nreg[694]), .B(n26574), .Z(n26577) );
  XNOR U28299 ( .A(n16275), .B(n26574), .Z(n26576) );
  XOR U28300 ( .A(n26578), .B(n26579), .Z(n16275) );
  XOR U28301 ( .A(n26580), .B(n26581), .Z(n26574) );
  AND U28302 ( .A(n26582), .B(n26583), .Z(n26581) );
  XOR U28303 ( .A(nreg[693]), .B(n26580), .Z(n26583) );
  XNOR U28304 ( .A(n16287), .B(n26580), .Z(n26582) );
  XOR U28305 ( .A(n26584), .B(n26585), .Z(n16287) );
  XOR U28306 ( .A(n26586), .B(n26587), .Z(n26580) );
  AND U28307 ( .A(n26588), .B(n26589), .Z(n26587) );
  XOR U28308 ( .A(nreg[692]), .B(n26586), .Z(n26589) );
  XNOR U28309 ( .A(n16299), .B(n26586), .Z(n26588) );
  XOR U28310 ( .A(n26590), .B(n26591), .Z(n16299) );
  XOR U28311 ( .A(n26592), .B(n26593), .Z(n26586) );
  AND U28312 ( .A(n26594), .B(n26595), .Z(n26593) );
  XOR U28313 ( .A(nreg[691]), .B(n26592), .Z(n26595) );
  XNOR U28314 ( .A(n16311), .B(n26592), .Z(n26594) );
  XOR U28315 ( .A(n26596), .B(n26597), .Z(n16311) );
  XOR U28316 ( .A(n26598), .B(n26599), .Z(n26592) );
  AND U28317 ( .A(n26600), .B(n26601), .Z(n26599) );
  XOR U28318 ( .A(nreg[690]), .B(n26598), .Z(n26601) );
  XNOR U28319 ( .A(n16323), .B(n26598), .Z(n26600) );
  XOR U28320 ( .A(n26602), .B(n26603), .Z(n16323) );
  XOR U28321 ( .A(n26604), .B(n26605), .Z(n26598) );
  AND U28322 ( .A(n26606), .B(n26607), .Z(n26605) );
  XOR U28323 ( .A(nreg[689]), .B(n26604), .Z(n26607) );
  XNOR U28324 ( .A(n16335), .B(n26604), .Z(n26606) );
  XOR U28325 ( .A(n26608), .B(n26609), .Z(n16335) );
  XOR U28326 ( .A(n26610), .B(n26611), .Z(n26604) );
  AND U28327 ( .A(n26612), .B(n26613), .Z(n26611) );
  XOR U28328 ( .A(nreg[688]), .B(n26610), .Z(n26613) );
  XNOR U28329 ( .A(n16347), .B(n26610), .Z(n26612) );
  XOR U28330 ( .A(n26614), .B(n26615), .Z(n16347) );
  XOR U28331 ( .A(n26616), .B(n26617), .Z(n26610) );
  AND U28332 ( .A(n26618), .B(n26619), .Z(n26617) );
  XOR U28333 ( .A(nreg[687]), .B(n26616), .Z(n26619) );
  XNOR U28334 ( .A(n16359), .B(n26616), .Z(n26618) );
  XOR U28335 ( .A(n26620), .B(n26621), .Z(n16359) );
  XOR U28336 ( .A(n26622), .B(n26623), .Z(n26616) );
  AND U28337 ( .A(n26624), .B(n26625), .Z(n26623) );
  XOR U28338 ( .A(nreg[686]), .B(n26622), .Z(n26625) );
  XNOR U28339 ( .A(n16371), .B(n26622), .Z(n26624) );
  XOR U28340 ( .A(n26626), .B(n26627), .Z(n16371) );
  XOR U28341 ( .A(n26628), .B(n26629), .Z(n26622) );
  AND U28342 ( .A(n26630), .B(n26631), .Z(n26629) );
  XOR U28343 ( .A(nreg[685]), .B(n26628), .Z(n26631) );
  XNOR U28344 ( .A(n16383), .B(n26628), .Z(n26630) );
  XOR U28345 ( .A(n26632), .B(n26633), .Z(n16383) );
  XOR U28346 ( .A(n26634), .B(n26635), .Z(n26628) );
  AND U28347 ( .A(n26636), .B(n26637), .Z(n26635) );
  XOR U28348 ( .A(nreg[684]), .B(n26634), .Z(n26637) );
  XNOR U28349 ( .A(n16395), .B(n26634), .Z(n26636) );
  XOR U28350 ( .A(n26638), .B(n26639), .Z(n16395) );
  XOR U28351 ( .A(n26640), .B(n26641), .Z(n26634) );
  AND U28352 ( .A(n26642), .B(n26643), .Z(n26641) );
  XOR U28353 ( .A(nreg[683]), .B(n26640), .Z(n26643) );
  XNOR U28354 ( .A(n16407), .B(n26640), .Z(n26642) );
  XOR U28355 ( .A(n26644), .B(n26645), .Z(n16407) );
  XOR U28356 ( .A(n26646), .B(n26647), .Z(n26640) );
  AND U28357 ( .A(n26648), .B(n26649), .Z(n26647) );
  XOR U28358 ( .A(nreg[682]), .B(n26646), .Z(n26649) );
  XNOR U28359 ( .A(n16419), .B(n26646), .Z(n26648) );
  XOR U28360 ( .A(n26650), .B(n26651), .Z(n16419) );
  XOR U28361 ( .A(n26652), .B(n26653), .Z(n26646) );
  AND U28362 ( .A(n26654), .B(n26655), .Z(n26653) );
  XOR U28363 ( .A(nreg[681]), .B(n26652), .Z(n26655) );
  XNOR U28364 ( .A(n16431), .B(n26652), .Z(n26654) );
  XOR U28365 ( .A(n26656), .B(n26657), .Z(n16431) );
  XOR U28366 ( .A(n26658), .B(n26659), .Z(n26652) );
  AND U28367 ( .A(n26660), .B(n26661), .Z(n26659) );
  XOR U28368 ( .A(nreg[680]), .B(n26658), .Z(n26661) );
  XNOR U28369 ( .A(n16443), .B(n26658), .Z(n26660) );
  XOR U28370 ( .A(n26662), .B(n26663), .Z(n16443) );
  XOR U28371 ( .A(n26664), .B(n26665), .Z(n26658) );
  AND U28372 ( .A(n26666), .B(n26667), .Z(n26665) );
  XOR U28373 ( .A(nreg[679]), .B(n26664), .Z(n26667) );
  XNOR U28374 ( .A(n16455), .B(n26664), .Z(n26666) );
  XOR U28375 ( .A(n26668), .B(n26669), .Z(n16455) );
  XOR U28376 ( .A(n26670), .B(n26671), .Z(n26664) );
  AND U28377 ( .A(n26672), .B(n26673), .Z(n26671) );
  XOR U28378 ( .A(nreg[678]), .B(n26670), .Z(n26673) );
  XNOR U28379 ( .A(n16467), .B(n26670), .Z(n26672) );
  XOR U28380 ( .A(n26674), .B(n26675), .Z(n16467) );
  XOR U28381 ( .A(n26676), .B(n26677), .Z(n26670) );
  AND U28382 ( .A(n26678), .B(n26679), .Z(n26677) );
  XOR U28383 ( .A(nreg[677]), .B(n26676), .Z(n26679) );
  XNOR U28384 ( .A(n16479), .B(n26676), .Z(n26678) );
  XOR U28385 ( .A(n26680), .B(n26681), .Z(n16479) );
  XOR U28386 ( .A(n26682), .B(n26683), .Z(n26676) );
  AND U28387 ( .A(n26684), .B(n26685), .Z(n26683) );
  XOR U28388 ( .A(nreg[676]), .B(n26682), .Z(n26685) );
  XNOR U28389 ( .A(n16491), .B(n26682), .Z(n26684) );
  XOR U28390 ( .A(n26686), .B(n26687), .Z(n16491) );
  XOR U28391 ( .A(n26688), .B(n26689), .Z(n26682) );
  AND U28392 ( .A(n26690), .B(n26691), .Z(n26689) );
  XOR U28393 ( .A(nreg[675]), .B(n26688), .Z(n26691) );
  XNOR U28394 ( .A(n16503), .B(n26688), .Z(n26690) );
  XOR U28395 ( .A(n26692), .B(n26693), .Z(n16503) );
  XOR U28396 ( .A(n26694), .B(n26695), .Z(n26688) );
  AND U28397 ( .A(n26696), .B(n26697), .Z(n26695) );
  XOR U28398 ( .A(nreg[674]), .B(n26694), .Z(n26697) );
  XNOR U28399 ( .A(n16515), .B(n26694), .Z(n26696) );
  XOR U28400 ( .A(n26698), .B(n26699), .Z(n16515) );
  XOR U28401 ( .A(n26700), .B(n26701), .Z(n26694) );
  AND U28402 ( .A(n26702), .B(n26703), .Z(n26701) );
  XOR U28403 ( .A(nreg[673]), .B(n26700), .Z(n26703) );
  XNOR U28404 ( .A(n16527), .B(n26700), .Z(n26702) );
  XOR U28405 ( .A(n26704), .B(n26705), .Z(n16527) );
  XOR U28406 ( .A(n26706), .B(n26707), .Z(n26700) );
  AND U28407 ( .A(n26708), .B(n26709), .Z(n26707) );
  XOR U28408 ( .A(nreg[672]), .B(n26706), .Z(n26709) );
  XNOR U28409 ( .A(n16539), .B(n26706), .Z(n26708) );
  XOR U28410 ( .A(n26710), .B(n26711), .Z(n16539) );
  XOR U28411 ( .A(n26712), .B(n26713), .Z(n26706) );
  AND U28412 ( .A(n26714), .B(n26715), .Z(n26713) );
  XOR U28413 ( .A(nreg[671]), .B(n26712), .Z(n26715) );
  XNOR U28414 ( .A(n16551), .B(n26712), .Z(n26714) );
  XOR U28415 ( .A(n26716), .B(n26717), .Z(n16551) );
  XOR U28416 ( .A(n26718), .B(n26719), .Z(n26712) );
  AND U28417 ( .A(n26720), .B(n26721), .Z(n26719) );
  XOR U28418 ( .A(nreg[670]), .B(n26718), .Z(n26721) );
  XNOR U28419 ( .A(n16563), .B(n26718), .Z(n26720) );
  XOR U28420 ( .A(n26722), .B(n26723), .Z(n16563) );
  XOR U28421 ( .A(n26724), .B(n26725), .Z(n26718) );
  AND U28422 ( .A(n26726), .B(n26727), .Z(n26725) );
  XOR U28423 ( .A(nreg[669]), .B(n26724), .Z(n26727) );
  XNOR U28424 ( .A(n16575), .B(n26724), .Z(n26726) );
  XOR U28425 ( .A(n26728), .B(n26729), .Z(n16575) );
  XOR U28426 ( .A(n26730), .B(n26731), .Z(n26724) );
  AND U28427 ( .A(n26732), .B(n26733), .Z(n26731) );
  XOR U28428 ( .A(nreg[668]), .B(n26730), .Z(n26733) );
  XNOR U28429 ( .A(n16587), .B(n26730), .Z(n26732) );
  XOR U28430 ( .A(n26734), .B(n26735), .Z(n16587) );
  XOR U28431 ( .A(n26736), .B(n26737), .Z(n26730) );
  AND U28432 ( .A(n26738), .B(n26739), .Z(n26737) );
  XOR U28433 ( .A(nreg[667]), .B(n26736), .Z(n26739) );
  XNOR U28434 ( .A(n16599), .B(n26736), .Z(n26738) );
  XOR U28435 ( .A(n26740), .B(n26741), .Z(n16599) );
  XOR U28436 ( .A(n26742), .B(n26743), .Z(n26736) );
  AND U28437 ( .A(n26744), .B(n26745), .Z(n26743) );
  XOR U28438 ( .A(nreg[666]), .B(n26742), .Z(n26745) );
  XNOR U28439 ( .A(n16611), .B(n26742), .Z(n26744) );
  XOR U28440 ( .A(n26746), .B(n26747), .Z(n16611) );
  XOR U28441 ( .A(n26748), .B(n26749), .Z(n26742) );
  AND U28442 ( .A(n26750), .B(n26751), .Z(n26749) );
  XOR U28443 ( .A(nreg[665]), .B(n26748), .Z(n26751) );
  XNOR U28444 ( .A(n16623), .B(n26748), .Z(n26750) );
  XOR U28445 ( .A(n26752), .B(n26753), .Z(n16623) );
  XOR U28446 ( .A(n26754), .B(n26755), .Z(n26748) );
  AND U28447 ( .A(n26756), .B(n26757), .Z(n26755) );
  XOR U28448 ( .A(nreg[664]), .B(n26754), .Z(n26757) );
  XNOR U28449 ( .A(n16635), .B(n26754), .Z(n26756) );
  XOR U28450 ( .A(n26758), .B(n26759), .Z(n16635) );
  XOR U28451 ( .A(n26760), .B(n26761), .Z(n26754) );
  AND U28452 ( .A(n26762), .B(n26763), .Z(n26761) );
  XOR U28453 ( .A(nreg[663]), .B(n26760), .Z(n26763) );
  XNOR U28454 ( .A(n16647), .B(n26760), .Z(n26762) );
  XOR U28455 ( .A(n26764), .B(n26765), .Z(n16647) );
  XOR U28456 ( .A(n26766), .B(n26767), .Z(n26760) );
  AND U28457 ( .A(n26768), .B(n26769), .Z(n26767) );
  XOR U28458 ( .A(nreg[662]), .B(n26766), .Z(n26769) );
  XNOR U28459 ( .A(n16659), .B(n26766), .Z(n26768) );
  XOR U28460 ( .A(n26770), .B(n26771), .Z(n16659) );
  XOR U28461 ( .A(n26772), .B(n26773), .Z(n26766) );
  AND U28462 ( .A(n26774), .B(n26775), .Z(n26773) );
  XOR U28463 ( .A(nreg[661]), .B(n26772), .Z(n26775) );
  XNOR U28464 ( .A(n16671), .B(n26772), .Z(n26774) );
  XOR U28465 ( .A(n26776), .B(n26777), .Z(n16671) );
  XOR U28466 ( .A(n26778), .B(n26779), .Z(n26772) );
  AND U28467 ( .A(n26780), .B(n26781), .Z(n26779) );
  XOR U28468 ( .A(nreg[660]), .B(n26778), .Z(n26781) );
  XNOR U28469 ( .A(n16683), .B(n26778), .Z(n26780) );
  XOR U28470 ( .A(n26782), .B(n26783), .Z(n16683) );
  XOR U28471 ( .A(n26784), .B(n26785), .Z(n26778) );
  AND U28472 ( .A(n26786), .B(n26787), .Z(n26785) );
  XOR U28473 ( .A(nreg[659]), .B(n26784), .Z(n26787) );
  XNOR U28474 ( .A(n16695), .B(n26784), .Z(n26786) );
  XOR U28475 ( .A(n26788), .B(n26789), .Z(n16695) );
  XOR U28476 ( .A(n26790), .B(n26791), .Z(n26784) );
  AND U28477 ( .A(n26792), .B(n26793), .Z(n26791) );
  XOR U28478 ( .A(nreg[658]), .B(n26790), .Z(n26793) );
  XNOR U28479 ( .A(n16707), .B(n26790), .Z(n26792) );
  XOR U28480 ( .A(n26794), .B(n26795), .Z(n16707) );
  XOR U28481 ( .A(n26796), .B(n26797), .Z(n26790) );
  AND U28482 ( .A(n26798), .B(n26799), .Z(n26797) );
  XOR U28483 ( .A(nreg[657]), .B(n26796), .Z(n26799) );
  XNOR U28484 ( .A(n16719), .B(n26796), .Z(n26798) );
  XOR U28485 ( .A(n26800), .B(n26801), .Z(n16719) );
  XOR U28486 ( .A(n26802), .B(n26803), .Z(n26796) );
  AND U28487 ( .A(n26804), .B(n26805), .Z(n26803) );
  XOR U28488 ( .A(nreg[656]), .B(n26802), .Z(n26805) );
  XNOR U28489 ( .A(n16731), .B(n26802), .Z(n26804) );
  XOR U28490 ( .A(n26806), .B(n26807), .Z(n16731) );
  XOR U28491 ( .A(n26808), .B(n26809), .Z(n26802) );
  AND U28492 ( .A(n26810), .B(n26811), .Z(n26809) );
  XOR U28493 ( .A(nreg[655]), .B(n26808), .Z(n26811) );
  XNOR U28494 ( .A(n16743), .B(n26808), .Z(n26810) );
  XOR U28495 ( .A(n26812), .B(n26813), .Z(n16743) );
  XOR U28496 ( .A(n26814), .B(n26815), .Z(n26808) );
  AND U28497 ( .A(n26816), .B(n26817), .Z(n26815) );
  XOR U28498 ( .A(nreg[654]), .B(n26814), .Z(n26817) );
  XNOR U28499 ( .A(n16755), .B(n26814), .Z(n26816) );
  XOR U28500 ( .A(n26818), .B(n26819), .Z(n16755) );
  XOR U28501 ( .A(n26820), .B(n26821), .Z(n26814) );
  AND U28502 ( .A(n26822), .B(n26823), .Z(n26821) );
  XOR U28503 ( .A(nreg[653]), .B(n26820), .Z(n26823) );
  XNOR U28504 ( .A(n16767), .B(n26820), .Z(n26822) );
  XOR U28505 ( .A(n26824), .B(n26825), .Z(n16767) );
  XOR U28506 ( .A(n26826), .B(n26827), .Z(n26820) );
  AND U28507 ( .A(n26828), .B(n26829), .Z(n26827) );
  XOR U28508 ( .A(nreg[652]), .B(n26826), .Z(n26829) );
  XNOR U28509 ( .A(n16779), .B(n26826), .Z(n26828) );
  XOR U28510 ( .A(n26830), .B(n26831), .Z(n16779) );
  XOR U28511 ( .A(n26832), .B(n26833), .Z(n26826) );
  AND U28512 ( .A(n26834), .B(n26835), .Z(n26833) );
  XOR U28513 ( .A(nreg[651]), .B(n26832), .Z(n26835) );
  XNOR U28514 ( .A(n16791), .B(n26832), .Z(n26834) );
  XOR U28515 ( .A(n26836), .B(n26837), .Z(n16791) );
  XOR U28516 ( .A(n26838), .B(n26839), .Z(n26832) );
  AND U28517 ( .A(n26840), .B(n26841), .Z(n26839) );
  XOR U28518 ( .A(nreg[650]), .B(n26838), .Z(n26841) );
  XNOR U28519 ( .A(n16803), .B(n26838), .Z(n26840) );
  XOR U28520 ( .A(n26842), .B(n26843), .Z(n16803) );
  XOR U28521 ( .A(n26844), .B(n26845), .Z(n26838) );
  AND U28522 ( .A(n26846), .B(n26847), .Z(n26845) );
  XOR U28523 ( .A(nreg[649]), .B(n26844), .Z(n26847) );
  XNOR U28524 ( .A(n16815), .B(n26844), .Z(n26846) );
  XOR U28525 ( .A(n26848), .B(n26849), .Z(n16815) );
  XOR U28526 ( .A(n26850), .B(n26851), .Z(n26844) );
  AND U28527 ( .A(n26852), .B(n26853), .Z(n26851) );
  XOR U28528 ( .A(nreg[648]), .B(n26850), .Z(n26853) );
  XNOR U28529 ( .A(n16827), .B(n26850), .Z(n26852) );
  XOR U28530 ( .A(n26854), .B(n26855), .Z(n16827) );
  XOR U28531 ( .A(n26856), .B(n26857), .Z(n26850) );
  AND U28532 ( .A(n26858), .B(n26859), .Z(n26857) );
  XOR U28533 ( .A(nreg[647]), .B(n26856), .Z(n26859) );
  XNOR U28534 ( .A(n16839), .B(n26856), .Z(n26858) );
  XOR U28535 ( .A(n26860), .B(n26861), .Z(n16839) );
  XOR U28536 ( .A(n26862), .B(n26863), .Z(n26856) );
  AND U28537 ( .A(n26864), .B(n26865), .Z(n26863) );
  XOR U28538 ( .A(nreg[646]), .B(n26862), .Z(n26865) );
  XNOR U28539 ( .A(n16851), .B(n26862), .Z(n26864) );
  XOR U28540 ( .A(n26866), .B(n26867), .Z(n16851) );
  XOR U28541 ( .A(n26868), .B(n26869), .Z(n26862) );
  AND U28542 ( .A(n26870), .B(n26871), .Z(n26869) );
  XOR U28543 ( .A(nreg[645]), .B(n26868), .Z(n26871) );
  XNOR U28544 ( .A(n16863), .B(n26868), .Z(n26870) );
  XOR U28545 ( .A(n26872), .B(n26873), .Z(n16863) );
  XOR U28546 ( .A(n26874), .B(n26875), .Z(n26868) );
  AND U28547 ( .A(n26876), .B(n26877), .Z(n26875) );
  XOR U28548 ( .A(nreg[644]), .B(n26874), .Z(n26877) );
  XNOR U28549 ( .A(n16875), .B(n26874), .Z(n26876) );
  XOR U28550 ( .A(n26878), .B(n26879), .Z(n16875) );
  XOR U28551 ( .A(n26880), .B(n26881), .Z(n26874) );
  AND U28552 ( .A(n26882), .B(n26883), .Z(n26881) );
  XOR U28553 ( .A(nreg[643]), .B(n26880), .Z(n26883) );
  XNOR U28554 ( .A(n16887), .B(n26880), .Z(n26882) );
  XOR U28555 ( .A(n26884), .B(n26885), .Z(n16887) );
  XOR U28556 ( .A(n26886), .B(n26887), .Z(n26880) );
  AND U28557 ( .A(n26888), .B(n26889), .Z(n26887) );
  XOR U28558 ( .A(nreg[642]), .B(n26886), .Z(n26889) );
  XNOR U28559 ( .A(n16899), .B(n26886), .Z(n26888) );
  XOR U28560 ( .A(n26890), .B(n26891), .Z(n16899) );
  XOR U28561 ( .A(n26892), .B(n26893), .Z(n26886) );
  AND U28562 ( .A(n26894), .B(n26895), .Z(n26893) );
  XOR U28563 ( .A(nreg[641]), .B(n26892), .Z(n26895) );
  XNOR U28564 ( .A(n16911), .B(n26892), .Z(n26894) );
  XOR U28565 ( .A(n26896), .B(n26897), .Z(n16911) );
  XOR U28566 ( .A(n26898), .B(n26899), .Z(n26892) );
  AND U28567 ( .A(n26900), .B(n26901), .Z(n26899) );
  XOR U28568 ( .A(nreg[640]), .B(n26898), .Z(n26901) );
  XNOR U28569 ( .A(n16923), .B(n26898), .Z(n26900) );
  XOR U28570 ( .A(n26902), .B(n26903), .Z(n16923) );
  XOR U28571 ( .A(n26904), .B(n26905), .Z(n26898) );
  AND U28572 ( .A(n26906), .B(n26907), .Z(n26905) );
  XOR U28573 ( .A(nreg[639]), .B(n26904), .Z(n26907) );
  XNOR U28574 ( .A(n16935), .B(n26904), .Z(n26906) );
  XOR U28575 ( .A(n26908), .B(n26909), .Z(n16935) );
  XOR U28576 ( .A(n26910), .B(n26911), .Z(n26904) );
  AND U28577 ( .A(n26912), .B(n26913), .Z(n26911) );
  XOR U28578 ( .A(nreg[638]), .B(n26910), .Z(n26913) );
  XNOR U28579 ( .A(n16947), .B(n26910), .Z(n26912) );
  XOR U28580 ( .A(n26914), .B(n26915), .Z(n16947) );
  XOR U28581 ( .A(n26916), .B(n26917), .Z(n26910) );
  AND U28582 ( .A(n26918), .B(n26919), .Z(n26917) );
  XOR U28583 ( .A(nreg[637]), .B(n26916), .Z(n26919) );
  XNOR U28584 ( .A(n16959), .B(n26916), .Z(n26918) );
  XOR U28585 ( .A(n26920), .B(n26921), .Z(n16959) );
  XOR U28586 ( .A(n26922), .B(n26923), .Z(n26916) );
  AND U28587 ( .A(n26924), .B(n26925), .Z(n26923) );
  XOR U28588 ( .A(nreg[636]), .B(n26922), .Z(n26925) );
  XNOR U28589 ( .A(n16971), .B(n26922), .Z(n26924) );
  XOR U28590 ( .A(n26926), .B(n26927), .Z(n16971) );
  XOR U28591 ( .A(n26928), .B(n26929), .Z(n26922) );
  AND U28592 ( .A(n26930), .B(n26931), .Z(n26929) );
  XOR U28593 ( .A(nreg[635]), .B(n26928), .Z(n26931) );
  XNOR U28594 ( .A(n16983), .B(n26928), .Z(n26930) );
  XOR U28595 ( .A(n26932), .B(n26933), .Z(n16983) );
  XOR U28596 ( .A(n26934), .B(n26935), .Z(n26928) );
  AND U28597 ( .A(n26936), .B(n26937), .Z(n26935) );
  XOR U28598 ( .A(nreg[634]), .B(n26934), .Z(n26937) );
  XNOR U28599 ( .A(n16995), .B(n26934), .Z(n26936) );
  XOR U28600 ( .A(n26938), .B(n26939), .Z(n16995) );
  XOR U28601 ( .A(n26940), .B(n26941), .Z(n26934) );
  AND U28602 ( .A(n26942), .B(n26943), .Z(n26941) );
  XOR U28603 ( .A(nreg[633]), .B(n26940), .Z(n26943) );
  XNOR U28604 ( .A(n17007), .B(n26940), .Z(n26942) );
  XOR U28605 ( .A(n26944), .B(n26945), .Z(n17007) );
  XOR U28606 ( .A(n26946), .B(n26947), .Z(n26940) );
  AND U28607 ( .A(n26948), .B(n26949), .Z(n26947) );
  XOR U28608 ( .A(nreg[632]), .B(n26946), .Z(n26949) );
  XNOR U28609 ( .A(n17019), .B(n26946), .Z(n26948) );
  XOR U28610 ( .A(n26950), .B(n26951), .Z(n17019) );
  XOR U28611 ( .A(n26952), .B(n26953), .Z(n26946) );
  AND U28612 ( .A(n26954), .B(n26955), .Z(n26953) );
  XOR U28613 ( .A(nreg[631]), .B(n26952), .Z(n26955) );
  XNOR U28614 ( .A(n17031), .B(n26952), .Z(n26954) );
  XOR U28615 ( .A(n26956), .B(n26957), .Z(n17031) );
  XOR U28616 ( .A(n26958), .B(n26959), .Z(n26952) );
  AND U28617 ( .A(n26960), .B(n26961), .Z(n26959) );
  XOR U28618 ( .A(nreg[630]), .B(n26958), .Z(n26961) );
  XNOR U28619 ( .A(n17043), .B(n26958), .Z(n26960) );
  XOR U28620 ( .A(n26962), .B(n26963), .Z(n17043) );
  XOR U28621 ( .A(n26964), .B(n26965), .Z(n26958) );
  AND U28622 ( .A(n26966), .B(n26967), .Z(n26965) );
  XOR U28623 ( .A(nreg[629]), .B(n26964), .Z(n26967) );
  XNOR U28624 ( .A(n17055), .B(n26964), .Z(n26966) );
  XOR U28625 ( .A(n26968), .B(n26969), .Z(n17055) );
  XOR U28626 ( .A(n26970), .B(n26971), .Z(n26964) );
  AND U28627 ( .A(n26972), .B(n26973), .Z(n26971) );
  XOR U28628 ( .A(nreg[628]), .B(n26970), .Z(n26973) );
  XNOR U28629 ( .A(n17067), .B(n26970), .Z(n26972) );
  XOR U28630 ( .A(n26974), .B(n26975), .Z(n17067) );
  XOR U28631 ( .A(n26976), .B(n26977), .Z(n26970) );
  AND U28632 ( .A(n26978), .B(n26979), .Z(n26977) );
  XOR U28633 ( .A(nreg[627]), .B(n26976), .Z(n26979) );
  XNOR U28634 ( .A(n17079), .B(n26976), .Z(n26978) );
  XOR U28635 ( .A(n26980), .B(n26981), .Z(n17079) );
  XOR U28636 ( .A(n26982), .B(n26983), .Z(n26976) );
  AND U28637 ( .A(n26984), .B(n26985), .Z(n26983) );
  XOR U28638 ( .A(nreg[626]), .B(n26982), .Z(n26985) );
  XNOR U28639 ( .A(n17091), .B(n26982), .Z(n26984) );
  XOR U28640 ( .A(n26986), .B(n26987), .Z(n17091) );
  XOR U28641 ( .A(n26988), .B(n26989), .Z(n26982) );
  AND U28642 ( .A(n26990), .B(n26991), .Z(n26989) );
  XOR U28643 ( .A(nreg[625]), .B(n26988), .Z(n26991) );
  XNOR U28644 ( .A(n17103), .B(n26988), .Z(n26990) );
  XOR U28645 ( .A(n26992), .B(n26993), .Z(n17103) );
  XOR U28646 ( .A(n26994), .B(n26995), .Z(n26988) );
  AND U28647 ( .A(n26996), .B(n26997), .Z(n26995) );
  XOR U28648 ( .A(nreg[624]), .B(n26994), .Z(n26997) );
  XNOR U28649 ( .A(n17115), .B(n26994), .Z(n26996) );
  XOR U28650 ( .A(n26998), .B(n26999), .Z(n17115) );
  XOR U28651 ( .A(n27000), .B(n27001), .Z(n26994) );
  AND U28652 ( .A(n27002), .B(n27003), .Z(n27001) );
  XOR U28653 ( .A(nreg[623]), .B(n27000), .Z(n27003) );
  XNOR U28654 ( .A(n17127), .B(n27000), .Z(n27002) );
  XOR U28655 ( .A(n27004), .B(n27005), .Z(n17127) );
  XOR U28656 ( .A(n27006), .B(n27007), .Z(n27000) );
  AND U28657 ( .A(n27008), .B(n27009), .Z(n27007) );
  XOR U28658 ( .A(nreg[622]), .B(n27006), .Z(n27009) );
  XNOR U28659 ( .A(n17139), .B(n27006), .Z(n27008) );
  XOR U28660 ( .A(n27010), .B(n27011), .Z(n17139) );
  XOR U28661 ( .A(n27012), .B(n27013), .Z(n27006) );
  AND U28662 ( .A(n27014), .B(n27015), .Z(n27013) );
  XOR U28663 ( .A(nreg[621]), .B(n27012), .Z(n27015) );
  XNOR U28664 ( .A(n17151), .B(n27012), .Z(n27014) );
  XOR U28665 ( .A(n27016), .B(n27017), .Z(n17151) );
  XOR U28666 ( .A(n27018), .B(n27019), .Z(n27012) );
  AND U28667 ( .A(n27020), .B(n27021), .Z(n27019) );
  XOR U28668 ( .A(nreg[620]), .B(n27018), .Z(n27021) );
  XNOR U28669 ( .A(n17163), .B(n27018), .Z(n27020) );
  XOR U28670 ( .A(n27022), .B(n27023), .Z(n17163) );
  XOR U28671 ( .A(n27024), .B(n27025), .Z(n27018) );
  AND U28672 ( .A(n27026), .B(n27027), .Z(n27025) );
  XOR U28673 ( .A(nreg[619]), .B(n27024), .Z(n27027) );
  XNOR U28674 ( .A(n17175), .B(n27024), .Z(n27026) );
  XOR U28675 ( .A(n27028), .B(n27029), .Z(n17175) );
  XOR U28676 ( .A(n27030), .B(n27031), .Z(n27024) );
  AND U28677 ( .A(n27032), .B(n27033), .Z(n27031) );
  XOR U28678 ( .A(nreg[618]), .B(n27030), .Z(n27033) );
  XNOR U28679 ( .A(n17187), .B(n27030), .Z(n27032) );
  XOR U28680 ( .A(n27034), .B(n27035), .Z(n17187) );
  XOR U28681 ( .A(n27036), .B(n27037), .Z(n27030) );
  AND U28682 ( .A(n27038), .B(n27039), .Z(n27037) );
  XOR U28683 ( .A(nreg[617]), .B(n27036), .Z(n27039) );
  XNOR U28684 ( .A(n17199), .B(n27036), .Z(n27038) );
  XOR U28685 ( .A(n27040), .B(n27041), .Z(n17199) );
  XOR U28686 ( .A(n27042), .B(n27043), .Z(n27036) );
  AND U28687 ( .A(n27044), .B(n27045), .Z(n27043) );
  XOR U28688 ( .A(nreg[616]), .B(n27042), .Z(n27045) );
  XNOR U28689 ( .A(n17211), .B(n27042), .Z(n27044) );
  XOR U28690 ( .A(n27046), .B(n27047), .Z(n17211) );
  XOR U28691 ( .A(n27048), .B(n27049), .Z(n27042) );
  AND U28692 ( .A(n27050), .B(n27051), .Z(n27049) );
  XOR U28693 ( .A(nreg[615]), .B(n27048), .Z(n27051) );
  XNOR U28694 ( .A(n17223), .B(n27048), .Z(n27050) );
  XOR U28695 ( .A(n27052), .B(n27053), .Z(n17223) );
  XOR U28696 ( .A(n27054), .B(n27055), .Z(n27048) );
  AND U28697 ( .A(n27056), .B(n27057), .Z(n27055) );
  XOR U28698 ( .A(nreg[614]), .B(n27054), .Z(n27057) );
  XNOR U28699 ( .A(n17235), .B(n27054), .Z(n27056) );
  XOR U28700 ( .A(n27058), .B(n27059), .Z(n17235) );
  XOR U28701 ( .A(n27060), .B(n27061), .Z(n27054) );
  AND U28702 ( .A(n27062), .B(n27063), .Z(n27061) );
  XOR U28703 ( .A(nreg[613]), .B(n27060), .Z(n27063) );
  XNOR U28704 ( .A(n17247), .B(n27060), .Z(n27062) );
  XOR U28705 ( .A(n27064), .B(n27065), .Z(n17247) );
  XOR U28706 ( .A(n27066), .B(n27067), .Z(n27060) );
  AND U28707 ( .A(n27068), .B(n27069), .Z(n27067) );
  XOR U28708 ( .A(nreg[612]), .B(n27066), .Z(n27069) );
  XNOR U28709 ( .A(n17259), .B(n27066), .Z(n27068) );
  XOR U28710 ( .A(n27070), .B(n27071), .Z(n17259) );
  XOR U28711 ( .A(n27072), .B(n27073), .Z(n27066) );
  AND U28712 ( .A(n27074), .B(n27075), .Z(n27073) );
  XOR U28713 ( .A(nreg[611]), .B(n27072), .Z(n27075) );
  XNOR U28714 ( .A(n17271), .B(n27072), .Z(n27074) );
  XOR U28715 ( .A(n27076), .B(n27077), .Z(n17271) );
  XOR U28716 ( .A(n27078), .B(n27079), .Z(n27072) );
  AND U28717 ( .A(n27080), .B(n27081), .Z(n27079) );
  XOR U28718 ( .A(nreg[610]), .B(n27078), .Z(n27081) );
  XNOR U28719 ( .A(n17283), .B(n27078), .Z(n27080) );
  XOR U28720 ( .A(n27082), .B(n27083), .Z(n17283) );
  XOR U28721 ( .A(n27084), .B(n27085), .Z(n27078) );
  AND U28722 ( .A(n27086), .B(n27087), .Z(n27085) );
  XOR U28723 ( .A(nreg[609]), .B(n27084), .Z(n27087) );
  XNOR U28724 ( .A(n17295), .B(n27084), .Z(n27086) );
  XOR U28725 ( .A(n27088), .B(n27089), .Z(n17295) );
  XOR U28726 ( .A(n27090), .B(n27091), .Z(n27084) );
  AND U28727 ( .A(n27092), .B(n27093), .Z(n27091) );
  XOR U28728 ( .A(nreg[608]), .B(n27090), .Z(n27093) );
  XNOR U28729 ( .A(n17307), .B(n27090), .Z(n27092) );
  XOR U28730 ( .A(n27094), .B(n27095), .Z(n17307) );
  XOR U28731 ( .A(n27096), .B(n27097), .Z(n27090) );
  AND U28732 ( .A(n27098), .B(n27099), .Z(n27097) );
  XOR U28733 ( .A(nreg[607]), .B(n27096), .Z(n27099) );
  XNOR U28734 ( .A(n17319), .B(n27096), .Z(n27098) );
  XOR U28735 ( .A(n27100), .B(n27101), .Z(n17319) );
  XOR U28736 ( .A(n27102), .B(n27103), .Z(n27096) );
  AND U28737 ( .A(n27104), .B(n27105), .Z(n27103) );
  XOR U28738 ( .A(nreg[606]), .B(n27102), .Z(n27105) );
  XNOR U28739 ( .A(n17331), .B(n27102), .Z(n27104) );
  XOR U28740 ( .A(n27106), .B(n27107), .Z(n17331) );
  XOR U28741 ( .A(n27108), .B(n27109), .Z(n27102) );
  AND U28742 ( .A(n27110), .B(n27111), .Z(n27109) );
  XOR U28743 ( .A(nreg[605]), .B(n27108), .Z(n27111) );
  XNOR U28744 ( .A(n17343), .B(n27108), .Z(n27110) );
  XOR U28745 ( .A(n27112), .B(n27113), .Z(n17343) );
  XOR U28746 ( .A(n27114), .B(n27115), .Z(n27108) );
  AND U28747 ( .A(n27116), .B(n27117), .Z(n27115) );
  XOR U28748 ( .A(nreg[604]), .B(n27114), .Z(n27117) );
  XNOR U28749 ( .A(n17355), .B(n27114), .Z(n27116) );
  XOR U28750 ( .A(n27118), .B(n27119), .Z(n17355) );
  XOR U28751 ( .A(n27120), .B(n27121), .Z(n27114) );
  AND U28752 ( .A(n27122), .B(n27123), .Z(n27121) );
  XOR U28753 ( .A(nreg[603]), .B(n27120), .Z(n27123) );
  XNOR U28754 ( .A(n17367), .B(n27120), .Z(n27122) );
  XOR U28755 ( .A(n27124), .B(n27125), .Z(n17367) );
  XOR U28756 ( .A(n27126), .B(n27127), .Z(n27120) );
  AND U28757 ( .A(n27128), .B(n27129), .Z(n27127) );
  XOR U28758 ( .A(nreg[602]), .B(n27126), .Z(n27129) );
  XNOR U28759 ( .A(n17379), .B(n27126), .Z(n27128) );
  XOR U28760 ( .A(n27130), .B(n27131), .Z(n17379) );
  XOR U28761 ( .A(n27132), .B(n27133), .Z(n27126) );
  AND U28762 ( .A(n27134), .B(n27135), .Z(n27133) );
  XOR U28763 ( .A(nreg[601]), .B(n27132), .Z(n27135) );
  XNOR U28764 ( .A(n17391), .B(n27132), .Z(n27134) );
  XOR U28765 ( .A(n27136), .B(n27137), .Z(n17391) );
  XOR U28766 ( .A(n27138), .B(n27139), .Z(n27132) );
  AND U28767 ( .A(n27140), .B(n27141), .Z(n27139) );
  XOR U28768 ( .A(nreg[600]), .B(n27138), .Z(n27141) );
  XNOR U28769 ( .A(n17403), .B(n27138), .Z(n27140) );
  XOR U28770 ( .A(n27142), .B(n27143), .Z(n17403) );
  XOR U28771 ( .A(n27144), .B(n27145), .Z(n27138) );
  AND U28772 ( .A(n27146), .B(n27147), .Z(n27145) );
  XOR U28773 ( .A(nreg[599]), .B(n27144), .Z(n27147) );
  XNOR U28774 ( .A(n17415), .B(n27144), .Z(n27146) );
  XOR U28775 ( .A(n27148), .B(n27149), .Z(n17415) );
  XOR U28776 ( .A(n27150), .B(n27151), .Z(n27144) );
  AND U28777 ( .A(n27152), .B(n27153), .Z(n27151) );
  XOR U28778 ( .A(nreg[598]), .B(n27150), .Z(n27153) );
  XNOR U28779 ( .A(n17427), .B(n27150), .Z(n27152) );
  XOR U28780 ( .A(n27154), .B(n27155), .Z(n17427) );
  XOR U28781 ( .A(n27156), .B(n27157), .Z(n27150) );
  AND U28782 ( .A(n27158), .B(n27159), .Z(n27157) );
  XOR U28783 ( .A(nreg[597]), .B(n27156), .Z(n27159) );
  XNOR U28784 ( .A(n17439), .B(n27156), .Z(n27158) );
  XOR U28785 ( .A(n27160), .B(n27161), .Z(n17439) );
  XOR U28786 ( .A(n27162), .B(n27163), .Z(n27156) );
  AND U28787 ( .A(n27164), .B(n27165), .Z(n27163) );
  XOR U28788 ( .A(nreg[596]), .B(n27162), .Z(n27165) );
  XNOR U28789 ( .A(n17451), .B(n27162), .Z(n27164) );
  XOR U28790 ( .A(n27166), .B(n27167), .Z(n17451) );
  XOR U28791 ( .A(n27168), .B(n27169), .Z(n27162) );
  AND U28792 ( .A(n27170), .B(n27171), .Z(n27169) );
  XOR U28793 ( .A(nreg[595]), .B(n27168), .Z(n27171) );
  XNOR U28794 ( .A(n17463), .B(n27168), .Z(n27170) );
  XOR U28795 ( .A(n27172), .B(n27173), .Z(n17463) );
  XOR U28796 ( .A(n27174), .B(n27175), .Z(n27168) );
  AND U28797 ( .A(n27176), .B(n27177), .Z(n27175) );
  XOR U28798 ( .A(nreg[594]), .B(n27174), .Z(n27177) );
  XNOR U28799 ( .A(n17475), .B(n27174), .Z(n27176) );
  XOR U28800 ( .A(n27178), .B(n27179), .Z(n17475) );
  XOR U28801 ( .A(n27180), .B(n27181), .Z(n27174) );
  AND U28802 ( .A(n27182), .B(n27183), .Z(n27181) );
  XOR U28803 ( .A(nreg[593]), .B(n27180), .Z(n27183) );
  XNOR U28804 ( .A(n17487), .B(n27180), .Z(n27182) );
  XOR U28805 ( .A(n27184), .B(n27185), .Z(n17487) );
  XOR U28806 ( .A(n27186), .B(n27187), .Z(n27180) );
  AND U28807 ( .A(n27188), .B(n27189), .Z(n27187) );
  XOR U28808 ( .A(nreg[592]), .B(n27186), .Z(n27189) );
  XNOR U28809 ( .A(n17499), .B(n27186), .Z(n27188) );
  XOR U28810 ( .A(n27190), .B(n27191), .Z(n17499) );
  XOR U28811 ( .A(n27192), .B(n27193), .Z(n27186) );
  AND U28812 ( .A(n27194), .B(n27195), .Z(n27193) );
  XOR U28813 ( .A(nreg[591]), .B(n27192), .Z(n27195) );
  XNOR U28814 ( .A(n17511), .B(n27192), .Z(n27194) );
  XOR U28815 ( .A(n27196), .B(n27197), .Z(n17511) );
  XOR U28816 ( .A(n27198), .B(n27199), .Z(n27192) );
  AND U28817 ( .A(n27200), .B(n27201), .Z(n27199) );
  XOR U28818 ( .A(nreg[590]), .B(n27198), .Z(n27201) );
  XNOR U28819 ( .A(n17523), .B(n27198), .Z(n27200) );
  XOR U28820 ( .A(n27202), .B(n27203), .Z(n17523) );
  XOR U28821 ( .A(n27204), .B(n27205), .Z(n27198) );
  AND U28822 ( .A(n27206), .B(n27207), .Z(n27205) );
  XOR U28823 ( .A(nreg[589]), .B(n27204), .Z(n27207) );
  XNOR U28824 ( .A(n17535), .B(n27204), .Z(n27206) );
  XOR U28825 ( .A(n27208), .B(n27209), .Z(n17535) );
  XOR U28826 ( .A(n27210), .B(n27211), .Z(n27204) );
  AND U28827 ( .A(n27212), .B(n27213), .Z(n27211) );
  XOR U28828 ( .A(nreg[588]), .B(n27210), .Z(n27213) );
  XNOR U28829 ( .A(n17547), .B(n27210), .Z(n27212) );
  XOR U28830 ( .A(n27214), .B(n27215), .Z(n17547) );
  XOR U28831 ( .A(n27216), .B(n27217), .Z(n27210) );
  AND U28832 ( .A(n27218), .B(n27219), .Z(n27217) );
  XOR U28833 ( .A(nreg[587]), .B(n27216), .Z(n27219) );
  XNOR U28834 ( .A(n17559), .B(n27216), .Z(n27218) );
  XOR U28835 ( .A(n27220), .B(n27221), .Z(n17559) );
  XOR U28836 ( .A(n27222), .B(n27223), .Z(n27216) );
  AND U28837 ( .A(n27224), .B(n27225), .Z(n27223) );
  XOR U28838 ( .A(nreg[586]), .B(n27222), .Z(n27225) );
  XNOR U28839 ( .A(n17571), .B(n27222), .Z(n27224) );
  XOR U28840 ( .A(n27226), .B(n27227), .Z(n17571) );
  XOR U28841 ( .A(n27228), .B(n27229), .Z(n27222) );
  AND U28842 ( .A(n27230), .B(n27231), .Z(n27229) );
  XOR U28843 ( .A(nreg[585]), .B(n27228), .Z(n27231) );
  XNOR U28844 ( .A(n17583), .B(n27228), .Z(n27230) );
  XOR U28845 ( .A(n27232), .B(n27233), .Z(n17583) );
  XOR U28846 ( .A(n27234), .B(n27235), .Z(n27228) );
  AND U28847 ( .A(n27236), .B(n27237), .Z(n27235) );
  XOR U28848 ( .A(nreg[584]), .B(n27234), .Z(n27237) );
  XNOR U28849 ( .A(n17595), .B(n27234), .Z(n27236) );
  XOR U28850 ( .A(n27238), .B(n27239), .Z(n17595) );
  XOR U28851 ( .A(n27240), .B(n27241), .Z(n27234) );
  AND U28852 ( .A(n27242), .B(n27243), .Z(n27241) );
  XOR U28853 ( .A(nreg[583]), .B(n27240), .Z(n27243) );
  XNOR U28854 ( .A(n17607), .B(n27240), .Z(n27242) );
  XOR U28855 ( .A(n27244), .B(n27245), .Z(n17607) );
  XOR U28856 ( .A(n27246), .B(n27247), .Z(n27240) );
  AND U28857 ( .A(n27248), .B(n27249), .Z(n27247) );
  XOR U28858 ( .A(nreg[582]), .B(n27246), .Z(n27249) );
  XNOR U28859 ( .A(n17619), .B(n27246), .Z(n27248) );
  XOR U28860 ( .A(n27250), .B(n27251), .Z(n17619) );
  XOR U28861 ( .A(n27252), .B(n27253), .Z(n27246) );
  AND U28862 ( .A(n27254), .B(n27255), .Z(n27253) );
  XOR U28863 ( .A(nreg[581]), .B(n27252), .Z(n27255) );
  XNOR U28864 ( .A(n17631), .B(n27252), .Z(n27254) );
  XOR U28865 ( .A(n27256), .B(n27257), .Z(n17631) );
  XOR U28866 ( .A(n27258), .B(n27259), .Z(n27252) );
  AND U28867 ( .A(n27260), .B(n27261), .Z(n27259) );
  XOR U28868 ( .A(nreg[580]), .B(n27258), .Z(n27261) );
  XNOR U28869 ( .A(n17643), .B(n27258), .Z(n27260) );
  XOR U28870 ( .A(n27262), .B(n27263), .Z(n17643) );
  XOR U28871 ( .A(n27264), .B(n27265), .Z(n27258) );
  AND U28872 ( .A(n27266), .B(n27267), .Z(n27265) );
  XOR U28873 ( .A(nreg[579]), .B(n27264), .Z(n27267) );
  XNOR U28874 ( .A(n17655), .B(n27264), .Z(n27266) );
  XOR U28875 ( .A(n27268), .B(n27269), .Z(n17655) );
  XOR U28876 ( .A(n27270), .B(n27271), .Z(n27264) );
  AND U28877 ( .A(n27272), .B(n27273), .Z(n27271) );
  XOR U28878 ( .A(nreg[578]), .B(n27270), .Z(n27273) );
  XNOR U28879 ( .A(n17667), .B(n27270), .Z(n27272) );
  XOR U28880 ( .A(n27274), .B(n27275), .Z(n17667) );
  XOR U28881 ( .A(n27276), .B(n27277), .Z(n27270) );
  AND U28882 ( .A(n27278), .B(n27279), .Z(n27277) );
  XOR U28883 ( .A(nreg[577]), .B(n27276), .Z(n27279) );
  XNOR U28884 ( .A(n17679), .B(n27276), .Z(n27278) );
  XOR U28885 ( .A(n27280), .B(n27281), .Z(n17679) );
  XOR U28886 ( .A(n27282), .B(n27283), .Z(n27276) );
  AND U28887 ( .A(n27284), .B(n27285), .Z(n27283) );
  XOR U28888 ( .A(nreg[576]), .B(n27282), .Z(n27285) );
  XNOR U28889 ( .A(n17691), .B(n27282), .Z(n27284) );
  XOR U28890 ( .A(n27286), .B(n27287), .Z(n17691) );
  XOR U28891 ( .A(n27288), .B(n27289), .Z(n27282) );
  AND U28892 ( .A(n27290), .B(n27291), .Z(n27289) );
  XOR U28893 ( .A(nreg[575]), .B(n27288), .Z(n27291) );
  XNOR U28894 ( .A(n17703), .B(n27288), .Z(n27290) );
  XOR U28895 ( .A(n27292), .B(n27293), .Z(n17703) );
  XOR U28896 ( .A(n27294), .B(n27295), .Z(n27288) );
  AND U28897 ( .A(n27296), .B(n27297), .Z(n27295) );
  XOR U28898 ( .A(nreg[574]), .B(n27294), .Z(n27297) );
  XNOR U28899 ( .A(n17715), .B(n27294), .Z(n27296) );
  XOR U28900 ( .A(n27298), .B(n27299), .Z(n17715) );
  XOR U28901 ( .A(n27300), .B(n27301), .Z(n27294) );
  AND U28902 ( .A(n27302), .B(n27303), .Z(n27301) );
  XOR U28903 ( .A(nreg[573]), .B(n27300), .Z(n27303) );
  XNOR U28904 ( .A(n17727), .B(n27300), .Z(n27302) );
  XOR U28905 ( .A(n27304), .B(n27305), .Z(n17727) );
  XOR U28906 ( .A(n27306), .B(n27307), .Z(n27300) );
  AND U28907 ( .A(n27308), .B(n27309), .Z(n27307) );
  XOR U28908 ( .A(nreg[572]), .B(n27306), .Z(n27309) );
  XNOR U28909 ( .A(n17739), .B(n27306), .Z(n27308) );
  XOR U28910 ( .A(n27310), .B(n27311), .Z(n17739) );
  XOR U28911 ( .A(n27312), .B(n27313), .Z(n27306) );
  AND U28912 ( .A(n27314), .B(n27315), .Z(n27313) );
  XOR U28913 ( .A(nreg[571]), .B(n27312), .Z(n27315) );
  XNOR U28914 ( .A(n17751), .B(n27312), .Z(n27314) );
  XOR U28915 ( .A(n27316), .B(n27317), .Z(n17751) );
  XOR U28916 ( .A(n27318), .B(n27319), .Z(n27312) );
  AND U28917 ( .A(n27320), .B(n27321), .Z(n27319) );
  XOR U28918 ( .A(nreg[570]), .B(n27318), .Z(n27321) );
  XNOR U28919 ( .A(n17763), .B(n27318), .Z(n27320) );
  XOR U28920 ( .A(n27322), .B(n27323), .Z(n17763) );
  XOR U28921 ( .A(n27324), .B(n27325), .Z(n27318) );
  AND U28922 ( .A(n27326), .B(n27327), .Z(n27325) );
  XOR U28923 ( .A(nreg[569]), .B(n27324), .Z(n27327) );
  XNOR U28924 ( .A(n17775), .B(n27324), .Z(n27326) );
  XOR U28925 ( .A(n27328), .B(n27329), .Z(n17775) );
  XOR U28926 ( .A(n27330), .B(n27331), .Z(n27324) );
  AND U28927 ( .A(n27332), .B(n27333), .Z(n27331) );
  XOR U28928 ( .A(nreg[568]), .B(n27330), .Z(n27333) );
  XNOR U28929 ( .A(n17787), .B(n27330), .Z(n27332) );
  XOR U28930 ( .A(n27334), .B(n27335), .Z(n17787) );
  XOR U28931 ( .A(n27336), .B(n27337), .Z(n27330) );
  AND U28932 ( .A(n27338), .B(n27339), .Z(n27337) );
  XOR U28933 ( .A(nreg[567]), .B(n27336), .Z(n27339) );
  XNOR U28934 ( .A(n17799), .B(n27336), .Z(n27338) );
  XOR U28935 ( .A(n27340), .B(n27341), .Z(n17799) );
  XOR U28936 ( .A(n27342), .B(n27343), .Z(n27336) );
  AND U28937 ( .A(n27344), .B(n27345), .Z(n27343) );
  XOR U28938 ( .A(nreg[566]), .B(n27342), .Z(n27345) );
  XNOR U28939 ( .A(n17811), .B(n27342), .Z(n27344) );
  XOR U28940 ( .A(n27346), .B(n27347), .Z(n17811) );
  XOR U28941 ( .A(n27348), .B(n27349), .Z(n27342) );
  AND U28942 ( .A(n27350), .B(n27351), .Z(n27349) );
  XOR U28943 ( .A(nreg[565]), .B(n27348), .Z(n27351) );
  XNOR U28944 ( .A(n17823), .B(n27348), .Z(n27350) );
  XOR U28945 ( .A(n27352), .B(n27353), .Z(n17823) );
  XOR U28946 ( .A(n27354), .B(n27355), .Z(n27348) );
  AND U28947 ( .A(n27356), .B(n27357), .Z(n27355) );
  XOR U28948 ( .A(nreg[564]), .B(n27354), .Z(n27357) );
  XNOR U28949 ( .A(n17835), .B(n27354), .Z(n27356) );
  XOR U28950 ( .A(n27358), .B(n27359), .Z(n17835) );
  XOR U28951 ( .A(n27360), .B(n27361), .Z(n27354) );
  AND U28952 ( .A(n27362), .B(n27363), .Z(n27361) );
  XOR U28953 ( .A(nreg[563]), .B(n27360), .Z(n27363) );
  XNOR U28954 ( .A(n17847), .B(n27360), .Z(n27362) );
  XOR U28955 ( .A(n27364), .B(n27365), .Z(n17847) );
  XOR U28956 ( .A(n27366), .B(n27367), .Z(n27360) );
  AND U28957 ( .A(n27368), .B(n27369), .Z(n27367) );
  XOR U28958 ( .A(nreg[562]), .B(n27366), .Z(n27369) );
  XNOR U28959 ( .A(n17859), .B(n27366), .Z(n27368) );
  XOR U28960 ( .A(n27370), .B(n27371), .Z(n17859) );
  XOR U28961 ( .A(n27372), .B(n27373), .Z(n27366) );
  AND U28962 ( .A(n27374), .B(n27375), .Z(n27373) );
  XOR U28963 ( .A(nreg[561]), .B(n27372), .Z(n27375) );
  XNOR U28964 ( .A(n17871), .B(n27372), .Z(n27374) );
  XOR U28965 ( .A(n27376), .B(n27377), .Z(n17871) );
  XOR U28966 ( .A(n27378), .B(n27379), .Z(n27372) );
  AND U28967 ( .A(n27380), .B(n27381), .Z(n27379) );
  XOR U28968 ( .A(nreg[560]), .B(n27378), .Z(n27381) );
  XNOR U28969 ( .A(n17883), .B(n27378), .Z(n27380) );
  XOR U28970 ( .A(n27382), .B(n27383), .Z(n17883) );
  XOR U28971 ( .A(n27384), .B(n27385), .Z(n27378) );
  AND U28972 ( .A(n27386), .B(n27387), .Z(n27385) );
  XOR U28973 ( .A(nreg[559]), .B(n27384), .Z(n27387) );
  XNOR U28974 ( .A(n17895), .B(n27384), .Z(n27386) );
  XOR U28975 ( .A(n27388), .B(n27389), .Z(n17895) );
  XOR U28976 ( .A(n27390), .B(n27391), .Z(n27384) );
  AND U28977 ( .A(n27392), .B(n27393), .Z(n27391) );
  XOR U28978 ( .A(nreg[558]), .B(n27390), .Z(n27393) );
  XNOR U28979 ( .A(n17907), .B(n27390), .Z(n27392) );
  XOR U28980 ( .A(n27394), .B(n27395), .Z(n17907) );
  XOR U28981 ( .A(n27396), .B(n27397), .Z(n27390) );
  AND U28982 ( .A(n27398), .B(n27399), .Z(n27397) );
  XOR U28983 ( .A(nreg[557]), .B(n27396), .Z(n27399) );
  XNOR U28984 ( .A(n17919), .B(n27396), .Z(n27398) );
  XOR U28985 ( .A(n27400), .B(n27401), .Z(n17919) );
  XOR U28986 ( .A(n27402), .B(n27403), .Z(n27396) );
  AND U28987 ( .A(n27404), .B(n27405), .Z(n27403) );
  XOR U28988 ( .A(nreg[556]), .B(n27402), .Z(n27405) );
  XNOR U28989 ( .A(n17931), .B(n27402), .Z(n27404) );
  XOR U28990 ( .A(n27406), .B(n27407), .Z(n17931) );
  XOR U28991 ( .A(n27408), .B(n27409), .Z(n27402) );
  AND U28992 ( .A(n27410), .B(n27411), .Z(n27409) );
  XOR U28993 ( .A(nreg[555]), .B(n27408), .Z(n27411) );
  XNOR U28994 ( .A(n17943), .B(n27408), .Z(n27410) );
  XOR U28995 ( .A(n27412), .B(n27413), .Z(n17943) );
  XOR U28996 ( .A(n27414), .B(n27415), .Z(n27408) );
  AND U28997 ( .A(n27416), .B(n27417), .Z(n27415) );
  XOR U28998 ( .A(nreg[554]), .B(n27414), .Z(n27417) );
  XNOR U28999 ( .A(n17955), .B(n27414), .Z(n27416) );
  XOR U29000 ( .A(n27418), .B(n27419), .Z(n17955) );
  XOR U29001 ( .A(n27420), .B(n27421), .Z(n27414) );
  AND U29002 ( .A(n27422), .B(n27423), .Z(n27421) );
  XOR U29003 ( .A(nreg[553]), .B(n27420), .Z(n27423) );
  XNOR U29004 ( .A(n17967), .B(n27420), .Z(n27422) );
  XOR U29005 ( .A(n27424), .B(n27425), .Z(n17967) );
  XOR U29006 ( .A(n27426), .B(n27427), .Z(n27420) );
  AND U29007 ( .A(n27428), .B(n27429), .Z(n27427) );
  XOR U29008 ( .A(nreg[552]), .B(n27426), .Z(n27429) );
  XNOR U29009 ( .A(n17979), .B(n27426), .Z(n27428) );
  XOR U29010 ( .A(n27430), .B(n27431), .Z(n17979) );
  XOR U29011 ( .A(n27432), .B(n27433), .Z(n27426) );
  AND U29012 ( .A(n27434), .B(n27435), .Z(n27433) );
  XOR U29013 ( .A(nreg[551]), .B(n27432), .Z(n27435) );
  XNOR U29014 ( .A(n17991), .B(n27432), .Z(n27434) );
  XOR U29015 ( .A(n27436), .B(n27437), .Z(n17991) );
  XOR U29016 ( .A(n27438), .B(n27439), .Z(n27432) );
  AND U29017 ( .A(n27440), .B(n27441), .Z(n27439) );
  XOR U29018 ( .A(nreg[550]), .B(n27438), .Z(n27441) );
  XNOR U29019 ( .A(n18003), .B(n27438), .Z(n27440) );
  XOR U29020 ( .A(n27442), .B(n27443), .Z(n18003) );
  XOR U29021 ( .A(n27444), .B(n27445), .Z(n27438) );
  AND U29022 ( .A(n27446), .B(n27447), .Z(n27445) );
  XOR U29023 ( .A(nreg[549]), .B(n27444), .Z(n27447) );
  XNOR U29024 ( .A(n18015), .B(n27444), .Z(n27446) );
  XOR U29025 ( .A(n27448), .B(n27449), .Z(n18015) );
  XOR U29026 ( .A(n27450), .B(n27451), .Z(n27444) );
  AND U29027 ( .A(n27452), .B(n27453), .Z(n27451) );
  XOR U29028 ( .A(nreg[548]), .B(n27450), .Z(n27453) );
  XNOR U29029 ( .A(n18027), .B(n27450), .Z(n27452) );
  XOR U29030 ( .A(n27454), .B(n27455), .Z(n18027) );
  XOR U29031 ( .A(n27456), .B(n27457), .Z(n27450) );
  AND U29032 ( .A(n27458), .B(n27459), .Z(n27457) );
  XOR U29033 ( .A(nreg[547]), .B(n27456), .Z(n27459) );
  XNOR U29034 ( .A(n18039), .B(n27456), .Z(n27458) );
  XOR U29035 ( .A(n27460), .B(n27461), .Z(n18039) );
  XOR U29036 ( .A(n27462), .B(n27463), .Z(n27456) );
  AND U29037 ( .A(n27464), .B(n27465), .Z(n27463) );
  XOR U29038 ( .A(nreg[546]), .B(n27462), .Z(n27465) );
  XNOR U29039 ( .A(n18051), .B(n27462), .Z(n27464) );
  XOR U29040 ( .A(n27466), .B(n27467), .Z(n18051) );
  XOR U29041 ( .A(n27468), .B(n27469), .Z(n27462) );
  AND U29042 ( .A(n27470), .B(n27471), .Z(n27469) );
  XOR U29043 ( .A(nreg[545]), .B(n27468), .Z(n27471) );
  XNOR U29044 ( .A(n18063), .B(n27468), .Z(n27470) );
  XOR U29045 ( .A(n27472), .B(n27473), .Z(n18063) );
  XOR U29046 ( .A(n27474), .B(n27475), .Z(n27468) );
  AND U29047 ( .A(n27476), .B(n27477), .Z(n27475) );
  XOR U29048 ( .A(nreg[544]), .B(n27474), .Z(n27477) );
  XNOR U29049 ( .A(n18075), .B(n27474), .Z(n27476) );
  XOR U29050 ( .A(n27478), .B(n27479), .Z(n18075) );
  XOR U29051 ( .A(n27480), .B(n27481), .Z(n27474) );
  AND U29052 ( .A(n27482), .B(n27483), .Z(n27481) );
  XOR U29053 ( .A(nreg[543]), .B(n27480), .Z(n27483) );
  XNOR U29054 ( .A(n18087), .B(n27480), .Z(n27482) );
  XOR U29055 ( .A(n27484), .B(n27485), .Z(n18087) );
  XOR U29056 ( .A(n27486), .B(n27487), .Z(n27480) );
  AND U29057 ( .A(n27488), .B(n27489), .Z(n27487) );
  XOR U29058 ( .A(nreg[542]), .B(n27486), .Z(n27489) );
  XNOR U29059 ( .A(n18099), .B(n27486), .Z(n27488) );
  XOR U29060 ( .A(n27490), .B(n27491), .Z(n18099) );
  XOR U29061 ( .A(n27492), .B(n27493), .Z(n27486) );
  AND U29062 ( .A(n27494), .B(n27495), .Z(n27493) );
  XOR U29063 ( .A(nreg[541]), .B(n27492), .Z(n27495) );
  XNOR U29064 ( .A(n18111), .B(n27492), .Z(n27494) );
  XOR U29065 ( .A(n27496), .B(n27497), .Z(n18111) );
  XOR U29066 ( .A(n27498), .B(n27499), .Z(n27492) );
  AND U29067 ( .A(n27500), .B(n27501), .Z(n27499) );
  XOR U29068 ( .A(nreg[540]), .B(n27498), .Z(n27501) );
  XNOR U29069 ( .A(n18123), .B(n27498), .Z(n27500) );
  XOR U29070 ( .A(n27502), .B(n27503), .Z(n18123) );
  XOR U29071 ( .A(n27504), .B(n27505), .Z(n27498) );
  AND U29072 ( .A(n27506), .B(n27507), .Z(n27505) );
  XOR U29073 ( .A(nreg[539]), .B(n27504), .Z(n27507) );
  XNOR U29074 ( .A(n18135), .B(n27504), .Z(n27506) );
  XOR U29075 ( .A(n27508), .B(n27509), .Z(n18135) );
  XOR U29076 ( .A(n27510), .B(n27511), .Z(n27504) );
  AND U29077 ( .A(n27512), .B(n27513), .Z(n27511) );
  XOR U29078 ( .A(nreg[538]), .B(n27510), .Z(n27513) );
  XNOR U29079 ( .A(n18147), .B(n27510), .Z(n27512) );
  XOR U29080 ( .A(n27514), .B(n27515), .Z(n18147) );
  XOR U29081 ( .A(n27516), .B(n27517), .Z(n27510) );
  AND U29082 ( .A(n27518), .B(n27519), .Z(n27517) );
  XOR U29083 ( .A(nreg[537]), .B(n27516), .Z(n27519) );
  XNOR U29084 ( .A(n18159), .B(n27516), .Z(n27518) );
  XOR U29085 ( .A(n27520), .B(n27521), .Z(n18159) );
  XOR U29086 ( .A(n27522), .B(n27523), .Z(n27516) );
  AND U29087 ( .A(n27524), .B(n27525), .Z(n27523) );
  XOR U29088 ( .A(nreg[536]), .B(n27522), .Z(n27525) );
  XNOR U29089 ( .A(n18171), .B(n27522), .Z(n27524) );
  XOR U29090 ( .A(n27526), .B(n27527), .Z(n18171) );
  XOR U29091 ( .A(n27528), .B(n27529), .Z(n27522) );
  AND U29092 ( .A(n27530), .B(n27531), .Z(n27529) );
  XOR U29093 ( .A(nreg[535]), .B(n27528), .Z(n27531) );
  XNOR U29094 ( .A(n18183), .B(n27528), .Z(n27530) );
  XOR U29095 ( .A(n27532), .B(n27533), .Z(n18183) );
  XOR U29096 ( .A(n27534), .B(n27535), .Z(n27528) );
  AND U29097 ( .A(n27536), .B(n27537), .Z(n27535) );
  XOR U29098 ( .A(nreg[534]), .B(n27534), .Z(n27537) );
  XNOR U29099 ( .A(n18195), .B(n27534), .Z(n27536) );
  XOR U29100 ( .A(n27538), .B(n27539), .Z(n18195) );
  XOR U29101 ( .A(n27540), .B(n27541), .Z(n27534) );
  AND U29102 ( .A(n27542), .B(n27543), .Z(n27541) );
  XOR U29103 ( .A(nreg[533]), .B(n27540), .Z(n27543) );
  XNOR U29104 ( .A(n18207), .B(n27540), .Z(n27542) );
  XOR U29105 ( .A(n27544), .B(n27545), .Z(n18207) );
  XOR U29106 ( .A(n27546), .B(n27547), .Z(n27540) );
  AND U29107 ( .A(n27548), .B(n27549), .Z(n27547) );
  XOR U29108 ( .A(nreg[532]), .B(n27546), .Z(n27549) );
  XNOR U29109 ( .A(n18219), .B(n27546), .Z(n27548) );
  XOR U29110 ( .A(n27550), .B(n27551), .Z(n18219) );
  XOR U29111 ( .A(n27552), .B(n27553), .Z(n27546) );
  AND U29112 ( .A(n27554), .B(n27555), .Z(n27553) );
  XOR U29113 ( .A(nreg[531]), .B(n27552), .Z(n27555) );
  XNOR U29114 ( .A(n18231), .B(n27552), .Z(n27554) );
  XOR U29115 ( .A(n27556), .B(n27557), .Z(n18231) );
  XOR U29116 ( .A(n27558), .B(n27559), .Z(n27552) );
  AND U29117 ( .A(n27560), .B(n27561), .Z(n27559) );
  XOR U29118 ( .A(nreg[530]), .B(n27558), .Z(n27561) );
  XNOR U29119 ( .A(n18243), .B(n27558), .Z(n27560) );
  XOR U29120 ( .A(n27562), .B(n27563), .Z(n18243) );
  XOR U29121 ( .A(n27564), .B(n27565), .Z(n27558) );
  AND U29122 ( .A(n27566), .B(n27567), .Z(n27565) );
  XOR U29123 ( .A(nreg[529]), .B(n27564), .Z(n27567) );
  XNOR U29124 ( .A(n18255), .B(n27564), .Z(n27566) );
  XOR U29125 ( .A(n27568), .B(n27569), .Z(n18255) );
  XOR U29126 ( .A(n27570), .B(n27571), .Z(n27564) );
  AND U29127 ( .A(n27572), .B(n27573), .Z(n27571) );
  XOR U29128 ( .A(nreg[528]), .B(n27570), .Z(n27573) );
  XNOR U29129 ( .A(n18267), .B(n27570), .Z(n27572) );
  XOR U29130 ( .A(n27574), .B(n27575), .Z(n18267) );
  XOR U29131 ( .A(n27576), .B(n27577), .Z(n27570) );
  AND U29132 ( .A(n27578), .B(n27579), .Z(n27577) );
  XOR U29133 ( .A(nreg[527]), .B(n27576), .Z(n27579) );
  XNOR U29134 ( .A(n18279), .B(n27576), .Z(n27578) );
  XOR U29135 ( .A(n27580), .B(n27581), .Z(n18279) );
  XOR U29136 ( .A(n27582), .B(n27583), .Z(n27576) );
  AND U29137 ( .A(n27584), .B(n27585), .Z(n27583) );
  XOR U29138 ( .A(nreg[526]), .B(n27582), .Z(n27585) );
  XNOR U29139 ( .A(n18291), .B(n27582), .Z(n27584) );
  XOR U29140 ( .A(n27586), .B(n27587), .Z(n18291) );
  XOR U29141 ( .A(n27588), .B(n27589), .Z(n27582) );
  AND U29142 ( .A(n27590), .B(n27591), .Z(n27589) );
  XOR U29143 ( .A(nreg[525]), .B(n27588), .Z(n27591) );
  XNOR U29144 ( .A(n18303), .B(n27588), .Z(n27590) );
  XOR U29145 ( .A(n27592), .B(n27593), .Z(n18303) );
  XOR U29146 ( .A(n27594), .B(n27595), .Z(n27588) );
  AND U29147 ( .A(n27596), .B(n27597), .Z(n27595) );
  XOR U29148 ( .A(nreg[524]), .B(n27594), .Z(n27597) );
  XNOR U29149 ( .A(n18315), .B(n27594), .Z(n27596) );
  XOR U29150 ( .A(n27598), .B(n27599), .Z(n18315) );
  XOR U29151 ( .A(n27600), .B(n27601), .Z(n27594) );
  AND U29152 ( .A(n27602), .B(n27603), .Z(n27601) );
  XOR U29153 ( .A(nreg[523]), .B(n27600), .Z(n27603) );
  XNOR U29154 ( .A(n18327), .B(n27600), .Z(n27602) );
  XOR U29155 ( .A(n27604), .B(n27605), .Z(n18327) );
  XOR U29156 ( .A(n27606), .B(n27607), .Z(n27600) );
  AND U29157 ( .A(n27608), .B(n27609), .Z(n27607) );
  XOR U29158 ( .A(nreg[522]), .B(n27606), .Z(n27609) );
  XNOR U29159 ( .A(n18339), .B(n27606), .Z(n27608) );
  XOR U29160 ( .A(n27610), .B(n27611), .Z(n18339) );
  XOR U29161 ( .A(n27612), .B(n27613), .Z(n27606) );
  AND U29162 ( .A(n27614), .B(n27615), .Z(n27613) );
  XOR U29163 ( .A(nreg[521]), .B(n27612), .Z(n27615) );
  XNOR U29164 ( .A(n18351), .B(n27612), .Z(n27614) );
  XOR U29165 ( .A(n27616), .B(n27617), .Z(n18351) );
  XOR U29166 ( .A(n27618), .B(n27619), .Z(n27612) );
  AND U29167 ( .A(n27620), .B(n27621), .Z(n27619) );
  XOR U29168 ( .A(nreg[520]), .B(n27618), .Z(n27621) );
  XNOR U29169 ( .A(n18363), .B(n27618), .Z(n27620) );
  XOR U29170 ( .A(n27622), .B(n27623), .Z(n18363) );
  XOR U29171 ( .A(n27624), .B(n27625), .Z(n27618) );
  AND U29172 ( .A(n27626), .B(n27627), .Z(n27625) );
  XOR U29173 ( .A(nreg[519]), .B(n27624), .Z(n27627) );
  XNOR U29174 ( .A(n18375), .B(n27624), .Z(n27626) );
  XOR U29175 ( .A(n27628), .B(n27629), .Z(n18375) );
  XOR U29176 ( .A(n27630), .B(n27631), .Z(n27624) );
  AND U29177 ( .A(n27632), .B(n27633), .Z(n27631) );
  XOR U29178 ( .A(nreg[518]), .B(n27630), .Z(n27633) );
  XNOR U29179 ( .A(n18387), .B(n27630), .Z(n27632) );
  XOR U29180 ( .A(n27634), .B(n27635), .Z(n18387) );
  XOR U29181 ( .A(n27636), .B(n27637), .Z(n27630) );
  AND U29182 ( .A(n27638), .B(n27639), .Z(n27637) );
  XOR U29183 ( .A(nreg[517]), .B(n27636), .Z(n27639) );
  XNOR U29184 ( .A(n18399), .B(n27636), .Z(n27638) );
  XOR U29185 ( .A(n27640), .B(n27641), .Z(n18399) );
  XOR U29186 ( .A(n27642), .B(n27643), .Z(n27636) );
  AND U29187 ( .A(n27644), .B(n27645), .Z(n27643) );
  XOR U29188 ( .A(nreg[516]), .B(n27642), .Z(n27645) );
  XNOR U29189 ( .A(n18411), .B(n27642), .Z(n27644) );
  XOR U29190 ( .A(n27646), .B(n27647), .Z(n18411) );
  XOR U29191 ( .A(n27648), .B(n27649), .Z(n27642) );
  AND U29192 ( .A(n27650), .B(n27651), .Z(n27649) );
  XOR U29193 ( .A(nreg[515]), .B(n27648), .Z(n27651) );
  XNOR U29194 ( .A(n18423), .B(n27648), .Z(n27650) );
  XOR U29195 ( .A(n27652), .B(n27653), .Z(n18423) );
  XOR U29196 ( .A(n27654), .B(n27655), .Z(n27648) );
  AND U29197 ( .A(n27656), .B(n27657), .Z(n27655) );
  XOR U29198 ( .A(nreg[514]), .B(n27654), .Z(n27657) );
  XNOR U29199 ( .A(n18435), .B(n27654), .Z(n27656) );
  XOR U29200 ( .A(n27658), .B(n27659), .Z(n18435) );
  XOR U29201 ( .A(n27660), .B(n27661), .Z(n27654) );
  AND U29202 ( .A(n27662), .B(n27663), .Z(n27661) );
  XOR U29203 ( .A(nreg[513]), .B(n27660), .Z(n27663) );
  XNOR U29204 ( .A(n18447), .B(n27660), .Z(n27662) );
  XOR U29205 ( .A(n27664), .B(n27665), .Z(n18447) );
  XOR U29206 ( .A(n27666), .B(n27667), .Z(n27660) );
  AND U29207 ( .A(n27668), .B(n27669), .Z(n27667) );
  XOR U29208 ( .A(nreg[512]), .B(n27666), .Z(n27669) );
  XNOR U29209 ( .A(n18459), .B(n27666), .Z(n27668) );
  XOR U29210 ( .A(n27670), .B(n27671), .Z(n18459) );
  XOR U29211 ( .A(n27672), .B(n27673), .Z(n27666) );
  AND U29212 ( .A(n27674), .B(n27675), .Z(n27673) );
  XOR U29213 ( .A(nreg[511]), .B(n27672), .Z(n27675) );
  XNOR U29214 ( .A(n18471), .B(n27672), .Z(n27674) );
  XOR U29215 ( .A(n27676), .B(n27677), .Z(n18471) );
  XOR U29216 ( .A(n27678), .B(n27679), .Z(n27672) );
  AND U29217 ( .A(n27680), .B(n27681), .Z(n27679) );
  XOR U29218 ( .A(nreg[510]), .B(n27678), .Z(n27681) );
  XNOR U29219 ( .A(n18483), .B(n27678), .Z(n27680) );
  XOR U29220 ( .A(n27682), .B(n27683), .Z(n18483) );
  XOR U29221 ( .A(n27684), .B(n27685), .Z(n27678) );
  AND U29222 ( .A(n27686), .B(n27687), .Z(n27685) );
  XOR U29223 ( .A(nreg[509]), .B(n27684), .Z(n27687) );
  XNOR U29224 ( .A(n18495), .B(n27684), .Z(n27686) );
  XOR U29225 ( .A(n27688), .B(n27689), .Z(n18495) );
  XOR U29226 ( .A(n27690), .B(n27691), .Z(n27684) );
  AND U29227 ( .A(n27692), .B(n27693), .Z(n27691) );
  XOR U29228 ( .A(nreg[508]), .B(n27690), .Z(n27693) );
  XNOR U29229 ( .A(n18507), .B(n27690), .Z(n27692) );
  XOR U29230 ( .A(n27694), .B(n27695), .Z(n18507) );
  XOR U29231 ( .A(n27696), .B(n27697), .Z(n27690) );
  AND U29232 ( .A(n27698), .B(n27699), .Z(n27697) );
  XOR U29233 ( .A(nreg[507]), .B(n27696), .Z(n27699) );
  XNOR U29234 ( .A(n18519), .B(n27696), .Z(n27698) );
  XOR U29235 ( .A(n27700), .B(n27701), .Z(n18519) );
  XOR U29236 ( .A(n27702), .B(n27703), .Z(n27696) );
  AND U29237 ( .A(n27704), .B(n27705), .Z(n27703) );
  XOR U29238 ( .A(nreg[506]), .B(n27702), .Z(n27705) );
  XNOR U29239 ( .A(n18531), .B(n27702), .Z(n27704) );
  XOR U29240 ( .A(n27706), .B(n27707), .Z(n18531) );
  XOR U29241 ( .A(n27708), .B(n27709), .Z(n27702) );
  AND U29242 ( .A(n27710), .B(n27711), .Z(n27709) );
  XOR U29243 ( .A(nreg[505]), .B(n27708), .Z(n27711) );
  XNOR U29244 ( .A(n18543), .B(n27708), .Z(n27710) );
  XOR U29245 ( .A(n27712), .B(n27713), .Z(n18543) );
  XOR U29246 ( .A(n27714), .B(n27715), .Z(n27708) );
  AND U29247 ( .A(n27716), .B(n27717), .Z(n27715) );
  XOR U29248 ( .A(nreg[504]), .B(n27714), .Z(n27717) );
  XNOR U29249 ( .A(n18555), .B(n27714), .Z(n27716) );
  XOR U29250 ( .A(n27718), .B(n27719), .Z(n18555) );
  XOR U29251 ( .A(n27720), .B(n27721), .Z(n27714) );
  AND U29252 ( .A(n27722), .B(n27723), .Z(n27721) );
  XOR U29253 ( .A(nreg[503]), .B(n27720), .Z(n27723) );
  XNOR U29254 ( .A(n18567), .B(n27720), .Z(n27722) );
  XOR U29255 ( .A(n27724), .B(n27725), .Z(n18567) );
  XOR U29256 ( .A(n27726), .B(n27727), .Z(n27720) );
  AND U29257 ( .A(n27728), .B(n27729), .Z(n27727) );
  XOR U29258 ( .A(nreg[502]), .B(n27726), .Z(n27729) );
  XNOR U29259 ( .A(n18579), .B(n27726), .Z(n27728) );
  XOR U29260 ( .A(n27730), .B(n27731), .Z(n18579) );
  XOR U29261 ( .A(n27732), .B(n27733), .Z(n27726) );
  AND U29262 ( .A(n27734), .B(n27735), .Z(n27733) );
  XOR U29263 ( .A(nreg[501]), .B(n27732), .Z(n27735) );
  XNOR U29264 ( .A(n18591), .B(n27732), .Z(n27734) );
  XOR U29265 ( .A(n27736), .B(n27737), .Z(n18591) );
  XOR U29266 ( .A(n27738), .B(n27739), .Z(n27732) );
  AND U29267 ( .A(n27740), .B(n27741), .Z(n27739) );
  XOR U29268 ( .A(nreg[500]), .B(n27738), .Z(n27741) );
  XNOR U29269 ( .A(n18603), .B(n27738), .Z(n27740) );
  XOR U29270 ( .A(n27742), .B(n27743), .Z(n18603) );
  XOR U29271 ( .A(n27744), .B(n27745), .Z(n27738) );
  AND U29272 ( .A(n27746), .B(n27747), .Z(n27745) );
  XOR U29273 ( .A(nreg[499]), .B(n27744), .Z(n27747) );
  XNOR U29274 ( .A(n18615), .B(n27744), .Z(n27746) );
  XOR U29275 ( .A(n27748), .B(n27749), .Z(n18615) );
  XOR U29276 ( .A(n27750), .B(n27751), .Z(n27744) );
  AND U29277 ( .A(n27752), .B(n27753), .Z(n27751) );
  XOR U29278 ( .A(nreg[498]), .B(n27750), .Z(n27753) );
  XNOR U29279 ( .A(n18627), .B(n27750), .Z(n27752) );
  XOR U29280 ( .A(n27754), .B(n27755), .Z(n18627) );
  XOR U29281 ( .A(n27756), .B(n27757), .Z(n27750) );
  AND U29282 ( .A(n27758), .B(n27759), .Z(n27757) );
  XOR U29283 ( .A(nreg[497]), .B(n27756), .Z(n27759) );
  XNOR U29284 ( .A(n18639), .B(n27756), .Z(n27758) );
  XOR U29285 ( .A(n27760), .B(n27761), .Z(n18639) );
  XOR U29286 ( .A(n27762), .B(n27763), .Z(n27756) );
  AND U29287 ( .A(n27764), .B(n27765), .Z(n27763) );
  XOR U29288 ( .A(nreg[496]), .B(n27762), .Z(n27765) );
  XNOR U29289 ( .A(n18651), .B(n27762), .Z(n27764) );
  XOR U29290 ( .A(n27766), .B(n27767), .Z(n18651) );
  XOR U29291 ( .A(n27768), .B(n27769), .Z(n27762) );
  AND U29292 ( .A(n27770), .B(n27771), .Z(n27769) );
  XOR U29293 ( .A(nreg[495]), .B(n27768), .Z(n27771) );
  XNOR U29294 ( .A(n18663), .B(n27768), .Z(n27770) );
  XOR U29295 ( .A(n27772), .B(n27773), .Z(n18663) );
  XOR U29296 ( .A(n27774), .B(n27775), .Z(n27768) );
  AND U29297 ( .A(n27776), .B(n27777), .Z(n27775) );
  XOR U29298 ( .A(nreg[494]), .B(n27774), .Z(n27777) );
  XNOR U29299 ( .A(n18675), .B(n27774), .Z(n27776) );
  XOR U29300 ( .A(n27778), .B(n27779), .Z(n18675) );
  XOR U29301 ( .A(n27780), .B(n27781), .Z(n27774) );
  AND U29302 ( .A(n27782), .B(n27783), .Z(n27781) );
  XOR U29303 ( .A(nreg[493]), .B(n27780), .Z(n27783) );
  XNOR U29304 ( .A(n18687), .B(n27780), .Z(n27782) );
  XOR U29305 ( .A(n27784), .B(n27785), .Z(n18687) );
  XOR U29306 ( .A(n27786), .B(n27787), .Z(n27780) );
  AND U29307 ( .A(n27788), .B(n27789), .Z(n27787) );
  XOR U29308 ( .A(nreg[492]), .B(n27786), .Z(n27789) );
  XNOR U29309 ( .A(n18699), .B(n27786), .Z(n27788) );
  XOR U29310 ( .A(n27790), .B(n27791), .Z(n18699) );
  XOR U29311 ( .A(n27792), .B(n27793), .Z(n27786) );
  AND U29312 ( .A(n27794), .B(n27795), .Z(n27793) );
  XOR U29313 ( .A(nreg[491]), .B(n27792), .Z(n27795) );
  XNOR U29314 ( .A(n18711), .B(n27792), .Z(n27794) );
  XOR U29315 ( .A(n27796), .B(n27797), .Z(n18711) );
  XOR U29316 ( .A(n27798), .B(n27799), .Z(n27792) );
  AND U29317 ( .A(n27800), .B(n27801), .Z(n27799) );
  XOR U29318 ( .A(nreg[490]), .B(n27798), .Z(n27801) );
  XNOR U29319 ( .A(n18723), .B(n27798), .Z(n27800) );
  XOR U29320 ( .A(n27802), .B(n27803), .Z(n18723) );
  XOR U29321 ( .A(n27804), .B(n27805), .Z(n27798) );
  AND U29322 ( .A(n27806), .B(n27807), .Z(n27805) );
  XOR U29323 ( .A(nreg[489]), .B(n27804), .Z(n27807) );
  XNOR U29324 ( .A(n18735), .B(n27804), .Z(n27806) );
  XOR U29325 ( .A(n27808), .B(n27809), .Z(n18735) );
  XOR U29326 ( .A(n27810), .B(n27811), .Z(n27804) );
  AND U29327 ( .A(n27812), .B(n27813), .Z(n27811) );
  XOR U29328 ( .A(nreg[488]), .B(n27810), .Z(n27813) );
  XNOR U29329 ( .A(n18747), .B(n27810), .Z(n27812) );
  XOR U29330 ( .A(n27814), .B(n27815), .Z(n18747) );
  XOR U29331 ( .A(n27816), .B(n27817), .Z(n27810) );
  AND U29332 ( .A(n27818), .B(n27819), .Z(n27817) );
  XOR U29333 ( .A(nreg[487]), .B(n27816), .Z(n27819) );
  XNOR U29334 ( .A(n18759), .B(n27816), .Z(n27818) );
  XOR U29335 ( .A(n27820), .B(n27821), .Z(n18759) );
  XOR U29336 ( .A(n27822), .B(n27823), .Z(n27816) );
  AND U29337 ( .A(n27824), .B(n27825), .Z(n27823) );
  XOR U29338 ( .A(nreg[486]), .B(n27822), .Z(n27825) );
  XNOR U29339 ( .A(n18771), .B(n27822), .Z(n27824) );
  XOR U29340 ( .A(n27826), .B(n27827), .Z(n18771) );
  XOR U29341 ( .A(n27828), .B(n27829), .Z(n27822) );
  AND U29342 ( .A(n27830), .B(n27831), .Z(n27829) );
  XOR U29343 ( .A(nreg[485]), .B(n27828), .Z(n27831) );
  XNOR U29344 ( .A(n18783), .B(n27828), .Z(n27830) );
  XOR U29345 ( .A(n27832), .B(n27833), .Z(n18783) );
  XOR U29346 ( .A(n27834), .B(n27835), .Z(n27828) );
  AND U29347 ( .A(n27836), .B(n27837), .Z(n27835) );
  XOR U29348 ( .A(nreg[484]), .B(n27834), .Z(n27837) );
  XNOR U29349 ( .A(n18795), .B(n27834), .Z(n27836) );
  XOR U29350 ( .A(n27838), .B(n27839), .Z(n18795) );
  XOR U29351 ( .A(n27840), .B(n27841), .Z(n27834) );
  AND U29352 ( .A(n27842), .B(n27843), .Z(n27841) );
  XOR U29353 ( .A(nreg[483]), .B(n27840), .Z(n27843) );
  XNOR U29354 ( .A(n18807), .B(n27840), .Z(n27842) );
  XOR U29355 ( .A(n27844), .B(n27845), .Z(n18807) );
  XOR U29356 ( .A(n27846), .B(n27847), .Z(n27840) );
  AND U29357 ( .A(n27848), .B(n27849), .Z(n27847) );
  XOR U29358 ( .A(nreg[482]), .B(n27846), .Z(n27849) );
  XNOR U29359 ( .A(n18819), .B(n27846), .Z(n27848) );
  XOR U29360 ( .A(n27850), .B(n27851), .Z(n18819) );
  XOR U29361 ( .A(n27852), .B(n27853), .Z(n27846) );
  AND U29362 ( .A(n27854), .B(n27855), .Z(n27853) );
  XOR U29363 ( .A(nreg[481]), .B(n27852), .Z(n27855) );
  XNOR U29364 ( .A(n18831), .B(n27852), .Z(n27854) );
  XOR U29365 ( .A(n27856), .B(n27857), .Z(n18831) );
  XOR U29366 ( .A(n27858), .B(n27859), .Z(n27852) );
  AND U29367 ( .A(n27860), .B(n27861), .Z(n27859) );
  XOR U29368 ( .A(nreg[480]), .B(n27858), .Z(n27861) );
  XNOR U29369 ( .A(n18843), .B(n27858), .Z(n27860) );
  XOR U29370 ( .A(n27862), .B(n27863), .Z(n18843) );
  XOR U29371 ( .A(n27864), .B(n27865), .Z(n27858) );
  AND U29372 ( .A(n27866), .B(n27867), .Z(n27865) );
  XOR U29373 ( .A(nreg[479]), .B(n27864), .Z(n27867) );
  XNOR U29374 ( .A(n18855), .B(n27864), .Z(n27866) );
  XOR U29375 ( .A(n27868), .B(n27869), .Z(n18855) );
  XOR U29376 ( .A(n27870), .B(n27871), .Z(n27864) );
  AND U29377 ( .A(n27872), .B(n27873), .Z(n27871) );
  XOR U29378 ( .A(nreg[478]), .B(n27870), .Z(n27873) );
  XNOR U29379 ( .A(n18867), .B(n27870), .Z(n27872) );
  XOR U29380 ( .A(n27874), .B(n27875), .Z(n18867) );
  XOR U29381 ( .A(n27876), .B(n27877), .Z(n27870) );
  AND U29382 ( .A(n27878), .B(n27879), .Z(n27877) );
  XOR U29383 ( .A(nreg[477]), .B(n27876), .Z(n27879) );
  XNOR U29384 ( .A(n18879), .B(n27876), .Z(n27878) );
  XOR U29385 ( .A(n27880), .B(n27881), .Z(n18879) );
  XOR U29386 ( .A(n27882), .B(n27883), .Z(n27876) );
  AND U29387 ( .A(n27884), .B(n27885), .Z(n27883) );
  XOR U29388 ( .A(nreg[476]), .B(n27882), .Z(n27885) );
  XNOR U29389 ( .A(n18891), .B(n27882), .Z(n27884) );
  XOR U29390 ( .A(n27886), .B(n27887), .Z(n18891) );
  XOR U29391 ( .A(n27888), .B(n27889), .Z(n27882) );
  AND U29392 ( .A(n27890), .B(n27891), .Z(n27889) );
  XOR U29393 ( .A(nreg[475]), .B(n27888), .Z(n27891) );
  XNOR U29394 ( .A(n18903), .B(n27888), .Z(n27890) );
  XOR U29395 ( .A(n27892), .B(n27893), .Z(n18903) );
  XOR U29396 ( .A(n27894), .B(n27895), .Z(n27888) );
  AND U29397 ( .A(n27896), .B(n27897), .Z(n27895) );
  XOR U29398 ( .A(nreg[474]), .B(n27894), .Z(n27897) );
  XNOR U29399 ( .A(n18915), .B(n27894), .Z(n27896) );
  XOR U29400 ( .A(n27898), .B(n27899), .Z(n18915) );
  XOR U29401 ( .A(n27900), .B(n27901), .Z(n27894) );
  AND U29402 ( .A(n27902), .B(n27903), .Z(n27901) );
  XOR U29403 ( .A(nreg[473]), .B(n27900), .Z(n27903) );
  XNOR U29404 ( .A(n18927), .B(n27900), .Z(n27902) );
  XOR U29405 ( .A(n27904), .B(n27905), .Z(n18927) );
  XOR U29406 ( .A(n27906), .B(n27907), .Z(n27900) );
  AND U29407 ( .A(n27908), .B(n27909), .Z(n27907) );
  XOR U29408 ( .A(nreg[472]), .B(n27906), .Z(n27909) );
  XNOR U29409 ( .A(n18939), .B(n27906), .Z(n27908) );
  XOR U29410 ( .A(n27910), .B(n27911), .Z(n18939) );
  XOR U29411 ( .A(n27912), .B(n27913), .Z(n27906) );
  AND U29412 ( .A(n27914), .B(n27915), .Z(n27913) );
  XOR U29413 ( .A(nreg[471]), .B(n27912), .Z(n27915) );
  XNOR U29414 ( .A(n18951), .B(n27912), .Z(n27914) );
  XOR U29415 ( .A(n27916), .B(n27917), .Z(n18951) );
  XOR U29416 ( .A(n27918), .B(n27919), .Z(n27912) );
  AND U29417 ( .A(n27920), .B(n27921), .Z(n27919) );
  XOR U29418 ( .A(nreg[470]), .B(n27918), .Z(n27921) );
  XNOR U29419 ( .A(n18963), .B(n27918), .Z(n27920) );
  XOR U29420 ( .A(n27922), .B(n27923), .Z(n18963) );
  XOR U29421 ( .A(n27924), .B(n27925), .Z(n27918) );
  AND U29422 ( .A(n27926), .B(n27927), .Z(n27925) );
  XOR U29423 ( .A(nreg[469]), .B(n27924), .Z(n27927) );
  XNOR U29424 ( .A(n18975), .B(n27924), .Z(n27926) );
  XOR U29425 ( .A(n27928), .B(n27929), .Z(n18975) );
  XOR U29426 ( .A(n27930), .B(n27931), .Z(n27924) );
  AND U29427 ( .A(n27932), .B(n27933), .Z(n27931) );
  XOR U29428 ( .A(nreg[468]), .B(n27930), .Z(n27933) );
  XNOR U29429 ( .A(n18987), .B(n27930), .Z(n27932) );
  XOR U29430 ( .A(n27934), .B(n27935), .Z(n18987) );
  XOR U29431 ( .A(n27936), .B(n27937), .Z(n27930) );
  AND U29432 ( .A(n27938), .B(n27939), .Z(n27937) );
  XOR U29433 ( .A(nreg[467]), .B(n27936), .Z(n27939) );
  XNOR U29434 ( .A(n18999), .B(n27936), .Z(n27938) );
  XOR U29435 ( .A(n27940), .B(n27941), .Z(n18999) );
  XOR U29436 ( .A(n27942), .B(n27943), .Z(n27936) );
  AND U29437 ( .A(n27944), .B(n27945), .Z(n27943) );
  XOR U29438 ( .A(nreg[466]), .B(n27942), .Z(n27945) );
  XNOR U29439 ( .A(n19011), .B(n27942), .Z(n27944) );
  XOR U29440 ( .A(n27946), .B(n27947), .Z(n19011) );
  XOR U29441 ( .A(n27948), .B(n27949), .Z(n27942) );
  AND U29442 ( .A(n27950), .B(n27951), .Z(n27949) );
  XOR U29443 ( .A(nreg[465]), .B(n27948), .Z(n27951) );
  XNOR U29444 ( .A(n19023), .B(n27948), .Z(n27950) );
  XOR U29445 ( .A(n27952), .B(n27953), .Z(n19023) );
  XOR U29446 ( .A(n27954), .B(n27955), .Z(n27948) );
  AND U29447 ( .A(n27956), .B(n27957), .Z(n27955) );
  XOR U29448 ( .A(nreg[464]), .B(n27954), .Z(n27957) );
  XNOR U29449 ( .A(n19035), .B(n27954), .Z(n27956) );
  XOR U29450 ( .A(n27958), .B(n27959), .Z(n19035) );
  XOR U29451 ( .A(n27960), .B(n27961), .Z(n27954) );
  AND U29452 ( .A(n27962), .B(n27963), .Z(n27961) );
  XOR U29453 ( .A(nreg[463]), .B(n27960), .Z(n27963) );
  XNOR U29454 ( .A(n19047), .B(n27960), .Z(n27962) );
  XOR U29455 ( .A(n27964), .B(n27965), .Z(n19047) );
  XOR U29456 ( .A(n27966), .B(n27967), .Z(n27960) );
  AND U29457 ( .A(n27968), .B(n27969), .Z(n27967) );
  XOR U29458 ( .A(nreg[462]), .B(n27966), .Z(n27969) );
  XNOR U29459 ( .A(n19059), .B(n27966), .Z(n27968) );
  XOR U29460 ( .A(n27970), .B(n27971), .Z(n19059) );
  XOR U29461 ( .A(n27972), .B(n27973), .Z(n27966) );
  AND U29462 ( .A(n27974), .B(n27975), .Z(n27973) );
  XOR U29463 ( .A(nreg[461]), .B(n27972), .Z(n27975) );
  XNOR U29464 ( .A(n19071), .B(n27972), .Z(n27974) );
  XOR U29465 ( .A(n27976), .B(n27977), .Z(n19071) );
  XOR U29466 ( .A(n27978), .B(n27979), .Z(n27972) );
  AND U29467 ( .A(n27980), .B(n27981), .Z(n27979) );
  XOR U29468 ( .A(nreg[460]), .B(n27978), .Z(n27981) );
  XNOR U29469 ( .A(n19083), .B(n27978), .Z(n27980) );
  XOR U29470 ( .A(n27982), .B(n27983), .Z(n19083) );
  XOR U29471 ( .A(n27984), .B(n27985), .Z(n27978) );
  AND U29472 ( .A(n27986), .B(n27987), .Z(n27985) );
  XOR U29473 ( .A(nreg[459]), .B(n27984), .Z(n27987) );
  XNOR U29474 ( .A(n19095), .B(n27984), .Z(n27986) );
  XOR U29475 ( .A(n27988), .B(n27989), .Z(n19095) );
  XOR U29476 ( .A(n27990), .B(n27991), .Z(n27984) );
  AND U29477 ( .A(n27992), .B(n27993), .Z(n27991) );
  XOR U29478 ( .A(nreg[458]), .B(n27990), .Z(n27993) );
  XNOR U29479 ( .A(n19107), .B(n27990), .Z(n27992) );
  XOR U29480 ( .A(n27994), .B(n27995), .Z(n19107) );
  XOR U29481 ( .A(n27996), .B(n27997), .Z(n27990) );
  AND U29482 ( .A(n27998), .B(n27999), .Z(n27997) );
  XOR U29483 ( .A(nreg[457]), .B(n27996), .Z(n27999) );
  XNOR U29484 ( .A(n19119), .B(n27996), .Z(n27998) );
  XOR U29485 ( .A(n28000), .B(n28001), .Z(n19119) );
  XOR U29486 ( .A(n28002), .B(n28003), .Z(n27996) );
  AND U29487 ( .A(n28004), .B(n28005), .Z(n28003) );
  XOR U29488 ( .A(nreg[456]), .B(n28002), .Z(n28005) );
  XNOR U29489 ( .A(n19131), .B(n28002), .Z(n28004) );
  XOR U29490 ( .A(n28006), .B(n28007), .Z(n19131) );
  XOR U29491 ( .A(n28008), .B(n28009), .Z(n28002) );
  AND U29492 ( .A(n28010), .B(n28011), .Z(n28009) );
  XOR U29493 ( .A(nreg[455]), .B(n28008), .Z(n28011) );
  XNOR U29494 ( .A(n19143), .B(n28008), .Z(n28010) );
  XOR U29495 ( .A(n28012), .B(n28013), .Z(n19143) );
  XOR U29496 ( .A(n28014), .B(n28015), .Z(n28008) );
  AND U29497 ( .A(n28016), .B(n28017), .Z(n28015) );
  XOR U29498 ( .A(nreg[454]), .B(n28014), .Z(n28017) );
  XNOR U29499 ( .A(n19155), .B(n28014), .Z(n28016) );
  XOR U29500 ( .A(n28018), .B(n28019), .Z(n19155) );
  XOR U29501 ( .A(n28020), .B(n28021), .Z(n28014) );
  AND U29502 ( .A(n28022), .B(n28023), .Z(n28021) );
  XOR U29503 ( .A(nreg[453]), .B(n28020), .Z(n28023) );
  XNOR U29504 ( .A(n19167), .B(n28020), .Z(n28022) );
  XOR U29505 ( .A(n28024), .B(n28025), .Z(n19167) );
  XOR U29506 ( .A(n28026), .B(n28027), .Z(n28020) );
  AND U29507 ( .A(n28028), .B(n28029), .Z(n28027) );
  XOR U29508 ( .A(nreg[452]), .B(n28026), .Z(n28029) );
  XNOR U29509 ( .A(n19179), .B(n28026), .Z(n28028) );
  XOR U29510 ( .A(n28030), .B(n28031), .Z(n19179) );
  XOR U29511 ( .A(n28032), .B(n28033), .Z(n28026) );
  AND U29512 ( .A(n28034), .B(n28035), .Z(n28033) );
  XOR U29513 ( .A(nreg[451]), .B(n28032), .Z(n28035) );
  XNOR U29514 ( .A(n19191), .B(n28032), .Z(n28034) );
  XOR U29515 ( .A(n28036), .B(n28037), .Z(n19191) );
  XOR U29516 ( .A(n28038), .B(n28039), .Z(n28032) );
  AND U29517 ( .A(n28040), .B(n28041), .Z(n28039) );
  XOR U29518 ( .A(nreg[450]), .B(n28038), .Z(n28041) );
  XNOR U29519 ( .A(n19203), .B(n28038), .Z(n28040) );
  XOR U29520 ( .A(n28042), .B(n28043), .Z(n19203) );
  XOR U29521 ( .A(n28044), .B(n28045), .Z(n28038) );
  AND U29522 ( .A(n28046), .B(n28047), .Z(n28045) );
  XOR U29523 ( .A(nreg[449]), .B(n28044), .Z(n28047) );
  XNOR U29524 ( .A(n19215), .B(n28044), .Z(n28046) );
  XOR U29525 ( .A(n28048), .B(n28049), .Z(n19215) );
  XOR U29526 ( .A(n28050), .B(n28051), .Z(n28044) );
  AND U29527 ( .A(n28052), .B(n28053), .Z(n28051) );
  XOR U29528 ( .A(nreg[448]), .B(n28050), .Z(n28053) );
  XNOR U29529 ( .A(n19227), .B(n28050), .Z(n28052) );
  XOR U29530 ( .A(n28054), .B(n28055), .Z(n19227) );
  XOR U29531 ( .A(n28056), .B(n28057), .Z(n28050) );
  AND U29532 ( .A(n28058), .B(n28059), .Z(n28057) );
  XOR U29533 ( .A(nreg[447]), .B(n28056), .Z(n28059) );
  XNOR U29534 ( .A(n19239), .B(n28056), .Z(n28058) );
  XOR U29535 ( .A(n28060), .B(n28061), .Z(n19239) );
  XOR U29536 ( .A(n28062), .B(n28063), .Z(n28056) );
  AND U29537 ( .A(n28064), .B(n28065), .Z(n28063) );
  XOR U29538 ( .A(nreg[446]), .B(n28062), .Z(n28065) );
  XNOR U29539 ( .A(n19251), .B(n28062), .Z(n28064) );
  XOR U29540 ( .A(n28066), .B(n28067), .Z(n19251) );
  XOR U29541 ( .A(n28068), .B(n28069), .Z(n28062) );
  AND U29542 ( .A(n28070), .B(n28071), .Z(n28069) );
  XOR U29543 ( .A(nreg[445]), .B(n28068), .Z(n28071) );
  XNOR U29544 ( .A(n19263), .B(n28068), .Z(n28070) );
  XOR U29545 ( .A(n28072), .B(n28073), .Z(n19263) );
  XOR U29546 ( .A(n28074), .B(n28075), .Z(n28068) );
  AND U29547 ( .A(n28076), .B(n28077), .Z(n28075) );
  XOR U29548 ( .A(nreg[444]), .B(n28074), .Z(n28077) );
  XNOR U29549 ( .A(n19275), .B(n28074), .Z(n28076) );
  XOR U29550 ( .A(n28078), .B(n28079), .Z(n19275) );
  XOR U29551 ( .A(n28080), .B(n28081), .Z(n28074) );
  AND U29552 ( .A(n28082), .B(n28083), .Z(n28081) );
  XOR U29553 ( .A(nreg[443]), .B(n28080), .Z(n28083) );
  XNOR U29554 ( .A(n19287), .B(n28080), .Z(n28082) );
  XOR U29555 ( .A(n28084), .B(n28085), .Z(n19287) );
  XOR U29556 ( .A(n28086), .B(n28087), .Z(n28080) );
  AND U29557 ( .A(n28088), .B(n28089), .Z(n28087) );
  XOR U29558 ( .A(nreg[442]), .B(n28086), .Z(n28089) );
  XNOR U29559 ( .A(n19299), .B(n28086), .Z(n28088) );
  XOR U29560 ( .A(n28090), .B(n28091), .Z(n19299) );
  XOR U29561 ( .A(n28092), .B(n28093), .Z(n28086) );
  AND U29562 ( .A(n28094), .B(n28095), .Z(n28093) );
  XOR U29563 ( .A(nreg[441]), .B(n28092), .Z(n28095) );
  XNOR U29564 ( .A(n19311), .B(n28092), .Z(n28094) );
  XOR U29565 ( .A(n28096), .B(n28097), .Z(n19311) );
  XOR U29566 ( .A(n28098), .B(n28099), .Z(n28092) );
  AND U29567 ( .A(n28100), .B(n28101), .Z(n28099) );
  XOR U29568 ( .A(nreg[440]), .B(n28098), .Z(n28101) );
  XNOR U29569 ( .A(n19323), .B(n28098), .Z(n28100) );
  XOR U29570 ( .A(n28102), .B(n28103), .Z(n19323) );
  XOR U29571 ( .A(n28104), .B(n28105), .Z(n28098) );
  AND U29572 ( .A(n28106), .B(n28107), .Z(n28105) );
  XOR U29573 ( .A(nreg[439]), .B(n28104), .Z(n28107) );
  XNOR U29574 ( .A(n19335), .B(n28104), .Z(n28106) );
  XOR U29575 ( .A(n28108), .B(n28109), .Z(n19335) );
  XOR U29576 ( .A(n28110), .B(n28111), .Z(n28104) );
  AND U29577 ( .A(n28112), .B(n28113), .Z(n28111) );
  XOR U29578 ( .A(nreg[438]), .B(n28110), .Z(n28113) );
  XNOR U29579 ( .A(n19347), .B(n28110), .Z(n28112) );
  XOR U29580 ( .A(n28114), .B(n28115), .Z(n19347) );
  XOR U29581 ( .A(n28116), .B(n28117), .Z(n28110) );
  AND U29582 ( .A(n28118), .B(n28119), .Z(n28117) );
  XOR U29583 ( .A(nreg[437]), .B(n28116), .Z(n28119) );
  XNOR U29584 ( .A(n19359), .B(n28116), .Z(n28118) );
  XOR U29585 ( .A(n28120), .B(n28121), .Z(n19359) );
  XOR U29586 ( .A(n28122), .B(n28123), .Z(n28116) );
  AND U29587 ( .A(n28124), .B(n28125), .Z(n28123) );
  XOR U29588 ( .A(nreg[436]), .B(n28122), .Z(n28125) );
  XNOR U29589 ( .A(n19371), .B(n28122), .Z(n28124) );
  XOR U29590 ( .A(n28126), .B(n28127), .Z(n19371) );
  XOR U29591 ( .A(n28128), .B(n28129), .Z(n28122) );
  AND U29592 ( .A(n28130), .B(n28131), .Z(n28129) );
  XOR U29593 ( .A(nreg[435]), .B(n28128), .Z(n28131) );
  XNOR U29594 ( .A(n19383), .B(n28128), .Z(n28130) );
  XOR U29595 ( .A(n28132), .B(n28133), .Z(n19383) );
  XOR U29596 ( .A(n28134), .B(n28135), .Z(n28128) );
  AND U29597 ( .A(n28136), .B(n28137), .Z(n28135) );
  XOR U29598 ( .A(nreg[434]), .B(n28134), .Z(n28137) );
  XNOR U29599 ( .A(n19395), .B(n28134), .Z(n28136) );
  XOR U29600 ( .A(n28138), .B(n28139), .Z(n19395) );
  XOR U29601 ( .A(n28140), .B(n28141), .Z(n28134) );
  AND U29602 ( .A(n28142), .B(n28143), .Z(n28141) );
  XOR U29603 ( .A(nreg[433]), .B(n28140), .Z(n28143) );
  XNOR U29604 ( .A(n19407), .B(n28140), .Z(n28142) );
  XOR U29605 ( .A(n28144), .B(n28145), .Z(n19407) );
  XOR U29606 ( .A(n28146), .B(n28147), .Z(n28140) );
  AND U29607 ( .A(n28148), .B(n28149), .Z(n28147) );
  XOR U29608 ( .A(nreg[432]), .B(n28146), .Z(n28149) );
  XNOR U29609 ( .A(n19419), .B(n28146), .Z(n28148) );
  XOR U29610 ( .A(n28150), .B(n28151), .Z(n19419) );
  XOR U29611 ( .A(n28152), .B(n28153), .Z(n28146) );
  AND U29612 ( .A(n28154), .B(n28155), .Z(n28153) );
  XOR U29613 ( .A(nreg[431]), .B(n28152), .Z(n28155) );
  XNOR U29614 ( .A(n19431), .B(n28152), .Z(n28154) );
  XOR U29615 ( .A(n28156), .B(n28157), .Z(n19431) );
  XOR U29616 ( .A(n28158), .B(n28159), .Z(n28152) );
  AND U29617 ( .A(n28160), .B(n28161), .Z(n28159) );
  XOR U29618 ( .A(nreg[430]), .B(n28158), .Z(n28161) );
  XNOR U29619 ( .A(n19443), .B(n28158), .Z(n28160) );
  XOR U29620 ( .A(n28162), .B(n28163), .Z(n19443) );
  XOR U29621 ( .A(n28164), .B(n28165), .Z(n28158) );
  AND U29622 ( .A(n28166), .B(n28167), .Z(n28165) );
  XOR U29623 ( .A(nreg[429]), .B(n28164), .Z(n28167) );
  XNOR U29624 ( .A(n19455), .B(n28164), .Z(n28166) );
  XOR U29625 ( .A(n28168), .B(n28169), .Z(n19455) );
  XOR U29626 ( .A(n28170), .B(n28171), .Z(n28164) );
  AND U29627 ( .A(n28172), .B(n28173), .Z(n28171) );
  XOR U29628 ( .A(nreg[428]), .B(n28170), .Z(n28173) );
  XNOR U29629 ( .A(n19467), .B(n28170), .Z(n28172) );
  XOR U29630 ( .A(n28174), .B(n28175), .Z(n19467) );
  XOR U29631 ( .A(n28176), .B(n28177), .Z(n28170) );
  AND U29632 ( .A(n28178), .B(n28179), .Z(n28177) );
  XOR U29633 ( .A(nreg[427]), .B(n28176), .Z(n28179) );
  XNOR U29634 ( .A(n19479), .B(n28176), .Z(n28178) );
  XOR U29635 ( .A(n28180), .B(n28181), .Z(n19479) );
  XOR U29636 ( .A(n28182), .B(n28183), .Z(n28176) );
  AND U29637 ( .A(n28184), .B(n28185), .Z(n28183) );
  XOR U29638 ( .A(nreg[426]), .B(n28182), .Z(n28185) );
  XNOR U29639 ( .A(n19491), .B(n28182), .Z(n28184) );
  XOR U29640 ( .A(n28186), .B(n28187), .Z(n19491) );
  XOR U29641 ( .A(n28188), .B(n28189), .Z(n28182) );
  AND U29642 ( .A(n28190), .B(n28191), .Z(n28189) );
  XOR U29643 ( .A(nreg[425]), .B(n28188), .Z(n28191) );
  XNOR U29644 ( .A(n19503), .B(n28188), .Z(n28190) );
  XOR U29645 ( .A(n28192), .B(n28193), .Z(n19503) );
  XOR U29646 ( .A(n28194), .B(n28195), .Z(n28188) );
  AND U29647 ( .A(n28196), .B(n28197), .Z(n28195) );
  XOR U29648 ( .A(nreg[424]), .B(n28194), .Z(n28197) );
  XNOR U29649 ( .A(n19515), .B(n28194), .Z(n28196) );
  XOR U29650 ( .A(n28198), .B(n28199), .Z(n19515) );
  XOR U29651 ( .A(n28200), .B(n28201), .Z(n28194) );
  AND U29652 ( .A(n28202), .B(n28203), .Z(n28201) );
  XOR U29653 ( .A(nreg[423]), .B(n28200), .Z(n28203) );
  XNOR U29654 ( .A(n19527), .B(n28200), .Z(n28202) );
  XOR U29655 ( .A(n28204), .B(n28205), .Z(n19527) );
  XOR U29656 ( .A(n28206), .B(n28207), .Z(n28200) );
  AND U29657 ( .A(n28208), .B(n28209), .Z(n28207) );
  XOR U29658 ( .A(nreg[422]), .B(n28206), .Z(n28209) );
  XNOR U29659 ( .A(n19539), .B(n28206), .Z(n28208) );
  XOR U29660 ( .A(n28210), .B(n28211), .Z(n19539) );
  XOR U29661 ( .A(n28212), .B(n28213), .Z(n28206) );
  AND U29662 ( .A(n28214), .B(n28215), .Z(n28213) );
  XOR U29663 ( .A(nreg[421]), .B(n28212), .Z(n28215) );
  XNOR U29664 ( .A(n19551), .B(n28212), .Z(n28214) );
  XOR U29665 ( .A(n28216), .B(n28217), .Z(n19551) );
  XOR U29666 ( .A(n28218), .B(n28219), .Z(n28212) );
  AND U29667 ( .A(n28220), .B(n28221), .Z(n28219) );
  XOR U29668 ( .A(nreg[420]), .B(n28218), .Z(n28221) );
  XNOR U29669 ( .A(n19563), .B(n28218), .Z(n28220) );
  XOR U29670 ( .A(n28222), .B(n28223), .Z(n19563) );
  XOR U29671 ( .A(n28224), .B(n28225), .Z(n28218) );
  AND U29672 ( .A(n28226), .B(n28227), .Z(n28225) );
  XOR U29673 ( .A(nreg[419]), .B(n28224), .Z(n28227) );
  XNOR U29674 ( .A(n19575), .B(n28224), .Z(n28226) );
  XOR U29675 ( .A(n28228), .B(n28229), .Z(n19575) );
  XOR U29676 ( .A(n28230), .B(n28231), .Z(n28224) );
  AND U29677 ( .A(n28232), .B(n28233), .Z(n28231) );
  XOR U29678 ( .A(nreg[418]), .B(n28230), .Z(n28233) );
  XNOR U29679 ( .A(n19587), .B(n28230), .Z(n28232) );
  XOR U29680 ( .A(n28234), .B(n28235), .Z(n19587) );
  XOR U29681 ( .A(n28236), .B(n28237), .Z(n28230) );
  AND U29682 ( .A(n28238), .B(n28239), .Z(n28237) );
  XOR U29683 ( .A(nreg[417]), .B(n28236), .Z(n28239) );
  XNOR U29684 ( .A(n19599), .B(n28236), .Z(n28238) );
  XOR U29685 ( .A(n28240), .B(n28241), .Z(n19599) );
  XOR U29686 ( .A(n28242), .B(n28243), .Z(n28236) );
  AND U29687 ( .A(n28244), .B(n28245), .Z(n28243) );
  XOR U29688 ( .A(nreg[416]), .B(n28242), .Z(n28245) );
  XNOR U29689 ( .A(n19611), .B(n28242), .Z(n28244) );
  XOR U29690 ( .A(n28246), .B(n28247), .Z(n19611) );
  XOR U29691 ( .A(n28248), .B(n28249), .Z(n28242) );
  AND U29692 ( .A(n28250), .B(n28251), .Z(n28249) );
  XOR U29693 ( .A(nreg[415]), .B(n28248), .Z(n28251) );
  XNOR U29694 ( .A(n19623), .B(n28248), .Z(n28250) );
  XOR U29695 ( .A(n28252), .B(n28253), .Z(n19623) );
  XOR U29696 ( .A(n28254), .B(n28255), .Z(n28248) );
  AND U29697 ( .A(n28256), .B(n28257), .Z(n28255) );
  XOR U29698 ( .A(nreg[414]), .B(n28254), .Z(n28257) );
  XNOR U29699 ( .A(n19635), .B(n28254), .Z(n28256) );
  XOR U29700 ( .A(n28258), .B(n28259), .Z(n19635) );
  XOR U29701 ( .A(n28260), .B(n28261), .Z(n28254) );
  AND U29702 ( .A(n28262), .B(n28263), .Z(n28261) );
  XOR U29703 ( .A(nreg[413]), .B(n28260), .Z(n28263) );
  XNOR U29704 ( .A(n19647), .B(n28260), .Z(n28262) );
  XOR U29705 ( .A(n28264), .B(n28265), .Z(n19647) );
  XOR U29706 ( .A(n28266), .B(n28267), .Z(n28260) );
  AND U29707 ( .A(n28268), .B(n28269), .Z(n28267) );
  XOR U29708 ( .A(nreg[412]), .B(n28266), .Z(n28269) );
  XNOR U29709 ( .A(n19659), .B(n28266), .Z(n28268) );
  XOR U29710 ( .A(n28270), .B(n28271), .Z(n19659) );
  XOR U29711 ( .A(n28272), .B(n28273), .Z(n28266) );
  AND U29712 ( .A(n28274), .B(n28275), .Z(n28273) );
  XOR U29713 ( .A(nreg[411]), .B(n28272), .Z(n28275) );
  XNOR U29714 ( .A(n19671), .B(n28272), .Z(n28274) );
  XOR U29715 ( .A(n28276), .B(n28277), .Z(n19671) );
  XOR U29716 ( .A(n28278), .B(n28279), .Z(n28272) );
  AND U29717 ( .A(n28280), .B(n28281), .Z(n28279) );
  XOR U29718 ( .A(nreg[410]), .B(n28278), .Z(n28281) );
  XNOR U29719 ( .A(n19683), .B(n28278), .Z(n28280) );
  XOR U29720 ( .A(n28282), .B(n28283), .Z(n19683) );
  XOR U29721 ( .A(n28284), .B(n28285), .Z(n28278) );
  AND U29722 ( .A(n28286), .B(n28287), .Z(n28285) );
  XOR U29723 ( .A(nreg[409]), .B(n28284), .Z(n28287) );
  XNOR U29724 ( .A(n19695), .B(n28284), .Z(n28286) );
  XOR U29725 ( .A(n28288), .B(n28289), .Z(n19695) );
  XOR U29726 ( .A(n28290), .B(n28291), .Z(n28284) );
  AND U29727 ( .A(n28292), .B(n28293), .Z(n28291) );
  XOR U29728 ( .A(nreg[408]), .B(n28290), .Z(n28293) );
  XNOR U29729 ( .A(n19707), .B(n28290), .Z(n28292) );
  XOR U29730 ( .A(n28294), .B(n28295), .Z(n19707) );
  XOR U29731 ( .A(n28296), .B(n28297), .Z(n28290) );
  AND U29732 ( .A(n28298), .B(n28299), .Z(n28297) );
  XOR U29733 ( .A(nreg[407]), .B(n28296), .Z(n28299) );
  XNOR U29734 ( .A(n19719), .B(n28296), .Z(n28298) );
  XOR U29735 ( .A(n28300), .B(n28301), .Z(n19719) );
  XOR U29736 ( .A(n28302), .B(n28303), .Z(n28296) );
  AND U29737 ( .A(n28304), .B(n28305), .Z(n28303) );
  XOR U29738 ( .A(nreg[406]), .B(n28302), .Z(n28305) );
  XNOR U29739 ( .A(n19731), .B(n28302), .Z(n28304) );
  XOR U29740 ( .A(n28306), .B(n28307), .Z(n19731) );
  XOR U29741 ( .A(n28308), .B(n28309), .Z(n28302) );
  AND U29742 ( .A(n28310), .B(n28311), .Z(n28309) );
  XOR U29743 ( .A(nreg[405]), .B(n28308), .Z(n28311) );
  XNOR U29744 ( .A(n19743), .B(n28308), .Z(n28310) );
  XOR U29745 ( .A(n28312), .B(n28313), .Z(n19743) );
  XOR U29746 ( .A(n28314), .B(n28315), .Z(n28308) );
  AND U29747 ( .A(n28316), .B(n28317), .Z(n28315) );
  XOR U29748 ( .A(nreg[404]), .B(n28314), .Z(n28317) );
  XNOR U29749 ( .A(n19755), .B(n28314), .Z(n28316) );
  XOR U29750 ( .A(n28318), .B(n28319), .Z(n19755) );
  XOR U29751 ( .A(n28320), .B(n28321), .Z(n28314) );
  AND U29752 ( .A(n28322), .B(n28323), .Z(n28321) );
  XOR U29753 ( .A(nreg[403]), .B(n28320), .Z(n28323) );
  XNOR U29754 ( .A(n19767), .B(n28320), .Z(n28322) );
  XOR U29755 ( .A(n28324), .B(n28325), .Z(n19767) );
  XOR U29756 ( .A(n28326), .B(n28327), .Z(n28320) );
  AND U29757 ( .A(n28328), .B(n28329), .Z(n28327) );
  XOR U29758 ( .A(nreg[402]), .B(n28326), .Z(n28329) );
  XNOR U29759 ( .A(n19779), .B(n28326), .Z(n28328) );
  XOR U29760 ( .A(n28330), .B(n28331), .Z(n19779) );
  XOR U29761 ( .A(n28332), .B(n28333), .Z(n28326) );
  AND U29762 ( .A(n28334), .B(n28335), .Z(n28333) );
  XOR U29763 ( .A(nreg[401]), .B(n28332), .Z(n28335) );
  XNOR U29764 ( .A(n19791), .B(n28332), .Z(n28334) );
  XOR U29765 ( .A(n28336), .B(n28337), .Z(n19791) );
  XOR U29766 ( .A(n28338), .B(n28339), .Z(n28332) );
  AND U29767 ( .A(n28340), .B(n28341), .Z(n28339) );
  XOR U29768 ( .A(nreg[400]), .B(n28338), .Z(n28341) );
  XNOR U29769 ( .A(n19803), .B(n28338), .Z(n28340) );
  XOR U29770 ( .A(n28342), .B(n28343), .Z(n19803) );
  XOR U29771 ( .A(n28344), .B(n28345), .Z(n28338) );
  AND U29772 ( .A(n28346), .B(n28347), .Z(n28345) );
  XOR U29773 ( .A(nreg[399]), .B(n28344), .Z(n28347) );
  XNOR U29774 ( .A(n19815), .B(n28344), .Z(n28346) );
  XOR U29775 ( .A(n28348), .B(n28349), .Z(n19815) );
  XOR U29776 ( .A(n28350), .B(n28351), .Z(n28344) );
  AND U29777 ( .A(n28352), .B(n28353), .Z(n28351) );
  XOR U29778 ( .A(nreg[398]), .B(n28350), .Z(n28353) );
  XNOR U29779 ( .A(n19827), .B(n28350), .Z(n28352) );
  XOR U29780 ( .A(n28354), .B(n28355), .Z(n19827) );
  XOR U29781 ( .A(n28356), .B(n28357), .Z(n28350) );
  AND U29782 ( .A(n28358), .B(n28359), .Z(n28357) );
  XOR U29783 ( .A(nreg[397]), .B(n28356), .Z(n28359) );
  XNOR U29784 ( .A(n19839), .B(n28356), .Z(n28358) );
  XOR U29785 ( .A(n28360), .B(n28361), .Z(n19839) );
  XOR U29786 ( .A(n28362), .B(n28363), .Z(n28356) );
  AND U29787 ( .A(n28364), .B(n28365), .Z(n28363) );
  XOR U29788 ( .A(nreg[396]), .B(n28362), .Z(n28365) );
  XNOR U29789 ( .A(n19851), .B(n28362), .Z(n28364) );
  XOR U29790 ( .A(n28366), .B(n28367), .Z(n19851) );
  XOR U29791 ( .A(n28368), .B(n28369), .Z(n28362) );
  AND U29792 ( .A(n28370), .B(n28371), .Z(n28369) );
  XOR U29793 ( .A(nreg[395]), .B(n28368), .Z(n28371) );
  XNOR U29794 ( .A(n19863), .B(n28368), .Z(n28370) );
  XOR U29795 ( .A(n28372), .B(n28373), .Z(n19863) );
  XOR U29796 ( .A(n28374), .B(n28375), .Z(n28368) );
  AND U29797 ( .A(n28376), .B(n28377), .Z(n28375) );
  XOR U29798 ( .A(nreg[394]), .B(n28374), .Z(n28377) );
  XNOR U29799 ( .A(n19875), .B(n28374), .Z(n28376) );
  XOR U29800 ( .A(n28378), .B(n28379), .Z(n19875) );
  XOR U29801 ( .A(n28380), .B(n28381), .Z(n28374) );
  AND U29802 ( .A(n28382), .B(n28383), .Z(n28381) );
  XOR U29803 ( .A(nreg[393]), .B(n28380), .Z(n28383) );
  XNOR U29804 ( .A(n19887), .B(n28380), .Z(n28382) );
  XOR U29805 ( .A(n28384), .B(n28385), .Z(n19887) );
  XOR U29806 ( .A(n28386), .B(n28387), .Z(n28380) );
  AND U29807 ( .A(n28388), .B(n28389), .Z(n28387) );
  XOR U29808 ( .A(nreg[392]), .B(n28386), .Z(n28389) );
  XNOR U29809 ( .A(n19899), .B(n28386), .Z(n28388) );
  XOR U29810 ( .A(n28390), .B(n28391), .Z(n19899) );
  XOR U29811 ( .A(n28392), .B(n28393), .Z(n28386) );
  AND U29812 ( .A(n28394), .B(n28395), .Z(n28393) );
  XOR U29813 ( .A(nreg[391]), .B(n28392), .Z(n28395) );
  XNOR U29814 ( .A(n19911), .B(n28392), .Z(n28394) );
  XOR U29815 ( .A(n28396), .B(n28397), .Z(n19911) );
  XOR U29816 ( .A(n28398), .B(n28399), .Z(n28392) );
  AND U29817 ( .A(n28400), .B(n28401), .Z(n28399) );
  XOR U29818 ( .A(nreg[390]), .B(n28398), .Z(n28401) );
  XNOR U29819 ( .A(n19923), .B(n28398), .Z(n28400) );
  XOR U29820 ( .A(n28402), .B(n28403), .Z(n19923) );
  XOR U29821 ( .A(n28404), .B(n28405), .Z(n28398) );
  AND U29822 ( .A(n28406), .B(n28407), .Z(n28405) );
  XOR U29823 ( .A(nreg[389]), .B(n28404), .Z(n28407) );
  XNOR U29824 ( .A(n19935), .B(n28404), .Z(n28406) );
  XOR U29825 ( .A(n28408), .B(n28409), .Z(n19935) );
  XOR U29826 ( .A(n28410), .B(n28411), .Z(n28404) );
  AND U29827 ( .A(n28412), .B(n28413), .Z(n28411) );
  XOR U29828 ( .A(nreg[388]), .B(n28410), .Z(n28413) );
  XNOR U29829 ( .A(n19947), .B(n28410), .Z(n28412) );
  XOR U29830 ( .A(n28414), .B(n28415), .Z(n19947) );
  XOR U29831 ( .A(n28416), .B(n28417), .Z(n28410) );
  AND U29832 ( .A(n28418), .B(n28419), .Z(n28417) );
  XOR U29833 ( .A(nreg[387]), .B(n28416), .Z(n28419) );
  XNOR U29834 ( .A(n19959), .B(n28416), .Z(n28418) );
  XOR U29835 ( .A(n28420), .B(n28421), .Z(n19959) );
  XOR U29836 ( .A(n28422), .B(n28423), .Z(n28416) );
  AND U29837 ( .A(n28424), .B(n28425), .Z(n28423) );
  XOR U29838 ( .A(nreg[386]), .B(n28422), .Z(n28425) );
  XNOR U29839 ( .A(n19971), .B(n28422), .Z(n28424) );
  XOR U29840 ( .A(n28426), .B(n28427), .Z(n19971) );
  XOR U29841 ( .A(n28428), .B(n28429), .Z(n28422) );
  AND U29842 ( .A(n28430), .B(n28431), .Z(n28429) );
  XOR U29843 ( .A(nreg[385]), .B(n28428), .Z(n28431) );
  XNOR U29844 ( .A(n19983), .B(n28428), .Z(n28430) );
  XOR U29845 ( .A(n28432), .B(n28433), .Z(n19983) );
  XOR U29846 ( .A(n28434), .B(n28435), .Z(n28428) );
  AND U29847 ( .A(n28436), .B(n28437), .Z(n28435) );
  XOR U29848 ( .A(nreg[384]), .B(n28434), .Z(n28437) );
  XNOR U29849 ( .A(n19995), .B(n28434), .Z(n28436) );
  XOR U29850 ( .A(n28438), .B(n28439), .Z(n19995) );
  XOR U29851 ( .A(n28440), .B(n28441), .Z(n28434) );
  AND U29852 ( .A(n28442), .B(n28443), .Z(n28441) );
  XOR U29853 ( .A(nreg[383]), .B(n28440), .Z(n28443) );
  XNOR U29854 ( .A(n20007), .B(n28440), .Z(n28442) );
  XOR U29855 ( .A(n28444), .B(n28445), .Z(n20007) );
  XOR U29856 ( .A(n28446), .B(n28447), .Z(n28440) );
  AND U29857 ( .A(n28448), .B(n28449), .Z(n28447) );
  XOR U29858 ( .A(nreg[382]), .B(n28446), .Z(n28449) );
  XNOR U29859 ( .A(n20019), .B(n28446), .Z(n28448) );
  XOR U29860 ( .A(n28450), .B(n28451), .Z(n20019) );
  XOR U29861 ( .A(n28452), .B(n28453), .Z(n28446) );
  AND U29862 ( .A(n28454), .B(n28455), .Z(n28453) );
  XOR U29863 ( .A(nreg[381]), .B(n28452), .Z(n28455) );
  XNOR U29864 ( .A(n20031), .B(n28452), .Z(n28454) );
  XOR U29865 ( .A(n28456), .B(n28457), .Z(n20031) );
  XOR U29866 ( .A(n28458), .B(n28459), .Z(n28452) );
  AND U29867 ( .A(n28460), .B(n28461), .Z(n28459) );
  XOR U29868 ( .A(nreg[380]), .B(n28458), .Z(n28461) );
  XNOR U29869 ( .A(n20043), .B(n28458), .Z(n28460) );
  XOR U29870 ( .A(n28462), .B(n28463), .Z(n20043) );
  XOR U29871 ( .A(n28464), .B(n28465), .Z(n28458) );
  AND U29872 ( .A(n28466), .B(n28467), .Z(n28465) );
  XOR U29873 ( .A(nreg[379]), .B(n28464), .Z(n28467) );
  XNOR U29874 ( .A(n20055), .B(n28464), .Z(n28466) );
  XOR U29875 ( .A(n28468), .B(n28469), .Z(n20055) );
  XOR U29876 ( .A(n28470), .B(n28471), .Z(n28464) );
  AND U29877 ( .A(n28472), .B(n28473), .Z(n28471) );
  XOR U29878 ( .A(nreg[378]), .B(n28470), .Z(n28473) );
  XNOR U29879 ( .A(n20067), .B(n28470), .Z(n28472) );
  XOR U29880 ( .A(n28474), .B(n28475), .Z(n20067) );
  XOR U29881 ( .A(n28476), .B(n28477), .Z(n28470) );
  AND U29882 ( .A(n28478), .B(n28479), .Z(n28477) );
  XOR U29883 ( .A(nreg[377]), .B(n28476), .Z(n28479) );
  XNOR U29884 ( .A(n20079), .B(n28476), .Z(n28478) );
  XOR U29885 ( .A(n28480), .B(n28481), .Z(n20079) );
  XOR U29886 ( .A(n28482), .B(n28483), .Z(n28476) );
  AND U29887 ( .A(n28484), .B(n28485), .Z(n28483) );
  XOR U29888 ( .A(nreg[376]), .B(n28482), .Z(n28485) );
  XNOR U29889 ( .A(n20091), .B(n28482), .Z(n28484) );
  XOR U29890 ( .A(n28486), .B(n28487), .Z(n20091) );
  XOR U29891 ( .A(n28488), .B(n28489), .Z(n28482) );
  AND U29892 ( .A(n28490), .B(n28491), .Z(n28489) );
  XOR U29893 ( .A(nreg[375]), .B(n28488), .Z(n28491) );
  XNOR U29894 ( .A(n20103), .B(n28488), .Z(n28490) );
  XOR U29895 ( .A(n28492), .B(n28493), .Z(n20103) );
  XOR U29896 ( .A(n28494), .B(n28495), .Z(n28488) );
  AND U29897 ( .A(n28496), .B(n28497), .Z(n28495) );
  XOR U29898 ( .A(nreg[374]), .B(n28494), .Z(n28497) );
  XNOR U29899 ( .A(n20115), .B(n28494), .Z(n28496) );
  XOR U29900 ( .A(n28498), .B(n28499), .Z(n20115) );
  XOR U29901 ( .A(n28500), .B(n28501), .Z(n28494) );
  AND U29902 ( .A(n28502), .B(n28503), .Z(n28501) );
  XOR U29903 ( .A(nreg[373]), .B(n28500), .Z(n28503) );
  XNOR U29904 ( .A(n20127), .B(n28500), .Z(n28502) );
  XOR U29905 ( .A(n28504), .B(n28505), .Z(n20127) );
  XOR U29906 ( .A(n28506), .B(n28507), .Z(n28500) );
  AND U29907 ( .A(n28508), .B(n28509), .Z(n28507) );
  XOR U29908 ( .A(nreg[372]), .B(n28506), .Z(n28509) );
  XNOR U29909 ( .A(n20139), .B(n28506), .Z(n28508) );
  XOR U29910 ( .A(n28510), .B(n28511), .Z(n20139) );
  XOR U29911 ( .A(n28512), .B(n28513), .Z(n28506) );
  AND U29912 ( .A(n28514), .B(n28515), .Z(n28513) );
  XOR U29913 ( .A(nreg[371]), .B(n28512), .Z(n28515) );
  XNOR U29914 ( .A(n20151), .B(n28512), .Z(n28514) );
  XOR U29915 ( .A(n28516), .B(n28517), .Z(n20151) );
  XOR U29916 ( .A(n28518), .B(n28519), .Z(n28512) );
  AND U29917 ( .A(n28520), .B(n28521), .Z(n28519) );
  XOR U29918 ( .A(nreg[370]), .B(n28518), .Z(n28521) );
  XNOR U29919 ( .A(n20163), .B(n28518), .Z(n28520) );
  XOR U29920 ( .A(n28522), .B(n28523), .Z(n20163) );
  XOR U29921 ( .A(n28524), .B(n28525), .Z(n28518) );
  AND U29922 ( .A(n28526), .B(n28527), .Z(n28525) );
  XOR U29923 ( .A(nreg[369]), .B(n28524), .Z(n28527) );
  XNOR U29924 ( .A(n20175), .B(n28524), .Z(n28526) );
  XOR U29925 ( .A(n28528), .B(n28529), .Z(n20175) );
  XOR U29926 ( .A(n28530), .B(n28531), .Z(n28524) );
  AND U29927 ( .A(n28532), .B(n28533), .Z(n28531) );
  XOR U29928 ( .A(nreg[368]), .B(n28530), .Z(n28533) );
  XNOR U29929 ( .A(n20187), .B(n28530), .Z(n28532) );
  XOR U29930 ( .A(n28534), .B(n28535), .Z(n20187) );
  XOR U29931 ( .A(n28536), .B(n28537), .Z(n28530) );
  AND U29932 ( .A(n28538), .B(n28539), .Z(n28537) );
  XOR U29933 ( .A(nreg[367]), .B(n28536), .Z(n28539) );
  XNOR U29934 ( .A(n20199), .B(n28536), .Z(n28538) );
  XOR U29935 ( .A(n28540), .B(n28541), .Z(n20199) );
  XOR U29936 ( .A(n28542), .B(n28543), .Z(n28536) );
  AND U29937 ( .A(n28544), .B(n28545), .Z(n28543) );
  XOR U29938 ( .A(nreg[366]), .B(n28542), .Z(n28545) );
  XNOR U29939 ( .A(n20211), .B(n28542), .Z(n28544) );
  XOR U29940 ( .A(n28546), .B(n28547), .Z(n20211) );
  XOR U29941 ( .A(n28548), .B(n28549), .Z(n28542) );
  AND U29942 ( .A(n28550), .B(n28551), .Z(n28549) );
  XOR U29943 ( .A(nreg[365]), .B(n28548), .Z(n28551) );
  XNOR U29944 ( .A(n20223), .B(n28548), .Z(n28550) );
  XOR U29945 ( .A(n28552), .B(n28553), .Z(n20223) );
  XOR U29946 ( .A(n28554), .B(n28555), .Z(n28548) );
  AND U29947 ( .A(n28556), .B(n28557), .Z(n28555) );
  XOR U29948 ( .A(nreg[364]), .B(n28554), .Z(n28557) );
  XNOR U29949 ( .A(n20235), .B(n28554), .Z(n28556) );
  XOR U29950 ( .A(n28558), .B(n28559), .Z(n20235) );
  XOR U29951 ( .A(n28560), .B(n28561), .Z(n28554) );
  AND U29952 ( .A(n28562), .B(n28563), .Z(n28561) );
  XOR U29953 ( .A(nreg[363]), .B(n28560), .Z(n28563) );
  XNOR U29954 ( .A(n20247), .B(n28560), .Z(n28562) );
  XOR U29955 ( .A(n28564), .B(n28565), .Z(n20247) );
  XOR U29956 ( .A(n28566), .B(n28567), .Z(n28560) );
  AND U29957 ( .A(n28568), .B(n28569), .Z(n28567) );
  XOR U29958 ( .A(nreg[362]), .B(n28566), .Z(n28569) );
  XNOR U29959 ( .A(n20259), .B(n28566), .Z(n28568) );
  XOR U29960 ( .A(n28570), .B(n28571), .Z(n20259) );
  XOR U29961 ( .A(n28572), .B(n28573), .Z(n28566) );
  AND U29962 ( .A(n28574), .B(n28575), .Z(n28573) );
  XOR U29963 ( .A(nreg[361]), .B(n28572), .Z(n28575) );
  XNOR U29964 ( .A(n20271), .B(n28572), .Z(n28574) );
  XOR U29965 ( .A(n28576), .B(n28577), .Z(n20271) );
  XOR U29966 ( .A(n28578), .B(n28579), .Z(n28572) );
  AND U29967 ( .A(n28580), .B(n28581), .Z(n28579) );
  XOR U29968 ( .A(nreg[360]), .B(n28578), .Z(n28581) );
  XNOR U29969 ( .A(n20283), .B(n28578), .Z(n28580) );
  XOR U29970 ( .A(n28582), .B(n28583), .Z(n20283) );
  XOR U29971 ( .A(n28584), .B(n28585), .Z(n28578) );
  AND U29972 ( .A(n28586), .B(n28587), .Z(n28585) );
  XOR U29973 ( .A(nreg[359]), .B(n28584), .Z(n28587) );
  XNOR U29974 ( .A(n20295), .B(n28584), .Z(n28586) );
  XOR U29975 ( .A(n28588), .B(n28589), .Z(n20295) );
  XOR U29976 ( .A(n28590), .B(n28591), .Z(n28584) );
  AND U29977 ( .A(n28592), .B(n28593), .Z(n28591) );
  XOR U29978 ( .A(nreg[358]), .B(n28590), .Z(n28593) );
  XNOR U29979 ( .A(n20307), .B(n28590), .Z(n28592) );
  XOR U29980 ( .A(n28594), .B(n28595), .Z(n20307) );
  XOR U29981 ( .A(n28596), .B(n28597), .Z(n28590) );
  AND U29982 ( .A(n28598), .B(n28599), .Z(n28597) );
  XOR U29983 ( .A(nreg[357]), .B(n28596), .Z(n28599) );
  XNOR U29984 ( .A(n20319), .B(n28596), .Z(n28598) );
  XOR U29985 ( .A(n28600), .B(n28601), .Z(n20319) );
  XOR U29986 ( .A(n28602), .B(n28603), .Z(n28596) );
  AND U29987 ( .A(n28604), .B(n28605), .Z(n28603) );
  XOR U29988 ( .A(nreg[356]), .B(n28602), .Z(n28605) );
  XNOR U29989 ( .A(n20331), .B(n28602), .Z(n28604) );
  XOR U29990 ( .A(n28606), .B(n28607), .Z(n20331) );
  XOR U29991 ( .A(n28608), .B(n28609), .Z(n28602) );
  AND U29992 ( .A(n28610), .B(n28611), .Z(n28609) );
  XOR U29993 ( .A(nreg[355]), .B(n28608), .Z(n28611) );
  XNOR U29994 ( .A(n20343), .B(n28608), .Z(n28610) );
  XOR U29995 ( .A(n28612), .B(n28613), .Z(n20343) );
  XOR U29996 ( .A(n28614), .B(n28615), .Z(n28608) );
  AND U29997 ( .A(n28616), .B(n28617), .Z(n28615) );
  XOR U29998 ( .A(nreg[354]), .B(n28614), .Z(n28617) );
  XNOR U29999 ( .A(n20355), .B(n28614), .Z(n28616) );
  XOR U30000 ( .A(n28618), .B(n28619), .Z(n20355) );
  XOR U30001 ( .A(n28620), .B(n28621), .Z(n28614) );
  AND U30002 ( .A(n28622), .B(n28623), .Z(n28621) );
  XOR U30003 ( .A(nreg[353]), .B(n28620), .Z(n28623) );
  XNOR U30004 ( .A(n20367), .B(n28620), .Z(n28622) );
  XOR U30005 ( .A(n28624), .B(n28625), .Z(n20367) );
  XOR U30006 ( .A(n28626), .B(n28627), .Z(n28620) );
  AND U30007 ( .A(n28628), .B(n28629), .Z(n28627) );
  XOR U30008 ( .A(nreg[352]), .B(n28626), .Z(n28629) );
  XNOR U30009 ( .A(n20379), .B(n28626), .Z(n28628) );
  XOR U30010 ( .A(n28630), .B(n28631), .Z(n20379) );
  XOR U30011 ( .A(n28632), .B(n28633), .Z(n28626) );
  AND U30012 ( .A(n28634), .B(n28635), .Z(n28633) );
  XOR U30013 ( .A(nreg[351]), .B(n28632), .Z(n28635) );
  XNOR U30014 ( .A(n20391), .B(n28632), .Z(n28634) );
  XOR U30015 ( .A(n28636), .B(n28637), .Z(n20391) );
  XOR U30016 ( .A(n28638), .B(n28639), .Z(n28632) );
  AND U30017 ( .A(n28640), .B(n28641), .Z(n28639) );
  XOR U30018 ( .A(nreg[350]), .B(n28638), .Z(n28641) );
  XNOR U30019 ( .A(n20403), .B(n28638), .Z(n28640) );
  XOR U30020 ( .A(n28642), .B(n28643), .Z(n20403) );
  XOR U30021 ( .A(n28644), .B(n28645), .Z(n28638) );
  AND U30022 ( .A(n28646), .B(n28647), .Z(n28645) );
  XOR U30023 ( .A(nreg[349]), .B(n28644), .Z(n28647) );
  XNOR U30024 ( .A(n20415), .B(n28644), .Z(n28646) );
  XOR U30025 ( .A(n28648), .B(n28649), .Z(n20415) );
  XOR U30026 ( .A(n28650), .B(n28651), .Z(n28644) );
  AND U30027 ( .A(n28652), .B(n28653), .Z(n28651) );
  XOR U30028 ( .A(nreg[348]), .B(n28650), .Z(n28653) );
  XNOR U30029 ( .A(n20427), .B(n28650), .Z(n28652) );
  XOR U30030 ( .A(n28654), .B(n28655), .Z(n20427) );
  XOR U30031 ( .A(n28656), .B(n28657), .Z(n28650) );
  AND U30032 ( .A(n28658), .B(n28659), .Z(n28657) );
  XOR U30033 ( .A(nreg[347]), .B(n28656), .Z(n28659) );
  XNOR U30034 ( .A(n20439), .B(n28656), .Z(n28658) );
  XOR U30035 ( .A(n28660), .B(n28661), .Z(n20439) );
  XOR U30036 ( .A(n28662), .B(n28663), .Z(n28656) );
  AND U30037 ( .A(n28664), .B(n28665), .Z(n28663) );
  XOR U30038 ( .A(nreg[346]), .B(n28662), .Z(n28665) );
  XNOR U30039 ( .A(n20451), .B(n28662), .Z(n28664) );
  XOR U30040 ( .A(n28666), .B(n28667), .Z(n20451) );
  XOR U30041 ( .A(n28668), .B(n28669), .Z(n28662) );
  AND U30042 ( .A(n28670), .B(n28671), .Z(n28669) );
  XOR U30043 ( .A(nreg[345]), .B(n28668), .Z(n28671) );
  XNOR U30044 ( .A(n20463), .B(n28668), .Z(n28670) );
  XOR U30045 ( .A(n28672), .B(n28673), .Z(n20463) );
  XOR U30046 ( .A(n28674), .B(n28675), .Z(n28668) );
  AND U30047 ( .A(n28676), .B(n28677), .Z(n28675) );
  XOR U30048 ( .A(nreg[344]), .B(n28674), .Z(n28677) );
  XNOR U30049 ( .A(n20475), .B(n28674), .Z(n28676) );
  XOR U30050 ( .A(n28678), .B(n28679), .Z(n20475) );
  XOR U30051 ( .A(n28680), .B(n28681), .Z(n28674) );
  AND U30052 ( .A(n28682), .B(n28683), .Z(n28681) );
  XOR U30053 ( .A(nreg[343]), .B(n28680), .Z(n28683) );
  XNOR U30054 ( .A(n20487), .B(n28680), .Z(n28682) );
  XOR U30055 ( .A(n28684), .B(n28685), .Z(n20487) );
  XOR U30056 ( .A(n28686), .B(n28687), .Z(n28680) );
  AND U30057 ( .A(n28688), .B(n28689), .Z(n28687) );
  XOR U30058 ( .A(nreg[342]), .B(n28686), .Z(n28689) );
  XNOR U30059 ( .A(n20499), .B(n28686), .Z(n28688) );
  XOR U30060 ( .A(n28690), .B(n28691), .Z(n20499) );
  XOR U30061 ( .A(n28692), .B(n28693), .Z(n28686) );
  AND U30062 ( .A(n28694), .B(n28695), .Z(n28693) );
  XOR U30063 ( .A(nreg[341]), .B(n28692), .Z(n28695) );
  XNOR U30064 ( .A(n20511), .B(n28692), .Z(n28694) );
  XOR U30065 ( .A(n28696), .B(n28697), .Z(n20511) );
  XOR U30066 ( .A(n28698), .B(n28699), .Z(n28692) );
  AND U30067 ( .A(n28700), .B(n28701), .Z(n28699) );
  XOR U30068 ( .A(nreg[340]), .B(n28698), .Z(n28701) );
  XNOR U30069 ( .A(n20523), .B(n28698), .Z(n28700) );
  XOR U30070 ( .A(n28702), .B(n28703), .Z(n20523) );
  XOR U30071 ( .A(n28704), .B(n28705), .Z(n28698) );
  AND U30072 ( .A(n28706), .B(n28707), .Z(n28705) );
  XOR U30073 ( .A(nreg[339]), .B(n28704), .Z(n28707) );
  XNOR U30074 ( .A(n20535), .B(n28704), .Z(n28706) );
  XOR U30075 ( .A(n28708), .B(n28709), .Z(n20535) );
  XOR U30076 ( .A(n28710), .B(n28711), .Z(n28704) );
  AND U30077 ( .A(n28712), .B(n28713), .Z(n28711) );
  XOR U30078 ( .A(nreg[338]), .B(n28710), .Z(n28713) );
  XNOR U30079 ( .A(n20547), .B(n28710), .Z(n28712) );
  XOR U30080 ( .A(n28714), .B(n28715), .Z(n20547) );
  XOR U30081 ( .A(n28716), .B(n28717), .Z(n28710) );
  AND U30082 ( .A(n28718), .B(n28719), .Z(n28717) );
  XOR U30083 ( .A(nreg[337]), .B(n28716), .Z(n28719) );
  XNOR U30084 ( .A(n20559), .B(n28716), .Z(n28718) );
  XOR U30085 ( .A(n28720), .B(n28721), .Z(n20559) );
  XOR U30086 ( .A(n28722), .B(n28723), .Z(n28716) );
  AND U30087 ( .A(n28724), .B(n28725), .Z(n28723) );
  XOR U30088 ( .A(nreg[336]), .B(n28722), .Z(n28725) );
  XNOR U30089 ( .A(n20571), .B(n28722), .Z(n28724) );
  XOR U30090 ( .A(n28726), .B(n28727), .Z(n20571) );
  XOR U30091 ( .A(n28728), .B(n28729), .Z(n28722) );
  AND U30092 ( .A(n28730), .B(n28731), .Z(n28729) );
  XOR U30093 ( .A(nreg[335]), .B(n28728), .Z(n28731) );
  XNOR U30094 ( .A(n20583), .B(n28728), .Z(n28730) );
  XOR U30095 ( .A(n28732), .B(n28733), .Z(n20583) );
  XOR U30096 ( .A(n28734), .B(n28735), .Z(n28728) );
  AND U30097 ( .A(n28736), .B(n28737), .Z(n28735) );
  XOR U30098 ( .A(nreg[334]), .B(n28734), .Z(n28737) );
  XNOR U30099 ( .A(n20595), .B(n28734), .Z(n28736) );
  XOR U30100 ( .A(n28738), .B(n28739), .Z(n20595) );
  XOR U30101 ( .A(n28740), .B(n28741), .Z(n28734) );
  AND U30102 ( .A(n28742), .B(n28743), .Z(n28741) );
  XOR U30103 ( .A(nreg[333]), .B(n28740), .Z(n28743) );
  XNOR U30104 ( .A(n20607), .B(n28740), .Z(n28742) );
  XOR U30105 ( .A(n28744), .B(n28745), .Z(n20607) );
  XOR U30106 ( .A(n28746), .B(n28747), .Z(n28740) );
  AND U30107 ( .A(n28748), .B(n28749), .Z(n28747) );
  XOR U30108 ( .A(nreg[332]), .B(n28746), .Z(n28749) );
  XNOR U30109 ( .A(n20619), .B(n28746), .Z(n28748) );
  XOR U30110 ( .A(n28750), .B(n28751), .Z(n20619) );
  XOR U30111 ( .A(n28752), .B(n28753), .Z(n28746) );
  AND U30112 ( .A(n28754), .B(n28755), .Z(n28753) );
  XOR U30113 ( .A(nreg[331]), .B(n28752), .Z(n28755) );
  XNOR U30114 ( .A(n20631), .B(n28752), .Z(n28754) );
  XOR U30115 ( .A(n28756), .B(n28757), .Z(n20631) );
  XOR U30116 ( .A(n28758), .B(n28759), .Z(n28752) );
  AND U30117 ( .A(n28760), .B(n28761), .Z(n28759) );
  XOR U30118 ( .A(nreg[330]), .B(n28758), .Z(n28761) );
  XNOR U30119 ( .A(n20643), .B(n28758), .Z(n28760) );
  XOR U30120 ( .A(n28762), .B(n28763), .Z(n20643) );
  XOR U30121 ( .A(n28764), .B(n28765), .Z(n28758) );
  AND U30122 ( .A(n28766), .B(n28767), .Z(n28765) );
  XOR U30123 ( .A(nreg[329]), .B(n28764), .Z(n28767) );
  XNOR U30124 ( .A(n20655), .B(n28764), .Z(n28766) );
  XOR U30125 ( .A(n28768), .B(n28769), .Z(n20655) );
  XOR U30126 ( .A(n28770), .B(n28771), .Z(n28764) );
  AND U30127 ( .A(n28772), .B(n28773), .Z(n28771) );
  XOR U30128 ( .A(nreg[328]), .B(n28770), .Z(n28773) );
  XNOR U30129 ( .A(n20667), .B(n28770), .Z(n28772) );
  XOR U30130 ( .A(n28774), .B(n28775), .Z(n20667) );
  XOR U30131 ( .A(n28776), .B(n28777), .Z(n28770) );
  AND U30132 ( .A(n28778), .B(n28779), .Z(n28777) );
  XOR U30133 ( .A(nreg[327]), .B(n28776), .Z(n28779) );
  XNOR U30134 ( .A(n20679), .B(n28776), .Z(n28778) );
  XOR U30135 ( .A(n28780), .B(n28781), .Z(n20679) );
  XOR U30136 ( .A(n28782), .B(n28783), .Z(n28776) );
  AND U30137 ( .A(n28784), .B(n28785), .Z(n28783) );
  XOR U30138 ( .A(nreg[326]), .B(n28782), .Z(n28785) );
  XNOR U30139 ( .A(n20691), .B(n28782), .Z(n28784) );
  XOR U30140 ( .A(n28786), .B(n28787), .Z(n20691) );
  XOR U30141 ( .A(n28788), .B(n28789), .Z(n28782) );
  AND U30142 ( .A(n28790), .B(n28791), .Z(n28789) );
  XOR U30143 ( .A(nreg[325]), .B(n28788), .Z(n28791) );
  XNOR U30144 ( .A(n20703), .B(n28788), .Z(n28790) );
  XOR U30145 ( .A(n28792), .B(n28793), .Z(n20703) );
  XOR U30146 ( .A(n28794), .B(n28795), .Z(n28788) );
  AND U30147 ( .A(n28796), .B(n28797), .Z(n28795) );
  XOR U30148 ( .A(nreg[324]), .B(n28794), .Z(n28797) );
  XNOR U30149 ( .A(n20715), .B(n28794), .Z(n28796) );
  XOR U30150 ( .A(n28798), .B(n28799), .Z(n20715) );
  XOR U30151 ( .A(n28800), .B(n28801), .Z(n28794) );
  AND U30152 ( .A(n28802), .B(n28803), .Z(n28801) );
  XOR U30153 ( .A(nreg[323]), .B(n28800), .Z(n28803) );
  XNOR U30154 ( .A(n20727), .B(n28800), .Z(n28802) );
  XOR U30155 ( .A(n28804), .B(n28805), .Z(n20727) );
  XOR U30156 ( .A(n28806), .B(n28807), .Z(n28800) );
  AND U30157 ( .A(n28808), .B(n28809), .Z(n28807) );
  XOR U30158 ( .A(nreg[322]), .B(n28806), .Z(n28809) );
  XNOR U30159 ( .A(n20739), .B(n28806), .Z(n28808) );
  XOR U30160 ( .A(n28810), .B(n28811), .Z(n20739) );
  XOR U30161 ( .A(n28812), .B(n28813), .Z(n28806) );
  AND U30162 ( .A(n28814), .B(n28815), .Z(n28813) );
  XOR U30163 ( .A(nreg[321]), .B(n28812), .Z(n28815) );
  XNOR U30164 ( .A(n20751), .B(n28812), .Z(n28814) );
  XOR U30165 ( .A(n28816), .B(n28817), .Z(n20751) );
  XOR U30166 ( .A(n28818), .B(n28819), .Z(n28812) );
  AND U30167 ( .A(n28820), .B(n28821), .Z(n28819) );
  XOR U30168 ( .A(nreg[320]), .B(n28818), .Z(n28821) );
  XNOR U30169 ( .A(n20763), .B(n28818), .Z(n28820) );
  XOR U30170 ( .A(n28822), .B(n28823), .Z(n20763) );
  XOR U30171 ( .A(n28824), .B(n28825), .Z(n28818) );
  AND U30172 ( .A(n28826), .B(n28827), .Z(n28825) );
  XOR U30173 ( .A(nreg[319]), .B(n28824), .Z(n28827) );
  XNOR U30174 ( .A(n20775), .B(n28824), .Z(n28826) );
  XOR U30175 ( .A(n28828), .B(n28829), .Z(n20775) );
  XOR U30176 ( .A(n28830), .B(n28831), .Z(n28824) );
  AND U30177 ( .A(n28832), .B(n28833), .Z(n28831) );
  XOR U30178 ( .A(nreg[318]), .B(n28830), .Z(n28833) );
  XNOR U30179 ( .A(n20787), .B(n28830), .Z(n28832) );
  XOR U30180 ( .A(n28834), .B(n28835), .Z(n20787) );
  XOR U30181 ( .A(n28836), .B(n28837), .Z(n28830) );
  AND U30182 ( .A(n28838), .B(n28839), .Z(n28837) );
  XOR U30183 ( .A(nreg[317]), .B(n28836), .Z(n28839) );
  XNOR U30184 ( .A(n20799), .B(n28836), .Z(n28838) );
  XOR U30185 ( .A(n28840), .B(n28841), .Z(n20799) );
  XOR U30186 ( .A(n28842), .B(n28843), .Z(n28836) );
  AND U30187 ( .A(n28844), .B(n28845), .Z(n28843) );
  XOR U30188 ( .A(nreg[316]), .B(n28842), .Z(n28845) );
  XNOR U30189 ( .A(n20811), .B(n28842), .Z(n28844) );
  XOR U30190 ( .A(n28846), .B(n28847), .Z(n20811) );
  XOR U30191 ( .A(n28848), .B(n28849), .Z(n28842) );
  AND U30192 ( .A(n28850), .B(n28851), .Z(n28849) );
  XOR U30193 ( .A(nreg[315]), .B(n28848), .Z(n28851) );
  XNOR U30194 ( .A(n20823), .B(n28848), .Z(n28850) );
  XOR U30195 ( .A(n28852), .B(n28853), .Z(n20823) );
  XOR U30196 ( .A(n28854), .B(n28855), .Z(n28848) );
  AND U30197 ( .A(n28856), .B(n28857), .Z(n28855) );
  XOR U30198 ( .A(nreg[314]), .B(n28854), .Z(n28857) );
  XNOR U30199 ( .A(n20835), .B(n28854), .Z(n28856) );
  XOR U30200 ( .A(n28858), .B(n28859), .Z(n20835) );
  XOR U30201 ( .A(n28860), .B(n28861), .Z(n28854) );
  AND U30202 ( .A(n28862), .B(n28863), .Z(n28861) );
  XOR U30203 ( .A(nreg[313]), .B(n28860), .Z(n28863) );
  XNOR U30204 ( .A(n20847), .B(n28860), .Z(n28862) );
  XOR U30205 ( .A(n28864), .B(n28865), .Z(n20847) );
  XOR U30206 ( .A(n28866), .B(n28867), .Z(n28860) );
  AND U30207 ( .A(n28868), .B(n28869), .Z(n28867) );
  XOR U30208 ( .A(nreg[312]), .B(n28866), .Z(n28869) );
  XNOR U30209 ( .A(n20859), .B(n28866), .Z(n28868) );
  XOR U30210 ( .A(n28870), .B(n28871), .Z(n20859) );
  XOR U30211 ( .A(n28872), .B(n28873), .Z(n28866) );
  AND U30212 ( .A(n28874), .B(n28875), .Z(n28873) );
  XOR U30213 ( .A(nreg[311]), .B(n28872), .Z(n28875) );
  XNOR U30214 ( .A(n20871), .B(n28872), .Z(n28874) );
  XOR U30215 ( .A(n28876), .B(n28877), .Z(n20871) );
  XOR U30216 ( .A(n28878), .B(n28879), .Z(n28872) );
  AND U30217 ( .A(n28880), .B(n28881), .Z(n28879) );
  XOR U30218 ( .A(nreg[310]), .B(n28878), .Z(n28881) );
  XNOR U30219 ( .A(n20883), .B(n28878), .Z(n28880) );
  XOR U30220 ( .A(n28882), .B(n28883), .Z(n20883) );
  XOR U30221 ( .A(n28884), .B(n28885), .Z(n28878) );
  AND U30222 ( .A(n28886), .B(n28887), .Z(n28885) );
  XOR U30223 ( .A(nreg[309]), .B(n28884), .Z(n28887) );
  XNOR U30224 ( .A(n20895), .B(n28884), .Z(n28886) );
  XOR U30225 ( .A(n28888), .B(n28889), .Z(n20895) );
  XOR U30226 ( .A(n28890), .B(n28891), .Z(n28884) );
  AND U30227 ( .A(n28892), .B(n28893), .Z(n28891) );
  XOR U30228 ( .A(nreg[308]), .B(n28890), .Z(n28893) );
  XNOR U30229 ( .A(n20907), .B(n28890), .Z(n28892) );
  XOR U30230 ( .A(n28894), .B(n28895), .Z(n20907) );
  XOR U30231 ( .A(n28896), .B(n28897), .Z(n28890) );
  AND U30232 ( .A(n28898), .B(n28899), .Z(n28897) );
  XOR U30233 ( .A(nreg[307]), .B(n28896), .Z(n28899) );
  XNOR U30234 ( .A(n20919), .B(n28896), .Z(n28898) );
  XOR U30235 ( .A(n28900), .B(n28901), .Z(n20919) );
  XOR U30236 ( .A(n28902), .B(n28903), .Z(n28896) );
  AND U30237 ( .A(n28904), .B(n28905), .Z(n28903) );
  XOR U30238 ( .A(nreg[306]), .B(n28902), .Z(n28905) );
  XNOR U30239 ( .A(n20931), .B(n28902), .Z(n28904) );
  XOR U30240 ( .A(n28906), .B(n28907), .Z(n20931) );
  XOR U30241 ( .A(n28908), .B(n28909), .Z(n28902) );
  AND U30242 ( .A(n28910), .B(n28911), .Z(n28909) );
  XOR U30243 ( .A(nreg[305]), .B(n28908), .Z(n28911) );
  XNOR U30244 ( .A(n20943), .B(n28908), .Z(n28910) );
  XOR U30245 ( .A(n28912), .B(n28913), .Z(n20943) );
  XOR U30246 ( .A(n28914), .B(n28915), .Z(n28908) );
  AND U30247 ( .A(n28916), .B(n28917), .Z(n28915) );
  XOR U30248 ( .A(nreg[304]), .B(n28914), .Z(n28917) );
  XNOR U30249 ( .A(n20955), .B(n28914), .Z(n28916) );
  XOR U30250 ( .A(n28918), .B(n28919), .Z(n20955) );
  XOR U30251 ( .A(n28920), .B(n28921), .Z(n28914) );
  AND U30252 ( .A(n28922), .B(n28923), .Z(n28921) );
  XOR U30253 ( .A(nreg[303]), .B(n28920), .Z(n28923) );
  XNOR U30254 ( .A(n20967), .B(n28920), .Z(n28922) );
  XOR U30255 ( .A(n28924), .B(n28925), .Z(n20967) );
  XOR U30256 ( .A(n28926), .B(n28927), .Z(n28920) );
  AND U30257 ( .A(n28928), .B(n28929), .Z(n28927) );
  XOR U30258 ( .A(nreg[302]), .B(n28926), .Z(n28929) );
  XNOR U30259 ( .A(n20979), .B(n28926), .Z(n28928) );
  XOR U30260 ( .A(n28930), .B(n28931), .Z(n20979) );
  XOR U30261 ( .A(n28932), .B(n28933), .Z(n28926) );
  AND U30262 ( .A(n28934), .B(n28935), .Z(n28933) );
  XOR U30263 ( .A(nreg[301]), .B(n28932), .Z(n28935) );
  XNOR U30264 ( .A(n20991), .B(n28932), .Z(n28934) );
  XOR U30265 ( .A(n28936), .B(n28937), .Z(n20991) );
  XOR U30266 ( .A(n28938), .B(n28939), .Z(n28932) );
  AND U30267 ( .A(n28940), .B(n28941), .Z(n28939) );
  XOR U30268 ( .A(nreg[300]), .B(n28938), .Z(n28941) );
  XNOR U30269 ( .A(n21003), .B(n28938), .Z(n28940) );
  XOR U30270 ( .A(n28942), .B(n28943), .Z(n21003) );
  XOR U30271 ( .A(n28944), .B(n28945), .Z(n28938) );
  AND U30272 ( .A(n28946), .B(n28947), .Z(n28945) );
  XOR U30273 ( .A(nreg[299]), .B(n28944), .Z(n28947) );
  XNOR U30274 ( .A(n21015), .B(n28944), .Z(n28946) );
  XOR U30275 ( .A(n28948), .B(n28949), .Z(n21015) );
  XOR U30276 ( .A(n28950), .B(n28951), .Z(n28944) );
  AND U30277 ( .A(n28952), .B(n28953), .Z(n28951) );
  XOR U30278 ( .A(nreg[298]), .B(n28950), .Z(n28953) );
  XNOR U30279 ( .A(n21027), .B(n28950), .Z(n28952) );
  XOR U30280 ( .A(n28954), .B(n28955), .Z(n21027) );
  XOR U30281 ( .A(n28956), .B(n28957), .Z(n28950) );
  AND U30282 ( .A(n28958), .B(n28959), .Z(n28957) );
  XOR U30283 ( .A(nreg[297]), .B(n28956), .Z(n28959) );
  XNOR U30284 ( .A(n21039), .B(n28956), .Z(n28958) );
  XOR U30285 ( .A(n28960), .B(n28961), .Z(n21039) );
  XOR U30286 ( .A(n28962), .B(n28963), .Z(n28956) );
  AND U30287 ( .A(n28964), .B(n28965), .Z(n28963) );
  XOR U30288 ( .A(nreg[296]), .B(n28962), .Z(n28965) );
  XNOR U30289 ( .A(n21051), .B(n28962), .Z(n28964) );
  XOR U30290 ( .A(n28966), .B(n28967), .Z(n21051) );
  XOR U30291 ( .A(n28968), .B(n28969), .Z(n28962) );
  AND U30292 ( .A(n28970), .B(n28971), .Z(n28969) );
  XOR U30293 ( .A(nreg[295]), .B(n28968), .Z(n28971) );
  XNOR U30294 ( .A(n21063), .B(n28968), .Z(n28970) );
  XOR U30295 ( .A(n28972), .B(n28973), .Z(n21063) );
  XOR U30296 ( .A(n28974), .B(n28975), .Z(n28968) );
  AND U30297 ( .A(n28976), .B(n28977), .Z(n28975) );
  XOR U30298 ( .A(nreg[294]), .B(n28974), .Z(n28977) );
  XNOR U30299 ( .A(n21075), .B(n28974), .Z(n28976) );
  XOR U30300 ( .A(n28978), .B(n28979), .Z(n21075) );
  XOR U30301 ( .A(n28980), .B(n28981), .Z(n28974) );
  AND U30302 ( .A(n28982), .B(n28983), .Z(n28981) );
  XOR U30303 ( .A(nreg[293]), .B(n28980), .Z(n28983) );
  XNOR U30304 ( .A(n21087), .B(n28980), .Z(n28982) );
  XOR U30305 ( .A(n28984), .B(n28985), .Z(n21087) );
  XOR U30306 ( .A(n28986), .B(n28987), .Z(n28980) );
  AND U30307 ( .A(n28988), .B(n28989), .Z(n28987) );
  XOR U30308 ( .A(nreg[292]), .B(n28986), .Z(n28989) );
  XNOR U30309 ( .A(n21099), .B(n28986), .Z(n28988) );
  XOR U30310 ( .A(n28990), .B(n28991), .Z(n21099) );
  XOR U30311 ( .A(n28992), .B(n28993), .Z(n28986) );
  AND U30312 ( .A(n28994), .B(n28995), .Z(n28993) );
  XOR U30313 ( .A(nreg[291]), .B(n28992), .Z(n28995) );
  XNOR U30314 ( .A(n21111), .B(n28992), .Z(n28994) );
  XOR U30315 ( .A(n28996), .B(n28997), .Z(n21111) );
  XOR U30316 ( .A(n28998), .B(n28999), .Z(n28992) );
  AND U30317 ( .A(n29000), .B(n29001), .Z(n28999) );
  XOR U30318 ( .A(nreg[290]), .B(n28998), .Z(n29001) );
  XNOR U30319 ( .A(n21123), .B(n28998), .Z(n29000) );
  XOR U30320 ( .A(n29002), .B(n29003), .Z(n21123) );
  XOR U30321 ( .A(n29004), .B(n29005), .Z(n28998) );
  AND U30322 ( .A(n29006), .B(n29007), .Z(n29005) );
  XOR U30323 ( .A(nreg[289]), .B(n29004), .Z(n29007) );
  XNOR U30324 ( .A(n21135), .B(n29004), .Z(n29006) );
  XOR U30325 ( .A(n29008), .B(n29009), .Z(n21135) );
  XOR U30326 ( .A(n29010), .B(n29011), .Z(n29004) );
  AND U30327 ( .A(n29012), .B(n29013), .Z(n29011) );
  XOR U30328 ( .A(nreg[288]), .B(n29010), .Z(n29013) );
  XNOR U30329 ( .A(n21147), .B(n29010), .Z(n29012) );
  XOR U30330 ( .A(n29014), .B(n29015), .Z(n21147) );
  XOR U30331 ( .A(n29016), .B(n29017), .Z(n29010) );
  AND U30332 ( .A(n29018), .B(n29019), .Z(n29017) );
  XOR U30333 ( .A(nreg[287]), .B(n29016), .Z(n29019) );
  XNOR U30334 ( .A(n21159), .B(n29016), .Z(n29018) );
  XOR U30335 ( .A(n29020), .B(n29021), .Z(n21159) );
  XOR U30336 ( .A(n29022), .B(n29023), .Z(n29016) );
  AND U30337 ( .A(n29024), .B(n29025), .Z(n29023) );
  XOR U30338 ( .A(nreg[286]), .B(n29022), .Z(n29025) );
  XNOR U30339 ( .A(n21171), .B(n29022), .Z(n29024) );
  XOR U30340 ( .A(n29026), .B(n29027), .Z(n21171) );
  XOR U30341 ( .A(n29028), .B(n29029), .Z(n29022) );
  AND U30342 ( .A(n29030), .B(n29031), .Z(n29029) );
  XOR U30343 ( .A(nreg[285]), .B(n29028), .Z(n29031) );
  XNOR U30344 ( .A(n21183), .B(n29028), .Z(n29030) );
  XOR U30345 ( .A(n29032), .B(n29033), .Z(n21183) );
  XOR U30346 ( .A(n29034), .B(n29035), .Z(n29028) );
  AND U30347 ( .A(n29036), .B(n29037), .Z(n29035) );
  XOR U30348 ( .A(nreg[284]), .B(n29034), .Z(n29037) );
  XNOR U30349 ( .A(n21195), .B(n29034), .Z(n29036) );
  XOR U30350 ( .A(n29038), .B(n29039), .Z(n21195) );
  XOR U30351 ( .A(n29040), .B(n29041), .Z(n29034) );
  AND U30352 ( .A(n29042), .B(n29043), .Z(n29041) );
  XOR U30353 ( .A(nreg[283]), .B(n29040), .Z(n29043) );
  XNOR U30354 ( .A(n21207), .B(n29040), .Z(n29042) );
  XOR U30355 ( .A(n29044), .B(n29045), .Z(n21207) );
  XOR U30356 ( .A(n29046), .B(n29047), .Z(n29040) );
  AND U30357 ( .A(n29048), .B(n29049), .Z(n29047) );
  XOR U30358 ( .A(nreg[282]), .B(n29046), .Z(n29049) );
  XNOR U30359 ( .A(n21219), .B(n29046), .Z(n29048) );
  XOR U30360 ( .A(n29050), .B(n29051), .Z(n21219) );
  XOR U30361 ( .A(n29052), .B(n29053), .Z(n29046) );
  AND U30362 ( .A(n29054), .B(n29055), .Z(n29053) );
  XOR U30363 ( .A(nreg[281]), .B(n29052), .Z(n29055) );
  XNOR U30364 ( .A(n21231), .B(n29052), .Z(n29054) );
  XOR U30365 ( .A(n29056), .B(n29057), .Z(n21231) );
  XOR U30366 ( .A(n29058), .B(n29059), .Z(n29052) );
  AND U30367 ( .A(n29060), .B(n29061), .Z(n29059) );
  XOR U30368 ( .A(nreg[280]), .B(n29058), .Z(n29061) );
  XNOR U30369 ( .A(n21243), .B(n29058), .Z(n29060) );
  XOR U30370 ( .A(n29062), .B(n29063), .Z(n21243) );
  XOR U30371 ( .A(n29064), .B(n29065), .Z(n29058) );
  AND U30372 ( .A(n29066), .B(n29067), .Z(n29065) );
  XOR U30373 ( .A(nreg[279]), .B(n29064), .Z(n29067) );
  XNOR U30374 ( .A(n21255), .B(n29064), .Z(n29066) );
  XOR U30375 ( .A(n29068), .B(n29069), .Z(n21255) );
  XOR U30376 ( .A(n29070), .B(n29071), .Z(n29064) );
  AND U30377 ( .A(n29072), .B(n29073), .Z(n29071) );
  XOR U30378 ( .A(nreg[278]), .B(n29070), .Z(n29073) );
  XNOR U30379 ( .A(n21267), .B(n29070), .Z(n29072) );
  XOR U30380 ( .A(n29074), .B(n29075), .Z(n21267) );
  XOR U30381 ( .A(n29076), .B(n29077), .Z(n29070) );
  AND U30382 ( .A(n29078), .B(n29079), .Z(n29077) );
  XOR U30383 ( .A(nreg[277]), .B(n29076), .Z(n29079) );
  XNOR U30384 ( .A(n21279), .B(n29076), .Z(n29078) );
  XOR U30385 ( .A(n29080), .B(n29081), .Z(n21279) );
  XOR U30386 ( .A(n29082), .B(n29083), .Z(n29076) );
  AND U30387 ( .A(n29084), .B(n29085), .Z(n29083) );
  XOR U30388 ( .A(nreg[276]), .B(n29082), .Z(n29085) );
  XNOR U30389 ( .A(n21291), .B(n29082), .Z(n29084) );
  XOR U30390 ( .A(n29086), .B(n29087), .Z(n21291) );
  XOR U30391 ( .A(n29088), .B(n29089), .Z(n29082) );
  AND U30392 ( .A(n29090), .B(n29091), .Z(n29089) );
  XOR U30393 ( .A(nreg[275]), .B(n29088), .Z(n29091) );
  XNOR U30394 ( .A(n21303), .B(n29088), .Z(n29090) );
  XOR U30395 ( .A(n29092), .B(n29093), .Z(n21303) );
  XOR U30396 ( .A(n29094), .B(n29095), .Z(n29088) );
  AND U30397 ( .A(n29096), .B(n29097), .Z(n29095) );
  XOR U30398 ( .A(nreg[274]), .B(n29094), .Z(n29097) );
  XNOR U30399 ( .A(n21315), .B(n29094), .Z(n29096) );
  XOR U30400 ( .A(n29098), .B(n29099), .Z(n21315) );
  XOR U30401 ( .A(n29100), .B(n29101), .Z(n29094) );
  AND U30402 ( .A(n29102), .B(n29103), .Z(n29101) );
  XOR U30403 ( .A(nreg[273]), .B(n29100), .Z(n29103) );
  XNOR U30404 ( .A(n21327), .B(n29100), .Z(n29102) );
  XOR U30405 ( .A(n29104), .B(n29105), .Z(n21327) );
  XOR U30406 ( .A(n29106), .B(n29107), .Z(n29100) );
  AND U30407 ( .A(n29108), .B(n29109), .Z(n29107) );
  XOR U30408 ( .A(nreg[272]), .B(n29106), .Z(n29109) );
  XNOR U30409 ( .A(n21339), .B(n29106), .Z(n29108) );
  XOR U30410 ( .A(n29110), .B(n29111), .Z(n21339) );
  XOR U30411 ( .A(n29112), .B(n29113), .Z(n29106) );
  AND U30412 ( .A(n29114), .B(n29115), .Z(n29113) );
  XOR U30413 ( .A(nreg[271]), .B(n29112), .Z(n29115) );
  XNOR U30414 ( .A(n21351), .B(n29112), .Z(n29114) );
  XOR U30415 ( .A(n29116), .B(n29117), .Z(n21351) );
  XOR U30416 ( .A(n29118), .B(n29119), .Z(n29112) );
  AND U30417 ( .A(n29120), .B(n29121), .Z(n29119) );
  XOR U30418 ( .A(nreg[270]), .B(n29118), .Z(n29121) );
  XNOR U30419 ( .A(n21363), .B(n29118), .Z(n29120) );
  XOR U30420 ( .A(n29122), .B(n29123), .Z(n21363) );
  XOR U30421 ( .A(n29124), .B(n29125), .Z(n29118) );
  AND U30422 ( .A(n29126), .B(n29127), .Z(n29125) );
  XOR U30423 ( .A(nreg[269]), .B(n29124), .Z(n29127) );
  XNOR U30424 ( .A(n21375), .B(n29124), .Z(n29126) );
  XOR U30425 ( .A(n29128), .B(n29129), .Z(n21375) );
  XOR U30426 ( .A(n29130), .B(n29131), .Z(n29124) );
  AND U30427 ( .A(n29132), .B(n29133), .Z(n29131) );
  XOR U30428 ( .A(nreg[268]), .B(n29130), .Z(n29133) );
  XNOR U30429 ( .A(n21387), .B(n29130), .Z(n29132) );
  XOR U30430 ( .A(n29134), .B(n29135), .Z(n21387) );
  XOR U30431 ( .A(n29136), .B(n29137), .Z(n29130) );
  AND U30432 ( .A(n29138), .B(n29139), .Z(n29137) );
  XOR U30433 ( .A(nreg[267]), .B(n29136), .Z(n29139) );
  XNOR U30434 ( .A(n21399), .B(n29136), .Z(n29138) );
  XOR U30435 ( .A(n29140), .B(n29141), .Z(n21399) );
  XOR U30436 ( .A(n29142), .B(n29143), .Z(n29136) );
  AND U30437 ( .A(n29144), .B(n29145), .Z(n29143) );
  XOR U30438 ( .A(nreg[266]), .B(n29142), .Z(n29145) );
  XNOR U30439 ( .A(n21411), .B(n29142), .Z(n29144) );
  XOR U30440 ( .A(n29146), .B(n29147), .Z(n21411) );
  XOR U30441 ( .A(n29148), .B(n29149), .Z(n29142) );
  AND U30442 ( .A(n29150), .B(n29151), .Z(n29149) );
  XOR U30443 ( .A(nreg[265]), .B(n29148), .Z(n29151) );
  XNOR U30444 ( .A(n21423), .B(n29148), .Z(n29150) );
  XOR U30445 ( .A(n29152), .B(n29153), .Z(n21423) );
  XOR U30446 ( .A(n29154), .B(n29155), .Z(n29148) );
  AND U30447 ( .A(n29156), .B(n29157), .Z(n29155) );
  XOR U30448 ( .A(nreg[264]), .B(n29154), .Z(n29157) );
  XNOR U30449 ( .A(n21435), .B(n29154), .Z(n29156) );
  XOR U30450 ( .A(n29158), .B(n29159), .Z(n21435) );
  XOR U30451 ( .A(n29160), .B(n29161), .Z(n29154) );
  AND U30452 ( .A(n29162), .B(n29163), .Z(n29161) );
  XOR U30453 ( .A(nreg[263]), .B(n29160), .Z(n29163) );
  XNOR U30454 ( .A(n21447), .B(n29160), .Z(n29162) );
  XOR U30455 ( .A(n29164), .B(n29165), .Z(n21447) );
  XOR U30456 ( .A(n29166), .B(n29167), .Z(n29160) );
  AND U30457 ( .A(n29168), .B(n29169), .Z(n29167) );
  XOR U30458 ( .A(nreg[262]), .B(n29166), .Z(n29169) );
  XNOR U30459 ( .A(n21459), .B(n29166), .Z(n29168) );
  XOR U30460 ( .A(n29170), .B(n29171), .Z(n21459) );
  XOR U30461 ( .A(n29172), .B(n29173), .Z(n29166) );
  AND U30462 ( .A(n29174), .B(n29175), .Z(n29173) );
  XOR U30463 ( .A(nreg[261]), .B(n29172), .Z(n29175) );
  XNOR U30464 ( .A(n21471), .B(n29172), .Z(n29174) );
  XOR U30465 ( .A(n29176), .B(n29177), .Z(n21471) );
  XOR U30466 ( .A(n29178), .B(n29179), .Z(n29172) );
  AND U30467 ( .A(n29180), .B(n29181), .Z(n29179) );
  XOR U30468 ( .A(nreg[260]), .B(n29178), .Z(n29181) );
  XNOR U30469 ( .A(n21483), .B(n29178), .Z(n29180) );
  XOR U30470 ( .A(n29182), .B(n29183), .Z(n21483) );
  XOR U30471 ( .A(n29184), .B(n29185), .Z(n29178) );
  AND U30472 ( .A(n29186), .B(n29187), .Z(n29185) );
  XOR U30473 ( .A(nreg[259]), .B(n29184), .Z(n29187) );
  XNOR U30474 ( .A(n21495), .B(n29184), .Z(n29186) );
  XOR U30475 ( .A(n29188), .B(n29189), .Z(n21495) );
  XOR U30476 ( .A(n29190), .B(n29191), .Z(n29184) );
  AND U30477 ( .A(n29192), .B(n29193), .Z(n29191) );
  XOR U30478 ( .A(nreg[258]), .B(n29190), .Z(n29193) );
  XNOR U30479 ( .A(n21507), .B(n29190), .Z(n29192) );
  XOR U30480 ( .A(n29194), .B(n29195), .Z(n21507) );
  XOR U30481 ( .A(n29196), .B(n29197), .Z(n29190) );
  AND U30482 ( .A(n29198), .B(n29199), .Z(n29197) );
  XOR U30483 ( .A(nreg[257]), .B(n29196), .Z(n29199) );
  XNOR U30484 ( .A(n21519), .B(n29196), .Z(n29198) );
  XOR U30485 ( .A(n29200), .B(n29201), .Z(n21519) );
  XOR U30486 ( .A(n29202), .B(n29203), .Z(n29196) );
  AND U30487 ( .A(n29204), .B(n29205), .Z(n29203) );
  XOR U30488 ( .A(nreg[256]), .B(n29202), .Z(n29205) );
  XNOR U30489 ( .A(n21531), .B(n29202), .Z(n29204) );
  XOR U30490 ( .A(n29206), .B(n29207), .Z(n21531) );
  XOR U30491 ( .A(n29208), .B(n29209), .Z(n29202) );
  AND U30492 ( .A(n29210), .B(n29211), .Z(n29209) );
  XOR U30493 ( .A(nreg[255]), .B(n29208), .Z(n29211) );
  XNOR U30494 ( .A(n21543), .B(n29208), .Z(n29210) );
  XOR U30495 ( .A(n29212), .B(n29213), .Z(n21543) );
  XOR U30496 ( .A(n29214), .B(n29215), .Z(n29208) );
  AND U30497 ( .A(n29216), .B(n29217), .Z(n29215) );
  XOR U30498 ( .A(nreg[254]), .B(n29214), .Z(n29217) );
  XNOR U30499 ( .A(n21555), .B(n29214), .Z(n29216) );
  XOR U30500 ( .A(n29218), .B(n29219), .Z(n21555) );
  XOR U30501 ( .A(n29220), .B(n29221), .Z(n29214) );
  AND U30502 ( .A(n29222), .B(n29223), .Z(n29221) );
  XOR U30503 ( .A(nreg[253]), .B(n29220), .Z(n29223) );
  XNOR U30504 ( .A(n21567), .B(n29220), .Z(n29222) );
  XOR U30505 ( .A(n29224), .B(n29225), .Z(n21567) );
  XOR U30506 ( .A(n29226), .B(n29227), .Z(n29220) );
  AND U30507 ( .A(n29228), .B(n29229), .Z(n29227) );
  XOR U30508 ( .A(nreg[252]), .B(n29226), .Z(n29229) );
  XNOR U30509 ( .A(n21579), .B(n29226), .Z(n29228) );
  XOR U30510 ( .A(n29230), .B(n29231), .Z(n21579) );
  XOR U30511 ( .A(n29232), .B(n29233), .Z(n29226) );
  AND U30512 ( .A(n29234), .B(n29235), .Z(n29233) );
  XOR U30513 ( .A(nreg[251]), .B(n29232), .Z(n29235) );
  XNOR U30514 ( .A(n21591), .B(n29232), .Z(n29234) );
  XOR U30515 ( .A(n29236), .B(n29237), .Z(n21591) );
  XOR U30516 ( .A(n29238), .B(n29239), .Z(n29232) );
  AND U30517 ( .A(n29240), .B(n29241), .Z(n29239) );
  XOR U30518 ( .A(nreg[250]), .B(n29238), .Z(n29241) );
  XNOR U30519 ( .A(n21603), .B(n29238), .Z(n29240) );
  XOR U30520 ( .A(n29242), .B(n29243), .Z(n21603) );
  XOR U30521 ( .A(n29244), .B(n29245), .Z(n29238) );
  AND U30522 ( .A(n29246), .B(n29247), .Z(n29245) );
  XOR U30523 ( .A(nreg[249]), .B(n29244), .Z(n29247) );
  XNOR U30524 ( .A(n21615), .B(n29244), .Z(n29246) );
  XOR U30525 ( .A(n29248), .B(n29249), .Z(n21615) );
  XOR U30526 ( .A(n29250), .B(n29251), .Z(n29244) );
  AND U30527 ( .A(n29252), .B(n29253), .Z(n29251) );
  XOR U30528 ( .A(nreg[248]), .B(n29250), .Z(n29253) );
  XNOR U30529 ( .A(n21627), .B(n29250), .Z(n29252) );
  XOR U30530 ( .A(n29254), .B(n29255), .Z(n21627) );
  XOR U30531 ( .A(n29256), .B(n29257), .Z(n29250) );
  AND U30532 ( .A(n29258), .B(n29259), .Z(n29257) );
  XOR U30533 ( .A(nreg[247]), .B(n29256), .Z(n29259) );
  XNOR U30534 ( .A(n21639), .B(n29256), .Z(n29258) );
  XOR U30535 ( .A(n29260), .B(n29261), .Z(n21639) );
  XOR U30536 ( .A(n29262), .B(n29263), .Z(n29256) );
  AND U30537 ( .A(n29264), .B(n29265), .Z(n29263) );
  XOR U30538 ( .A(nreg[246]), .B(n29262), .Z(n29265) );
  XNOR U30539 ( .A(n21651), .B(n29262), .Z(n29264) );
  XOR U30540 ( .A(n29266), .B(n29267), .Z(n21651) );
  XOR U30541 ( .A(n29268), .B(n29269), .Z(n29262) );
  AND U30542 ( .A(n29270), .B(n29271), .Z(n29269) );
  XOR U30543 ( .A(nreg[245]), .B(n29268), .Z(n29271) );
  XNOR U30544 ( .A(n21663), .B(n29268), .Z(n29270) );
  XOR U30545 ( .A(n29272), .B(n29273), .Z(n21663) );
  XOR U30546 ( .A(n29274), .B(n29275), .Z(n29268) );
  AND U30547 ( .A(n29276), .B(n29277), .Z(n29275) );
  XOR U30548 ( .A(nreg[244]), .B(n29274), .Z(n29277) );
  XNOR U30549 ( .A(n21675), .B(n29274), .Z(n29276) );
  XOR U30550 ( .A(n29278), .B(n29279), .Z(n21675) );
  XOR U30551 ( .A(n29280), .B(n29281), .Z(n29274) );
  AND U30552 ( .A(n29282), .B(n29283), .Z(n29281) );
  XOR U30553 ( .A(nreg[243]), .B(n29280), .Z(n29283) );
  XNOR U30554 ( .A(n21687), .B(n29280), .Z(n29282) );
  XOR U30555 ( .A(n29284), .B(n29285), .Z(n21687) );
  XOR U30556 ( .A(n29286), .B(n29287), .Z(n29280) );
  AND U30557 ( .A(n29288), .B(n29289), .Z(n29287) );
  XOR U30558 ( .A(nreg[242]), .B(n29286), .Z(n29289) );
  XNOR U30559 ( .A(n21699), .B(n29286), .Z(n29288) );
  XOR U30560 ( .A(n29290), .B(n29291), .Z(n21699) );
  XOR U30561 ( .A(n29292), .B(n29293), .Z(n29286) );
  AND U30562 ( .A(n29294), .B(n29295), .Z(n29293) );
  XOR U30563 ( .A(nreg[241]), .B(n29292), .Z(n29295) );
  XNOR U30564 ( .A(n21711), .B(n29292), .Z(n29294) );
  XOR U30565 ( .A(n29296), .B(n29297), .Z(n21711) );
  XOR U30566 ( .A(n29298), .B(n29299), .Z(n29292) );
  AND U30567 ( .A(n29300), .B(n29301), .Z(n29299) );
  XOR U30568 ( .A(nreg[240]), .B(n29298), .Z(n29301) );
  XNOR U30569 ( .A(n21723), .B(n29298), .Z(n29300) );
  XOR U30570 ( .A(n29302), .B(n29303), .Z(n21723) );
  XOR U30571 ( .A(n29304), .B(n29305), .Z(n29298) );
  AND U30572 ( .A(n29306), .B(n29307), .Z(n29305) );
  XOR U30573 ( .A(nreg[239]), .B(n29304), .Z(n29307) );
  XNOR U30574 ( .A(n21735), .B(n29304), .Z(n29306) );
  XOR U30575 ( .A(n29308), .B(n29309), .Z(n21735) );
  XOR U30576 ( .A(n29310), .B(n29311), .Z(n29304) );
  AND U30577 ( .A(n29312), .B(n29313), .Z(n29311) );
  XOR U30578 ( .A(nreg[238]), .B(n29310), .Z(n29313) );
  XNOR U30579 ( .A(n21747), .B(n29310), .Z(n29312) );
  XOR U30580 ( .A(n29314), .B(n29315), .Z(n21747) );
  XOR U30581 ( .A(n29316), .B(n29317), .Z(n29310) );
  AND U30582 ( .A(n29318), .B(n29319), .Z(n29317) );
  XOR U30583 ( .A(nreg[237]), .B(n29316), .Z(n29319) );
  XNOR U30584 ( .A(n21759), .B(n29316), .Z(n29318) );
  XOR U30585 ( .A(n29320), .B(n29321), .Z(n21759) );
  XOR U30586 ( .A(n29322), .B(n29323), .Z(n29316) );
  AND U30587 ( .A(n29324), .B(n29325), .Z(n29323) );
  XOR U30588 ( .A(nreg[236]), .B(n29322), .Z(n29325) );
  XNOR U30589 ( .A(n21771), .B(n29322), .Z(n29324) );
  XOR U30590 ( .A(n29326), .B(n29327), .Z(n21771) );
  XOR U30591 ( .A(n29328), .B(n29329), .Z(n29322) );
  AND U30592 ( .A(n29330), .B(n29331), .Z(n29329) );
  XOR U30593 ( .A(nreg[235]), .B(n29328), .Z(n29331) );
  XNOR U30594 ( .A(n21783), .B(n29328), .Z(n29330) );
  XOR U30595 ( .A(n29332), .B(n29333), .Z(n21783) );
  XOR U30596 ( .A(n29334), .B(n29335), .Z(n29328) );
  AND U30597 ( .A(n29336), .B(n29337), .Z(n29335) );
  XOR U30598 ( .A(nreg[234]), .B(n29334), .Z(n29337) );
  XNOR U30599 ( .A(n21795), .B(n29334), .Z(n29336) );
  XOR U30600 ( .A(n29338), .B(n29339), .Z(n21795) );
  XOR U30601 ( .A(n29340), .B(n29341), .Z(n29334) );
  AND U30602 ( .A(n29342), .B(n29343), .Z(n29341) );
  XOR U30603 ( .A(nreg[233]), .B(n29340), .Z(n29343) );
  XNOR U30604 ( .A(n21807), .B(n29340), .Z(n29342) );
  XOR U30605 ( .A(n29344), .B(n29345), .Z(n21807) );
  XOR U30606 ( .A(n29346), .B(n29347), .Z(n29340) );
  AND U30607 ( .A(n29348), .B(n29349), .Z(n29347) );
  XOR U30608 ( .A(nreg[232]), .B(n29346), .Z(n29349) );
  XNOR U30609 ( .A(n21819), .B(n29346), .Z(n29348) );
  XOR U30610 ( .A(n29350), .B(n29351), .Z(n21819) );
  XOR U30611 ( .A(n29352), .B(n29353), .Z(n29346) );
  AND U30612 ( .A(n29354), .B(n29355), .Z(n29353) );
  XOR U30613 ( .A(nreg[231]), .B(n29352), .Z(n29355) );
  XNOR U30614 ( .A(n21831), .B(n29352), .Z(n29354) );
  XOR U30615 ( .A(n29356), .B(n29357), .Z(n21831) );
  XOR U30616 ( .A(n29358), .B(n29359), .Z(n29352) );
  AND U30617 ( .A(n29360), .B(n29361), .Z(n29359) );
  XOR U30618 ( .A(nreg[230]), .B(n29358), .Z(n29361) );
  XNOR U30619 ( .A(n21843), .B(n29358), .Z(n29360) );
  XOR U30620 ( .A(n29362), .B(n29363), .Z(n21843) );
  XOR U30621 ( .A(n29364), .B(n29365), .Z(n29358) );
  AND U30622 ( .A(n29366), .B(n29367), .Z(n29365) );
  XOR U30623 ( .A(nreg[229]), .B(n29364), .Z(n29367) );
  XNOR U30624 ( .A(n21855), .B(n29364), .Z(n29366) );
  XOR U30625 ( .A(n29368), .B(n29369), .Z(n21855) );
  XOR U30626 ( .A(n29370), .B(n29371), .Z(n29364) );
  AND U30627 ( .A(n29372), .B(n29373), .Z(n29371) );
  XOR U30628 ( .A(nreg[228]), .B(n29370), .Z(n29373) );
  XNOR U30629 ( .A(n21867), .B(n29370), .Z(n29372) );
  XOR U30630 ( .A(n29374), .B(n29375), .Z(n21867) );
  XOR U30631 ( .A(n29376), .B(n29377), .Z(n29370) );
  AND U30632 ( .A(n29378), .B(n29379), .Z(n29377) );
  XOR U30633 ( .A(nreg[227]), .B(n29376), .Z(n29379) );
  XNOR U30634 ( .A(n21879), .B(n29376), .Z(n29378) );
  XOR U30635 ( .A(n29380), .B(n29381), .Z(n21879) );
  XOR U30636 ( .A(n29382), .B(n29383), .Z(n29376) );
  AND U30637 ( .A(n29384), .B(n29385), .Z(n29383) );
  XOR U30638 ( .A(nreg[226]), .B(n29382), .Z(n29385) );
  XNOR U30639 ( .A(n21891), .B(n29382), .Z(n29384) );
  XOR U30640 ( .A(n29386), .B(n29387), .Z(n21891) );
  XOR U30641 ( .A(n29388), .B(n29389), .Z(n29382) );
  AND U30642 ( .A(n29390), .B(n29391), .Z(n29389) );
  XOR U30643 ( .A(nreg[225]), .B(n29388), .Z(n29391) );
  XNOR U30644 ( .A(n21903), .B(n29388), .Z(n29390) );
  XOR U30645 ( .A(n29392), .B(n29393), .Z(n21903) );
  XOR U30646 ( .A(n29394), .B(n29395), .Z(n29388) );
  AND U30647 ( .A(n29396), .B(n29397), .Z(n29395) );
  XOR U30648 ( .A(nreg[224]), .B(n29394), .Z(n29397) );
  XNOR U30649 ( .A(n21915), .B(n29394), .Z(n29396) );
  XOR U30650 ( .A(n29398), .B(n29399), .Z(n21915) );
  XOR U30651 ( .A(n29400), .B(n29401), .Z(n29394) );
  AND U30652 ( .A(n29402), .B(n29403), .Z(n29401) );
  XOR U30653 ( .A(nreg[223]), .B(n29400), .Z(n29403) );
  XNOR U30654 ( .A(n21927), .B(n29400), .Z(n29402) );
  XOR U30655 ( .A(n29404), .B(n29405), .Z(n21927) );
  XOR U30656 ( .A(n29406), .B(n29407), .Z(n29400) );
  AND U30657 ( .A(n29408), .B(n29409), .Z(n29407) );
  XOR U30658 ( .A(nreg[222]), .B(n29406), .Z(n29409) );
  XNOR U30659 ( .A(n21939), .B(n29406), .Z(n29408) );
  XOR U30660 ( .A(n29410), .B(n29411), .Z(n21939) );
  XOR U30661 ( .A(n29412), .B(n29413), .Z(n29406) );
  AND U30662 ( .A(n29414), .B(n29415), .Z(n29413) );
  XOR U30663 ( .A(nreg[221]), .B(n29412), .Z(n29415) );
  XNOR U30664 ( .A(n21951), .B(n29412), .Z(n29414) );
  XOR U30665 ( .A(n29416), .B(n29417), .Z(n21951) );
  XOR U30666 ( .A(n29418), .B(n29419), .Z(n29412) );
  AND U30667 ( .A(n29420), .B(n29421), .Z(n29419) );
  XOR U30668 ( .A(nreg[220]), .B(n29418), .Z(n29421) );
  XNOR U30669 ( .A(n21963), .B(n29418), .Z(n29420) );
  XOR U30670 ( .A(n29422), .B(n29423), .Z(n21963) );
  XOR U30671 ( .A(n29424), .B(n29425), .Z(n29418) );
  AND U30672 ( .A(n29426), .B(n29427), .Z(n29425) );
  XOR U30673 ( .A(nreg[219]), .B(n29424), .Z(n29427) );
  XNOR U30674 ( .A(n21975), .B(n29424), .Z(n29426) );
  XOR U30675 ( .A(n29428), .B(n29429), .Z(n21975) );
  XOR U30676 ( .A(n29430), .B(n29431), .Z(n29424) );
  AND U30677 ( .A(n29432), .B(n29433), .Z(n29431) );
  XOR U30678 ( .A(nreg[218]), .B(n29430), .Z(n29433) );
  XNOR U30679 ( .A(n21987), .B(n29430), .Z(n29432) );
  XOR U30680 ( .A(n29434), .B(n29435), .Z(n21987) );
  XOR U30681 ( .A(n29436), .B(n29437), .Z(n29430) );
  AND U30682 ( .A(n29438), .B(n29439), .Z(n29437) );
  XOR U30683 ( .A(nreg[217]), .B(n29436), .Z(n29439) );
  XNOR U30684 ( .A(n21999), .B(n29436), .Z(n29438) );
  XOR U30685 ( .A(n29440), .B(n29441), .Z(n21999) );
  XOR U30686 ( .A(n29442), .B(n29443), .Z(n29436) );
  AND U30687 ( .A(n29444), .B(n29445), .Z(n29443) );
  XOR U30688 ( .A(nreg[216]), .B(n29442), .Z(n29445) );
  XNOR U30689 ( .A(n22011), .B(n29442), .Z(n29444) );
  XOR U30690 ( .A(n29446), .B(n29447), .Z(n22011) );
  XOR U30691 ( .A(n29448), .B(n29449), .Z(n29442) );
  AND U30692 ( .A(n29450), .B(n29451), .Z(n29449) );
  XOR U30693 ( .A(nreg[215]), .B(n29448), .Z(n29451) );
  XNOR U30694 ( .A(n22023), .B(n29448), .Z(n29450) );
  XOR U30695 ( .A(n29452), .B(n29453), .Z(n22023) );
  XOR U30696 ( .A(n29454), .B(n29455), .Z(n29448) );
  AND U30697 ( .A(n29456), .B(n29457), .Z(n29455) );
  XOR U30698 ( .A(nreg[214]), .B(n29454), .Z(n29457) );
  XNOR U30699 ( .A(n22035), .B(n29454), .Z(n29456) );
  XOR U30700 ( .A(n29458), .B(n29459), .Z(n22035) );
  XOR U30701 ( .A(n29460), .B(n29461), .Z(n29454) );
  AND U30702 ( .A(n29462), .B(n29463), .Z(n29461) );
  XOR U30703 ( .A(nreg[213]), .B(n29460), .Z(n29463) );
  XNOR U30704 ( .A(n22047), .B(n29460), .Z(n29462) );
  XOR U30705 ( .A(n29464), .B(n29465), .Z(n22047) );
  XOR U30706 ( .A(n29466), .B(n29467), .Z(n29460) );
  AND U30707 ( .A(n29468), .B(n29469), .Z(n29467) );
  XOR U30708 ( .A(nreg[212]), .B(n29466), .Z(n29469) );
  XNOR U30709 ( .A(n22059), .B(n29466), .Z(n29468) );
  XOR U30710 ( .A(n29470), .B(n29471), .Z(n22059) );
  XOR U30711 ( .A(n29472), .B(n29473), .Z(n29466) );
  AND U30712 ( .A(n29474), .B(n29475), .Z(n29473) );
  XOR U30713 ( .A(nreg[211]), .B(n29472), .Z(n29475) );
  XNOR U30714 ( .A(n22071), .B(n29472), .Z(n29474) );
  XOR U30715 ( .A(n29476), .B(n29477), .Z(n22071) );
  XOR U30716 ( .A(n29478), .B(n29479), .Z(n29472) );
  AND U30717 ( .A(n29480), .B(n29481), .Z(n29479) );
  XOR U30718 ( .A(nreg[210]), .B(n29478), .Z(n29481) );
  XNOR U30719 ( .A(n22083), .B(n29478), .Z(n29480) );
  XOR U30720 ( .A(n29482), .B(n29483), .Z(n22083) );
  XOR U30721 ( .A(n29484), .B(n29485), .Z(n29478) );
  AND U30722 ( .A(n29486), .B(n29487), .Z(n29485) );
  XOR U30723 ( .A(nreg[209]), .B(n29484), .Z(n29487) );
  XNOR U30724 ( .A(n22095), .B(n29484), .Z(n29486) );
  XOR U30725 ( .A(n29488), .B(n29489), .Z(n22095) );
  XOR U30726 ( .A(n29490), .B(n29491), .Z(n29484) );
  AND U30727 ( .A(n29492), .B(n29493), .Z(n29491) );
  XOR U30728 ( .A(nreg[208]), .B(n29490), .Z(n29493) );
  XNOR U30729 ( .A(n22107), .B(n29490), .Z(n29492) );
  XOR U30730 ( .A(n29494), .B(n29495), .Z(n22107) );
  XOR U30731 ( .A(n29496), .B(n29497), .Z(n29490) );
  AND U30732 ( .A(n29498), .B(n29499), .Z(n29497) );
  XOR U30733 ( .A(nreg[207]), .B(n29496), .Z(n29499) );
  XNOR U30734 ( .A(n22119), .B(n29496), .Z(n29498) );
  XOR U30735 ( .A(n29500), .B(n29501), .Z(n22119) );
  XOR U30736 ( .A(n29502), .B(n29503), .Z(n29496) );
  AND U30737 ( .A(n29504), .B(n29505), .Z(n29503) );
  XOR U30738 ( .A(nreg[206]), .B(n29502), .Z(n29505) );
  XNOR U30739 ( .A(n22131), .B(n29502), .Z(n29504) );
  XOR U30740 ( .A(n29506), .B(n29507), .Z(n22131) );
  XOR U30741 ( .A(n29508), .B(n29509), .Z(n29502) );
  AND U30742 ( .A(n29510), .B(n29511), .Z(n29509) );
  XOR U30743 ( .A(nreg[205]), .B(n29508), .Z(n29511) );
  XNOR U30744 ( .A(n22143), .B(n29508), .Z(n29510) );
  XOR U30745 ( .A(n29512), .B(n29513), .Z(n22143) );
  XOR U30746 ( .A(n29514), .B(n29515), .Z(n29508) );
  AND U30747 ( .A(n29516), .B(n29517), .Z(n29515) );
  XOR U30748 ( .A(nreg[204]), .B(n29514), .Z(n29517) );
  XNOR U30749 ( .A(n22155), .B(n29514), .Z(n29516) );
  XOR U30750 ( .A(n29518), .B(n29519), .Z(n22155) );
  XOR U30751 ( .A(n29520), .B(n29521), .Z(n29514) );
  AND U30752 ( .A(n29522), .B(n29523), .Z(n29521) );
  XOR U30753 ( .A(nreg[203]), .B(n29520), .Z(n29523) );
  XNOR U30754 ( .A(n22167), .B(n29520), .Z(n29522) );
  XOR U30755 ( .A(n29524), .B(n29525), .Z(n22167) );
  XOR U30756 ( .A(n29526), .B(n29527), .Z(n29520) );
  AND U30757 ( .A(n29528), .B(n29529), .Z(n29527) );
  XOR U30758 ( .A(nreg[202]), .B(n29526), .Z(n29529) );
  XNOR U30759 ( .A(n22179), .B(n29526), .Z(n29528) );
  XOR U30760 ( .A(n29530), .B(n29531), .Z(n22179) );
  XOR U30761 ( .A(n29532), .B(n29533), .Z(n29526) );
  AND U30762 ( .A(n29534), .B(n29535), .Z(n29533) );
  XOR U30763 ( .A(nreg[201]), .B(n29532), .Z(n29535) );
  XNOR U30764 ( .A(n22191), .B(n29532), .Z(n29534) );
  XOR U30765 ( .A(n29536), .B(n29537), .Z(n22191) );
  XOR U30766 ( .A(n29538), .B(n29539), .Z(n29532) );
  AND U30767 ( .A(n29540), .B(n29541), .Z(n29539) );
  XOR U30768 ( .A(nreg[200]), .B(n29538), .Z(n29541) );
  XNOR U30769 ( .A(n22203), .B(n29538), .Z(n29540) );
  XOR U30770 ( .A(n29542), .B(n29543), .Z(n22203) );
  XOR U30771 ( .A(n29544), .B(n29545), .Z(n29538) );
  AND U30772 ( .A(n29546), .B(n29547), .Z(n29545) );
  XOR U30773 ( .A(nreg[199]), .B(n29544), .Z(n29547) );
  XNOR U30774 ( .A(n22215), .B(n29544), .Z(n29546) );
  XOR U30775 ( .A(n29548), .B(n29549), .Z(n22215) );
  XOR U30776 ( .A(n29550), .B(n29551), .Z(n29544) );
  AND U30777 ( .A(n29552), .B(n29553), .Z(n29551) );
  XOR U30778 ( .A(nreg[198]), .B(n29550), .Z(n29553) );
  XNOR U30779 ( .A(n22227), .B(n29550), .Z(n29552) );
  XOR U30780 ( .A(n29554), .B(n29555), .Z(n22227) );
  XOR U30781 ( .A(n29556), .B(n29557), .Z(n29550) );
  AND U30782 ( .A(n29558), .B(n29559), .Z(n29557) );
  XOR U30783 ( .A(nreg[197]), .B(n29556), .Z(n29559) );
  XNOR U30784 ( .A(n22239), .B(n29556), .Z(n29558) );
  XOR U30785 ( .A(n29560), .B(n29561), .Z(n22239) );
  XOR U30786 ( .A(n29562), .B(n29563), .Z(n29556) );
  AND U30787 ( .A(n29564), .B(n29565), .Z(n29563) );
  XOR U30788 ( .A(nreg[196]), .B(n29562), .Z(n29565) );
  XNOR U30789 ( .A(n22251), .B(n29562), .Z(n29564) );
  XOR U30790 ( .A(n29566), .B(n29567), .Z(n22251) );
  XOR U30791 ( .A(n29568), .B(n29569), .Z(n29562) );
  AND U30792 ( .A(n29570), .B(n29571), .Z(n29569) );
  XOR U30793 ( .A(nreg[195]), .B(n29568), .Z(n29571) );
  XNOR U30794 ( .A(n22263), .B(n29568), .Z(n29570) );
  XOR U30795 ( .A(n29572), .B(n29573), .Z(n22263) );
  XOR U30796 ( .A(n29574), .B(n29575), .Z(n29568) );
  AND U30797 ( .A(n29576), .B(n29577), .Z(n29575) );
  XOR U30798 ( .A(nreg[194]), .B(n29574), .Z(n29577) );
  XNOR U30799 ( .A(n22275), .B(n29574), .Z(n29576) );
  XOR U30800 ( .A(n29578), .B(n29579), .Z(n22275) );
  XOR U30801 ( .A(n29580), .B(n29581), .Z(n29574) );
  AND U30802 ( .A(n29582), .B(n29583), .Z(n29581) );
  XOR U30803 ( .A(nreg[193]), .B(n29580), .Z(n29583) );
  XNOR U30804 ( .A(n22287), .B(n29580), .Z(n29582) );
  XOR U30805 ( .A(n29584), .B(n29585), .Z(n22287) );
  XOR U30806 ( .A(n29586), .B(n29587), .Z(n29580) );
  AND U30807 ( .A(n29588), .B(n29589), .Z(n29587) );
  XOR U30808 ( .A(nreg[192]), .B(n29586), .Z(n29589) );
  XNOR U30809 ( .A(n22299), .B(n29586), .Z(n29588) );
  XOR U30810 ( .A(n29590), .B(n29591), .Z(n22299) );
  XOR U30811 ( .A(n29592), .B(n29593), .Z(n29586) );
  AND U30812 ( .A(n29594), .B(n29595), .Z(n29593) );
  XOR U30813 ( .A(nreg[191]), .B(n29592), .Z(n29595) );
  XNOR U30814 ( .A(n22311), .B(n29592), .Z(n29594) );
  XOR U30815 ( .A(n29596), .B(n29597), .Z(n22311) );
  XOR U30816 ( .A(n29598), .B(n29599), .Z(n29592) );
  AND U30817 ( .A(n29600), .B(n29601), .Z(n29599) );
  XOR U30818 ( .A(nreg[190]), .B(n29598), .Z(n29601) );
  XNOR U30819 ( .A(n22323), .B(n29598), .Z(n29600) );
  XOR U30820 ( .A(n29602), .B(n29603), .Z(n22323) );
  XOR U30821 ( .A(n29604), .B(n29605), .Z(n29598) );
  AND U30822 ( .A(n29606), .B(n29607), .Z(n29605) );
  XOR U30823 ( .A(nreg[189]), .B(n29604), .Z(n29607) );
  XNOR U30824 ( .A(n22335), .B(n29604), .Z(n29606) );
  XOR U30825 ( .A(n29608), .B(n29609), .Z(n22335) );
  XOR U30826 ( .A(n29610), .B(n29611), .Z(n29604) );
  AND U30827 ( .A(n29612), .B(n29613), .Z(n29611) );
  XOR U30828 ( .A(nreg[188]), .B(n29610), .Z(n29613) );
  XNOR U30829 ( .A(n22347), .B(n29610), .Z(n29612) );
  XOR U30830 ( .A(n29614), .B(n29615), .Z(n22347) );
  XOR U30831 ( .A(n29616), .B(n29617), .Z(n29610) );
  AND U30832 ( .A(n29618), .B(n29619), .Z(n29617) );
  XOR U30833 ( .A(nreg[187]), .B(n29616), .Z(n29619) );
  XNOR U30834 ( .A(n22359), .B(n29616), .Z(n29618) );
  XOR U30835 ( .A(n29620), .B(n29621), .Z(n22359) );
  XOR U30836 ( .A(n29622), .B(n29623), .Z(n29616) );
  AND U30837 ( .A(n29624), .B(n29625), .Z(n29623) );
  XOR U30838 ( .A(nreg[186]), .B(n29622), .Z(n29625) );
  XNOR U30839 ( .A(n22371), .B(n29622), .Z(n29624) );
  XOR U30840 ( .A(n29626), .B(n29627), .Z(n22371) );
  XOR U30841 ( .A(n29628), .B(n29629), .Z(n29622) );
  AND U30842 ( .A(n29630), .B(n29631), .Z(n29629) );
  XOR U30843 ( .A(nreg[185]), .B(n29628), .Z(n29631) );
  XNOR U30844 ( .A(n22383), .B(n29628), .Z(n29630) );
  XOR U30845 ( .A(n29632), .B(n29633), .Z(n22383) );
  XOR U30846 ( .A(n29634), .B(n29635), .Z(n29628) );
  AND U30847 ( .A(n29636), .B(n29637), .Z(n29635) );
  XOR U30848 ( .A(nreg[184]), .B(n29634), .Z(n29637) );
  XNOR U30849 ( .A(n22395), .B(n29634), .Z(n29636) );
  XOR U30850 ( .A(n29638), .B(n29639), .Z(n22395) );
  XOR U30851 ( .A(n29640), .B(n29641), .Z(n29634) );
  AND U30852 ( .A(n29642), .B(n29643), .Z(n29641) );
  XOR U30853 ( .A(nreg[183]), .B(n29640), .Z(n29643) );
  XNOR U30854 ( .A(n22407), .B(n29640), .Z(n29642) );
  XOR U30855 ( .A(n29644), .B(n29645), .Z(n22407) );
  XOR U30856 ( .A(n29646), .B(n29647), .Z(n29640) );
  AND U30857 ( .A(n29648), .B(n29649), .Z(n29647) );
  XOR U30858 ( .A(nreg[182]), .B(n29646), .Z(n29649) );
  XNOR U30859 ( .A(n22419), .B(n29646), .Z(n29648) );
  XOR U30860 ( .A(n29650), .B(n29651), .Z(n22419) );
  XOR U30861 ( .A(n29652), .B(n29653), .Z(n29646) );
  AND U30862 ( .A(n29654), .B(n29655), .Z(n29653) );
  XOR U30863 ( .A(nreg[181]), .B(n29652), .Z(n29655) );
  XNOR U30864 ( .A(n22431), .B(n29652), .Z(n29654) );
  XOR U30865 ( .A(n29656), .B(n29657), .Z(n22431) );
  XOR U30866 ( .A(n29658), .B(n29659), .Z(n29652) );
  AND U30867 ( .A(n29660), .B(n29661), .Z(n29659) );
  XOR U30868 ( .A(nreg[180]), .B(n29658), .Z(n29661) );
  XNOR U30869 ( .A(n22443), .B(n29658), .Z(n29660) );
  XOR U30870 ( .A(n29662), .B(n29663), .Z(n22443) );
  XOR U30871 ( .A(n29664), .B(n29665), .Z(n29658) );
  AND U30872 ( .A(n29666), .B(n29667), .Z(n29665) );
  XOR U30873 ( .A(nreg[179]), .B(n29664), .Z(n29667) );
  XNOR U30874 ( .A(n22455), .B(n29664), .Z(n29666) );
  XOR U30875 ( .A(n29668), .B(n29669), .Z(n22455) );
  XOR U30876 ( .A(n29670), .B(n29671), .Z(n29664) );
  AND U30877 ( .A(n29672), .B(n29673), .Z(n29671) );
  XOR U30878 ( .A(nreg[178]), .B(n29670), .Z(n29673) );
  XNOR U30879 ( .A(n22467), .B(n29670), .Z(n29672) );
  XOR U30880 ( .A(n29674), .B(n29675), .Z(n22467) );
  XOR U30881 ( .A(n29676), .B(n29677), .Z(n29670) );
  AND U30882 ( .A(n29678), .B(n29679), .Z(n29677) );
  XOR U30883 ( .A(nreg[177]), .B(n29676), .Z(n29679) );
  XNOR U30884 ( .A(n22479), .B(n29676), .Z(n29678) );
  XOR U30885 ( .A(n29680), .B(n29681), .Z(n22479) );
  XOR U30886 ( .A(n29682), .B(n29683), .Z(n29676) );
  AND U30887 ( .A(n29684), .B(n29685), .Z(n29683) );
  XOR U30888 ( .A(nreg[176]), .B(n29682), .Z(n29685) );
  XNOR U30889 ( .A(n22491), .B(n29682), .Z(n29684) );
  XOR U30890 ( .A(n29686), .B(n29687), .Z(n22491) );
  XOR U30891 ( .A(n29688), .B(n29689), .Z(n29682) );
  AND U30892 ( .A(n29690), .B(n29691), .Z(n29689) );
  XOR U30893 ( .A(nreg[175]), .B(n29688), .Z(n29691) );
  XNOR U30894 ( .A(n22503), .B(n29688), .Z(n29690) );
  XOR U30895 ( .A(n29692), .B(n29693), .Z(n22503) );
  XOR U30896 ( .A(n29694), .B(n29695), .Z(n29688) );
  AND U30897 ( .A(n29696), .B(n29697), .Z(n29695) );
  XOR U30898 ( .A(nreg[174]), .B(n29694), .Z(n29697) );
  XNOR U30899 ( .A(n22515), .B(n29694), .Z(n29696) );
  XOR U30900 ( .A(n29698), .B(n29699), .Z(n22515) );
  XOR U30901 ( .A(n29700), .B(n29701), .Z(n29694) );
  AND U30902 ( .A(n29702), .B(n29703), .Z(n29701) );
  XOR U30903 ( .A(nreg[173]), .B(n29700), .Z(n29703) );
  XNOR U30904 ( .A(n22527), .B(n29700), .Z(n29702) );
  XOR U30905 ( .A(n29704), .B(n29705), .Z(n22527) );
  XOR U30906 ( .A(n29706), .B(n29707), .Z(n29700) );
  AND U30907 ( .A(n29708), .B(n29709), .Z(n29707) );
  XOR U30908 ( .A(nreg[172]), .B(n29706), .Z(n29709) );
  XNOR U30909 ( .A(n22539), .B(n29706), .Z(n29708) );
  XOR U30910 ( .A(n29710), .B(n29711), .Z(n22539) );
  XOR U30911 ( .A(n29712), .B(n29713), .Z(n29706) );
  AND U30912 ( .A(n29714), .B(n29715), .Z(n29713) );
  XOR U30913 ( .A(nreg[171]), .B(n29712), .Z(n29715) );
  XNOR U30914 ( .A(n22551), .B(n29712), .Z(n29714) );
  XOR U30915 ( .A(n29716), .B(n29717), .Z(n22551) );
  XOR U30916 ( .A(n29718), .B(n29719), .Z(n29712) );
  AND U30917 ( .A(n29720), .B(n29721), .Z(n29719) );
  XOR U30918 ( .A(nreg[170]), .B(n29718), .Z(n29721) );
  XNOR U30919 ( .A(n22563), .B(n29718), .Z(n29720) );
  XOR U30920 ( .A(n29722), .B(n29723), .Z(n22563) );
  XOR U30921 ( .A(n29724), .B(n29725), .Z(n29718) );
  AND U30922 ( .A(n29726), .B(n29727), .Z(n29725) );
  XOR U30923 ( .A(nreg[169]), .B(n29724), .Z(n29727) );
  XNOR U30924 ( .A(n22575), .B(n29724), .Z(n29726) );
  XOR U30925 ( .A(n29728), .B(n29729), .Z(n22575) );
  XOR U30926 ( .A(n29730), .B(n29731), .Z(n29724) );
  AND U30927 ( .A(n29732), .B(n29733), .Z(n29731) );
  XOR U30928 ( .A(nreg[168]), .B(n29730), .Z(n29733) );
  XNOR U30929 ( .A(n22587), .B(n29730), .Z(n29732) );
  XOR U30930 ( .A(n29734), .B(n29735), .Z(n22587) );
  XOR U30931 ( .A(n29736), .B(n29737), .Z(n29730) );
  AND U30932 ( .A(n29738), .B(n29739), .Z(n29737) );
  XOR U30933 ( .A(nreg[167]), .B(n29736), .Z(n29739) );
  XNOR U30934 ( .A(n22599), .B(n29736), .Z(n29738) );
  XOR U30935 ( .A(n29740), .B(n29741), .Z(n22599) );
  XOR U30936 ( .A(n29742), .B(n29743), .Z(n29736) );
  AND U30937 ( .A(n29744), .B(n29745), .Z(n29743) );
  XOR U30938 ( .A(nreg[166]), .B(n29742), .Z(n29745) );
  XNOR U30939 ( .A(n22611), .B(n29742), .Z(n29744) );
  XOR U30940 ( .A(n29746), .B(n29747), .Z(n22611) );
  XOR U30941 ( .A(n29748), .B(n29749), .Z(n29742) );
  AND U30942 ( .A(n29750), .B(n29751), .Z(n29749) );
  XOR U30943 ( .A(nreg[165]), .B(n29748), .Z(n29751) );
  XNOR U30944 ( .A(n22623), .B(n29748), .Z(n29750) );
  XOR U30945 ( .A(n29752), .B(n29753), .Z(n22623) );
  XOR U30946 ( .A(n29754), .B(n29755), .Z(n29748) );
  AND U30947 ( .A(n29756), .B(n29757), .Z(n29755) );
  XOR U30948 ( .A(nreg[164]), .B(n29754), .Z(n29757) );
  XNOR U30949 ( .A(n22635), .B(n29754), .Z(n29756) );
  XOR U30950 ( .A(n29758), .B(n29759), .Z(n22635) );
  XOR U30951 ( .A(n29760), .B(n29761), .Z(n29754) );
  AND U30952 ( .A(n29762), .B(n29763), .Z(n29761) );
  XOR U30953 ( .A(nreg[163]), .B(n29760), .Z(n29763) );
  XNOR U30954 ( .A(n22647), .B(n29760), .Z(n29762) );
  XOR U30955 ( .A(n29764), .B(n29765), .Z(n22647) );
  XOR U30956 ( .A(n29766), .B(n29767), .Z(n29760) );
  AND U30957 ( .A(n29768), .B(n29769), .Z(n29767) );
  XOR U30958 ( .A(nreg[162]), .B(n29766), .Z(n29769) );
  XNOR U30959 ( .A(n22659), .B(n29766), .Z(n29768) );
  XOR U30960 ( .A(n29770), .B(n29771), .Z(n22659) );
  XOR U30961 ( .A(n29772), .B(n29773), .Z(n29766) );
  AND U30962 ( .A(n29774), .B(n29775), .Z(n29773) );
  XOR U30963 ( .A(nreg[161]), .B(n29772), .Z(n29775) );
  XNOR U30964 ( .A(n22671), .B(n29772), .Z(n29774) );
  XOR U30965 ( .A(n29776), .B(n29777), .Z(n22671) );
  XOR U30966 ( .A(n29778), .B(n29779), .Z(n29772) );
  AND U30967 ( .A(n29780), .B(n29781), .Z(n29779) );
  XOR U30968 ( .A(nreg[160]), .B(n29778), .Z(n29781) );
  XNOR U30969 ( .A(n22683), .B(n29778), .Z(n29780) );
  XOR U30970 ( .A(n29782), .B(n29783), .Z(n22683) );
  XOR U30971 ( .A(n29784), .B(n29785), .Z(n29778) );
  AND U30972 ( .A(n29786), .B(n29787), .Z(n29785) );
  XOR U30973 ( .A(nreg[159]), .B(n29784), .Z(n29787) );
  XNOR U30974 ( .A(n22695), .B(n29784), .Z(n29786) );
  XOR U30975 ( .A(n29788), .B(n29789), .Z(n22695) );
  XOR U30976 ( .A(n29790), .B(n29791), .Z(n29784) );
  AND U30977 ( .A(n29792), .B(n29793), .Z(n29791) );
  XOR U30978 ( .A(nreg[158]), .B(n29790), .Z(n29793) );
  XNOR U30979 ( .A(n22707), .B(n29790), .Z(n29792) );
  XOR U30980 ( .A(n29794), .B(n29795), .Z(n22707) );
  XOR U30981 ( .A(n29796), .B(n29797), .Z(n29790) );
  AND U30982 ( .A(n29798), .B(n29799), .Z(n29797) );
  XOR U30983 ( .A(nreg[157]), .B(n29796), .Z(n29799) );
  XNOR U30984 ( .A(n22719), .B(n29796), .Z(n29798) );
  XOR U30985 ( .A(n29800), .B(n29801), .Z(n22719) );
  XOR U30986 ( .A(n29802), .B(n29803), .Z(n29796) );
  AND U30987 ( .A(n29804), .B(n29805), .Z(n29803) );
  XOR U30988 ( .A(nreg[156]), .B(n29802), .Z(n29805) );
  XNOR U30989 ( .A(n22731), .B(n29802), .Z(n29804) );
  XOR U30990 ( .A(n29806), .B(n29807), .Z(n22731) );
  XOR U30991 ( .A(n29808), .B(n29809), .Z(n29802) );
  AND U30992 ( .A(n29810), .B(n29811), .Z(n29809) );
  XOR U30993 ( .A(nreg[155]), .B(n29808), .Z(n29811) );
  XNOR U30994 ( .A(n22743), .B(n29808), .Z(n29810) );
  XOR U30995 ( .A(n29812), .B(n29813), .Z(n22743) );
  XOR U30996 ( .A(n29814), .B(n29815), .Z(n29808) );
  AND U30997 ( .A(n29816), .B(n29817), .Z(n29815) );
  XOR U30998 ( .A(nreg[154]), .B(n29814), .Z(n29817) );
  XNOR U30999 ( .A(n22755), .B(n29814), .Z(n29816) );
  XOR U31000 ( .A(n29818), .B(n29819), .Z(n22755) );
  XOR U31001 ( .A(n29820), .B(n29821), .Z(n29814) );
  AND U31002 ( .A(n29822), .B(n29823), .Z(n29821) );
  XOR U31003 ( .A(nreg[153]), .B(n29820), .Z(n29823) );
  XNOR U31004 ( .A(n22767), .B(n29820), .Z(n29822) );
  XOR U31005 ( .A(n29824), .B(n29825), .Z(n22767) );
  XOR U31006 ( .A(n29826), .B(n29827), .Z(n29820) );
  AND U31007 ( .A(n29828), .B(n29829), .Z(n29827) );
  XOR U31008 ( .A(nreg[152]), .B(n29826), .Z(n29829) );
  XNOR U31009 ( .A(n22779), .B(n29826), .Z(n29828) );
  XOR U31010 ( .A(n29830), .B(n29831), .Z(n22779) );
  XOR U31011 ( .A(n29832), .B(n29833), .Z(n29826) );
  AND U31012 ( .A(n29834), .B(n29835), .Z(n29833) );
  XOR U31013 ( .A(nreg[151]), .B(n29832), .Z(n29835) );
  XNOR U31014 ( .A(n22791), .B(n29832), .Z(n29834) );
  XOR U31015 ( .A(n29836), .B(n29837), .Z(n22791) );
  XOR U31016 ( .A(n29838), .B(n29839), .Z(n29832) );
  AND U31017 ( .A(n29840), .B(n29841), .Z(n29839) );
  XOR U31018 ( .A(nreg[150]), .B(n29838), .Z(n29841) );
  XNOR U31019 ( .A(n22803), .B(n29838), .Z(n29840) );
  XOR U31020 ( .A(n29842), .B(n29843), .Z(n22803) );
  XOR U31021 ( .A(n29844), .B(n29845), .Z(n29838) );
  AND U31022 ( .A(n29846), .B(n29847), .Z(n29845) );
  XOR U31023 ( .A(nreg[149]), .B(n29844), .Z(n29847) );
  XNOR U31024 ( .A(n22815), .B(n29844), .Z(n29846) );
  XOR U31025 ( .A(n29848), .B(n29849), .Z(n22815) );
  XOR U31026 ( .A(n29850), .B(n29851), .Z(n29844) );
  AND U31027 ( .A(n29852), .B(n29853), .Z(n29851) );
  XOR U31028 ( .A(nreg[148]), .B(n29850), .Z(n29853) );
  XNOR U31029 ( .A(n22827), .B(n29850), .Z(n29852) );
  XOR U31030 ( .A(n29854), .B(n29855), .Z(n22827) );
  XOR U31031 ( .A(n29856), .B(n29857), .Z(n29850) );
  AND U31032 ( .A(n29858), .B(n29859), .Z(n29857) );
  XOR U31033 ( .A(nreg[147]), .B(n29856), .Z(n29859) );
  XNOR U31034 ( .A(n22839), .B(n29856), .Z(n29858) );
  XOR U31035 ( .A(n29860), .B(n29861), .Z(n22839) );
  XOR U31036 ( .A(n29862), .B(n29863), .Z(n29856) );
  AND U31037 ( .A(n29864), .B(n29865), .Z(n29863) );
  XOR U31038 ( .A(nreg[146]), .B(n29862), .Z(n29865) );
  XNOR U31039 ( .A(n22851), .B(n29862), .Z(n29864) );
  XOR U31040 ( .A(n29866), .B(n29867), .Z(n22851) );
  XOR U31041 ( .A(n29868), .B(n29869), .Z(n29862) );
  AND U31042 ( .A(n29870), .B(n29871), .Z(n29869) );
  XOR U31043 ( .A(nreg[145]), .B(n29868), .Z(n29871) );
  XNOR U31044 ( .A(n22863), .B(n29868), .Z(n29870) );
  XOR U31045 ( .A(n29872), .B(n29873), .Z(n22863) );
  XOR U31046 ( .A(n29874), .B(n29875), .Z(n29868) );
  AND U31047 ( .A(n29876), .B(n29877), .Z(n29875) );
  XOR U31048 ( .A(nreg[144]), .B(n29874), .Z(n29877) );
  XNOR U31049 ( .A(n22875), .B(n29874), .Z(n29876) );
  XOR U31050 ( .A(n29878), .B(n29879), .Z(n22875) );
  XOR U31051 ( .A(n29880), .B(n29881), .Z(n29874) );
  AND U31052 ( .A(n29882), .B(n29883), .Z(n29881) );
  XOR U31053 ( .A(nreg[143]), .B(n29880), .Z(n29883) );
  XNOR U31054 ( .A(n22887), .B(n29880), .Z(n29882) );
  XOR U31055 ( .A(n29884), .B(n29885), .Z(n22887) );
  XOR U31056 ( .A(n29886), .B(n29887), .Z(n29880) );
  AND U31057 ( .A(n29888), .B(n29889), .Z(n29887) );
  XOR U31058 ( .A(nreg[142]), .B(n29886), .Z(n29889) );
  XNOR U31059 ( .A(n22899), .B(n29886), .Z(n29888) );
  XOR U31060 ( .A(n29890), .B(n29891), .Z(n22899) );
  XOR U31061 ( .A(n29892), .B(n29893), .Z(n29886) );
  AND U31062 ( .A(n29894), .B(n29895), .Z(n29893) );
  XOR U31063 ( .A(nreg[141]), .B(n29892), .Z(n29895) );
  XNOR U31064 ( .A(n22911), .B(n29892), .Z(n29894) );
  XOR U31065 ( .A(n29896), .B(n29897), .Z(n22911) );
  XOR U31066 ( .A(n29898), .B(n29899), .Z(n29892) );
  AND U31067 ( .A(n29900), .B(n29901), .Z(n29899) );
  XOR U31068 ( .A(nreg[140]), .B(n29898), .Z(n29901) );
  XNOR U31069 ( .A(n22923), .B(n29898), .Z(n29900) );
  XOR U31070 ( .A(n29902), .B(n29903), .Z(n22923) );
  XOR U31071 ( .A(n29904), .B(n29905), .Z(n29898) );
  AND U31072 ( .A(n29906), .B(n29907), .Z(n29905) );
  XOR U31073 ( .A(nreg[139]), .B(n29904), .Z(n29907) );
  XNOR U31074 ( .A(n22935), .B(n29904), .Z(n29906) );
  XOR U31075 ( .A(n29908), .B(n29909), .Z(n22935) );
  XOR U31076 ( .A(n29910), .B(n29911), .Z(n29904) );
  AND U31077 ( .A(n29912), .B(n29913), .Z(n29911) );
  XOR U31078 ( .A(nreg[138]), .B(n29910), .Z(n29913) );
  XNOR U31079 ( .A(n22947), .B(n29910), .Z(n29912) );
  XOR U31080 ( .A(n29914), .B(n29915), .Z(n22947) );
  XOR U31081 ( .A(n29916), .B(n29917), .Z(n29910) );
  AND U31082 ( .A(n29918), .B(n29919), .Z(n29917) );
  XOR U31083 ( .A(nreg[137]), .B(n29916), .Z(n29919) );
  XNOR U31084 ( .A(n22959), .B(n29916), .Z(n29918) );
  XOR U31085 ( .A(n29920), .B(n29921), .Z(n22959) );
  XOR U31086 ( .A(n29922), .B(n29923), .Z(n29916) );
  AND U31087 ( .A(n29924), .B(n29925), .Z(n29923) );
  XOR U31088 ( .A(nreg[136]), .B(n29922), .Z(n29925) );
  XNOR U31089 ( .A(n22971), .B(n29922), .Z(n29924) );
  XOR U31090 ( .A(n29926), .B(n29927), .Z(n22971) );
  XOR U31091 ( .A(n29928), .B(n29929), .Z(n29922) );
  AND U31092 ( .A(n29930), .B(n29931), .Z(n29929) );
  XOR U31093 ( .A(nreg[135]), .B(n29928), .Z(n29931) );
  XNOR U31094 ( .A(n22983), .B(n29928), .Z(n29930) );
  XOR U31095 ( .A(n29932), .B(n29933), .Z(n22983) );
  XOR U31096 ( .A(n29934), .B(n29935), .Z(n29928) );
  AND U31097 ( .A(n29936), .B(n29937), .Z(n29935) );
  XOR U31098 ( .A(nreg[134]), .B(n29934), .Z(n29937) );
  XNOR U31099 ( .A(n22995), .B(n29934), .Z(n29936) );
  XOR U31100 ( .A(n29938), .B(n29939), .Z(n22995) );
  XOR U31101 ( .A(n29940), .B(n29941), .Z(n29934) );
  AND U31102 ( .A(n29942), .B(n29943), .Z(n29941) );
  XOR U31103 ( .A(nreg[133]), .B(n29940), .Z(n29943) );
  XNOR U31104 ( .A(n23007), .B(n29940), .Z(n29942) );
  XOR U31105 ( .A(n29944), .B(n29945), .Z(n23007) );
  XOR U31106 ( .A(n29946), .B(n29947), .Z(n29940) );
  AND U31107 ( .A(n29948), .B(n29949), .Z(n29947) );
  XOR U31108 ( .A(nreg[132]), .B(n29946), .Z(n29949) );
  XNOR U31109 ( .A(n23019), .B(n29946), .Z(n29948) );
  XOR U31110 ( .A(n29950), .B(n29951), .Z(n23019) );
  XOR U31111 ( .A(n29952), .B(n29953), .Z(n29946) );
  AND U31112 ( .A(n29954), .B(n29955), .Z(n29953) );
  XOR U31113 ( .A(nreg[131]), .B(n29952), .Z(n29955) );
  XNOR U31114 ( .A(n23031), .B(n29952), .Z(n29954) );
  XOR U31115 ( .A(n29956), .B(n29957), .Z(n23031) );
  XOR U31116 ( .A(n29958), .B(n29959), .Z(n29952) );
  AND U31117 ( .A(n29960), .B(n29961), .Z(n29959) );
  XOR U31118 ( .A(nreg[130]), .B(n29958), .Z(n29961) );
  XNOR U31119 ( .A(n23043), .B(n29958), .Z(n29960) );
  XOR U31120 ( .A(n29962), .B(n29963), .Z(n23043) );
  XOR U31121 ( .A(n29964), .B(n29965), .Z(n29958) );
  AND U31122 ( .A(n29966), .B(n29967), .Z(n29965) );
  XOR U31123 ( .A(nreg[129]), .B(n29964), .Z(n29967) );
  XNOR U31124 ( .A(n23055), .B(n29964), .Z(n29966) );
  XOR U31125 ( .A(n29968), .B(n29969), .Z(n23055) );
  XOR U31126 ( .A(n29970), .B(n29971), .Z(n29964) );
  AND U31127 ( .A(n29972), .B(n29973), .Z(n29971) );
  XOR U31128 ( .A(nreg[128]), .B(n29970), .Z(n29973) );
  XNOR U31129 ( .A(n23067), .B(n29970), .Z(n29972) );
  XOR U31130 ( .A(n29974), .B(n29975), .Z(n23067) );
  XOR U31131 ( .A(n29976), .B(n29977), .Z(n29970) );
  AND U31132 ( .A(n29978), .B(n29979), .Z(n29977) );
  XOR U31133 ( .A(nreg[127]), .B(n29976), .Z(n29979) );
  XNOR U31134 ( .A(n23079), .B(n29976), .Z(n29978) );
  XOR U31135 ( .A(n29980), .B(n29981), .Z(n23079) );
  XOR U31136 ( .A(n29982), .B(n29983), .Z(n29976) );
  AND U31137 ( .A(n29984), .B(n29985), .Z(n29983) );
  XOR U31138 ( .A(nreg[126]), .B(n29982), .Z(n29985) );
  XNOR U31139 ( .A(n23091), .B(n29982), .Z(n29984) );
  XOR U31140 ( .A(n29986), .B(n29987), .Z(n23091) );
  XOR U31141 ( .A(n29988), .B(n29989), .Z(n29982) );
  AND U31142 ( .A(n29990), .B(n29991), .Z(n29989) );
  XOR U31143 ( .A(nreg[125]), .B(n29988), .Z(n29991) );
  XNOR U31144 ( .A(n23103), .B(n29988), .Z(n29990) );
  XOR U31145 ( .A(n29992), .B(n29993), .Z(n23103) );
  XOR U31146 ( .A(n29994), .B(n29995), .Z(n29988) );
  AND U31147 ( .A(n29996), .B(n29997), .Z(n29995) );
  XOR U31148 ( .A(nreg[124]), .B(n29994), .Z(n29997) );
  XNOR U31149 ( .A(n23115), .B(n29994), .Z(n29996) );
  XOR U31150 ( .A(n29998), .B(n29999), .Z(n23115) );
  XOR U31151 ( .A(n30000), .B(n30001), .Z(n29994) );
  AND U31152 ( .A(n30002), .B(n30003), .Z(n30001) );
  XOR U31153 ( .A(nreg[123]), .B(n30000), .Z(n30003) );
  XNOR U31154 ( .A(n23127), .B(n30000), .Z(n30002) );
  XOR U31155 ( .A(n30004), .B(n30005), .Z(n23127) );
  XOR U31156 ( .A(n30006), .B(n30007), .Z(n30000) );
  AND U31157 ( .A(n30008), .B(n30009), .Z(n30007) );
  XOR U31158 ( .A(nreg[122]), .B(n30006), .Z(n30009) );
  XNOR U31159 ( .A(n23139), .B(n30006), .Z(n30008) );
  XOR U31160 ( .A(n30010), .B(n30011), .Z(n23139) );
  XOR U31161 ( .A(n30012), .B(n30013), .Z(n30006) );
  AND U31162 ( .A(n30014), .B(n30015), .Z(n30013) );
  XOR U31163 ( .A(nreg[121]), .B(n30012), .Z(n30015) );
  XNOR U31164 ( .A(n23151), .B(n30012), .Z(n30014) );
  XOR U31165 ( .A(n30016), .B(n30017), .Z(n23151) );
  XOR U31166 ( .A(n30018), .B(n30019), .Z(n30012) );
  AND U31167 ( .A(n30020), .B(n30021), .Z(n30019) );
  XOR U31168 ( .A(nreg[120]), .B(n30018), .Z(n30021) );
  XNOR U31169 ( .A(n23163), .B(n30018), .Z(n30020) );
  XOR U31170 ( .A(n30022), .B(n30023), .Z(n23163) );
  XOR U31171 ( .A(n30024), .B(n30025), .Z(n30018) );
  AND U31172 ( .A(n30026), .B(n30027), .Z(n30025) );
  XOR U31173 ( .A(nreg[119]), .B(n30024), .Z(n30027) );
  XNOR U31174 ( .A(n23175), .B(n30024), .Z(n30026) );
  XOR U31175 ( .A(n30028), .B(n30029), .Z(n23175) );
  XOR U31176 ( .A(n30030), .B(n30031), .Z(n30024) );
  AND U31177 ( .A(n30032), .B(n30033), .Z(n30031) );
  XOR U31178 ( .A(nreg[118]), .B(n30030), .Z(n30033) );
  XNOR U31179 ( .A(n23187), .B(n30030), .Z(n30032) );
  XOR U31180 ( .A(n30034), .B(n30035), .Z(n23187) );
  XOR U31181 ( .A(n30036), .B(n30037), .Z(n30030) );
  AND U31182 ( .A(n30038), .B(n30039), .Z(n30037) );
  XOR U31183 ( .A(nreg[117]), .B(n30036), .Z(n30039) );
  XNOR U31184 ( .A(n23199), .B(n30036), .Z(n30038) );
  XOR U31185 ( .A(n30040), .B(n30041), .Z(n23199) );
  XOR U31186 ( .A(n30042), .B(n30043), .Z(n30036) );
  AND U31187 ( .A(n30044), .B(n30045), .Z(n30043) );
  XOR U31188 ( .A(nreg[116]), .B(n30042), .Z(n30045) );
  XNOR U31189 ( .A(n23211), .B(n30042), .Z(n30044) );
  XOR U31190 ( .A(n30046), .B(n30047), .Z(n23211) );
  XOR U31191 ( .A(n30048), .B(n30049), .Z(n30042) );
  AND U31192 ( .A(n30050), .B(n30051), .Z(n30049) );
  XOR U31193 ( .A(nreg[115]), .B(n30048), .Z(n30051) );
  XNOR U31194 ( .A(n23223), .B(n30048), .Z(n30050) );
  XOR U31195 ( .A(n30052), .B(n30053), .Z(n23223) );
  XOR U31196 ( .A(n30054), .B(n30055), .Z(n30048) );
  AND U31197 ( .A(n30056), .B(n30057), .Z(n30055) );
  XOR U31198 ( .A(nreg[114]), .B(n30054), .Z(n30057) );
  XNOR U31199 ( .A(n23235), .B(n30054), .Z(n30056) );
  XOR U31200 ( .A(n30058), .B(n30059), .Z(n23235) );
  XOR U31201 ( .A(n30060), .B(n30061), .Z(n30054) );
  AND U31202 ( .A(n30062), .B(n30063), .Z(n30061) );
  XOR U31203 ( .A(nreg[113]), .B(n30060), .Z(n30063) );
  XNOR U31204 ( .A(n23247), .B(n30060), .Z(n30062) );
  XOR U31205 ( .A(n30064), .B(n30065), .Z(n23247) );
  XOR U31206 ( .A(n30066), .B(n30067), .Z(n30060) );
  AND U31207 ( .A(n30068), .B(n30069), .Z(n30067) );
  XOR U31208 ( .A(nreg[112]), .B(n30066), .Z(n30069) );
  XNOR U31209 ( .A(n23259), .B(n30066), .Z(n30068) );
  XOR U31210 ( .A(n30070), .B(n30071), .Z(n23259) );
  XOR U31211 ( .A(n30072), .B(n30073), .Z(n30066) );
  AND U31212 ( .A(n30074), .B(n30075), .Z(n30073) );
  XOR U31213 ( .A(nreg[111]), .B(n30072), .Z(n30075) );
  XNOR U31214 ( .A(n23271), .B(n30072), .Z(n30074) );
  XOR U31215 ( .A(n30076), .B(n30077), .Z(n23271) );
  XOR U31216 ( .A(n30078), .B(n30079), .Z(n30072) );
  AND U31217 ( .A(n30080), .B(n30081), .Z(n30079) );
  XOR U31218 ( .A(nreg[110]), .B(n30078), .Z(n30081) );
  XNOR U31219 ( .A(n23283), .B(n30078), .Z(n30080) );
  XOR U31220 ( .A(n30082), .B(n30083), .Z(n23283) );
  XOR U31221 ( .A(n30084), .B(n30085), .Z(n30078) );
  AND U31222 ( .A(n30086), .B(n30087), .Z(n30085) );
  XOR U31223 ( .A(nreg[109]), .B(n30084), .Z(n30087) );
  XNOR U31224 ( .A(n23295), .B(n30084), .Z(n30086) );
  XOR U31225 ( .A(n30088), .B(n30089), .Z(n23295) );
  XOR U31226 ( .A(n30090), .B(n30091), .Z(n30084) );
  AND U31227 ( .A(n30092), .B(n30093), .Z(n30091) );
  XOR U31228 ( .A(nreg[108]), .B(n30090), .Z(n30093) );
  XNOR U31229 ( .A(n23307), .B(n30090), .Z(n30092) );
  XOR U31230 ( .A(n30094), .B(n30095), .Z(n23307) );
  XOR U31231 ( .A(n30096), .B(n30097), .Z(n30090) );
  AND U31232 ( .A(n30098), .B(n30099), .Z(n30097) );
  XOR U31233 ( .A(nreg[107]), .B(n30096), .Z(n30099) );
  XNOR U31234 ( .A(n23319), .B(n30096), .Z(n30098) );
  XOR U31235 ( .A(n30100), .B(n30101), .Z(n23319) );
  XOR U31236 ( .A(n30102), .B(n30103), .Z(n30096) );
  AND U31237 ( .A(n30104), .B(n30105), .Z(n30103) );
  XOR U31238 ( .A(nreg[106]), .B(n30102), .Z(n30105) );
  XNOR U31239 ( .A(n23331), .B(n30102), .Z(n30104) );
  XOR U31240 ( .A(n30106), .B(n30107), .Z(n23331) );
  XOR U31241 ( .A(n30108), .B(n30109), .Z(n30102) );
  AND U31242 ( .A(n30110), .B(n30111), .Z(n30109) );
  XOR U31243 ( .A(nreg[105]), .B(n30108), .Z(n30111) );
  XNOR U31244 ( .A(n23343), .B(n30108), .Z(n30110) );
  XOR U31245 ( .A(n30112), .B(n30113), .Z(n23343) );
  XOR U31246 ( .A(n30114), .B(n30115), .Z(n30108) );
  AND U31247 ( .A(n30116), .B(n30117), .Z(n30115) );
  XOR U31248 ( .A(nreg[104]), .B(n30114), .Z(n30117) );
  XNOR U31249 ( .A(n23355), .B(n30114), .Z(n30116) );
  XOR U31250 ( .A(n30118), .B(n30119), .Z(n23355) );
  XOR U31251 ( .A(n30120), .B(n30121), .Z(n30114) );
  AND U31252 ( .A(n30122), .B(n30123), .Z(n30121) );
  XOR U31253 ( .A(nreg[103]), .B(n30120), .Z(n30123) );
  XNOR U31254 ( .A(n23367), .B(n30120), .Z(n30122) );
  XOR U31255 ( .A(n30124), .B(n30125), .Z(n23367) );
  XOR U31256 ( .A(n30126), .B(n30127), .Z(n30120) );
  AND U31257 ( .A(n30128), .B(n30129), .Z(n30127) );
  XOR U31258 ( .A(nreg[102]), .B(n30126), .Z(n30129) );
  XNOR U31259 ( .A(n23379), .B(n30126), .Z(n30128) );
  XOR U31260 ( .A(n30130), .B(n30131), .Z(n23379) );
  XOR U31261 ( .A(n30132), .B(n30133), .Z(n30126) );
  AND U31262 ( .A(n30134), .B(n30135), .Z(n30133) );
  XOR U31263 ( .A(nreg[101]), .B(n30132), .Z(n30135) );
  XNOR U31264 ( .A(n23391), .B(n30132), .Z(n30134) );
  XOR U31265 ( .A(n30136), .B(n30137), .Z(n23391) );
  XOR U31266 ( .A(n30138), .B(n30139), .Z(n30132) );
  AND U31267 ( .A(n30140), .B(n30141), .Z(n30139) );
  XOR U31268 ( .A(nreg[100]), .B(n30138), .Z(n30141) );
  XNOR U31269 ( .A(n23403), .B(n30138), .Z(n30140) );
  XOR U31270 ( .A(n30142), .B(n30143), .Z(n23403) );
  XOR U31271 ( .A(n30144), .B(n30145), .Z(n30138) );
  AND U31272 ( .A(n30146), .B(n30147), .Z(n30145) );
  XOR U31273 ( .A(nreg[99]), .B(n30144), .Z(n30147) );
  XNOR U31274 ( .A(n23415), .B(n30144), .Z(n30146) );
  XOR U31275 ( .A(n30148), .B(n30149), .Z(n23415) );
  XOR U31276 ( .A(n30150), .B(n30151), .Z(n30144) );
  AND U31277 ( .A(n30152), .B(n30153), .Z(n30151) );
  XOR U31278 ( .A(nreg[98]), .B(n30150), .Z(n30153) );
  XNOR U31279 ( .A(n23427), .B(n30150), .Z(n30152) );
  XOR U31280 ( .A(n30154), .B(n30155), .Z(n23427) );
  XOR U31281 ( .A(n30156), .B(n30157), .Z(n30150) );
  AND U31282 ( .A(n30158), .B(n30159), .Z(n30157) );
  XOR U31283 ( .A(nreg[97]), .B(n30156), .Z(n30159) );
  XNOR U31284 ( .A(n23439), .B(n30156), .Z(n30158) );
  XOR U31285 ( .A(n30160), .B(n30161), .Z(n23439) );
  XOR U31286 ( .A(n30162), .B(n30163), .Z(n30156) );
  AND U31287 ( .A(n30164), .B(n30165), .Z(n30163) );
  XOR U31288 ( .A(nreg[96]), .B(n30162), .Z(n30165) );
  XNOR U31289 ( .A(n23451), .B(n30162), .Z(n30164) );
  XOR U31290 ( .A(n30166), .B(n30167), .Z(n23451) );
  XOR U31291 ( .A(n30168), .B(n30169), .Z(n30162) );
  AND U31292 ( .A(n30170), .B(n30171), .Z(n30169) );
  XOR U31293 ( .A(nreg[95]), .B(n30168), .Z(n30171) );
  XNOR U31294 ( .A(n23463), .B(n30168), .Z(n30170) );
  XOR U31295 ( .A(n30172), .B(n30173), .Z(n23463) );
  XOR U31296 ( .A(n30174), .B(n30175), .Z(n30168) );
  AND U31297 ( .A(n30176), .B(n30177), .Z(n30175) );
  XOR U31298 ( .A(nreg[94]), .B(n30174), .Z(n30177) );
  XNOR U31299 ( .A(n23475), .B(n30174), .Z(n30176) );
  XOR U31300 ( .A(n30178), .B(n30179), .Z(n23475) );
  XOR U31301 ( .A(n30180), .B(n30181), .Z(n30174) );
  AND U31302 ( .A(n30182), .B(n30183), .Z(n30181) );
  XOR U31303 ( .A(nreg[93]), .B(n30180), .Z(n30183) );
  XNOR U31304 ( .A(n23487), .B(n30180), .Z(n30182) );
  XOR U31305 ( .A(n30184), .B(n30185), .Z(n23487) );
  XOR U31306 ( .A(n30186), .B(n30187), .Z(n30180) );
  AND U31307 ( .A(n30188), .B(n30189), .Z(n30187) );
  XOR U31308 ( .A(nreg[92]), .B(n30186), .Z(n30189) );
  XNOR U31309 ( .A(n23499), .B(n30186), .Z(n30188) );
  XOR U31310 ( .A(n30190), .B(n30191), .Z(n23499) );
  XOR U31311 ( .A(n30192), .B(n30193), .Z(n30186) );
  AND U31312 ( .A(n30194), .B(n30195), .Z(n30193) );
  XOR U31313 ( .A(nreg[91]), .B(n30192), .Z(n30195) );
  XNOR U31314 ( .A(n23511), .B(n30192), .Z(n30194) );
  XOR U31315 ( .A(n30196), .B(n30197), .Z(n23511) );
  XOR U31316 ( .A(n30198), .B(n30199), .Z(n30192) );
  AND U31317 ( .A(n30200), .B(n30201), .Z(n30199) );
  XOR U31318 ( .A(nreg[90]), .B(n30198), .Z(n30201) );
  XNOR U31319 ( .A(n23523), .B(n30198), .Z(n30200) );
  XOR U31320 ( .A(n30202), .B(n30203), .Z(n23523) );
  XOR U31321 ( .A(n30204), .B(n30205), .Z(n30198) );
  AND U31322 ( .A(n30206), .B(n30207), .Z(n30205) );
  XOR U31323 ( .A(nreg[89]), .B(n30204), .Z(n30207) );
  XNOR U31324 ( .A(n23535), .B(n30204), .Z(n30206) );
  XOR U31325 ( .A(n30208), .B(n30209), .Z(n23535) );
  XOR U31326 ( .A(n30210), .B(n30211), .Z(n30204) );
  AND U31327 ( .A(n30212), .B(n30213), .Z(n30211) );
  XOR U31328 ( .A(nreg[88]), .B(n30210), .Z(n30213) );
  XNOR U31329 ( .A(n23547), .B(n30210), .Z(n30212) );
  XOR U31330 ( .A(n30214), .B(n30215), .Z(n23547) );
  XOR U31331 ( .A(n30216), .B(n30217), .Z(n30210) );
  AND U31332 ( .A(n30218), .B(n30219), .Z(n30217) );
  XOR U31333 ( .A(nreg[87]), .B(n30216), .Z(n30219) );
  XNOR U31334 ( .A(n23559), .B(n30216), .Z(n30218) );
  XOR U31335 ( .A(n30220), .B(n30221), .Z(n23559) );
  XOR U31336 ( .A(n30222), .B(n30223), .Z(n30216) );
  AND U31337 ( .A(n30224), .B(n30225), .Z(n30223) );
  XOR U31338 ( .A(nreg[86]), .B(n30222), .Z(n30225) );
  XNOR U31339 ( .A(n23571), .B(n30222), .Z(n30224) );
  XOR U31340 ( .A(n30226), .B(n30227), .Z(n23571) );
  XOR U31341 ( .A(n30228), .B(n30229), .Z(n30222) );
  AND U31342 ( .A(n30230), .B(n30231), .Z(n30229) );
  XOR U31343 ( .A(nreg[85]), .B(n30228), .Z(n30231) );
  XNOR U31344 ( .A(n23583), .B(n30228), .Z(n30230) );
  XOR U31345 ( .A(n30232), .B(n30233), .Z(n23583) );
  XOR U31346 ( .A(n30234), .B(n30235), .Z(n30228) );
  AND U31347 ( .A(n30236), .B(n30237), .Z(n30235) );
  XOR U31348 ( .A(nreg[84]), .B(n30234), .Z(n30237) );
  XNOR U31349 ( .A(n23595), .B(n30234), .Z(n30236) );
  XOR U31350 ( .A(n30238), .B(n30239), .Z(n23595) );
  XOR U31351 ( .A(n30240), .B(n30241), .Z(n30234) );
  AND U31352 ( .A(n30242), .B(n30243), .Z(n30241) );
  XOR U31353 ( .A(nreg[83]), .B(n30240), .Z(n30243) );
  XNOR U31354 ( .A(n23607), .B(n30240), .Z(n30242) );
  XOR U31355 ( .A(n30244), .B(n30245), .Z(n23607) );
  XOR U31356 ( .A(n30246), .B(n30247), .Z(n30240) );
  AND U31357 ( .A(n30248), .B(n30249), .Z(n30247) );
  XOR U31358 ( .A(nreg[82]), .B(n30246), .Z(n30249) );
  XNOR U31359 ( .A(n23619), .B(n30246), .Z(n30248) );
  XOR U31360 ( .A(n30250), .B(n30251), .Z(n23619) );
  XOR U31361 ( .A(n30252), .B(n30253), .Z(n30246) );
  AND U31362 ( .A(n30254), .B(n30255), .Z(n30253) );
  XOR U31363 ( .A(nreg[81]), .B(n30252), .Z(n30255) );
  XNOR U31364 ( .A(n23631), .B(n30252), .Z(n30254) );
  XOR U31365 ( .A(n30256), .B(n30257), .Z(n23631) );
  XOR U31366 ( .A(n30258), .B(n30259), .Z(n30252) );
  AND U31367 ( .A(n30260), .B(n30261), .Z(n30259) );
  XOR U31368 ( .A(nreg[80]), .B(n30258), .Z(n30261) );
  XNOR U31369 ( .A(n23643), .B(n30258), .Z(n30260) );
  XOR U31370 ( .A(n30262), .B(n30263), .Z(n23643) );
  XOR U31371 ( .A(n30264), .B(n30265), .Z(n30258) );
  AND U31372 ( .A(n30266), .B(n30267), .Z(n30265) );
  XOR U31373 ( .A(nreg[79]), .B(n30264), .Z(n30267) );
  XNOR U31374 ( .A(n23655), .B(n30264), .Z(n30266) );
  XOR U31375 ( .A(n30268), .B(n30269), .Z(n23655) );
  XOR U31376 ( .A(n30270), .B(n30271), .Z(n30264) );
  AND U31377 ( .A(n30272), .B(n30273), .Z(n30271) );
  XOR U31378 ( .A(nreg[78]), .B(n30270), .Z(n30273) );
  XNOR U31379 ( .A(n23667), .B(n30270), .Z(n30272) );
  XOR U31380 ( .A(n30274), .B(n30275), .Z(n23667) );
  XOR U31381 ( .A(n30276), .B(n30277), .Z(n30270) );
  AND U31382 ( .A(n30278), .B(n30279), .Z(n30277) );
  XOR U31383 ( .A(nreg[77]), .B(n30276), .Z(n30279) );
  XNOR U31384 ( .A(n23679), .B(n30276), .Z(n30278) );
  XOR U31385 ( .A(n30280), .B(n30281), .Z(n23679) );
  XOR U31386 ( .A(n30282), .B(n30283), .Z(n30276) );
  AND U31387 ( .A(n30284), .B(n30285), .Z(n30283) );
  XOR U31388 ( .A(nreg[76]), .B(n30282), .Z(n30285) );
  XNOR U31389 ( .A(n23691), .B(n30282), .Z(n30284) );
  XOR U31390 ( .A(n30286), .B(n30287), .Z(n23691) );
  XOR U31391 ( .A(n30288), .B(n30289), .Z(n30282) );
  AND U31392 ( .A(n30290), .B(n30291), .Z(n30289) );
  XOR U31393 ( .A(nreg[75]), .B(n30288), .Z(n30291) );
  XNOR U31394 ( .A(n23703), .B(n30288), .Z(n30290) );
  XOR U31395 ( .A(n30292), .B(n30293), .Z(n23703) );
  XOR U31396 ( .A(n30294), .B(n30295), .Z(n30288) );
  AND U31397 ( .A(n30296), .B(n30297), .Z(n30295) );
  XOR U31398 ( .A(nreg[74]), .B(n30294), .Z(n30297) );
  XNOR U31399 ( .A(n23715), .B(n30294), .Z(n30296) );
  XOR U31400 ( .A(n30298), .B(n30299), .Z(n23715) );
  XOR U31401 ( .A(n30300), .B(n30301), .Z(n30294) );
  AND U31402 ( .A(n30302), .B(n30303), .Z(n30301) );
  XOR U31403 ( .A(nreg[73]), .B(n30300), .Z(n30303) );
  XNOR U31404 ( .A(n23727), .B(n30300), .Z(n30302) );
  XOR U31405 ( .A(n30304), .B(n30305), .Z(n23727) );
  XOR U31406 ( .A(n30306), .B(n30307), .Z(n30300) );
  AND U31407 ( .A(n30308), .B(n30309), .Z(n30307) );
  XOR U31408 ( .A(nreg[72]), .B(n30306), .Z(n30309) );
  XNOR U31409 ( .A(n23739), .B(n30306), .Z(n30308) );
  XOR U31410 ( .A(n30310), .B(n30311), .Z(n23739) );
  XOR U31411 ( .A(n30312), .B(n30313), .Z(n30306) );
  AND U31412 ( .A(n30314), .B(n30315), .Z(n30313) );
  XOR U31413 ( .A(nreg[71]), .B(n30312), .Z(n30315) );
  XNOR U31414 ( .A(n23751), .B(n30312), .Z(n30314) );
  XOR U31415 ( .A(n30316), .B(n30317), .Z(n23751) );
  XOR U31416 ( .A(n30318), .B(n30319), .Z(n30312) );
  AND U31417 ( .A(n30320), .B(n30321), .Z(n30319) );
  XOR U31418 ( .A(nreg[70]), .B(n30318), .Z(n30321) );
  XNOR U31419 ( .A(n23763), .B(n30318), .Z(n30320) );
  XOR U31420 ( .A(n30322), .B(n30323), .Z(n23763) );
  XOR U31421 ( .A(n30324), .B(n30325), .Z(n30318) );
  AND U31422 ( .A(n30326), .B(n30327), .Z(n30325) );
  XOR U31423 ( .A(nreg[69]), .B(n30324), .Z(n30327) );
  XNOR U31424 ( .A(n23775), .B(n30324), .Z(n30326) );
  XOR U31425 ( .A(n30328), .B(n30329), .Z(n23775) );
  XOR U31426 ( .A(n30330), .B(n30331), .Z(n30324) );
  AND U31427 ( .A(n30332), .B(n30333), .Z(n30331) );
  XOR U31428 ( .A(nreg[68]), .B(n30330), .Z(n30333) );
  XNOR U31429 ( .A(n23787), .B(n30330), .Z(n30332) );
  XOR U31430 ( .A(n30334), .B(n30335), .Z(n23787) );
  XOR U31431 ( .A(n30336), .B(n30337), .Z(n30330) );
  AND U31432 ( .A(n30338), .B(n30339), .Z(n30337) );
  XOR U31433 ( .A(nreg[67]), .B(n30336), .Z(n30339) );
  XNOR U31434 ( .A(n23799), .B(n30336), .Z(n30338) );
  XOR U31435 ( .A(n30340), .B(n30341), .Z(n23799) );
  XOR U31436 ( .A(n30342), .B(n30343), .Z(n30336) );
  AND U31437 ( .A(n30344), .B(n30345), .Z(n30343) );
  XOR U31438 ( .A(nreg[66]), .B(n30342), .Z(n30345) );
  XNOR U31439 ( .A(n23811), .B(n30342), .Z(n30344) );
  XOR U31440 ( .A(n30346), .B(n30347), .Z(n23811) );
  XOR U31441 ( .A(n30348), .B(n30349), .Z(n30342) );
  AND U31442 ( .A(n30350), .B(n30351), .Z(n30349) );
  XOR U31443 ( .A(nreg[65]), .B(n30348), .Z(n30351) );
  XNOR U31444 ( .A(n23823), .B(n30348), .Z(n30350) );
  XOR U31445 ( .A(n30352), .B(n30353), .Z(n23823) );
  XOR U31446 ( .A(n30354), .B(n30355), .Z(n30348) );
  AND U31447 ( .A(n30356), .B(n30357), .Z(n30355) );
  XOR U31448 ( .A(nreg[64]), .B(n30354), .Z(n30357) );
  XNOR U31449 ( .A(n23835), .B(n30354), .Z(n30356) );
  XOR U31450 ( .A(n30358), .B(n30359), .Z(n23835) );
  XOR U31451 ( .A(n30360), .B(n30361), .Z(n30354) );
  AND U31452 ( .A(n30362), .B(n30363), .Z(n30361) );
  XOR U31453 ( .A(nreg[63]), .B(n30360), .Z(n30363) );
  XNOR U31454 ( .A(n23847), .B(n30360), .Z(n30362) );
  XOR U31455 ( .A(n30364), .B(n30365), .Z(n23847) );
  XOR U31456 ( .A(n30366), .B(n30367), .Z(n30360) );
  AND U31457 ( .A(n30368), .B(n30369), .Z(n30367) );
  XOR U31458 ( .A(nreg[62]), .B(n30366), .Z(n30369) );
  XNOR U31459 ( .A(n23859), .B(n30366), .Z(n30368) );
  XOR U31460 ( .A(n30370), .B(n30371), .Z(n23859) );
  XOR U31461 ( .A(n30372), .B(n30373), .Z(n30366) );
  AND U31462 ( .A(n30374), .B(n30375), .Z(n30373) );
  XOR U31463 ( .A(nreg[61]), .B(n30372), .Z(n30375) );
  XNOR U31464 ( .A(n23871), .B(n30372), .Z(n30374) );
  XOR U31465 ( .A(n30376), .B(n30377), .Z(n23871) );
  XOR U31466 ( .A(n30378), .B(n30379), .Z(n30372) );
  AND U31467 ( .A(n30380), .B(n30381), .Z(n30379) );
  XOR U31468 ( .A(nreg[60]), .B(n30378), .Z(n30381) );
  XNOR U31469 ( .A(n23883), .B(n30378), .Z(n30380) );
  XOR U31470 ( .A(n30382), .B(n30383), .Z(n23883) );
  XOR U31471 ( .A(n30384), .B(n30385), .Z(n30378) );
  AND U31472 ( .A(n30386), .B(n30387), .Z(n30385) );
  XOR U31473 ( .A(nreg[59]), .B(n30384), .Z(n30387) );
  XNOR U31474 ( .A(n23895), .B(n30384), .Z(n30386) );
  XOR U31475 ( .A(n30388), .B(n30389), .Z(n23895) );
  XOR U31476 ( .A(n30390), .B(n30391), .Z(n30384) );
  AND U31477 ( .A(n30392), .B(n30393), .Z(n30391) );
  XOR U31478 ( .A(nreg[58]), .B(n30390), .Z(n30393) );
  XNOR U31479 ( .A(n23907), .B(n30390), .Z(n30392) );
  XOR U31480 ( .A(n30394), .B(n30395), .Z(n23907) );
  XOR U31481 ( .A(n30396), .B(n30397), .Z(n30390) );
  AND U31482 ( .A(n30398), .B(n30399), .Z(n30397) );
  XOR U31483 ( .A(nreg[57]), .B(n30396), .Z(n30399) );
  XNOR U31484 ( .A(n23919), .B(n30396), .Z(n30398) );
  XOR U31485 ( .A(n30400), .B(n30401), .Z(n23919) );
  XOR U31486 ( .A(n30402), .B(n30403), .Z(n30396) );
  AND U31487 ( .A(n30404), .B(n30405), .Z(n30403) );
  XOR U31488 ( .A(nreg[56]), .B(n30402), .Z(n30405) );
  XNOR U31489 ( .A(n23931), .B(n30402), .Z(n30404) );
  XOR U31490 ( .A(n30406), .B(n30407), .Z(n23931) );
  XOR U31491 ( .A(n30408), .B(n30409), .Z(n30402) );
  AND U31492 ( .A(n30410), .B(n30411), .Z(n30409) );
  XOR U31493 ( .A(nreg[55]), .B(n30408), .Z(n30411) );
  XNOR U31494 ( .A(n23943), .B(n30408), .Z(n30410) );
  XOR U31495 ( .A(n30412), .B(n30413), .Z(n23943) );
  XOR U31496 ( .A(n30414), .B(n30415), .Z(n30408) );
  AND U31497 ( .A(n30416), .B(n30417), .Z(n30415) );
  XOR U31498 ( .A(nreg[54]), .B(n30414), .Z(n30417) );
  XNOR U31499 ( .A(n23955), .B(n30414), .Z(n30416) );
  XOR U31500 ( .A(n30418), .B(n30419), .Z(n23955) );
  XOR U31501 ( .A(n30420), .B(n30421), .Z(n30414) );
  AND U31502 ( .A(n30422), .B(n30423), .Z(n30421) );
  XOR U31503 ( .A(nreg[53]), .B(n30420), .Z(n30423) );
  XNOR U31504 ( .A(n23967), .B(n30420), .Z(n30422) );
  XOR U31505 ( .A(n30424), .B(n30425), .Z(n23967) );
  XOR U31506 ( .A(n30426), .B(n30427), .Z(n30420) );
  AND U31507 ( .A(n30428), .B(n30429), .Z(n30427) );
  XOR U31508 ( .A(nreg[52]), .B(n30426), .Z(n30429) );
  XNOR U31509 ( .A(n23979), .B(n30426), .Z(n30428) );
  XOR U31510 ( .A(n30430), .B(n30431), .Z(n23979) );
  XOR U31511 ( .A(n30432), .B(n30433), .Z(n30426) );
  AND U31512 ( .A(n30434), .B(n30435), .Z(n30433) );
  XOR U31513 ( .A(nreg[51]), .B(n30432), .Z(n30435) );
  XNOR U31514 ( .A(n23991), .B(n30432), .Z(n30434) );
  XOR U31515 ( .A(n30436), .B(n30437), .Z(n23991) );
  XOR U31516 ( .A(n30438), .B(n30439), .Z(n30432) );
  AND U31517 ( .A(n30440), .B(n30441), .Z(n30439) );
  XOR U31518 ( .A(nreg[50]), .B(n30438), .Z(n30441) );
  XNOR U31519 ( .A(n24003), .B(n30438), .Z(n30440) );
  XOR U31520 ( .A(n30442), .B(n30443), .Z(n24003) );
  XOR U31521 ( .A(n30444), .B(n30445), .Z(n30438) );
  AND U31522 ( .A(n30446), .B(n30447), .Z(n30445) );
  XOR U31523 ( .A(nreg[49]), .B(n30444), .Z(n30447) );
  XNOR U31524 ( .A(n24015), .B(n30444), .Z(n30446) );
  XOR U31525 ( .A(n30448), .B(n30449), .Z(n24015) );
  XOR U31526 ( .A(n30450), .B(n30451), .Z(n30444) );
  AND U31527 ( .A(n30452), .B(n30453), .Z(n30451) );
  XOR U31528 ( .A(nreg[48]), .B(n30450), .Z(n30453) );
  XNOR U31529 ( .A(n24027), .B(n30450), .Z(n30452) );
  XOR U31530 ( .A(n30454), .B(n30455), .Z(n24027) );
  XOR U31531 ( .A(n30456), .B(n30457), .Z(n30450) );
  AND U31532 ( .A(n30458), .B(n30459), .Z(n30457) );
  XOR U31533 ( .A(nreg[47]), .B(n30456), .Z(n30459) );
  XNOR U31534 ( .A(n24039), .B(n30456), .Z(n30458) );
  XOR U31535 ( .A(n30460), .B(n30461), .Z(n24039) );
  XOR U31536 ( .A(n30462), .B(n30463), .Z(n30456) );
  AND U31537 ( .A(n30464), .B(n30465), .Z(n30463) );
  XOR U31538 ( .A(nreg[46]), .B(n30462), .Z(n30465) );
  XNOR U31539 ( .A(n24051), .B(n30462), .Z(n30464) );
  XOR U31540 ( .A(n30466), .B(n30467), .Z(n24051) );
  XOR U31541 ( .A(n30468), .B(n30469), .Z(n30462) );
  AND U31542 ( .A(n30470), .B(n30471), .Z(n30469) );
  XOR U31543 ( .A(nreg[45]), .B(n30468), .Z(n30471) );
  XNOR U31544 ( .A(n24063), .B(n30468), .Z(n30470) );
  XOR U31545 ( .A(n30472), .B(n30473), .Z(n24063) );
  XOR U31546 ( .A(n30474), .B(n30475), .Z(n30468) );
  AND U31547 ( .A(n30476), .B(n30477), .Z(n30475) );
  XOR U31548 ( .A(nreg[44]), .B(n30474), .Z(n30477) );
  XNOR U31549 ( .A(n24075), .B(n30474), .Z(n30476) );
  XOR U31550 ( .A(n30478), .B(n30479), .Z(n24075) );
  XOR U31551 ( .A(n30480), .B(n30481), .Z(n30474) );
  AND U31552 ( .A(n30482), .B(n30483), .Z(n30481) );
  XOR U31553 ( .A(nreg[43]), .B(n30480), .Z(n30483) );
  XNOR U31554 ( .A(n24087), .B(n30480), .Z(n30482) );
  XOR U31555 ( .A(n30484), .B(n30485), .Z(n24087) );
  XOR U31556 ( .A(n30486), .B(n30487), .Z(n30480) );
  AND U31557 ( .A(n30488), .B(n30489), .Z(n30487) );
  XOR U31558 ( .A(nreg[42]), .B(n30486), .Z(n30489) );
  XNOR U31559 ( .A(n24099), .B(n30486), .Z(n30488) );
  XOR U31560 ( .A(n30490), .B(n30491), .Z(n24099) );
  XOR U31561 ( .A(n30492), .B(n30493), .Z(n30486) );
  AND U31562 ( .A(n30494), .B(n30495), .Z(n30493) );
  XOR U31563 ( .A(nreg[41]), .B(n30492), .Z(n30495) );
  XNOR U31564 ( .A(n24111), .B(n30492), .Z(n30494) );
  XOR U31565 ( .A(n30496), .B(n30497), .Z(n24111) );
  XOR U31566 ( .A(n30498), .B(n30499), .Z(n30492) );
  AND U31567 ( .A(n30500), .B(n30501), .Z(n30499) );
  XOR U31568 ( .A(nreg[40]), .B(n30498), .Z(n30501) );
  XNOR U31569 ( .A(n24123), .B(n30498), .Z(n30500) );
  XOR U31570 ( .A(n30502), .B(n30503), .Z(n24123) );
  XOR U31571 ( .A(n30504), .B(n30505), .Z(n30498) );
  AND U31572 ( .A(n30506), .B(n30507), .Z(n30505) );
  XOR U31573 ( .A(nreg[39]), .B(n30504), .Z(n30507) );
  XNOR U31574 ( .A(n24135), .B(n30504), .Z(n30506) );
  XOR U31575 ( .A(n30508), .B(n30509), .Z(n24135) );
  XOR U31576 ( .A(n30510), .B(n30511), .Z(n30504) );
  AND U31577 ( .A(n30512), .B(n30513), .Z(n30511) );
  XOR U31578 ( .A(nreg[38]), .B(n30510), .Z(n30513) );
  XNOR U31579 ( .A(n24147), .B(n30510), .Z(n30512) );
  XOR U31580 ( .A(n30514), .B(n30515), .Z(n24147) );
  XOR U31581 ( .A(n30516), .B(n30517), .Z(n30510) );
  AND U31582 ( .A(n30518), .B(n30519), .Z(n30517) );
  XOR U31583 ( .A(nreg[37]), .B(n30516), .Z(n30519) );
  XNOR U31584 ( .A(n24159), .B(n30516), .Z(n30518) );
  XOR U31585 ( .A(n30520), .B(n30521), .Z(n24159) );
  XOR U31586 ( .A(n30522), .B(n30523), .Z(n30516) );
  AND U31587 ( .A(n30524), .B(n30525), .Z(n30523) );
  XOR U31588 ( .A(nreg[36]), .B(n30522), .Z(n30525) );
  XNOR U31589 ( .A(n24171), .B(n30522), .Z(n30524) );
  XOR U31590 ( .A(n30526), .B(n30527), .Z(n24171) );
  XOR U31591 ( .A(n30528), .B(n30529), .Z(n30522) );
  AND U31592 ( .A(n30530), .B(n30531), .Z(n30529) );
  XOR U31593 ( .A(nreg[35]), .B(n30528), .Z(n30531) );
  XNOR U31594 ( .A(n24183), .B(n30528), .Z(n30530) );
  XOR U31595 ( .A(n30532), .B(n30533), .Z(n24183) );
  XOR U31596 ( .A(n30534), .B(n30535), .Z(n30528) );
  AND U31597 ( .A(n30536), .B(n30537), .Z(n30535) );
  XOR U31598 ( .A(nreg[34]), .B(n30534), .Z(n30537) );
  XNOR U31599 ( .A(n24195), .B(n30534), .Z(n30536) );
  XOR U31600 ( .A(n30538), .B(n30539), .Z(n24195) );
  XOR U31601 ( .A(n30540), .B(n30541), .Z(n30534) );
  AND U31602 ( .A(n30542), .B(n30543), .Z(n30541) );
  XOR U31603 ( .A(nreg[33]), .B(n30540), .Z(n30543) );
  XNOR U31604 ( .A(n24207), .B(n30540), .Z(n30542) );
  XOR U31605 ( .A(n30544), .B(n30545), .Z(n24207) );
  XOR U31606 ( .A(n30546), .B(n30547), .Z(n30540) );
  AND U31607 ( .A(n30548), .B(n30549), .Z(n30547) );
  XOR U31608 ( .A(nreg[32]), .B(n30546), .Z(n30549) );
  XNOR U31609 ( .A(n24219), .B(n30546), .Z(n30548) );
  XOR U31610 ( .A(n30550), .B(n30551), .Z(n24219) );
  XOR U31611 ( .A(n30552), .B(n30553), .Z(n30546) );
  AND U31612 ( .A(n30554), .B(n30555), .Z(n30553) );
  XOR U31613 ( .A(nreg[31]), .B(n30552), .Z(n30555) );
  XNOR U31614 ( .A(n24231), .B(n30552), .Z(n30554) );
  XOR U31615 ( .A(n30556), .B(n30557), .Z(n24231) );
  XOR U31616 ( .A(n30558), .B(n30559), .Z(n30552) );
  AND U31617 ( .A(n30560), .B(n30561), .Z(n30559) );
  XOR U31618 ( .A(nreg[30]), .B(n30558), .Z(n30561) );
  XNOR U31619 ( .A(n24243), .B(n30558), .Z(n30560) );
  XOR U31620 ( .A(n30562), .B(n30563), .Z(n24243) );
  XOR U31621 ( .A(n30564), .B(n30565), .Z(n30558) );
  AND U31622 ( .A(n30566), .B(n30567), .Z(n30565) );
  XOR U31623 ( .A(nreg[29]), .B(n30564), .Z(n30567) );
  XNOR U31624 ( .A(n24255), .B(n30564), .Z(n30566) );
  XOR U31625 ( .A(n30568), .B(n30569), .Z(n24255) );
  XOR U31626 ( .A(n30570), .B(n30571), .Z(n30564) );
  AND U31627 ( .A(n30572), .B(n30573), .Z(n30571) );
  XOR U31628 ( .A(nreg[28]), .B(n30570), .Z(n30573) );
  XNOR U31629 ( .A(n24267), .B(n30570), .Z(n30572) );
  XOR U31630 ( .A(n30574), .B(n30575), .Z(n24267) );
  XOR U31631 ( .A(n30576), .B(n30577), .Z(n30570) );
  AND U31632 ( .A(n30578), .B(n30579), .Z(n30577) );
  XOR U31633 ( .A(nreg[27]), .B(n30576), .Z(n30579) );
  XNOR U31634 ( .A(n24279), .B(n30576), .Z(n30578) );
  XOR U31635 ( .A(n30580), .B(n30581), .Z(n24279) );
  XOR U31636 ( .A(n30582), .B(n30583), .Z(n30576) );
  AND U31637 ( .A(n30584), .B(n30585), .Z(n30583) );
  XOR U31638 ( .A(nreg[26]), .B(n30582), .Z(n30585) );
  XNOR U31639 ( .A(n24291), .B(n30582), .Z(n30584) );
  XOR U31640 ( .A(n30586), .B(n30587), .Z(n24291) );
  XOR U31641 ( .A(n30588), .B(n30589), .Z(n30582) );
  AND U31642 ( .A(n30590), .B(n30591), .Z(n30589) );
  XOR U31643 ( .A(nreg[25]), .B(n30588), .Z(n30591) );
  XNOR U31644 ( .A(n24303), .B(n30588), .Z(n30590) );
  XOR U31645 ( .A(n30592), .B(n30593), .Z(n24303) );
  XOR U31646 ( .A(n30594), .B(n30595), .Z(n30588) );
  AND U31647 ( .A(n30596), .B(n30597), .Z(n30595) );
  XOR U31648 ( .A(nreg[24]), .B(n30594), .Z(n30597) );
  XNOR U31649 ( .A(n24315), .B(n30594), .Z(n30596) );
  XOR U31650 ( .A(n30598), .B(n30599), .Z(n24315) );
  XOR U31651 ( .A(n30600), .B(n30601), .Z(n30594) );
  AND U31652 ( .A(n30602), .B(n30603), .Z(n30601) );
  XOR U31653 ( .A(nreg[23]), .B(n30600), .Z(n30603) );
  XNOR U31654 ( .A(n24327), .B(n30600), .Z(n30602) );
  XOR U31655 ( .A(n30604), .B(n30605), .Z(n24327) );
  XOR U31656 ( .A(n30606), .B(n30607), .Z(n30600) );
  AND U31657 ( .A(n30608), .B(n30609), .Z(n30607) );
  XOR U31658 ( .A(nreg[22]), .B(n30606), .Z(n30609) );
  XNOR U31659 ( .A(n24339), .B(n30606), .Z(n30608) );
  XOR U31660 ( .A(n30610), .B(n30611), .Z(n24339) );
  XOR U31661 ( .A(n30612), .B(n30613), .Z(n30606) );
  AND U31662 ( .A(n30614), .B(n30615), .Z(n30613) );
  XOR U31663 ( .A(nreg[21]), .B(n30612), .Z(n30615) );
  XNOR U31664 ( .A(n24351), .B(n30612), .Z(n30614) );
  XOR U31665 ( .A(n30616), .B(n30617), .Z(n24351) );
  XOR U31666 ( .A(n30618), .B(n30619), .Z(n30612) );
  AND U31667 ( .A(n30620), .B(n30621), .Z(n30619) );
  XOR U31668 ( .A(nreg[20]), .B(n30618), .Z(n30621) );
  XNOR U31669 ( .A(n24363), .B(n30618), .Z(n30620) );
  XOR U31670 ( .A(n30622), .B(n30623), .Z(n24363) );
  XOR U31671 ( .A(n30624), .B(n30625), .Z(n30618) );
  AND U31672 ( .A(n30626), .B(n30627), .Z(n30625) );
  XOR U31673 ( .A(nreg[19]), .B(n30624), .Z(n30627) );
  XNOR U31674 ( .A(n24375), .B(n30624), .Z(n30626) );
  XOR U31675 ( .A(n30628), .B(n30629), .Z(n24375) );
  XOR U31676 ( .A(n30630), .B(n30631), .Z(n30624) );
  AND U31677 ( .A(n30632), .B(n30633), .Z(n30631) );
  XOR U31678 ( .A(nreg[18]), .B(n30630), .Z(n30633) );
  XNOR U31679 ( .A(n24387), .B(n30630), .Z(n30632) );
  XOR U31680 ( .A(n30634), .B(n30635), .Z(n24387) );
  XOR U31681 ( .A(n30636), .B(n30637), .Z(n30630) );
  AND U31682 ( .A(n30638), .B(n30639), .Z(n30637) );
  XOR U31683 ( .A(nreg[17]), .B(n30636), .Z(n30639) );
  XNOR U31684 ( .A(n24399), .B(n30636), .Z(n30638) );
  XOR U31685 ( .A(n30640), .B(n30641), .Z(n24399) );
  XOR U31686 ( .A(n30642), .B(n30643), .Z(n30636) );
  AND U31687 ( .A(n30644), .B(n30645), .Z(n30643) );
  XOR U31688 ( .A(nreg[16]), .B(n30642), .Z(n30645) );
  XNOR U31689 ( .A(n24411), .B(n30642), .Z(n30644) );
  XOR U31690 ( .A(n30646), .B(n30647), .Z(n24411) );
  XOR U31691 ( .A(n30648), .B(n30649), .Z(n30642) );
  AND U31692 ( .A(n30650), .B(n30651), .Z(n30649) );
  XOR U31693 ( .A(nreg[15]), .B(n30648), .Z(n30651) );
  XNOR U31694 ( .A(n24423), .B(n30648), .Z(n30650) );
  XOR U31695 ( .A(n30652), .B(n30653), .Z(n24423) );
  XOR U31696 ( .A(n30654), .B(n30655), .Z(n30648) );
  AND U31697 ( .A(n30656), .B(n30657), .Z(n30655) );
  XOR U31698 ( .A(nreg[14]), .B(n30654), .Z(n30657) );
  XNOR U31699 ( .A(n24435), .B(n30654), .Z(n30656) );
  XOR U31700 ( .A(n30658), .B(n30659), .Z(n24435) );
  XOR U31701 ( .A(n30660), .B(n30661), .Z(n30654) );
  AND U31702 ( .A(n30662), .B(n30663), .Z(n30661) );
  XOR U31703 ( .A(nreg[13]), .B(n30660), .Z(n30663) );
  XNOR U31704 ( .A(n24447), .B(n30660), .Z(n30662) );
  XOR U31705 ( .A(n30664), .B(n30665), .Z(n24447) );
  XOR U31706 ( .A(n30666), .B(n30667), .Z(n30660) );
  AND U31707 ( .A(n30668), .B(n30669), .Z(n30667) );
  XOR U31708 ( .A(nreg[12]), .B(n30666), .Z(n30669) );
  XNOR U31709 ( .A(n24459), .B(n30666), .Z(n30668) );
  XOR U31710 ( .A(n30670), .B(n30671), .Z(n24459) );
  XOR U31711 ( .A(n30672), .B(n30673), .Z(n30666) );
  AND U31712 ( .A(n30674), .B(n30675), .Z(n30673) );
  XOR U31713 ( .A(nreg[11]), .B(n30672), .Z(n30675) );
  XNOR U31714 ( .A(n24471), .B(n30672), .Z(n30674) );
  XOR U31715 ( .A(n30676), .B(n30677), .Z(n24471) );
  XOR U31716 ( .A(n30678), .B(n30679), .Z(n30672) );
  AND U31717 ( .A(n30680), .B(n30681), .Z(n30679) );
  XOR U31718 ( .A(nreg[10]), .B(n30678), .Z(n30681) );
  XNOR U31719 ( .A(n24483), .B(n30678), .Z(n30680) );
  XOR U31720 ( .A(n30682), .B(n30683), .Z(n24483) );
  XOR U31721 ( .A(n30684), .B(n30685), .Z(n30678) );
  AND U31722 ( .A(n30686), .B(n30687), .Z(n30685) );
  XOR U31723 ( .A(nreg[9]), .B(n30684), .Z(n30687) );
  XNOR U31724 ( .A(n24495), .B(n30684), .Z(n30686) );
  XOR U31725 ( .A(n30688), .B(n30689), .Z(n24495) );
  XOR U31726 ( .A(n30690), .B(n30691), .Z(n30684) );
  AND U31727 ( .A(n30692), .B(n30693), .Z(n30691) );
  XOR U31728 ( .A(nreg[8]), .B(n30690), .Z(n30693) );
  XNOR U31729 ( .A(n24507), .B(n30690), .Z(n30692) );
  XOR U31730 ( .A(n30694), .B(n30695), .Z(n24507) );
  XOR U31731 ( .A(n30696), .B(n30697), .Z(n30690) );
  AND U31732 ( .A(n30698), .B(n30699), .Z(n30697) );
  XOR U31733 ( .A(nreg[7]), .B(n30696), .Z(n30699) );
  XNOR U31734 ( .A(n24519), .B(n30696), .Z(n30698) );
  XOR U31735 ( .A(n30700), .B(n30701), .Z(n24519) );
  XOR U31736 ( .A(n30702), .B(n30703), .Z(n30696) );
  AND U31737 ( .A(n30704), .B(n30705), .Z(n30703) );
  XOR U31738 ( .A(nreg[6]), .B(n30702), .Z(n30705) );
  XNOR U31739 ( .A(n24531), .B(n30702), .Z(n30704) );
  XOR U31740 ( .A(n30706), .B(n30707), .Z(n24531) );
  XOR U31741 ( .A(n30708), .B(n30709), .Z(n30702) );
  AND U31742 ( .A(n30710), .B(n30711), .Z(n30709) );
  XOR U31743 ( .A(nreg[5]), .B(n30708), .Z(n30711) );
  XNOR U31744 ( .A(n24543), .B(n30708), .Z(n30710) );
  XOR U31745 ( .A(n30712), .B(n30713), .Z(n24543) );
  XOR U31746 ( .A(n30714), .B(n30715), .Z(n30708) );
  AND U31747 ( .A(n30716), .B(n30717), .Z(n30715) );
  XOR U31748 ( .A(nreg[4]), .B(n30714), .Z(n30717) );
  XNOR U31749 ( .A(n24555), .B(n30714), .Z(n30716) );
  XOR U31750 ( .A(n30718), .B(n30719), .Z(n24555) );
  XOR U31751 ( .A(n30720), .B(n30721), .Z(n30714) );
  AND U31752 ( .A(n30722), .B(n30723), .Z(n30721) );
  XOR U31753 ( .A(nreg[3]), .B(n30720), .Z(n30723) );
  XNOR U31754 ( .A(n24567), .B(n30720), .Z(n30722) );
  XOR U31755 ( .A(n30724), .B(n30725), .Z(n24567) );
  XNOR U31756 ( .A(n30726), .B(n30727), .Z(n30720) );
  AND U31757 ( .A(n30728), .B(n30729), .Z(n30727) );
  XNOR U31758 ( .A(nreg[2]), .B(n30726), .Z(n30729) );
  XNOR U31759 ( .A(n24579), .B(n30726), .Z(n30728) );
  XOR U31760 ( .A(n30730), .B(n30731), .Z(n24579) );
  XOR U31761 ( .A(n30732), .B(n30733), .Z(n30726) );
  NAND U31762 ( .A(n30734), .B(n30735), .Z(n30732) );
  XNOR U31763 ( .A(nreg[1]), .B(n30736), .Z(n30735) );
  IV U31764 ( .A(n30733), .Z(n30736) );
  XNOR U31765 ( .A(n24592), .B(n30733), .Z(n30734) );
  ANDN U31766 ( .A(nreg[0]), .B(n24589), .Z(n30733) );
  XOR U31767 ( .A(n30737), .B(n30738), .Z(n12309) );
  XOR U31768 ( .A(n30739), .B(\modmult_1/zin[0][1024] ), .Z(n30737) );
  NAND U31769 ( .A(n30738), .B(n12315), .Z(n30739) );
  XNOR U31770 ( .A(n30740), .B(\modmult_1/zin[0][1023] ), .Z(n12315) );
  IV U31771 ( .A(n30738), .Z(n30740) );
  XOR U31772 ( .A(n30741), .B(n30742), .Z(n30738) );
  ANDN U31773 ( .A(n30743), .B(n24605), .Z(n30742) );
  XOR U31774 ( .A(n30744), .B(\modmult_1/zin[0][1022] ), .Z(n24605) );
  IV U31775 ( .A(n30741), .Z(n30744) );
  XNOR U31776 ( .A(n30741), .B(n24604), .Z(n30743) );
  XOR U31777 ( .A(n30745), .B(n30746), .Z(n24604) );
  ANDN U31778 ( .A(\modmult_1/xin[1023] ), .B(n30745), .Z(n30746) );
  XOR U31779 ( .A(n30747), .B(mreg[1023]), .Z(n30745) );
  NAND U31780 ( .A(n30748), .B(mul_pow), .Z(n30747) );
  XOR U31781 ( .A(mreg[1023]), .B(creg[1023]), .Z(n30748) );
  XOR U31782 ( .A(n30749), .B(n30750), .Z(n30741) );
  ANDN U31783 ( .A(n30751), .B(n24611), .Z(n30750) );
  XOR U31784 ( .A(n30752), .B(\modmult_1/zin[0][1021] ), .Z(n24611) );
  IV U31785 ( .A(n30749), .Z(n30752) );
  XNOR U31786 ( .A(n30749), .B(n24610), .Z(n30751) );
  XOR U31787 ( .A(n30753), .B(n30754), .Z(n24610) );
  AND U31788 ( .A(\modmult_1/xin[1023] ), .B(n30755), .Z(n30754) );
  IV U31789 ( .A(n30753), .Z(n30755) );
  XOR U31790 ( .A(n30756), .B(mreg[1022]), .Z(n30753) );
  NAND U31791 ( .A(n30757), .B(mul_pow), .Z(n30756) );
  XOR U31792 ( .A(mreg[1022]), .B(creg[1022]), .Z(n30757) );
  XOR U31793 ( .A(n30758), .B(n30759), .Z(n30749) );
  ANDN U31794 ( .A(n30760), .B(n24617), .Z(n30759) );
  XOR U31795 ( .A(n30761), .B(\modmult_1/zin[0][1020] ), .Z(n24617) );
  IV U31796 ( .A(n30758), .Z(n30761) );
  XNOR U31797 ( .A(n30758), .B(n24616), .Z(n30760) );
  XOR U31798 ( .A(n30762), .B(n30763), .Z(n24616) );
  AND U31799 ( .A(\modmult_1/xin[1023] ), .B(n30764), .Z(n30763) );
  IV U31800 ( .A(n30762), .Z(n30764) );
  XOR U31801 ( .A(n30765), .B(mreg[1021]), .Z(n30762) );
  NAND U31802 ( .A(n30766), .B(mul_pow), .Z(n30765) );
  XOR U31803 ( .A(mreg[1021]), .B(creg[1021]), .Z(n30766) );
  XOR U31804 ( .A(n30767), .B(n30768), .Z(n30758) );
  ANDN U31805 ( .A(n30769), .B(n24623), .Z(n30768) );
  XOR U31806 ( .A(n30770), .B(\modmult_1/zin[0][1019] ), .Z(n24623) );
  IV U31807 ( .A(n30767), .Z(n30770) );
  XNOR U31808 ( .A(n30767), .B(n24622), .Z(n30769) );
  XOR U31809 ( .A(n30771), .B(n30772), .Z(n24622) );
  AND U31810 ( .A(\modmult_1/xin[1023] ), .B(n30773), .Z(n30772) );
  IV U31811 ( .A(n30771), .Z(n30773) );
  XOR U31812 ( .A(n30774), .B(mreg[1020]), .Z(n30771) );
  NAND U31813 ( .A(n30775), .B(mul_pow), .Z(n30774) );
  XOR U31814 ( .A(mreg[1020]), .B(creg[1020]), .Z(n30775) );
  XOR U31815 ( .A(n30776), .B(n30777), .Z(n30767) );
  ANDN U31816 ( .A(n30778), .B(n24629), .Z(n30777) );
  XOR U31817 ( .A(n30779), .B(\modmult_1/zin[0][1018] ), .Z(n24629) );
  IV U31818 ( .A(n30776), .Z(n30779) );
  XNOR U31819 ( .A(n30776), .B(n24628), .Z(n30778) );
  XOR U31820 ( .A(n30780), .B(n30781), .Z(n24628) );
  AND U31821 ( .A(\modmult_1/xin[1023] ), .B(n30782), .Z(n30781) );
  IV U31822 ( .A(n30780), .Z(n30782) );
  XOR U31823 ( .A(n30783), .B(mreg[1019]), .Z(n30780) );
  NAND U31824 ( .A(n30784), .B(mul_pow), .Z(n30783) );
  XOR U31825 ( .A(mreg[1019]), .B(creg[1019]), .Z(n30784) );
  XOR U31826 ( .A(n30785), .B(n30786), .Z(n30776) );
  ANDN U31827 ( .A(n30787), .B(n24635), .Z(n30786) );
  XOR U31828 ( .A(n30788), .B(\modmult_1/zin[0][1017] ), .Z(n24635) );
  IV U31829 ( .A(n30785), .Z(n30788) );
  XNOR U31830 ( .A(n30785), .B(n24634), .Z(n30787) );
  XOR U31831 ( .A(n30789), .B(n30790), .Z(n24634) );
  AND U31832 ( .A(\modmult_1/xin[1023] ), .B(n30791), .Z(n30790) );
  IV U31833 ( .A(n30789), .Z(n30791) );
  XOR U31834 ( .A(n30792), .B(mreg[1018]), .Z(n30789) );
  NAND U31835 ( .A(n30793), .B(mul_pow), .Z(n30792) );
  XOR U31836 ( .A(mreg[1018]), .B(creg[1018]), .Z(n30793) );
  XOR U31837 ( .A(n30794), .B(n30795), .Z(n30785) );
  ANDN U31838 ( .A(n30796), .B(n24641), .Z(n30795) );
  XOR U31839 ( .A(n30797), .B(\modmult_1/zin[0][1016] ), .Z(n24641) );
  IV U31840 ( .A(n30794), .Z(n30797) );
  XNOR U31841 ( .A(n30794), .B(n24640), .Z(n30796) );
  XOR U31842 ( .A(n30798), .B(n30799), .Z(n24640) );
  AND U31843 ( .A(\modmult_1/xin[1023] ), .B(n30800), .Z(n30799) );
  IV U31844 ( .A(n30798), .Z(n30800) );
  XOR U31845 ( .A(n30801), .B(mreg[1017]), .Z(n30798) );
  NAND U31846 ( .A(n30802), .B(mul_pow), .Z(n30801) );
  XOR U31847 ( .A(mreg[1017]), .B(creg[1017]), .Z(n30802) );
  XOR U31848 ( .A(n30803), .B(n30804), .Z(n30794) );
  ANDN U31849 ( .A(n30805), .B(n24647), .Z(n30804) );
  XOR U31850 ( .A(n30806), .B(\modmult_1/zin[0][1015] ), .Z(n24647) );
  IV U31851 ( .A(n30803), .Z(n30806) );
  XNOR U31852 ( .A(n30803), .B(n24646), .Z(n30805) );
  XOR U31853 ( .A(n30807), .B(n30808), .Z(n24646) );
  AND U31854 ( .A(\modmult_1/xin[1023] ), .B(n30809), .Z(n30808) );
  IV U31855 ( .A(n30807), .Z(n30809) );
  XOR U31856 ( .A(n30810), .B(mreg[1016]), .Z(n30807) );
  NAND U31857 ( .A(n30811), .B(mul_pow), .Z(n30810) );
  XOR U31858 ( .A(mreg[1016]), .B(creg[1016]), .Z(n30811) );
  XOR U31859 ( .A(n30812), .B(n30813), .Z(n30803) );
  ANDN U31860 ( .A(n30814), .B(n24653), .Z(n30813) );
  XOR U31861 ( .A(n30815), .B(\modmult_1/zin[0][1014] ), .Z(n24653) );
  IV U31862 ( .A(n30812), .Z(n30815) );
  XNOR U31863 ( .A(n30812), .B(n24652), .Z(n30814) );
  XOR U31864 ( .A(n30816), .B(n30817), .Z(n24652) );
  AND U31865 ( .A(\modmult_1/xin[1023] ), .B(n30818), .Z(n30817) );
  IV U31866 ( .A(n30816), .Z(n30818) );
  XOR U31867 ( .A(n30819), .B(mreg[1015]), .Z(n30816) );
  NAND U31868 ( .A(n30820), .B(mul_pow), .Z(n30819) );
  XOR U31869 ( .A(mreg[1015]), .B(creg[1015]), .Z(n30820) );
  XOR U31870 ( .A(n30821), .B(n30822), .Z(n30812) );
  ANDN U31871 ( .A(n30823), .B(n24659), .Z(n30822) );
  XOR U31872 ( .A(n30824), .B(\modmult_1/zin[0][1013] ), .Z(n24659) );
  IV U31873 ( .A(n30821), .Z(n30824) );
  XNOR U31874 ( .A(n30821), .B(n24658), .Z(n30823) );
  XOR U31875 ( .A(n30825), .B(n30826), .Z(n24658) );
  AND U31876 ( .A(\modmult_1/xin[1023] ), .B(n30827), .Z(n30826) );
  IV U31877 ( .A(n30825), .Z(n30827) );
  XOR U31878 ( .A(n30828), .B(mreg[1014]), .Z(n30825) );
  NAND U31879 ( .A(n30829), .B(mul_pow), .Z(n30828) );
  XOR U31880 ( .A(mreg[1014]), .B(creg[1014]), .Z(n30829) );
  XOR U31881 ( .A(n30830), .B(n30831), .Z(n30821) );
  ANDN U31882 ( .A(n30832), .B(n24665), .Z(n30831) );
  XOR U31883 ( .A(n30833), .B(\modmult_1/zin[0][1012] ), .Z(n24665) );
  IV U31884 ( .A(n30830), .Z(n30833) );
  XNOR U31885 ( .A(n30830), .B(n24664), .Z(n30832) );
  XOR U31886 ( .A(n30834), .B(n30835), .Z(n24664) );
  AND U31887 ( .A(\modmult_1/xin[1023] ), .B(n30836), .Z(n30835) );
  IV U31888 ( .A(n30834), .Z(n30836) );
  XOR U31889 ( .A(n30837), .B(mreg[1013]), .Z(n30834) );
  NAND U31890 ( .A(n30838), .B(mul_pow), .Z(n30837) );
  XOR U31891 ( .A(mreg[1013]), .B(creg[1013]), .Z(n30838) );
  XOR U31892 ( .A(n30839), .B(n30840), .Z(n30830) );
  ANDN U31893 ( .A(n30841), .B(n24671), .Z(n30840) );
  XOR U31894 ( .A(n30842), .B(\modmult_1/zin[0][1011] ), .Z(n24671) );
  IV U31895 ( .A(n30839), .Z(n30842) );
  XNOR U31896 ( .A(n30839), .B(n24670), .Z(n30841) );
  XOR U31897 ( .A(n30843), .B(n30844), .Z(n24670) );
  AND U31898 ( .A(\modmult_1/xin[1023] ), .B(n30845), .Z(n30844) );
  IV U31899 ( .A(n30843), .Z(n30845) );
  XOR U31900 ( .A(n30846), .B(mreg[1012]), .Z(n30843) );
  NAND U31901 ( .A(n30847), .B(mul_pow), .Z(n30846) );
  XOR U31902 ( .A(mreg[1012]), .B(creg[1012]), .Z(n30847) );
  XOR U31903 ( .A(n30848), .B(n30849), .Z(n30839) );
  ANDN U31904 ( .A(n30850), .B(n24677), .Z(n30849) );
  XOR U31905 ( .A(n30851), .B(\modmult_1/zin[0][1010] ), .Z(n24677) );
  IV U31906 ( .A(n30848), .Z(n30851) );
  XNOR U31907 ( .A(n30848), .B(n24676), .Z(n30850) );
  XOR U31908 ( .A(n30852), .B(n30853), .Z(n24676) );
  AND U31909 ( .A(\modmult_1/xin[1023] ), .B(n30854), .Z(n30853) );
  IV U31910 ( .A(n30852), .Z(n30854) );
  XOR U31911 ( .A(n30855), .B(mreg[1011]), .Z(n30852) );
  NAND U31912 ( .A(n30856), .B(mul_pow), .Z(n30855) );
  XOR U31913 ( .A(mreg[1011]), .B(creg[1011]), .Z(n30856) );
  XOR U31914 ( .A(n30857), .B(n30858), .Z(n30848) );
  ANDN U31915 ( .A(n30859), .B(n24683), .Z(n30858) );
  XOR U31916 ( .A(n30860), .B(\modmult_1/zin[0][1009] ), .Z(n24683) );
  IV U31917 ( .A(n30857), .Z(n30860) );
  XNOR U31918 ( .A(n30857), .B(n24682), .Z(n30859) );
  XOR U31919 ( .A(n30861), .B(n30862), .Z(n24682) );
  AND U31920 ( .A(\modmult_1/xin[1023] ), .B(n30863), .Z(n30862) );
  IV U31921 ( .A(n30861), .Z(n30863) );
  XOR U31922 ( .A(n30864), .B(mreg[1010]), .Z(n30861) );
  NAND U31923 ( .A(n30865), .B(mul_pow), .Z(n30864) );
  XOR U31924 ( .A(mreg[1010]), .B(creg[1010]), .Z(n30865) );
  XOR U31925 ( .A(n30866), .B(n30867), .Z(n30857) );
  ANDN U31926 ( .A(n30868), .B(n24689), .Z(n30867) );
  XOR U31927 ( .A(n30869), .B(\modmult_1/zin[0][1008] ), .Z(n24689) );
  IV U31928 ( .A(n30866), .Z(n30869) );
  XNOR U31929 ( .A(n30866), .B(n24688), .Z(n30868) );
  XOR U31930 ( .A(n30870), .B(n30871), .Z(n24688) );
  AND U31931 ( .A(\modmult_1/xin[1023] ), .B(n30872), .Z(n30871) );
  IV U31932 ( .A(n30870), .Z(n30872) );
  XOR U31933 ( .A(n30873), .B(mreg[1009]), .Z(n30870) );
  NAND U31934 ( .A(n30874), .B(mul_pow), .Z(n30873) );
  XOR U31935 ( .A(mreg[1009]), .B(creg[1009]), .Z(n30874) );
  XOR U31936 ( .A(n30875), .B(n30876), .Z(n30866) );
  ANDN U31937 ( .A(n30877), .B(n24695), .Z(n30876) );
  XOR U31938 ( .A(n30878), .B(\modmult_1/zin[0][1007] ), .Z(n24695) );
  IV U31939 ( .A(n30875), .Z(n30878) );
  XNOR U31940 ( .A(n30875), .B(n24694), .Z(n30877) );
  XOR U31941 ( .A(n30879), .B(n30880), .Z(n24694) );
  AND U31942 ( .A(\modmult_1/xin[1023] ), .B(n30881), .Z(n30880) );
  IV U31943 ( .A(n30879), .Z(n30881) );
  XOR U31944 ( .A(n30882), .B(mreg[1008]), .Z(n30879) );
  NAND U31945 ( .A(n30883), .B(mul_pow), .Z(n30882) );
  XOR U31946 ( .A(mreg[1008]), .B(creg[1008]), .Z(n30883) );
  XOR U31947 ( .A(n30884), .B(n30885), .Z(n30875) );
  ANDN U31948 ( .A(n30886), .B(n24701), .Z(n30885) );
  XOR U31949 ( .A(n30887), .B(\modmult_1/zin[0][1006] ), .Z(n24701) );
  IV U31950 ( .A(n30884), .Z(n30887) );
  XNOR U31951 ( .A(n30884), .B(n24700), .Z(n30886) );
  XOR U31952 ( .A(n30888), .B(n30889), .Z(n24700) );
  AND U31953 ( .A(\modmult_1/xin[1023] ), .B(n30890), .Z(n30889) );
  IV U31954 ( .A(n30888), .Z(n30890) );
  XOR U31955 ( .A(n30891), .B(mreg[1007]), .Z(n30888) );
  NAND U31956 ( .A(n30892), .B(mul_pow), .Z(n30891) );
  XOR U31957 ( .A(mreg[1007]), .B(creg[1007]), .Z(n30892) );
  XOR U31958 ( .A(n30893), .B(n30894), .Z(n30884) );
  ANDN U31959 ( .A(n30895), .B(n24707), .Z(n30894) );
  XOR U31960 ( .A(n30896), .B(\modmult_1/zin[0][1005] ), .Z(n24707) );
  IV U31961 ( .A(n30893), .Z(n30896) );
  XNOR U31962 ( .A(n30893), .B(n24706), .Z(n30895) );
  XOR U31963 ( .A(n30897), .B(n30898), .Z(n24706) );
  AND U31964 ( .A(\modmult_1/xin[1023] ), .B(n30899), .Z(n30898) );
  IV U31965 ( .A(n30897), .Z(n30899) );
  XOR U31966 ( .A(n30900), .B(mreg[1006]), .Z(n30897) );
  NAND U31967 ( .A(n30901), .B(mul_pow), .Z(n30900) );
  XOR U31968 ( .A(mreg[1006]), .B(creg[1006]), .Z(n30901) );
  XOR U31969 ( .A(n30902), .B(n30903), .Z(n30893) );
  ANDN U31970 ( .A(n30904), .B(n24713), .Z(n30903) );
  XOR U31971 ( .A(n30905), .B(\modmult_1/zin[0][1004] ), .Z(n24713) );
  IV U31972 ( .A(n30902), .Z(n30905) );
  XNOR U31973 ( .A(n30902), .B(n24712), .Z(n30904) );
  XOR U31974 ( .A(n30906), .B(n30907), .Z(n24712) );
  AND U31975 ( .A(\modmult_1/xin[1023] ), .B(n30908), .Z(n30907) );
  IV U31976 ( .A(n30906), .Z(n30908) );
  XOR U31977 ( .A(n30909), .B(mreg[1005]), .Z(n30906) );
  NAND U31978 ( .A(n30910), .B(mul_pow), .Z(n30909) );
  XOR U31979 ( .A(mreg[1005]), .B(creg[1005]), .Z(n30910) );
  XOR U31980 ( .A(n30911), .B(n30912), .Z(n30902) );
  ANDN U31981 ( .A(n30913), .B(n24719), .Z(n30912) );
  XOR U31982 ( .A(n30914), .B(\modmult_1/zin[0][1003] ), .Z(n24719) );
  IV U31983 ( .A(n30911), .Z(n30914) );
  XNOR U31984 ( .A(n30911), .B(n24718), .Z(n30913) );
  XOR U31985 ( .A(n30915), .B(n30916), .Z(n24718) );
  AND U31986 ( .A(\modmult_1/xin[1023] ), .B(n30917), .Z(n30916) );
  IV U31987 ( .A(n30915), .Z(n30917) );
  XOR U31988 ( .A(n30918), .B(mreg[1004]), .Z(n30915) );
  NAND U31989 ( .A(n30919), .B(mul_pow), .Z(n30918) );
  XOR U31990 ( .A(mreg[1004]), .B(creg[1004]), .Z(n30919) );
  XOR U31991 ( .A(n30920), .B(n30921), .Z(n30911) );
  ANDN U31992 ( .A(n30922), .B(n24725), .Z(n30921) );
  XOR U31993 ( .A(n30923), .B(\modmult_1/zin[0][1002] ), .Z(n24725) );
  IV U31994 ( .A(n30920), .Z(n30923) );
  XNOR U31995 ( .A(n30920), .B(n24724), .Z(n30922) );
  XOR U31996 ( .A(n30924), .B(n30925), .Z(n24724) );
  AND U31997 ( .A(\modmult_1/xin[1023] ), .B(n30926), .Z(n30925) );
  IV U31998 ( .A(n30924), .Z(n30926) );
  XOR U31999 ( .A(n30927), .B(mreg[1003]), .Z(n30924) );
  NAND U32000 ( .A(n30928), .B(mul_pow), .Z(n30927) );
  XOR U32001 ( .A(mreg[1003]), .B(creg[1003]), .Z(n30928) );
  XOR U32002 ( .A(n30929), .B(n30930), .Z(n30920) );
  ANDN U32003 ( .A(n30931), .B(n24731), .Z(n30930) );
  XOR U32004 ( .A(n30932), .B(\modmult_1/zin[0][1001] ), .Z(n24731) );
  IV U32005 ( .A(n30929), .Z(n30932) );
  XNOR U32006 ( .A(n30929), .B(n24730), .Z(n30931) );
  XOR U32007 ( .A(n30933), .B(n30934), .Z(n24730) );
  AND U32008 ( .A(\modmult_1/xin[1023] ), .B(n30935), .Z(n30934) );
  IV U32009 ( .A(n30933), .Z(n30935) );
  XOR U32010 ( .A(n30936), .B(mreg[1002]), .Z(n30933) );
  NAND U32011 ( .A(n30937), .B(mul_pow), .Z(n30936) );
  XOR U32012 ( .A(mreg[1002]), .B(creg[1002]), .Z(n30937) );
  XOR U32013 ( .A(n30938), .B(n30939), .Z(n30929) );
  ANDN U32014 ( .A(n30940), .B(n24737), .Z(n30939) );
  XOR U32015 ( .A(n30941), .B(\modmult_1/zin[0][1000] ), .Z(n24737) );
  IV U32016 ( .A(n30938), .Z(n30941) );
  XNOR U32017 ( .A(n30938), .B(n24736), .Z(n30940) );
  XOR U32018 ( .A(n30942), .B(n30943), .Z(n24736) );
  AND U32019 ( .A(\modmult_1/xin[1023] ), .B(n30944), .Z(n30943) );
  IV U32020 ( .A(n30942), .Z(n30944) );
  XOR U32021 ( .A(n30945), .B(mreg[1001]), .Z(n30942) );
  NAND U32022 ( .A(n30946), .B(mul_pow), .Z(n30945) );
  XOR U32023 ( .A(mreg[1001]), .B(creg[1001]), .Z(n30946) );
  XOR U32024 ( .A(n30947), .B(n30948), .Z(n30938) );
  ANDN U32025 ( .A(n30949), .B(n24743), .Z(n30948) );
  XOR U32026 ( .A(n30950), .B(\modmult_1/zin[0][999] ), .Z(n24743) );
  IV U32027 ( .A(n30947), .Z(n30950) );
  XNOR U32028 ( .A(n30947), .B(n24742), .Z(n30949) );
  XOR U32029 ( .A(n30951), .B(n30952), .Z(n24742) );
  AND U32030 ( .A(\modmult_1/xin[1023] ), .B(n30953), .Z(n30952) );
  IV U32031 ( .A(n30951), .Z(n30953) );
  XOR U32032 ( .A(n30954), .B(mreg[1000]), .Z(n30951) );
  NAND U32033 ( .A(n30955), .B(mul_pow), .Z(n30954) );
  XOR U32034 ( .A(mreg[1000]), .B(creg[1000]), .Z(n30955) );
  XOR U32035 ( .A(n30956), .B(n30957), .Z(n30947) );
  ANDN U32036 ( .A(n30958), .B(n24749), .Z(n30957) );
  XOR U32037 ( .A(n30959), .B(\modmult_1/zin[0][998] ), .Z(n24749) );
  IV U32038 ( .A(n30956), .Z(n30959) );
  XNOR U32039 ( .A(n30956), .B(n24748), .Z(n30958) );
  XOR U32040 ( .A(n30960), .B(n30961), .Z(n24748) );
  AND U32041 ( .A(\modmult_1/xin[1023] ), .B(n30962), .Z(n30961) );
  IV U32042 ( .A(n30960), .Z(n30962) );
  XOR U32043 ( .A(n30963), .B(mreg[999]), .Z(n30960) );
  NAND U32044 ( .A(n30964), .B(mul_pow), .Z(n30963) );
  XOR U32045 ( .A(mreg[999]), .B(creg[999]), .Z(n30964) );
  XOR U32046 ( .A(n30965), .B(n30966), .Z(n30956) );
  ANDN U32047 ( .A(n30967), .B(n24755), .Z(n30966) );
  XOR U32048 ( .A(n30968), .B(\modmult_1/zin[0][997] ), .Z(n24755) );
  IV U32049 ( .A(n30965), .Z(n30968) );
  XNOR U32050 ( .A(n30965), .B(n24754), .Z(n30967) );
  XOR U32051 ( .A(n30969), .B(n30970), .Z(n24754) );
  AND U32052 ( .A(\modmult_1/xin[1023] ), .B(n30971), .Z(n30970) );
  IV U32053 ( .A(n30969), .Z(n30971) );
  XOR U32054 ( .A(n30972), .B(mreg[998]), .Z(n30969) );
  NAND U32055 ( .A(n30973), .B(mul_pow), .Z(n30972) );
  XOR U32056 ( .A(mreg[998]), .B(creg[998]), .Z(n30973) );
  XOR U32057 ( .A(n30974), .B(n30975), .Z(n30965) );
  ANDN U32058 ( .A(n30976), .B(n24761), .Z(n30975) );
  XOR U32059 ( .A(n30977), .B(\modmult_1/zin[0][996] ), .Z(n24761) );
  IV U32060 ( .A(n30974), .Z(n30977) );
  XNOR U32061 ( .A(n30974), .B(n24760), .Z(n30976) );
  XOR U32062 ( .A(n30978), .B(n30979), .Z(n24760) );
  AND U32063 ( .A(\modmult_1/xin[1023] ), .B(n30980), .Z(n30979) );
  IV U32064 ( .A(n30978), .Z(n30980) );
  XOR U32065 ( .A(n30981), .B(mreg[997]), .Z(n30978) );
  NAND U32066 ( .A(n30982), .B(mul_pow), .Z(n30981) );
  XOR U32067 ( .A(mreg[997]), .B(creg[997]), .Z(n30982) );
  XOR U32068 ( .A(n30983), .B(n30984), .Z(n30974) );
  ANDN U32069 ( .A(n30985), .B(n24767), .Z(n30984) );
  XOR U32070 ( .A(n30986), .B(\modmult_1/zin[0][995] ), .Z(n24767) );
  IV U32071 ( .A(n30983), .Z(n30986) );
  XNOR U32072 ( .A(n30983), .B(n24766), .Z(n30985) );
  XOR U32073 ( .A(n30987), .B(n30988), .Z(n24766) );
  AND U32074 ( .A(\modmult_1/xin[1023] ), .B(n30989), .Z(n30988) );
  IV U32075 ( .A(n30987), .Z(n30989) );
  XOR U32076 ( .A(n30990), .B(mreg[996]), .Z(n30987) );
  NAND U32077 ( .A(n30991), .B(mul_pow), .Z(n30990) );
  XOR U32078 ( .A(mreg[996]), .B(creg[996]), .Z(n30991) );
  XOR U32079 ( .A(n30992), .B(n30993), .Z(n30983) );
  ANDN U32080 ( .A(n30994), .B(n24773), .Z(n30993) );
  XOR U32081 ( .A(n30995), .B(\modmult_1/zin[0][994] ), .Z(n24773) );
  IV U32082 ( .A(n30992), .Z(n30995) );
  XNOR U32083 ( .A(n30992), .B(n24772), .Z(n30994) );
  XOR U32084 ( .A(n30996), .B(n30997), .Z(n24772) );
  AND U32085 ( .A(\modmult_1/xin[1023] ), .B(n30998), .Z(n30997) );
  IV U32086 ( .A(n30996), .Z(n30998) );
  XOR U32087 ( .A(n30999), .B(mreg[995]), .Z(n30996) );
  NAND U32088 ( .A(n31000), .B(mul_pow), .Z(n30999) );
  XOR U32089 ( .A(mreg[995]), .B(creg[995]), .Z(n31000) );
  XOR U32090 ( .A(n31001), .B(n31002), .Z(n30992) );
  ANDN U32091 ( .A(n31003), .B(n24779), .Z(n31002) );
  XOR U32092 ( .A(n31004), .B(\modmult_1/zin[0][993] ), .Z(n24779) );
  IV U32093 ( .A(n31001), .Z(n31004) );
  XNOR U32094 ( .A(n31001), .B(n24778), .Z(n31003) );
  XOR U32095 ( .A(n31005), .B(n31006), .Z(n24778) );
  AND U32096 ( .A(\modmult_1/xin[1023] ), .B(n31007), .Z(n31006) );
  IV U32097 ( .A(n31005), .Z(n31007) );
  XOR U32098 ( .A(n31008), .B(mreg[994]), .Z(n31005) );
  NAND U32099 ( .A(n31009), .B(mul_pow), .Z(n31008) );
  XOR U32100 ( .A(mreg[994]), .B(creg[994]), .Z(n31009) );
  XOR U32101 ( .A(n31010), .B(n31011), .Z(n31001) );
  ANDN U32102 ( .A(n31012), .B(n24785), .Z(n31011) );
  XOR U32103 ( .A(n31013), .B(\modmult_1/zin[0][992] ), .Z(n24785) );
  IV U32104 ( .A(n31010), .Z(n31013) );
  XNOR U32105 ( .A(n31010), .B(n24784), .Z(n31012) );
  XOR U32106 ( .A(n31014), .B(n31015), .Z(n24784) );
  AND U32107 ( .A(\modmult_1/xin[1023] ), .B(n31016), .Z(n31015) );
  IV U32108 ( .A(n31014), .Z(n31016) );
  XOR U32109 ( .A(n31017), .B(mreg[993]), .Z(n31014) );
  NAND U32110 ( .A(n31018), .B(mul_pow), .Z(n31017) );
  XOR U32111 ( .A(mreg[993]), .B(creg[993]), .Z(n31018) );
  XOR U32112 ( .A(n31019), .B(n31020), .Z(n31010) );
  ANDN U32113 ( .A(n31021), .B(n24791), .Z(n31020) );
  XOR U32114 ( .A(n31022), .B(\modmult_1/zin[0][991] ), .Z(n24791) );
  IV U32115 ( .A(n31019), .Z(n31022) );
  XNOR U32116 ( .A(n31019), .B(n24790), .Z(n31021) );
  XOR U32117 ( .A(n31023), .B(n31024), .Z(n24790) );
  AND U32118 ( .A(\modmult_1/xin[1023] ), .B(n31025), .Z(n31024) );
  IV U32119 ( .A(n31023), .Z(n31025) );
  XOR U32120 ( .A(n31026), .B(mreg[992]), .Z(n31023) );
  NAND U32121 ( .A(n31027), .B(mul_pow), .Z(n31026) );
  XOR U32122 ( .A(mreg[992]), .B(creg[992]), .Z(n31027) );
  XOR U32123 ( .A(n31028), .B(n31029), .Z(n31019) );
  ANDN U32124 ( .A(n31030), .B(n24797), .Z(n31029) );
  XOR U32125 ( .A(n31031), .B(\modmult_1/zin[0][990] ), .Z(n24797) );
  IV U32126 ( .A(n31028), .Z(n31031) );
  XNOR U32127 ( .A(n31028), .B(n24796), .Z(n31030) );
  XOR U32128 ( .A(n31032), .B(n31033), .Z(n24796) );
  AND U32129 ( .A(\modmult_1/xin[1023] ), .B(n31034), .Z(n31033) );
  IV U32130 ( .A(n31032), .Z(n31034) );
  XOR U32131 ( .A(n31035), .B(mreg[991]), .Z(n31032) );
  NAND U32132 ( .A(n31036), .B(mul_pow), .Z(n31035) );
  XOR U32133 ( .A(mreg[991]), .B(creg[991]), .Z(n31036) );
  XOR U32134 ( .A(n31037), .B(n31038), .Z(n31028) );
  ANDN U32135 ( .A(n31039), .B(n24803), .Z(n31038) );
  XOR U32136 ( .A(n31040), .B(\modmult_1/zin[0][989] ), .Z(n24803) );
  IV U32137 ( .A(n31037), .Z(n31040) );
  XNOR U32138 ( .A(n31037), .B(n24802), .Z(n31039) );
  XOR U32139 ( .A(n31041), .B(n31042), .Z(n24802) );
  AND U32140 ( .A(\modmult_1/xin[1023] ), .B(n31043), .Z(n31042) );
  IV U32141 ( .A(n31041), .Z(n31043) );
  XOR U32142 ( .A(n31044), .B(mreg[990]), .Z(n31041) );
  NAND U32143 ( .A(n31045), .B(mul_pow), .Z(n31044) );
  XOR U32144 ( .A(mreg[990]), .B(creg[990]), .Z(n31045) );
  XOR U32145 ( .A(n31046), .B(n31047), .Z(n31037) );
  ANDN U32146 ( .A(n31048), .B(n24809), .Z(n31047) );
  XOR U32147 ( .A(n31049), .B(\modmult_1/zin[0][988] ), .Z(n24809) );
  IV U32148 ( .A(n31046), .Z(n31049) );
  XNOR U32149 ( .A(n31046), .B(n24808), .Z(n31048) );
  XOR U32150 ( .A(n31050), .B(n31051), .Z(n24808) );
  AND U32151 ( .A(\modmult_1/xin[1023] ), .B(n31052), .Z(n31051) );
  IV U32152 ( .A(n31050), .Z(n31052) );
  XOR U32153 ( .A(n31053), .B(mreg[989]), .Z(n31050) );
  NAND U32154 ( .A(n31054), .B(mul_pow), .Z(n31053) );
  XOR U32155 ( .A(mreg[989]), .B(creg[989]), .Z(n31054) );
  XOR U32156 ( .A(n31055), .B(n31056), .Z(n31046) );
  ANDN U32157 ( .A(n31057), .B(n24815), .Z(n31056) );
  XOR U32158 ( .A(n31058), .B(\modmult_1/zin[0][987] ), .Z(n24815) );
  IV U32159 ( .A(n31055), .Z(n31058) );
  XNOR U32160 ( .A(n31055), .B(n24814), .Z(n31057) );
  XOR U32161 ( .A(n31059), .B(n31060), .Z(n24814) );
  AND U32162 ( .A(\modmult_1/xin[1023] ), .B(n31061), .Z(n31060) );
  IV U32163 ( .A(n31059), .Z(n31061) );
  XOR U32164 ( .A(n31062), .B(mreg[988]), .Z(n31059) );
  NAND U32165 ( .A(n31063), .B(mul_pow), .Z(n31062) );
  XOR U32166 ( .A(mreg[988]), .B(creg[988]), .Z(n31063) );
  XOR U32167 ( .A(n31064), .B(n31065), .Z(n31055) );
  ANDN U32168 ( .A(n31066), .B(n24821), .Z(n31065) );
  XOR U32169 ( .A(n31067), .B(\modmult_1/zin[0][986] ), .Z(n24821) );
  IV U32170 ( .A(n31064), .Z(n31067) );
  XNOR U32171 ( .A(n31064), .B(n24820), .Z(n31066) );
  XOR U32172 ( .A(n31068), .B(n31069), .Z(n24820) );
  AND U32173 ( .A(\modmult_1/xin[1023] ), .B(n31070), .Z(n31069) );
  IV U32174 ( .A(n31068), .Z(n31070) );
  XOR U32175 ( .A(n31071), .B(mreg[987]), .Z(n31068) );
  NAND U32176 ( .A(n31072), .B(mul_pow), .Z(n31071) );
  XOR U32177 ( .A(mreg[987]), .B(creg[987]), .Z(n31072) );
  XOR U32178 ( .A(n31073), .B(n31074), .Z(n31064) );
  ANDN U32179 ( .A(n31075), .B(n24827), .Z(n31074) );
  XOR U32180 ( .A(n31076), .B(\modmult_1/zin[0][985] ), .Z(n24827) );
  IV U32181 ( .A(n31073), .Z(n31076) );
  XNOR U32182 ( .A(n31073), .B(n24826), .Z(n31075) );
  XOR U32183 ( .A(n31077), .B(n31078), .Z(n24826) );
  AND U32184 ( .A(\modmult_1/xin[1023] ), .B(n31079), .Z(n31078) );
  IV U32185 ( .A(n31077), .Z(n31079) );
  XOR U32186 ( .A(n31080), .B(mreg[986]), .Z(n31077) );
  NAND U32187 ( .A(n31081), .B(mul_pow), .Z(n31080) );
  XOR U32188 ( .A(mreg[986]), .B(creg[986]), .Z(n31081) );
  XOR U32189 ( .A(n31082), .B(n31083), .Z(n31073) );
  ANDN U32190 ( .A(n31084), .B(n24833), .Z(n31083) );
  XOR U32191 ( .A(n31085), .B(\modmult_1/zin[0][984] ), .Z(n24833) );
  IV U32192 ( .A(n31082), .Z(n31085) );
  XNOR U32193 ( .A(n31082), .B(n24832), .Z(n31084) );
  XOR U32194 ( .A(n31086), .B(n31087), .Z(n24832) );
  AND U32195 ( .A(\modmult_1/xin[1023] ), .B(n31088), .Z(n31087) );
  IV U32196 ( .A(n31086), .Z(n31088) );
  XOR U32197 ( .A(n31089), .B(mreg[985]), .Z(n31086) );
  NAND U32198 ( .A(n31090), .B(mul_pow), .Z(n31089) );
  XOR U32199 ( .A(mreg[985]), .B(creg[985]), .Z(n31090) );
  XOR U32200 ( .A(n31091), .B(n31092), .Z(n31082) );
  ANDN U32201 ( .A(n31093), .B(n24839), .Z(n31092) );
  XOR U32202 ( .A(n31094), .B(\modmult_1/zin[0][983] ), .Z(n24839) );
  IV U32203 ( .A(n31091), .Z(n31094) );
  XNOR U32204 ( .A(n31091), .B(n24838), .Z(n31093) );
  XOR U32205 ( .A(n31095), .B(n31096), .Z(n24838) );
  AND U32206 ( .A(\modmult_1/xin[1023] ), .B(n31097), .Z(n31096) );
  IV U32207 ( .A(n31095), .Z(n31097) );
  XOR U32208 ( .A(n31098), .B(mreg[984]), .Z(n31095) );
  NAND U32209 ( .A(n31099), .B(mul_pow), .Z(n31098) );
  XOR U32210 ( .A(mreg[984]), .B(creg[984]), .Z(n31099) );
  XOR U32211 ( .A(n31100), .B(n31101), .Z(n31091) );
  ANDN U32212 ( .A(n31102), .B(n24845), .Z(n31101) );
  XOR U32213 ( .A(n31103), .B(\modmult_1/zin[0][982] ), .Z(n24845) );
  IV U32214 ( .A(n31100), .Z(n31103) );
  XNOR U32215 ( .A(n31100), .B(n24844), .Z(n31102) );
  XOR U32216 ( .A(n31104), .B(n31105), .Z(n24844) );
  AND U32217 ( .A(\modmult_1/xin[1023] ), .B(n31106), .Z(n31105) );
  IV U32218 ( .A(n31104), .Z(n31106) );
  XOR U32219 ( .A(n31107), .B(mreg[983]), .Z(n31104) );
  NAND U32220 ( .A(n31108), .B(mul_pow), .Z(n31107) );
  XOR U32221 ( .A(mreg[983]), .B(creg[983]), .Z(n31108) );
  XOR U32222 ( .A(n31109), .B(n31110), .Z(n31100) );
  ANDN U32223 ( .A(n31111), .B(n24851), .Z(n31110) );
  XOR U32224 ( .A(n31112), .B(\modmult_1/zin[0][981] ), .Z(n24851) );
  IV U32225 ( .A(n31109), .Z(n31112) );
  XNOR U32226 ( .A(n31109), .B(n24850), .Z(n31111) );
  XOR U32227 ( .A(n31113), .B(n31114), .Z(n24850) );
  AND U32228 ( .A(\modmult_1/xin[1023] ), .B(n31115), .Z(n31114) );
  IV U32229 ( .A(n31113), .Z(n31115) );
  XOR U32230 ( .A(n31116), .B(mreg[982]), .Z(n31113) );
  NAND U32231 ( .A(n31117), .B(mul_pow), .Z(n31116) );
  XOR U32232 ( .A(mreg[982]), .B(creg[982]), .Z(n31117) );
  XOR U32233 ( .A(n31118), .B(n31119), .Z(n31109) );
  ANDN U32234 ( .A(n31120), .B(n24857), .Z(n31119) );
  XOR U32235 ( .A(n31121), .B(\modmult_1/zin[0][980] ), .Z(n24857) );
  IV U32236 ( .A(n31118), .Z(n31121) );
  XNOR U32237 ( .A(n31118), .B(n24856), .Z(n31120) );
  XOR U32238 ( .A(n31122), .B(n31123), .Z(n24856) );
  AND U32239 ( .A(\modmult_1/xin[1023] ), .B(n31124), .Z(n31123) );
  IV U32240 ( .A(n31122), .Z(n31124) );
  XOR U32241 ( .A(n31125), .B(mreg[981]), .Z(n31122) );
  NAND U32242 ( .A(n31126), .B(mul_pow), .Z(n31125) );
  XOR U32243 ( .A(mreg[981]), .B(creg[981]), .Z(n31126) );
  XOR U32244 ( .A(n31127), .B(n31128), .Z(n31118) );
  ANDN U32245 ( .A(n31129), .B(n24863), .Z(n31128) );
  XOR U32246 ( .A(n31130), .B(\modmult_1/zin[0][979] ), .Z(n24863) );
  IV U32247 ( .A(n31127), .Z(n31130) );
  XNOR U32248 ( .A(n31127), .B(n24862), .Z(n31129) );
  XOR U32249 ( .A(n31131), .B(n31132), .Z(n24862) );
  AND U32250 ( .A(\modmult_1/xin[1023] ), .B(n31133), .Z(n31132) );
  IV U32251 ( .A(n31131), .Z(n31133) );
  XOR U32252 ( .A(n31134), .B(mreg[980]), .Z(n31131) );
  NAND U32253 ( .A(n31135), .B(mul_pow), .Z(n31134) );
  XOR U32254 ( .A(mreg[980]), .B(creg[980]), .Z(n31135) );
  XOR U32255 ( .A(n31136), .B(n31137), .Z(n31127) );
  ANDN U32256 ( .A(n31138), .B(n24869), .Z(n31137) );
  XOR U32257 ( .A(n31139), .B(\modmult_1/zin[0][978] ), .Z(n24869) );
  IV U32258 ( .A(n31136), .Z(n31139) );
  XNOR U32259 ( .A(n31136), .B(n24868), .Z(n31138) );
  XOR U32260 ( .A(n31140), .B(n31141), .Z(n24868) );
  AND U32261 ( .A(\modmult_1/xin[1023] ), .B(n31142), .Z(n31141) );
  IV U32262 ( .A(n31140), .Z(n31142) );
  XOR U32263 ( .A(n31143), .B(mreg[979]), .Z(n31140) );
  NAND U32264 ( .A(n31144), .B(mul_pow), .Z(n31143) );
  XOR U32265 ( .A(mreg[979]), .B(creg[979]), .Z(n31144) );
  XOR U32266 ( .A(n31145), .B(n31146), .Z(n31136) );
  ANDN U32267 ( .A(n31147), .B(n24875), .Z(n31146) );
  XOR U32268 ( .A(n31148), .B(\modmult_1/zin[0][977] ), .Z(n24875) );
  IV U32269 ( .A(n31145), .Z(n31148) );
  XNOR U32270 ( .A(n31145), .B(n24874), .Z(n31147) );
  XOR U32271 ( .A(n31149), .B(n31150), .Z(n24874) );
  AND U32272 ( .A(\modmult_1/xin[1023] ), .B(n31151), .Z(n31150) );
  IV U32273 ( .A(n31149), .Z(n31151) );
  XOR U32274 ( .A(n31152), .B(mreg[978]), .Z(n31149) );
  NAND U32275 ( .A(n31153), .B(mul_pow), .Z(n31152) );
  XOR U32276 ( .A(mreg[978]), .B(creg[978]), .Z(n31153) );
  XOR U32277 ( .A(n31154), .B(n31155), .Z(n31145) );
  ANDN U32278 ( .A(n31156), .B(n24881), .Z(n31155) );
  XOR U32279 ( .A(n31157), .B(\modmult_1/zin[0][976] ), .Z(n24881) );
  IV U32280 ( .A(n31154), .Z(n31157) );
  XNOR U32281 ( .A(n31154), .B(n24880), .Z(n31156) );
  XOR U32282 ( .A(n31158), .B(n31159), .Z(n24880) );
  AND U32283 ( .A(\modmult_1/xin[1023] ), .B(n31160), .Z(n31159) );
  IV U32284 ( .A(n31158), .Z(n31160) );
  XOR U32285 ( .A(n31161), .B(mreg[977]), .Z(n31158) );
  NAND U32286 ( .A(n31162), .B(mul_pow), .Z(n31161) );
  XOR U32287 ( .A(mreg[977]), .B(creg[977]), .Z(n31162) );
  XOR U32288 ( .A(n31163), .B(n31164), .Z(n31154) );
  ANDN U32289 ( .A(n31165), .B(n24887), .Z(n31164) );
  XOR U32290 ( .A(n31166), .B(\modmult_1/zin[0][975] ), .Z(n24887) );
  IV U32291 ( .A(n31163), .Z(n31166) );
  XNOR U32292 ( .A(n31163), .B(n24886), .Z(n31165) );
  XOR U32293 ( .A(n31167), .B(n31168), .Z(n24886) );
  AND U32294 ( .A(\modmult_1/xin[1023] ), .B(n31169), .Z(n31168) );
  IV U32295 ( .A(n31167), .Z(n31169) );
  XOR U32296 ( .A(n31170), .B(mreg[976]), .Z(n31167) );
  NAND U32297 ( .A(n31171), .B(mul_pow), .Z(n31170) );
  XOR U32298 ( .A(mreg[976]), .B(creg[976]), .Z(n31171) );
  XOR U32299 ( .A(n31172), .B(n31173), .Z(n31163) );
  ANDN U32300 ( .A(n31174), .B(n24893), .Z(n31173) );
  XOR U32301 ( .A(n31175), .B(\modmult_1/zin[0][974] ), .Z(n24893) );
  IV U32302 ( .A(n31172), .Z(n31175) );
  XNOR U32303 ( .A(n31172), .B(n24892), .Z(n31174) );
  XOR U32304 ( .A(n31176), .B(n31177), .Z(n24892) );
  AND U32305 ( .A(\modmult_1/xin[1023] ), .B(n31178), .Z(n31177) );
  IV U32306 ( .A(n31176), .Z(n31178) );
  XOR U32307 ( .A(n31179), .B(mreg[975]), .Z(n31176) );
  NAND U32308 ( .A(n31180), .B(mul_pow), .Z(n31179) );
  XOR U32309 ( .A(mreg[975]), .B(creg[975]), .Z(n31180) );
  XOR U32310 ( .A(n31181), .B(n31182), .Z(n31172) );
  ANDN U32311 ( .A(n31183), .B(n24899), .Z(n31182) );
  XOR U32312 ( .A(n31184), .B(\modmult_1/zin[0][973] ), .Z(n24899) );
  IV U32313 ( .A(n31181), .Z(n31184) );
  XNOR U32314 ( .A(n31181), .B(n24898), .Z(n31183) );
  XOR U32315 ( .A(n31185), .B(n31186), .Z(n24898) );
  AND U32316 ( .A(\modmult_1/xin[1023] ), .B(n31187), .Z(n31186) );
  IV U32317 ( .A(n31185), .Z(n31187) );
  XOR U32318 ( .A(n31188), .B(mreg[974]), .Z(n31185) );
  NAND U32319 ( .A(n31189), .B(mul_pow), .Z(n31188) );
  XOR U32320 ( .A(mreg[974]), .B(creg[974]), .Z(n31189) );
  XOR U32321 ( .A(n31190), .B(n31191), .Z(n31181) );
  ANDN U32322 ( .A(n31192), .B(n24905), .Z(n31191) );
  XOR U32323 ( .A(n31193), .B(\modmult_1/zin[0][972] ), .Z(n24905) );
  IV U32324 ( .A(n31190), .Z(n31193) );
  XNOR U32325 ( .A(n31190), .B(n24904), .Z(n31192) );
  XOR U32326 ( .A(n31194), .B(n31195), .Z(n24904) );
  AND U32327 ( .A(\modmult_1/xin[1023] ), .B(n31196), .Z(n31195) );
  IV U32328 ( .A(n31194), .Z(n31196) );
  XOR U32329 ( .A(n31197), .B(mreg[973]), .Z(n31194) );
  NAND U32330 ( .A(n31198), .B(mul_pow), .Z(n31197) );
  XOR U32331 ( .A(mreg[973]), .B(creg[973]), .Z(n31198) );
  XOR U32332 ( .A(n31199), .B(n31200), .Z(n31190) );
  ANDN U32333 ( .A(n31201), .B(n24911), .Z(n31200) );
  XOR U32334 ( .A(n31202), .B(\modmult_1/zin[0][971] ), .Z(n24911) );
  IV U32335 ( .A(n31199), .Z(n31202) );
  XNOR U32336 ( .A(n31199), .B(n24910), .Z(n31201) );
  XOR U32337 ( .A(n31203), .B(n31204), .Z(n24910) );
  AND U32338 ( .A(\modmult_1/xin[1023] ), .B(n31205), .Z(n31204) );
  IV U32339 ( .A(n31203), .Z(n31205) );
  XOR U32340 ( .A(n31206), .B(mreg[972]), .Z(n31203) );
  NAND U32341 ( .A(n31207), .B(mul_pow), .Z(n31206) );
  XOR U32342 ( .A(mreg[972]), .B(creg[972]), .Z(n31207) );
  XOR U32343 ( .A(n31208), .B(n31209), .Z(n31199) );
  ANDN U32344 ( .A(n31210), .B(n24917), .Z(n31209) );
  XOR U32345 ( .A(n31211), .B(\modmult_1/zin[0][970] ), .Z(n24917) );
  IV U32346 ( .A(n31208), .Z(n31211) );
  XNOR U32347 ( .A(n31208), .B(n24916), .Z(n31210) );
  XOR U32348 ( .A(n31212), .B(n31213), .Z(n24916) );
  AND U32349 ( .A(\modmult_1/xin[1023] ), .B(n31214), .Z(n31213) );
  IV U32350 ( .A(n31212), .Z(n31214) );
  XOR U32351 ( .A(n31215), .B(mreg[971]), .Z(n31212) );
  NAND U32352 ( .A(n31216), .B(mul_pow), .Z(n31215) );
  XOR U32353 ( .A(mreg[971]), .B(creg[971]), .Z(n31216) );
  XOR U32354 ( .A(n31217), .B(n31218), .Z(n31208) );
  ANDN U32355 ( .A(n31219), .B(n24923), .Z(n31218) );
  XOR U32356 ( .A(n31220), .B(\modmult_1/zin[0][969] ), .Z(n24923) );
  IV U32357 ( .A(n31217), .Z(n31220) );
  XNOR U32358 ( .A(n31217), .B(n24922), .Z(n31219) );
  XOR U32359 ( .A(n31221), .B(n31222), .Z(n24922) );
  AND U32360 ( .A(\modmult_1/xin[1023] ), .B(n31223), .Z(n31222) );
  IV U32361 ( .A(n31221), .Z(n31223) );
  XOR U32362 ( .A(n31224), .B(mreg[970]), .Z(n31221) );
  NAND U32363 ( .A(n31225), .B(mul_pow), .Z(n31224) );
  XOR U32364 ( .A(mreg[970]), .B(creg[970]), .Z(n31225) );
  XOR U32365 ( .A(n31226), .B(n31227), .Z(n31217) );
  ANDN U32366 ( .A(n31228), .B(n24929), .Z(n31227) );
  XOR U32367 ( .A(n31229), .B(\modmult_1/zin[0][968] ), .Z(n24929) );
  IV U32368 ( .A(n31226), .Z(n31229) );
  XNOR U32369 ( .A(n31226), .B(n24928), .Z(n31228) );
  XOR U32370 ( .A(n31230), .B(n31231), .Z(n24928) );
  AND U32371 ( .A(\modmult_1/xin[1023] ), .B(n31232), .Z(n31231) );
  IV U32372 ( .A(n31230), .Z(n31232) );
  XOR U32373 ( .A(n31233), .B(mreg[969]), .Z(n31230) );
  NAND U32374 ( .A(n31234), .B(mul_pow), .Z(n31233) );
  XOR U32375 ( .A(mreg[969]), .B(creg[969]), .Z(n31234) );
  XOR U32376 ( .A(n31235), .B(n31236), .Z(n31226) );
  ANDN U32377 ( .A(n31237), .B(n24935), .Z(n31236) );
  XOR U32378 ( .A(n31238), .B(\modmult_1/zin[0][967] ), .Z(n24935) );
  IV U32379 ( .A(n31235), .Z(n31238) );
  XNOR U32380 ( .A(n31235), .B(n24934), .Z(n31237) );
  XOR U32381 ( .A(n31239), .B(n31240), .Z(n24934) );
  AND U32382 ( .A(\modmult_1/xin[1023] ), .B(n31241), .Z(n31240) );
  IV U32383 ( .A(n31239), .Z(n31241) );
  XOR U32384 ( .A(n31242), .B(mreg[968]), .Z(n31239) );
  NAND U32385 ( .A(n31243), .B(mul_pow), .Z(n31242) );
  XOR U32386 ( .A(mreg[968]), .B(creg[968]), .Z(n31243) );
  XOR U32387 ( .A(n31244), .B(n31245), .Z(n31235) );
  ANDN U32388 ( .A(n31246), .B(n24941), .Z(n31245) );
  XOR U32389 ( .A(n31247), .B(\modmult_1/zin[0][966] ), .Z(n24941) );
  IV U32390 ( .A(n31244), .Z(n31247) );
  XNOR U32391 ( .A(n31244), .B(n24940), .Z(n31246) );
  XOR U32392 ( .A(n31248), .B(n31249), .Z(n24940) );
  AND U32393 ( .A(\modmult_1/xin[1023] ), .B(n31250), .Z(n31249) );
  IV U32394 ( .A(n31248), .Z(n31250) );
  XOR U32395 ( .A(n31251), .B(mreg[967]), .Z(n31248) );
  NAND U32396 ( .A(n31252), .B(mul_pow), .Z(n31251) );
  XOR U32397 ( .A(mreg[967]), .B(creg[967]), .Z(n31252) );
  XOR U32398 ( .A(n31253), .B(n31254), .Z(n31244) );
  ANDN U32399 ( .A(n31255), .B(n24947), .Z(n31254) );
  XOR U32400 ( .A(n31256), .B(\modmult_1/zin[0][965] ), .Z(n24947) );
  IV U32401 ( .A(n31253), .Z(n31256) );
  XNOR U32402 ( .A(n31253), .B(n24946), .Z(n31255) );
  XOR U32403 ( .A(n31257), .B(n31258), .Z(n24946) );
  AND U32404 ( .A(\modmult_1/xin[1023] ), .B(n31259), .Z(n31258) );
  IV U32405 ( .A(n31257), .Z(n31259) );
  XOR U32406 ( .A(n31260), .B(mreg[966]), .Z(n31257) );
  NAND U32407 ( .A(n31261), .B(mul_pow), .Z(n31260) );
  XOR U32408 ( .A(mreg[966]), .B(creg[966]), .Z(n31261) );
  XOR U32409 ( .A(n31262), .B(n31263), .Z(n31253) );
  ANDN U32410 ( .A(n31264), .B(n24953), .Z(n31263) );
  XOR U32411 ( .A(n31265), .B(\modmult_1/zin[0][964] ), .Z(n24953) );
  IV U32412 ( .A(n31262), .Z(n31265) );
  XNOR U32413 ( .A(n31262), .B(n24952), .Z(n31264) );
  XOR U32414 ( .A(n31266), .B(n31267), .Z(n24952) );
  AND U32415 ( .A(\modmult_1/xin[1023] ), .B(n31268), .Z(n31267) );
  IV U32416 ( .A(n31266), .Z(n31268) );
  XOR U32417 ( .A(n31269), .B(mreg[965]), .Z(n31266) );
  NAND U32418 ( .A(n31270), .B(mul_pow), .Z(n31269) );
  XOR U32419 ( .A(mreg[965]), .B(creg[965]), .Z(n31270) );
  XOR U32420 ( .A(n31271), .B(n31272), .Z(n31262) );
  ANDN U32421 ( .A(n31273), .B(n24959), .Z(n31272) );
  XOR U32422 ( .A(n31274), .B(\modmult_1/zin[0][963] ), .Z(n24959) );
  IV U32423 ( .A(n31271), .Z(n31274) );
  XNOR U32424 ( .A(n31271), .B(n24958), .Z(n31273) );
  XOR U32425 ( .A(n31275), .B(n31276), .Z(n24958) );
  AND U32426 ( .A(\modmult_1/xin[1023] ), .B(n31277), .Z(n31276) );
  IV U32427 ( .A(n31275), .Z(n31277) );
  XOR U32428 ( .A(n31278), .B(mreg[964]), .Z(n31275) );
  NAND U32429 ( .A(n31279), .B(mul_pow), .Z(n31278) );
  XOR U32430 ( .A(mreg[964]), .B(creg[964]), .Z(n31279) );
  XOR U32431 ( .A(n31280), .B(n31281), .Z(n31271) );
  ANDN U32432 ( .A(n31282), .B(n24965), .Z(n31281) );
  XOR U32433 ( .A(n31283), .B(\modmult_1/zin[0][962] ), .Z(n24965) );
  IV U32434 ( .A(n31280), .Z(n31283) );
  XNOR U32435 ( .A(n31280), .B(n24964), .Z(n31282) );
  XOR U32436 ( .A(n31284), .B(n31285), .Z(n24964) );
  AND U32437 ( .A(\modmult_1/xin[1023] ), .B(n31286), .Z(n31285) );
  IV U32438 ( .A(n31284), .Z(n31286) );
  XOR U32439 ( .A(n31287), .B(mreg[963]), .Z(n31284) );
  NAND U32440 ( .A(n31288), .B(mul_pow), .Z(n31287) );
  XOR U32441 ( .A(mreg[963]), .B(creg[963]), .Z(n31288) );
  XOR U32442 ( .A(n31289), .B(n31290), .Z(n31280) );
  ANDN U32443 ( .A(n31291), .B(n24971), .Z(n31290) );
  XOR U32444 ( .A(n31292), .B(\modmult_1/zin[0][961] ), .Z(n24971) );
  IV U32445 ( .A(n31289), .Z(n31292) );
  XNOR U32446 ( .A(n31289), .B(n24970), .Z(n31291) );
  XOR U32447 ( .A(n31293), .B(n31294), .Z(n24970) );
  AND U32448 ( .A(\modmult_1/xin[1023] ), .B(n31295), .Z(n31294) );
  IV U32449 ( .A(n31293), .Z(n31295) );
  XOR U32450 ( .A(n31296), .B(mreg[962]), .Z(n31293) );
  NAND U32451 ( .A(n31297), .B(mul_pow), .Z(n31296) );
  XOR U32452 ( .A(mreg[962]), .B(creg[962]), .Z(n31297) );
  XOR U32453 ( .A(n31298), .B(n31299), .Z(n31289) );
  ANDN U32454 ( .A(n31300), .B(n24977), .Z(n31299) );
  XOR U32455 ( .A(n31301), .B(\modmult_1/zin[0][960] ), .Z(n24977) );
  IV U32456 ( .A(n31298), .Z(n31301) );
  XNOR U32457 ( .A(n31298), .B(n24976), .Z(n31300) );
  XOR U32458 ( .A(n31302), .B(n31303), .Z(n24976) );
  AND U32459 ( .A(\modmult_1/xin[1023] ), .B(n31304), .Z(n31303) );
  IV U32460 ( .A(n31302), .Z(n31304) );
  XOR U32461 ( .A(n31305), .B(mreg[961]), .Z(n31302) );
  NAND U32462 ( .A(n31306), .B(mul_pow), .Z(n31305) );
  XOR U32463 ( .A(mreg[961]), .B(creg[961]), .Z(n31306) );
  XOR U32464 ( .A(n31307), .B(n31308), .Z(n31298) );
  ANDN U32465 ( .A(n31309), .B(n24983), .Z(n31308) );
  XOR U32466 ( .A(n31310), .B(\modmult_1/zin[0][959] ), .Z(n24983) );
  IV U32467 ( .A(n31307), .Z(n31310) );
  XNOR U32468 ( .A(n31307), .B(n24982), .Z(n31309) );
  XOR U32469 ( .A(n31311), .B(n31312), .Z(n24982) );
  AND U32470 ( .A(\modmult_1/xin[1023] ), .B(n31313), .Z(n31312) );
  IV U32471 ( .A(n31311), .Z(n31313) );
  XOR U32472 ( .A(n31314), .B(mreg[960]), .Z(n31311) );
  NAND U32473 ( .A(n31315), .B(mul_pow), .Z(n31314) );
  XOR U32474 ( .A(mreg[960]), .B(creg[960]), .Z(n31315) );
  XOR U32475 ( .A(n31316), .B(n31317), .Z(n31307) );
  ANDN U32476 ( .A(n31318), .B(n24989), .Z(n31317) );
  XOR U32477 ( .A(n31319), .B(\modmult_1/zin[0][958] ), .Z(n24989) );
  IV U32478 ( .A(n31316), .Z(n31319) );
  XNOR U32479 ( .A(n31316), .B(n24988), .Z(n31318) );
  XOR U32480 ( .A(n31320), .B(n31321), .Z(n24988) );
  AND U32481 ( .A(\modmult_1/xin[1023] ), .B(n31322), .Z(n31321) );
  IV U32482 ( .A(n31320), .Z(n31322) );
  XOR U32483 ( .A(n31323), .B(mreg[959]), .Z(n31320) );
  NAND U32484 ( .A(n31324), .B(mul_pow), .Z(n31323) );
  XOR U32485 ( .A(mreg[959]), .B(creg[959]), .Z(n31324) );
  XOR U32486 ( .A(n31325), .B(n31326), .Z(n31316) );
  ANDN U32487 ( .A(n31327), .B(n24995), .Z(n31326) );
  XOR U32488 ( .A(n31328), .B(\modmult_1/zin[0][957] ), .Z(n24995) );
  IV U32489 ( .A(n31325), .Z(n31328) );
  XNOR U32490 ( .A(n31325), .B(n24994), .Z(n31327) );
  XOR U32491 ( .A(n31329), .B(n31330), .Z(n24994) );
  AND U32492 ( .A(\modmult_1/xin[1023] ), .B(n31331), .Z(n31330) );
  IV U32493 ( .A(n31329), .Z(n31331) );
  XOR U32494 ( .A(n31332), .B(mreg[958]), .Z(n31329) );
  NAND U32495 ( .A(n31333), .B(mul_pow), .Z(n31332) );
  XOR U32496 ( .A(mreg[958]), .B(creg[958]), .Z(n31333) );
  XOR U32497 ( .A(n31334), .B(n31335), .Z(n31325) );
  ANDN U32498 ( .A(n31336), .B(n25001), .Z(n31335) );
  XOR U32499 ( .A(n31337), .B(\modmult_1/zin[0][956] ), .Z(n25001) );
  IV U32500 ( .A(n31334), .Z(n31337) );
  XNOR U32501 ( .A(n31334), .B(n25000), .Z(n31336) );
  XOR U32502 ( .A(n31338), .B(n31339), .Z(n25000) );
  AND U32503 ( .A(\modmult_1/xin[1023] ), .B(n31340), .Z(n31339) );
  IV U32504 ( .A(n31338), .Z(n31340) );
  XOR U32505 ( .A(n31341), .B(mreg[957]), .Z(n31338) );
  NAND U32506 ( .A(n31342), .B(mul_pow), .Z(n31341) );
  XOR U32507 ( .A(mreg[957]), .B(creg[957]), .Z(n31342) );
  XOR U32508 ( .A(n31343), .B(n31344), .Z(n31334) );
  ANDN U32509 ( .A(n31345), .B(n25007), .Z(n31344) );
  XOR U32510 ( .A(n31346), .B(\modmult_1/zin[0][955] ), .Z(n25007) );
  IV U32511 ( .A(n31343), .Z(n31346) );
  XNOR U32512 ( .A(n31343), .B(n25006), .Z(n31345) );
  XOR U32513 ( .A(n31347), .B(n31348), .Z(n25006) );
  AND U32514 ( .A(\modmult_1/xin[1023] ), .B(n31349), .Z(n31348) );
  IV U32515 ( .A(n31347), .Z(n31349) );
  XOR U32516 ( .A(n31350), .B(mreg[956]), .Z(n31347) );
  NAND U32517 ( .A(n31351), .B(mul_pow), .Z(n31350) );
  XOR U32518 ( .A(mreg[956]), .B(creg[956]), .Z(n31351) );
  XOR U32519 ( .A(n31352), .B(n31353), .Z(n31343) );
  ANDN U32520 ( .A(n31354), .B(n25013), .Z(n31353) );
  XOR U32521 ( .A(n31355), .B(\modmult_1/zin[0][954] ), .Z(n25013) );
  IV U32522 ( .A(n31352), .Z(n31355) );
  XNOR U32523 ( .A(n31352), .B(n25012), .Z(n31354) );
  XOR U32524 ( .A(n31356), .B(n31357), .Z(n25012) );
  AND U32525 ( .A(\modmult_1/xin[1023] ), .B(n31358), .Z(n31357) );
  IV U32526 ( .A(n31356), .Z(n31358) );
  XOR U32527 ( .A(n31359), .B(mreg[955]), .Z(n31356) );
  NAND U32528 ( .A(n31360), .B(mul_pow), .Z(n31359) );
  XOR U32529 ( .A(mreg[955]), .B(creg[955]), .Z(n31360) );
  XOR U32530 ( .A(n31361), .B(n31362), .Z(n31352) );
  ANDN U32531 ( .A(n31363), .B(n25019), .Z(n31362) );
  XOR U32532 ( .A(n31364), .B(\modmult_1/zin[0][953] ), .Z(n25019) );
  IV U32533 ( .A(n31361), .Z(n31364) );
  XNOR U32534 ( .A(n31361), .B(n25018), .Z(n31363) );
  XOR U32535 ( .A(n31365), .B(n31366), .Z(n25018) );
  AND U32536 ( .A(\modmult_1/xin[1023] ), .B(n31367), .Z(n31366) );
  IV U32537 ( .A(n31365), .Z(n31367) );
  XOR U32538 ( .A(n31368), .B(mreg[954]), .Z(n31365) );
  NAND U32539 ( .A(n31369), .B(mul_pow), .Z(n31368) );
  XOR U32540 ( .A(mreg[954]), .B(creg[954]), .Z(n31369) );
  XOR U32541 ( .A(n31370), .B(n31371), .Z(n31361) );
  ANDN U32542 ( .A(n31372), .B(n25025), .Z(n31371) );
  XOR U32543 ( .A(n31373), .B(\modmult_1/zin[0][952] ), .Z(n25025) );
  IV U32544 ( .A(n31370), .Z(n31373) );
  XNOR U32545 ( .A(n31370), .B(n25024), .Z(n31372) );
  XOR U32546 ( .A(n31374), .B(n31375), .Z(n25024) );
  AND U32547 ( .A(\modmult_1/xin[1023] ), .B(n31376), .Z(n31375) );
  IV U32548 ( .A(n31374), .Z(n31376) );
  XOR U32549 ( .A(n31377), .B(mreg[953]), .Z(n31374) );
  NAND U32550 ( .A(n31378), .B(mul_pow), .Z(n31377) );
  XOR U32551 ( .A(mreg[953]), .B(creg[953]), .Z(n31378) );
  XOR U32552 ( .A(n31379), .B(n31380), .Z(n31370) );
  ANDN U32553 ( .A(n31381), .B(n25031), .Z(n31380) );
  XOR U32554 ( .A(n31382), .B(\modmult_1/zin[0][951] ), .Z(n25031) );
  IV U32555 ( .A(n31379), .Z(n31382) );
  XNOR U32556 ( .A(n31379), .B(n25030), .Z(n31381) );
  XOR U32557 ( .A(n31383), .B(n31384), .Z(n25030) );
  AND U32558 ( .A(\modmult_1/xin[1023] ), .B(n31385), .Z(n31384) );
  IV U32559 ( .A(n31383), .Z(n31385) );
  XOR U32560 ( .A(n31386), .B(mreg[952]), .Z(n31383) );
  NAND U32561 ( .A(n31387), .B(mul_pow), .Z(n31386) );
  XOR U32562 ( .A(mreg[952]), .B(creg[952]), .Z(n31387) );
  XOR U32563 ( .A(n31388), .B(n31389), .Z(n31379) );
  ANDN U32564 ( .A(n31390), .B(n25037), .Z(n31389) );
  XOR U32565 ( .A(n31391), .B(\modmult_1/zin[0][950] ), .Z(n25037) );
  IV U32566 ( .A(n31388), .Z(n31391) );
  XNOR U32567 ( .A(n31388), .B(n25036), .Z(n31390) );
  XOR U32568 ( .A(n31392), .B(n31393), .Z(n25036) );
  AND U32569 ( .A(\modmult_1/xin[1023] ), .B(n31394), .Z(n31393) );
  IV U32570 ( .A(n31392), .Z(n31394) );
  XOR U32571 ( .A(n31395), .B(mreg[951]), .Z(n31392) );
  NAND U32572 ( .A(n31396), .B(mul_pow), .Z(n31395) );
  XOR U32573 ( .A(mreg[951]), .B(creg[951]), .Z(n31396) );
  XOR U32574 ( .A(n31397), .B(n31398), .Z(n31388) );
  ANDN U32575 ( .A(n31399), .B(n25043), .Z(n31398) );
  XOR U32576 ( .A(n31400), .B(\modmult_1/zin[0][949] ), .Z(n25043) );
  IV U32577 ( .A(n31397), .Z(n31400) );
  XNOR U32578 ( .A(n31397), .B(n25042), .Z(n31399) );
  XOR U32579 ( .A(n31401), .B(n31402), .Z(n25042) );
  AND U32580 ( .A(\modmult_1/xin[1023] ), .B(n31403), .Z(n31402) );
  IV U32581 ( .A(n31401), .Z(n31403) );
  XOR U32582 ( .A(n31404), .B(mreg[950]), .Z(n31401) );
  NAND U32583 ( .A(n31405), .B(mul_pow), .Z(n31404) );
  XOR U32584 ( .A(mreg[950]), .B(creg[950]), .Z(n31405) );
  XOR U32585 ( .A(n31406), .B(n31407), .Z(n31397) );
  ANDN U32586 ( .A(n31408), .B(n25049), .Z(n31407) );
  XOR U32587 ( .A(n31409), .B(\modmult_1/zin[0][948] ), .Z(n25049) );
  IV U32588 ( .A(n31406), .Z(n31409) );
  XNOR U32589 ( .A(n31406), .B(n25048), .Z(n31408) );
  XOR U32590 ( .A(n31410), .B(n31411), .Z(n25048) );
  AND U32591 ( .A(\modmult_1/xin[1023] ), .B(n31412), .Z(n31411) );
  IV U32592 ( .A(n31410), .Z(n31412) );
  XOR U32593 ( .A(n31413), .B(mreg[949]), .Z(n31410) );
  NAND U32594 ( .A(n31414), .B(mul_pow), .Z(n31413) );
  XOR U32595 ( .A(mreg[949]), .B(creg[949]), .Z(n31414) );
  XOR U32596 ( .A(n31415), .B(n31416), .Z(n31406) );
  ANDN U32597 ( .A(n31417), .B(n25055), .Z(n31416) );
  XOR U32598 ( .A(n31418), .B(\modmult_1/zin[0][947] ), .Z(n25055) );
  IV U32599 ( .A(n31415), .Z(n31418) );
  XNOR U32600 ( .A(n31415), .B(n25054), .Z(n31417) );
  XOR U32601 ( .A(n31419), .B(n31420), .Z(n25054) );
  AND U32602 ( .A(\modmult_1/xin[1023] ), .B(n31421), .Z(n31420) );
  IV U32603 ( .A(n31419), .Z(n31421) );
  XOR U32604 ( .A(n31422), .B(mreg[948]), .Z(n31419) );
  NAND U32605 ( .A(n31423), .B(mul_pow), .Z(n31422) );
  XOR U32606 ( .A(mreg[948]), .B(creg[948]), .Z(n31423) );
  XOR U32607 ( .A(n31424), .B(n31425), .Z(n31415) );
  ANDN U32608 ( .A(n31426), .B(n25061), .Z(n31425) );
  XOR U32609 ( .A(n31427), .B(\modmult_1/zin[0][946] ), .Z(n25061) );
  IV U32610 ( .A(n31424), .Z(n31427) );
  XNOR U32611 ( .A(n31424), .B(n25060), .Z(n31426) );
  XOR U32612 ( .A(n31428), .B(n31429), .Z(n25060) );
  AND U32613 ( .A(\modmult_1/xin[1023] ), .B(n31430), .Z(n31429) );
  IV U32614 ( .A(n31428), .Z(n31430) );
  XOR U32615 ( .A(n31431), .B(mreg[947]), .Z(n31428) );
  NAND U32616 ( .A(n31432), .B(mul_pow), .Z(n31431) );
  XOR U32617 ( .A(mreg[947]), .B(creg[947]), .Z(n31432) );
  XOR U32618 ( .A(n31433), .B(n31434), .Z(n31424) );
  ANDN U32619 ( .A(n31435), .B(n25067), .Z(n31434) );
  XOR U32620 ( .A(n31436), .B(\modmult_1/zin[0][945] ), .Z(n25067) );
  IV U32621 ( .A(n31433), .Z(n31436) );
  XNOR U32622 ( .A(n31433), .B(n25066), .Z(n31435) );
  XOR U32623 ( .A(n31437), .B(n31438), .Z(n25066) );
  AND U32624 ( .A(\modmult_1/xin[1023] ), .B(n31439), .Z(n31438) );
  IV U32625 ( .A(n31437), .Z(n31439) );
  XOR U32626 ( .A(n31440), .B(mreg[946]), .Z(n31437) );
  NAND U32627 ( .A(n31441), .B(mul_pow), .Z(n31440) );
  XOR U32628 ( .A(mreg[946]), .B(creg[946]), .Z(n31441) );
  XOR U32629 ( .A(n31442), .B(n31443), .Z(n31433) );
  ANDN U32630 ( .A(n31444), .B(n25073), .Z(n31443) );
  XOR U32631 ( .A(n31445), .B(\modmult_1/zin[0][944] ), .Z(n25073) );
  IV U32632 ( .A(n31442), .Z(n31445) );
  XNOR U32633 ( .A(n31442), .B(n25072), .Z(n31444) );
  XOR U32634 ( .A(n31446), .B(n31447), .Z(n25072) );
  AND U32635 ( .A(\modmult_1/xin[1023] ), .B(n31448), .Z(n31447) );
  IV U32636 ( .A(n31446), .Z(n31448) );
  XOR U32637 ( .A(n31449), .B(mreg[945]), .Z(n31446) );
  NAND U32638 ( .A(n31450), .B(mul_pow), .Z(n31449) );
  XOR U32639 ( .A(mreg[945]), .B(creg[945]), .Z(n31450) );
  XOR U32640 ( .A(n31451), .B(n31452), .Z(n31442) );
  ANDN U32641 ( .A(n31453), .B(n25079), .Z(n31452) );
  XOR U32642 ( .A(n31454), .B(\modmult_1/zin[0][943] ), .Z(n25079) );
  IV U32643 ( .A(n31451), .Z(n31454) );
  XNOR U32644 ( .A(n31451), .B(n25078), .Z(n31453) );
  XOR U32645 ( .A(n31455), .B(n31456), .Z(n25078) );
  AND U32646 ( .A(\modmult_1/xin[1023] ), .B(n31457), .Z(n31456) );
  IV U32647 ( .A(n31455), .Z(n31457) );
  XOR U32648 ( .A(n31458), .B(mreg[944]), .Z(n31455) );
  NAND U32649 ( .A(n31459), .B(mul_pow), .Z(n31458) );
  XOR U32650 ( .A(mreg[944]), .B(creg[944]), .Z(n31459) );
  XOR U32651 ( .A(n31460), .B(n31461), .Z(n31451) );
  ANDN U32652 ( .A(n31462), .B(n25085), .Z(n31461) );
  XOR U32653 ( .A(n31463), .B(\modmult_1/zin[0][942] ), .Z(n25085) );
  IV U32654 ( .A(n31460), .Z(n31463) );
  XNOR U32655 ( .A(n31460), .B(n25084), .Z(n31462) );
  XOR U32656 ( .A(n31464), .B(n31465), .Z(n25084) );
  AND U32657 ( .A(\modmult_1/xin[1023] ), .B(n31466), .Z(n31465) );
  IV U32658 ( .A(n31464), .Z(n31466) );
  XOR U32659 ( .A(n31467), .B(mreg[943]), .Z(n31464) );
  NAND U32660 ( .A(n31468), .B(mul_pow), .Z(n31467) );
  XOR U32661 ( .A(mreg[943]), .B(creg[943]), .Z(n31468) );
  XOR U32662 ( .A(n31469), .B(n31470), .Z(n31460) );
  ANDN U32663 ( .A(n31471), .B(n25091), .Z(n31470) );
  XOR U32664 ( .A(n31472), .B(\modmult_1/zin[0][941] ), .Z(n25091) );
  IV U32665 ( .A(n31469), .Z(n31472) );
  XNOR U32666 ( .A(n31469), .B(n25090), .Z(n31471) );
  XOR U32667 ( .A(n31473), .B(n31474), .Z(n25090) );
  AND U32668 ( .A(\modmult_1/xin[1023] ), .B(n31475), .Z(n31474) );
  IV U32669 ( .A(n31473), .Z(n31475) );
  XOR U32670 ( .A(n31476), .B(mreg[942]), .Z(n31473) );
  NAND U32671 ( .A(n31477), .B(mul_pow), .Z(n31476) );
  XOR U32672 ( .A(mreg[942]), .B(creg[942]), .Z(n31477) );
  XOR U32673 ( .A(n31478), .B(n31479), .Z(n31469) );
  ANDN U32674 ( .A(n31480), .B(n25097), .Z(n31479) );
  XOR U32675 ( .A(n31481), .B(\modmult_1/zin[0][940] ), .Z(n25097) );
  IV U32676 ( .A(n31478), .Z(n31481) );
  XNOR U32677 ( .A(n31478), .B(n25096), .Z(n31480) );
  XOR U32678 ( .A(n31482), .B(n31483), .Z(n25096) );
  AND U32679 ( .A(\modmult_1/xin[1023] ), .B(n31484), .Z(n31483) );
  IV U32680 ( .A(n31482), .Z(n31484) );
  XOR U32681 ( .A(n31485), .B(mreg[941]), .Z(n31482) );
  NAND U32682 ( .A(n31486), .B(mul_pow), .Z(n31485) );
  XOR U32683 ( .A(mreg[941]), .B(creg[941]), .Z(n31486) );
  XOR U32684 ( .A(n31487), .B(n31488), .Z(n31478) );
  ANDN U32685 ( .A(n31489), .B(n25103), .Z(n31488) );
  XOR U32686 ( .A(n31490), .B(\modmult_1/zin[0][939] ), .Z(n25103) );
  IV U32687 ( .A(n31487), .Z(n31490) );
  XNOR U32688 ( .A(n31487), .B(n25102), .Z(n31489) );
  XOR U32689 ( .A(n31491), .B(n31492), .Z(n25102) );
  AND U32690 ( .A(\modmult_1/xin[1023] ), .B(n31493), .Z(n31492) );
  IV U32691 ( .A(n31491), .Z(n31493) );
  XOR U32692 ( .A(n31494), .B(mreg[940]), .Z(n31491) );
  NAND U32693 ( .A(n31495), .B(mul_pow), .Z(n31494) );
  XOR U32694 ( .A(mreg[940]), .B(creg[940]), .Z(n31495) );
  XOR U32695 ( .A(n31496), .B(n31497), .Z(n31487) );
  ANDN U32696 ( .A(n31498), .B(n25109), .Z(n31497) );
  XOR U32697 ( .A(n31499), .B(\modmult_1/zin[0][938] ), .Z(n25109) );
  IV U32698 ( .A(n31496), .Z(n31499) );
  XNOR U32699 ( .A(n31496), .B(n25108), .Z(n31498) );
  XOR U32700 ( .A(n31500), .B(n31501), .Z(n25108) );
  AND U32701 ( .A(\modmult_1/xin[1023] ), .B(n31502), .Z(n31501) );
  IV U32702 ( .A(n31500), .Z(n31502) );
  XOR U32703 ( .A(n31503), .B(mreg[939]), .Z(n31500) );
  NAND U32704 ( .A(n31504), .B(mul_pow), .Z(n31503) );
  XOR U32705 ( .A(mreg[939]), .B(creg[939]), .Z(n31504) );
  XOR U32706 ( .A(n31505), .B(n31506), .Z(n31496) );
  ANDN U32707 ( .A(n31507), .B(n25115), .Z(n31506) );
  XOR U32708 ( .A(n31508), .B(\modmult_1/zin[0][937] ), .Z(n25115) );
  IV U32709 ( .A(n31505), .Z(n31508) );
  XNOR U32710 ( .A(n31505), .B(n25114), .Z(n31507) );
  XOR U32711 ( .A(n31509), .B(n31510), .Z(n25114) );
  AND U32712 ( .A(\modmult_1/xin[1023] ), .B(n31511), .Z(n31510) );
  IV U32713 ( .A(n31509), .Z(n31511) );
  XOR U32714 ( .A(n31512), .B(mreg[938]), .Z(n31509) );
  NAND U32715 ( .A(n31513), .B(mul_pow), .Z(n31512) );
  XOR U32716 ( .A(mreg[938]), .B(creg[938]), .Z(n31513) );
  XOR U32717 ( .A(n31514), .B(n31515), .Z(n31505) );
  ANDN U32718 ( .A(n31516), .B(n25121), .Z(n31515) );
  XOR U32719 ( .A(n31517), .B(\modmult_1/zin[0][936] ), .Z(n25121) );
  IV U32720 ( .A(n31514), .Z(n31517) );
  XNOR U32721 ( .A(n31514), .B(n25120), .Z(n31516) );
  XOR U32722 ( .A(n31518), .B(n31519), .Z(n25120) );
  AND U32723 ( .A(\modmult_1/xin[1023] ), .B(n31520), .Z(n31519) );
  IV U32724 ( .A(n31518), .Z(n31520) );
  XOR U32725 ( .A(n31521), .B(mreg[937]), .Z(n31518) );
  NAND U32726 ( .A(n31522), .B(mul_pow), .Z(n31521) );
  XOR U32727 ( .A(mreg[937]), .B(creg[937]), .Z(n31522) );
  XOR U32728 ( .A(n31523), .B(n31524), .Z(n31514) );
  ANDN U32729 ( .A(n31525), .B(n25127), .Z(n31524) );
  XOR U32730 ( .A(n31526), .B(\modmult_1/zin[0][935] ), .Z(n25127) );
  IV U32731 ( .A(n31523), .Z(n31526) );
  XNOR U32732 ( .A(n31523), .B(n25126), .Z(n31525) );
  XOR U32733 ( .A(n31527), .B(n31528), .Z(n25126) );
  AND U32734 ( .A(\modmult_1/xin[1023] ), .B(n31529), .Z(n31528) );
  IV U32735 ( .A(n31527), .Z(n31529) );
  XOR U32736 ( .A(n31530), .B(mreg[936]), .Z(n31527) );
  NAND U32737 ( .A(n31531), .B(mul_pow), .Z(n31530) );
  XOR U32738 ( .A(mreg[936]), .B(creg[936]), .Z(n31531) );
  XOR U32739 ( .A(n31532), .B(n31533), .Z(n31523) );
  ANDN U32740 ( .A(n31534), .B(n25133), .Z(n31533) );
  XOR U32741 ( .A(n31535), .B(\modmult_1/zin[0][934] ), .Z(n25133) );
  IV U32742 ( .A(n31532), .Z(n31535) );
  XNOR U32743 ( .A(n31532), .B(n25132), .Z(n31534) );
  XOR U32744 ( .A(n31536), .B(n31537), .Z(n25132) );
  AND U32745 ( .A(\modmult_1/xin[1023] ), .B(n31538), .Z(n31537) );
  IV U32746 ( .A(n31536), .Z(n31538) );
  XOR U32747 ( .A(n31539), .B(mreg[935]), .Z(n31536) );
  NAND U32748 ( .A(n31540), .B(mul_pow), .Z(n31539) );
  XOR U32749 ( .A(mreg[935]), .B(creg[935]), .Z(n31540) );
  XOR U32750 ( .A(n31541), .B(n31542), .Z(n31532) );
  ANDN U32751 ( .A(n31543), .B(n25139), .Z(n31542) );
  XOR U32752 ( .A(n31544), .B(\modmult_1/zin[0][933] ), .Z(n25139) );
  IV U32753 ( .A(n31541), .Z(n31544) );
  XNOR U32754 ( .A(n31541), .B(n25138), .Z(n31543) );
  XOR U32755 ( .A(n31545), .B(n31546), .Z(n25138) );
  AND U32756 ( .A(\modmult_1/xin[1023] ), .B(n31547), .Z(n31546) );
  IV U32757 ( .A(n31545), .Z(n31547) );
  XOR U32758 ( .A(n31548), .B(mreg[934]), .Z(n31545) );
  NAND U32759 ( .A(n31549), .B(mul_pow), .Z(n31548) );
  XOR U32760 ( .A(mreg[934]), .B(creg[934]), .Z(n31549) );
  XOR U32761 ( .A(n31550), .B(n31551), .Z(n31541) );
  ANDN U32762 ( .A(n31552), .B(n25145), .Z(n31551) );
  XOR U32763 ( .A(n31553), .B(\modmult_1/zin[0][932] ), .Z(n25145) );
  IV U32764 ( .A(n31550), .Z(n31553) );
  XNOR U32765 ( .A(n31550), .B(n25144), .Z(n31552) );
  XOR U32766 ( .A(n31554), .B(n31555), .Z(n25144) );
  AND U32767 ( .A(\modmult_1/xin[1023] ), .B(n31556), .Z(n31555) );
  IV U32768 ( .A(n31554), .Z(n31556) );
  XOR U32769 ( .A(n31557), .B(mreg[933]), .Z(n31554) );
  NAND U32770 ( .A(n31558), .B(mul_pow), .Z(n31557) );
  XOR U32771 ( .A(mreg[933]), .B(creg[933]), .Z(n31558) );
  XOR U32772 ( .A(n31559), .B(n31560), .Z(n31550) );
  ANDN U32773 ( .A(n31561), .B(n25151), .Z(n31560) );
  XOR U32774 ( .A(n31562), .B(\modmult_1/zin[0][931] ), .Z(n25151) );
  IV U32775 ( .A(n31559), .Z(n31562) );
  XNOR U32776 ( .A(n31559), .B(n25150), .Z(n31561) );
  XOR U32777 ( .A(n31563), .B(n31564), .Z(n25150) );
  AND U32778 ( .A(\modmult_1/xin[1023] ), .B(n31565), .Z(n31564) );
  IV U32779 ( .A(n31563), .Z(n31565) );
  XOR U32780 ( .A(n31566), .B(mreg[932]), .Z(n31563) );
  NAND U32781 ( .A(n31567), .B(mul_pow), .Z(n31566) );
  XOR U32782 ( .A(mreg[932]), .B(creg[932]), .Z(n31567) );
  XOR U32783 ( .A(n31568), .B(n31569), .Z(n31559) );
  ANDN U32784 ( .A(n31570), .B(n25157), .Z(n31569) );
  XOR U32785 ( .A(n31571), .B(\modmult_1/zin[0][930] ), .Z(n25157) );
  IV U32786 ( .A(n31568), .Z(n31571) );
  XNOR U32787 ( .A(n31568), .B(n25156), .Z(n31570) );
  XOR U32788 ( .A(n31572), .B(n31573), .Z(n25156) );
  AND U32789 ( .A(\modmult_1/xin[1023] ), .B(n31574), .Z(n31573) );
  IV U32790 ( .A(n31572), .Z(n31574) );
  XOR U32791 ( .A(n31575), .B(mreg[931]), .Z(n31572) );
  NAND U32792 ( .A(n31576), .B(mul_pow), .Z(n31575) );
  XOR U32793 ( .A(mreg[931]), .B(creg[931]), .Z(n31576) );
  XOR U32794 ( .A(n31577), .B(n31578), .Z(n31568) );
  ANDN U32795 ( .A(n31579), .B(n25163), .Z(n31578) );
  XOR U32796 ( .A(n31580), .B(\modmult_1/zin[0][929] ), .Z(n25163) );
  IV U32797 ( .A(n31577), .Z(n31580) );
  XNOR U32798 ( .A(n31577), .B(n25162), .Z(n31579) );
  XOR U32799 ( .A(n31581), .B(n31582), .Z(n25162) );
  AND U32800 ( .A(\modmult_1/xin[1023] ), .B(n31583), .Z(n31582) );
  IV U32801 ( .A(n31581), .Z(n31583) );
  XOR U32802 ( .A(n31584), .B(mreg[930]), .Z(n31581) );
  NAND U32803 ( .A(n31585), .B(mul_pow), .Z(n31584) );
  XOR U32804 ( .A(mreg[930]), .B(creg[930]), .Z(n31585) );
  XOR U32805 ( .A(n31586), .B(n31587), .Z(n31577) );
  ANDN U32806 ( .A(n31588), .B(n25169), .Z(n31587) );
  XOR U32807 ( .A(n31589), .B(\modmult_1/zin[0][928] ), .Z(n25169) );
  IV U32808 ( .A(n31586), .Z(n31589) );
  XNOR U32809 ( .A(n31586), .B(n25168), .Z(n31588) );
  XOR U32810 ( .A(n31590), .B(n31591), .Z(n25168) );
  AND U32811 ( .A(\modmult_1/xin[1023] ), .B(n31592), .Z(n31591) );
  IV U32812 ( .A(n31590), .Z(n31592) );
  XOR U32813 ( .A(n31593), .B(mreg[929]), .Z(n31590) );
  NAND U32814 ( .A(n31594), .B(mul_pow), .Z(n31593) );
  XOR U32815 ( .A(mreg[929]), .B(creg[929]), .Z(n31594) );
  XOR U32816 ( .A(n31595), .B(n31596), .Z(n31586) );
  ANDN U32817 ( .A(n31597), .B(n25175), .Z(n31596) );
  XOR U32818 ( .A(n31598), .B(\modmult_1/zin[0][927] ), .Z(n25175) );
  IV U32819 ( .A(n31595), .Z(n31598) );
  XNOR U32820 ( .A(n31595), .B(n25174), .Z(n31597) );
  XOR U32821 ( .A(n31599), .B(n31600), .Z(n25174) );
  AND U32822 ( .A(\modmult_1/xin[1023] ), .B(n31601), .Z(n31600) );
  IV U32823 ( .A(n31599), .Z(n31601) );
  XOR U32824 ( .A(n31602), .B(mreg[928]), .Z(n31599) );
  NAND U32825 ( .A(n31603), .B(mul_pow), .Z(n31602) );
  XOR U32826 ( .A(mreg[928]), .B(creg[928]), .Z(n31603) );
  XOR U32827 ( .A(n31604), .B(n31605), .Z(n31595) );
  ANDN U32828 ( .A(n31606), .B(n25181), .Z(n31605) );
  XOR U32829 ( .A(n31607), .B(\modmult_1/zin[0][926] ), .Z(n25181) );
  IV U32830 ( .A(n31604), .Z(n31607) );
  XNOR U32831 ( .A(n31604), .B(n25180), .Z(n31606) );
  XOR U32832 ( .A(n31608), .B(n31609), .Z(n25180) );
  AND U32833 ( .A(\modmult_1/xin[1023] ), .B(n31610), .Z(n31609) );
  IV U32834 ( .A(n31608), .Z(n31610) );
  XOR U32835 ( .A(n31611), .B(mreg[927]), .Z(n31608) );
  NAND U32836 ( .A(n31612), .B(mul_pow), .Z(n31611) );
  XOR U32837 ( .A(mreg[927]), .B(creg[927]), .Z(n31612) );
  XOR U32838 ( .A(n31613), .B(n31614), .Z(n31604) );
  ANDN U32839 ( .A(n31615), .B(n25187), .Z(n31614) );
  XOR U32840 ( .A(n31616), .B(\modmult_1/zin[0][925] ), .Z(n25187) );
  IV U32841 ( .A(n31613), .Z(n31616) );
  XNOR U32842 ( .A(n31613), .B(n25186), .Z(n31615) );
  XOR U32843 ( .A(n31617), .B(n31618), .Z(n25186) );
  AND U32844 ( .A(\modmult_1/xin[1023] ), .B(n31619), .Z(n31618) );
  IV U32845 ( .A(n31617), .Z(n31619) );
  XOR U32846 ( .A(n31620), .B(mreg[926]), .Z(n31617) );
  NAND U32847 ( .A(n31621), .B(mul_pow), .Z(n31620) );
  XOR U32848 ( .A(mreg[926]), .B(creg[926]), .Z(n31621) );
  XOR U32849 ( .A(n31622), .B(n31623), .Z(n31613) );
  ANDN U32850 ( .A(n31624), .B(n25193), .Z(n31623) );
  XOR U32851 ( .A(n31625), .B(\modmult_1/zin[0][924] ), .Z(n25193) );
  IV U32852 ( .A(n31622), .Z(n31625) );
  XNOR U32853 ( .A(n31622), .B(n25192), .Z(n31624) );
  XOR U32854 ( .A(n31626), .B(n31627), .Z(n25192) );
  AND U32855 ( .A(\modmult_1/xin[1023] ), .B(n31628), .Z(n31627) );
  IV U32856 ( .A(n31626), .Z(n31628) );
  XOR U32857 ( .A(n31629), .B(mreg[925]), .Z(n31626) );
  NAND U32858 ( .A(n31630), .B(mul_pow), .Z(n31629) );
  XOR U32859 ( .A(mreg[925]), .B(creg[925]), .Z(n31630) );
  XOR U32860 ( .A(n31631), .B(n31632), .Z(n31622) );
  ANDN U32861 ( .A(n31633), .B(n25199), .Z(n31632) );
  XOR U32862 ( .A(n31634), .B(\modmult_1/zin[0][923] ), .Z(n25199) );
  IV U32863 ( .A(n31631), .Z(n31634) );
  XNOR U32864 ( .A(n31631), .B(n25198), .Z(n31633) );
  XOR U32865 ( .A(n31635), .B(n31636), .Z(n25198) );
  AND U32866 ( .A(\modmult_1/xin[1023] ), .B(n31637), .Z(n31636) );
  IV U32867 ( .A(n31635), .Z(n31637) );
  XOR U32868 ( .A(n31638), .B(mreg[924]), .Z(n31635) );
  NAND U32869 ( .A(n31639), .B(mul_pow), .Z(n31638) );
  XOR U32870 ( .A(mreg[924]), .B(creg[924]), .Z(n31639) );
  XOR U32871 ( .A(n31640), .B(n31641), .Z(n31631) );
  ANDN U32872 ( .A(n31642), .B(n25205), .Z(n31641) );
  XOR U32873 ( .A(n31643), .B(\modmult_1/zin[0][922] ), .Z(n25205) );
  IV U32874 ( .A(n31640), .Z(n31643) );
  XNOR U32875 ( .A(n31640), .B(n25204), .Z(n31642) );
  XOR U32876 ( .A(n31644), .B(n31645), .Z(n25204) );
  AND U32877 ( .A(\modmult_1/xin[1023] ), .B(n31646), .Z(n31645) );
  IV U32878 ( .A(n31644), .Z(n31646) );
  XOR U32879 ( .A(n31647), .B(mreg[923]), .Z(n31644) );
  NAND U32880 ( .A(n31648), .B(mul_pow), .Z(n31647) );
  XOR U32881 ( .A(mreg[923]), .B(creg[923]), .Z(n31648) );
  XOR U32882 ( .A(n31649), .B(n31650), .Z(n31640) );
  ANDN U32883 ( .A(n31651), .B(n25211), .Z(n31650) );
  XOR U32884 ( .A(n31652), .B(\modmult_1/zin[0][921] ), .Z(n25211) );
  IV U32885 ( .A(n31649), .Z(n31652) );
  XNOR U32886 ( .A(n31649), .B(n25210), .Z(n31651) );
  XOR U32887 ( .A(n31653), .B(n31654), .Z(n25210) );
  AND U32888 ( .A(\modmult_1/xin[1023] ), .B(n31655), .Z(n31654) );
  IV U32889 ( .A(n31653), .Z(n31655) );
  XOR U32890 ( .A(n31656), .B(mreg[922]), .Z(n31653) );
  NAND U32891 ( .A(n31657), .B(mul_pow), .Z(n31656) );
  XOR U32892 ( .A(mreg[922]), .B(creg[922]), .Z(n31657) );
  XOR U32893 ( .A(n31658), .B(n31659), .Z(n31649) );
  ANDN U32894 ( .A(n31660), .B(n25217), .Z(n31659) );
  XOR U32895 ( .A(n31661), .B(\modmult_1/zin[0][920] ), .Z(n25217) );
  IV U32896 ( .A(n31658), .Z(n31661) );
  XNOR U32897 ( .A(n31658), .B(n25216), .Z(n31660) );
  XOR U32898 ( .A(n31662), .B(n31663), .Z(n25216) );
  AND U32899 ( .A(\modmult_1/xin[1023] ), .B(n31664), .Z(n31663) );
  IV U32900 ( .A(n31662), .Z(n31664) );
  XOR U32901 ( .A(n31665), .B(mreg[921]), .Z(n31662) );
  NAND U32902 ( .A(n31666), .B(mul_pow), .Z(n31665) );
  XOR U32903 ( .A(mreg[921]), .B(creg[921]), .Z(n31666) );
  XOR U32904 ( .A(n31667), .B(n31668), .Z(n31658) );
  ANDN U32905 ( .A(n31669), .B(n25223), .Z(n31668) );
  XOR U32906 ( .A(n31670), .B(\modmult_1/zin[0][919] ), .Z(n25223) );
  IV U32907 ( .A(n31667), .Z(n31670) );
  XNOR U32908 ( .A(n31667), .B(n25222), .Z(n31669) );
  XOR U32909 ( .A(n31671), .B(n31672), .Z(n25222) );
  AND U32910 ( .A(\modmult_1/xin[1023] ), .B(n31673), .Z(n31672) );
  IV U32911 ( .A(n31671), .Z(n31673) );
  XOR U32912 ( .A(n31674), .B(mreg[920]), .Z(n31671) );
  NAND U32913 ( .A(n31675), .B(mul_pow), .Z(n31674) );
  XOR U32914 ( .A(mreg[920]), .B(creg[920]), .Z(n31675) );
  XOR U32915 ( .A(n31676), .B(n31677), .Z(n31667) );
  ANDN U32916 ( .A(n31678), .B(n25229), .Z(n31677) );
  XOR U32917 ( .A(n31679), .B(\modmult_1/zin[0][918] ), .Z(n25229) );
  IV U32918 ( .A(n31676), .Z(n31679) );
  XNOR U32919 ( .A(n31676), .B(n25228), .Z(n31678) );
  XOR U32920 ( .A(n31680), .B(n31681), .Z(n25228) );
  AND U32921 ( .A(\modmult_1/xin[1023] ), .B(n31682), .Z(n31681) );
  IV U32922 ( .A(n31680), .Z(n31682) );
  XOR U32923 ( .A(n31683), .B(mreg[919]), .Z(n31680) );
  NAND U32924 ( .A(n31684), .B(mul_pow), .Z(n31683) );
  XOR U32925 ( .A(mreg[919]), .B(creg[919]), .Z(n31684) );
  XOR U32926 ( .A(n31685), .B(n31686), .Z(n31676) );
  ANDN U32927 ( .A(n31687), .B(n25235), .Z(n31686) );
  XOR U32928 ( .A(n31688), .B(\modmult_1/zin[0][917] ), .Z(n25235) );
  IV U32929 ( .A(n31685), .Z(n31688) );
  XNOR U32930 ( .A(n31685), .B(n25234), .Z(n31687) );
  XOR U32931 ( .A(n31689), .B(n31690), .Z(n25234) );
  AND U32932 ( .A(\modmult_1/xin[1023] ), .B(n31691), .Z(n31690) );
  IV U32933 ( .A(n31689), .Z(n31691) );
  XOR U32934 ( .A(n31692), .B(mreg[918]), .Z(n31689) );
  NAND U32935 ( .A(n31693), .B(mul_pow), .Z(n31692) );
  XOR U32936 ( .A(mreg[918]), .B(creg[918]), .Z(n31693) );
  XOR U32937 ( .A(n31694), .B(n31695), .Z(n31685) );
  ANDN U32938 ( .A(n31696), .B(n25241), .Z(n31695) );
  XOR U32939 ( .A(n31697), .B(\modmult_1/zin[0][916] ), .Z(n25241) );
  IV U32940 ( .A(n31694), .Z(n31697) );
  XNOR U32941 ( .A(n31694), .B(n25240), .Z(n31696) );
  XOR U32942 ( .A(n31698), .B(n31699), .Z(n25240) );
  AND U32943 ( .A(\modmult_1/xin[1023] ), .B(n31700), .Z(n31699) );
  IV U32944 ( .A(n31698), .Z(n31700) );
  XOR U32945 ( .A(n31701), .B(mreg[917]), .Z(n31698) );
  NAND U32946 ( .A(n31702), .B(mul_pow), .Z(n31701) );
  XOR U32947 ( .A(mreg[917]), .B(creg[917]), .Z(n31702) );
  XOR U32948 ( .A(n31703), .B(n31704), .Z(n31694) );
  ANDN U32949 ( .A(n31705), .B(n25247), .Z(n31704) );
  XOR U32950 ( .A(n31706), .B(\modmult_1/zin[0][915] ), .Z(n25247) );
  IV U32951 ( .A(n31703), .Z(n31706) );
  XNOR U32952 ( .A(n31703), .B(n25246), .Z(n31705) );
  XOR U32953 ( .A(n31707), .B(n31708), .Z(n25246) );
  AND U32954 ( .A(\modmult_1/xin[1023] ), .B(n31709), .Z(n31708) );
  IV U32955 ( .A(n31707), .Z(n31709) );
  XOR U32956 ( .A(n31710), .B(mreg[916]), .Z(n31707) );
  NAND U32957 ( .A(n31711), .B(mul_pow), .Z(n31710) );
  XOR U32958 ( .A(mreg[916]), .B(creg[916]), .Z(n31711) );
  XOR U32959 ( .A(n31712), .B(n31713), .Z(n31703) );
  ANDN U32960 ( .A(n31714), .B(n25253), .Z(n31713) );
  XOR U32961 ( .A(n31715), .B(\modmult_1/zin[0][914] ), .Z(n25253) );
  IV U32962 ( .A(n31712), .Z(n31715) );
  XNOR U32963 ( .A(n31712), .B(n25252), .Z(n31714) );
  XOR U32964 ( .A(n31716), .B(n31717), .Z(n25252) );
  AND U32965 ( .A(\modmult_1/xin[1023] ), .B(n31718), .Z(n31717) );
  IV U32966 ( .A(n31716), .Z(n31718) );
  XOR U32967 ( .A(n31719), .B(mreg[915]), .Z(n31716) );
  NAND U32968 ( .A(n31720), .B(mul_pow), .Z(n31719) );
  XOR U32969 ( .A(mreg[915]), .B(creg[915]), .Z(n31720) );
  XOR U32970 ( .A(n31721), .B(n31722), .Z(n31712) );
  ANDN U32971 ( .A(n31723), .B(n25259), .Z(n31722) );
  XOR U32972 ( .A(n31724), .B(\modmult_1/zin[0][913] ), .Z(n25259) );
  IV U32973 ( .A(n31721), .Z(n31724) );
  XNOR U32974 ( .A(n31721), .B(n25258), .Z(n31723) );
  XOR U32975 ( .A(n31725), .B(n31726), .Z(n25258) );
  AND U32976 ( .A(\modmult_1/xin[1023] ), .B(n31727), .Z(n31726) );
  IV U32977 ( .A(n31725), .Z(n31727) );
  XOR U32978 ( .A(n31728), .B(mreg[914]), .Z(n31725) );
  NAND U32979 ( .A(n31729), .B(mul_pow), .Z(n31728) );
  XOR U32980 ( .A(mreg[914]), .B(creg[914]), .Z(n31729) );
  XOR U32981 ( .A(n31730), .B(n31731), .Z(n31721) );
  ANDN U32982 ( .A(n31732), .B(n25265), .Z(n31731) );
  XOR U32983 ( .A(n31733), .B(\modmult_1/zin[0][912] ), .Z(n25265) );
  IV U32984 ( .A(n31730), .Z(n31733) );
  XNOR U32985 ( .A(n31730), .B(n25264), .Z(n31732) );
  XOR U32986 ( .A(n31734), .B(n31735), .Z(n25264) );
  AND U32987 ( .A(\modmult_1/xin[1023] ), .B(n31736), .Z(n31735) );
  IV U32988 ( .A(n31734), .Z(n31736) );
  XOR U32989 ( .A(n31737), .B(mreg[913]), .Z(n31734) );
  NAND U32990 ( .A(n31738), .B(mul_pow), .Z(n31737) );
  XOR U32991 ( .A(mreg[913]), .B(creg[913]), .Z(n31738) );
  XOR U32992 ( .A(n31739), .B(n31740), .Z(n31730) );
  ANDN U32993 ( .A(n31741), .B(n25271), .Z(n31740) );
  XOR U32994 ( .A(n31742), .B(\modmult_1/zin[0][911] ), .Z(n25271) );
  IV U32995 ( .A(n31739), .Z(n31742) );
  XNOR U32996 ( .A(n31739), .B(n25270), .Z(n31741) );
  XOR U32997 ( .A(n31743), .B(n31744), .Z(n25270) );
  AND U32998 ( .A(\modmult_1/xin[1023] ), .B(n31745), .Z(n31744) );
  IV U32999 ( .A(n31743), .Z(n31745) );
  XOR U33000 ( .A(n31746), .B(mreg[912]), .Z(n31743) );
  NAND U33001 ( .A(n31747), .B(mul_pow), .Z(n31746) );
  XOR U33002 ( .A(mreg[912]), .B(creg[912]), .Z(n31747) );
  XOR U33003 ( .A(n31748), .B(n31749), .Z(n31739) );
  ANDN U33004 ( .A(n31750), .B(n25277), .Z(n31749) );
  XOR U33005 ( .A(n31751), .B(\modmult_1/zin[0][910] ), .Z(n25277) );
  IV U33006 ( .A(n31748), .Z(n31751) );
  XNOR U33007 ( .A(n31748), .B(n25276), .Z(n31750) );
  XOR U33008 ( .A(n31752), .B(n31753), .Z(n25276) );
  AND U33009 ( .A(\modmult_1/xin[1023] ), .B(n31754), .Z(n31753) );
  IV U33010 ( .A(n31752), .Z(n31754) );
  XOR U33011 ( .A(n31755), .B(mreg[911]), .Z(n31752) );
  NAND U33012 ( .A(n31756), .B(mul_pow), .Z(n31755) );
  XOR U33013 ( .A(mreg[911]), .B(creg[911]), .Z(n31756) );
  XOR U33014 ( .A(n31757), .B(n31758), .Z(n31748) );
  ANDN U33015 ( .A(n31759), .B(n25283), .Z(n31758) );
  XOR U33016 ( .A(n31760), .B(\modmult_1/zin[0][909] ), .Z(n25283) );
  IV U33017 ( .A(n31757), .Z(n31760) );
  XNOR U33018 ( .A(n31757), .B(n25282), .Z(n31759) );
  XOR U33019 ( .A(n31761), .B(n31762), .Z(n25282) );
  AND U33020 ( .A(\modmult_1/xin[1023] ), .B(n31763), .Z(n31762) );
  IV U33021 ( .A(n31761), .Z(n31763) );
  XOR U33022 ( .A(n31764), .B(mreg[910]), .Z(n31761) );
  NAND U33023 ( .A(n31765), .B(mul_pow), .Z(n31764) );
  XOR U33024 ( .A(mreg[910]), .B(creg[910]), .Z(n31765) );
  XOR U33025 ( .A(n31766), .B(n31767), .Z(n31757) );
  ANDN U33026 ( .A(n31768), .B(n25289), .Z(n31767) );
  XOR U33027 ( .A(n31769), .B(\modmult_1/zin[0][908] ), .Z(n25289) );
  IV U33028 ( .A(n31766), .Z(n31769) );
  XNOR U33029 ( .A(n31766), .B(n25288), .Z(n31768) );
  XOR U33030 ( .A(n31770), .B(n31771), .Z(n25288) );
  AND U33031 ( .A(\modmult_1/xin[1023] ), .B(n31772), .Z(n31771) );
  IV U33032 ( .A(n31770), .Z(n31772) );
  XOR U33033 ( .A(n31773), .B(mreg[909]), .Z(n31770) );
  NAND U33034 ( .A(n31774), .B(mul_pow), .Z(n31773) );
  XOR U33035 ( .A(mreg[909]), .B(creg[909]), .Z(n31774) );
  XOR U33036 ( .A(n31775), .B(n31776), .Z(n31766) );
  ANDN U33037 ( .A(n31777), .B(n25295), .Z(n31776) );
  XOR U33038 ( .A(n31778), .B(\modmult_1/zin[0][907] ), .Z(n25295) );
  IV U33039 ( .A(n31775), .Z(n31778) );
  XNOR U33040 ( .A(n31775), .B(n25294), .Z(n31777) );
  XOR U33041 ( .A(n31779), .B(n31780), .Z(n25294) );
  AND U33042 ( .A(\modmult_1/xin[1023] ), .B(n31781), .Z(n31780) );
  IV U33043 ( .A(n31779), .Z(n31781) );
  XOR U33044 ( .A(n31782), .B(mreg[908]), .Z(n31779) );
  NAND U33045 ( .A(n31783), .B(mul_pow), .Z(n31782) );
  XOR U33046 ( .A(mreg[908]), .B(creg[908]), .Z(n31783) );
  XOR U33047 ( .A(n31784), .B(n31785), .Z(n31775) );
  ANDN U33048 ( .A(n31786), .B(n25301), .Z(n31785) );
  XOR U33049 ( .A(n31787), .B(\modmult_1/zin[0][906] ), .Z(n25301) );
  IV U33050 ( .A(n31784), .Z(n31787) );
  XNOR U33051 ( .A(n31784), .B(n25300), .Z(n31786) );
  XOR U33052 ( .A(n31788), .B(n31789), .Z(n25300) );
  AND U33053 ( .A(\modmult_1/xin[1023] ), .B(n31790), .Z(n31789) );
  IV U33054 ( .A(n31788), .Z(n31790) );
  XOR U33055 ( .A(n31791), .B(mreg[907]), .Z(n31788) );
  NAND U33056 ( .A(n31792), .B(mul_pow), .Z(n31791) );
  XOR U33057 ( .A(mreg[907]), .B(creg[907]), .Z(n31792) );
  XOR U33058 ( .A(n31793), .B(n31794), .Z(n31784) );
  ANDN U33059 ( .A(n31795), .B(n25307), .Z(n31794) );
  XOR U33060 ( .A(n31796), .B(\modmult_1/zin[0][905] ), .Z(n25307) );
  IV U33061 ( .A(n31793), .Z(n31796) );
  XNOR U33062 ( .A(n31793), .B(n25306), .Z(n31795) );
  XOR U33063 ( .A(n31797), .B(n31798), .Z(n25306) );
  AND U33064 ( .A(\modmult_1/xin[1023] ), .B(n31799), .Z(n31798) );
  IV U33065 ( .A(n31797), .Z(n31799) );
  XOR U33066 ( .A(n31800), .B(mreg[906]), .Z(n31797) );
  NAND U33067 ( .A(n31801), .B(mul_pow), .Z(n31800) );
  XOR U33068 ( .A(mreg[906]), .B(creg[906]), .Z(n31801) );
  XOR U33069 ( .A(n31802), .B(n31803), .Z(n31793) );
  ANDN U33070 ( .A(n31804), .B(n25313), .Z(n31803) );
  XOR U33071 ( .A(n31805), .B(\modmult_1/zin[0][904] ), .Z(n25313) );
  IV U33072 ( .A(n31802), .Z(n31805) );
  XNOR U33073 ( .A(n31802), .B(n25312), .Z(n31804) );
  XOR U33074 ( .A(n31806), .B(n31807), .Z(n25312) );
  AND U33075 ( .A(\modmult_1/xin[1023] ), .B(n31808), .Z(n31807) );
  IV U33076 ( .A(n31806), .Z(n31808) );
  XOR U33077 ( .A(n31809), .B(mreg[905]), .Z(n31806) );
  NAND U33078 ( .A(n31810), .B(mul_pow), .Z(n31809) );
  XOR U33079 ( .A(mreg[905]), .B(creg[905]), .Z(n31810) );
  XOR U33080 ( .A(n31811), .B(n31812), .Z(n31802) );
  ANDN U33081 ( .A(n31813), .B(n25319), .Z(n31812) );
  XOR U33082 ( .A(n31814), .B(\modmult_1/zin[0][903] ), .Z(n25319) );
  IV U33083 ( .A(n31811), .Z(n31814) );
  XNOR U33084 ( .A(n31811), .B(n25318), .Z(n31813) );
  XOR U33085 ( .A(n31815), .B(n31816), .Z(n25318) );
  AND U33086 ( .A(\modmult_1/xin[1023] ), .B(n31817), .Z(n31816) );
  IV U33087 ( .A(n31815), .Z(n31817) );
  XOR U33088 ( .A(n31818), .B(mreg[904]), .Z(n31815) );
  NAND U33089 ( .A(n31819), .B(mul_pow), .Z(n31818) );
  XOR U33090 ( .A(mreg[904]), .B(creg[904]), .Z(n31819) );
  XOR U33091 ( .A(n31820), .B(n31821), .Z(n31811) );
  ANDN U33092 ( .A(n31822), .B(n25325), .Z(n31821) );
  XOR U33093 ( .A(n31823), .B(\modmult_1/zin[0][902] ), .Z(n25325) );
  IV U33094 ( .A(n31820), .Z(n31823) );
  XNOR U33095 ( .A(n31820), .B(n25324), .Z(n31822) );
  XOR U33096 ( .A(n31824), .B(n31825), .Z(n25324) );
  AND U33097 ( .A(\modmult_1/xin[1023] ), .B(n31826), .Z(n31825) );
  IV U33098 ( .A(n31824), .Z(n31826) );
  XOR U33099 ( .A(n31827), .B(mreg[903]), .Z(n31824) );
  NAND U33100 ( .A(n31828), .B(mul_pow), .Z(n31827) );
  XOR U33101 ( .A(mreg[903]), .B(creg[903]), .Z(n31828) );
  XOR U33102 ( .A(n31829), .B(n31830), .Z(n31820) );
  ANDN U33103 ( .A(n31831), .B(n25331), .Z(n31830) );
  XOR U33104 ( .A(n31832), .B(\modmult_1/zin[0][901] ), .Z(n25331) );
  IV U33105 ( .A(n31829), .Z(n31832) );
  XNOR U33106 ( .A(n31829), .B(n25330), .Z(n31831) );
  XOR U33107 ( .A(n31833), .B(n31834), .Z(n25330) );
  AND U33108 ( .A(\modmult_1/xin[1023] ), .B(n31835), .Z(n31834) );
  IV U33109 ( .A(n31833), .Z(n31835) );
  XOR U33110 ( .A(n31836), .B(mreg[902]), .Z(n31833) );
  NAND U33111 ( .A(n31837), .B(mul_pow), .Z(n31836) );
  XOR U33112 ( .A(mreg[902]), .B(creg[902]), .Z(n31837) );
  XOR U33113 ( .A(n31838), .B(n31839), .Z(n31829) );
  ANDN U33114 ( .A(n31840), .B(n25337), .Z(n31839) );
  XOR U33115 ( .A(n31841), .B(\modmult_1/zin[0][900] ), .Z(n25337) );
  IV U33116 ( .A(n31838), .Z(n31841) );
  XNOR U33117 ( .A(n31838), .B(n25336), .Z(n31840) );
  XOR U33118 ( .A(n31842), .B(n31843), .Z(n25336) );
  AND U33119 ( .A(\modmult_1/xin[1023] ), .B(n31844), .Z(n31843) );
  IV U33120 ( .A(n31842), .Z(n31844) );
  XOR U33121 ( .A(n31845), .B(mreg[901]), .Z(n31842) );
  NAND U33122 ( .A(n31846), .B(mul_pow), .Z(n31845) );
  XOR U33123 ( .A(mreg[901]), .B(creg[901]), .Z(n31846) );
  XOR U33124 ( .A(n31847), .B(n31848), .Z(n31838) );
  ANDN U33125 ( .A(n31849), .B(n25343), .Z(n31848) );
  XOR U33126 ( .A(n31850), .B(\modmult_1/zin[0][899] ), .Z(n25343) );
  IV U33127 ( .A(n31847), .Z(n31850) );
  XNOR U33128 ( .A(n31847), .B(n25342), .Z(n31849) );
  XOR U33129 ( .A(n31851), .B(n31852), .Z(n25342) );
  AND U33130 ( .A(\modmult_1/xin[1023] ), .B(n31853), .Z(n31852) );
  IV U33131 ( .A(n31851), .Z(n31853) );
  XOR U33132 ( .A(n31854), .B(mreg[900]), .Z(n31851) );
  NAND U33133 ( .A(n31855), .B(mul_pow), .Z(n31854) );
  XOR U33134 ( .A(mreg[900]), .B(creg[900]), .Z(n31855) );
  XOR U33135 ( .A(n31856), .B(n31857), .Z(n31847) );
  ANDN U33136 ( .A(n31858), .B(n25349), .Z(n31857) );
  XOR U33137 ( .A(n31859), .B(\modmult_1/zin[0][898] ), .Z(n25349) );
  IV U33138 ( .A(n31856), .Z(n31859) );
  XNOR U33139 ( .A(n31856), .B(n25348), .Z(n31858) );
  XOR U33140 ( .A(n31860), .B(n31861), .Z(n25348) );
  AND U33141 ( .A(\modmult_1/xin[1023] ), .B(n31862), .Z(n31861) );
  IV U33142 ( .A(n31860), .Z(n31862) );
  XOR U33143 ( .A(n31863), .B(mreg[899]), .Z(n31860) );
  NAND U33144 ( .A(n31864), .B(mul_pow), .Z(n31863) );
  XOR U33145 ( .A(mreg[899]), .B(creg[899]), .Z(n31864) );
  XOR U33146 ( .A(n31865), .B(n31866), .Z(n31856) );
  ANDN U33147 ( .A(n31867), .B(n25355), .Z(n31866) );
  XOR U33148 ( .A(n31868), .B(\modmult_1/zin[0][897] ), .Z(n25355) );
  IV U33149 ( .A(n31865), .Z(n31868) );
  XNOR U33150 ( .A(n31865), .B(n25354), .Z(n31867) );
  XOR U33151 ( .A(n31869), .B(n31870), .Z(n25354) );
  AND U33152 ( .A(\modmult_1/xin[1023] ), .B(n31871), .Z(n31870) );
  IV U33153 ( .A(n31869), .Z(n31871) );
  XOR U33154 ( .A(n31872), .B(mreg[898]), .Z(n31869) );
  NAND U33155 ( .A(n31873), .B(mul_pow), .Z(n31872) );
  XOR U33156 ( .A(mreg[898]), .B(creg[898]), .Z(n31873) );
  XOR U33157 ( .A(n31874), .B(n31875), .Z(n31865) );
  ANDN U33158 ( .A(n31876), .B(n25361), .Z(n31875) );
  XOR U33159 ( .A(n31877), .B(\modmult_1/zin[0][896] ), .Z(n25361) );
  IV U33160 ( .A(n31874), .Z(n31877) );
  XNOR U33161 ( .A(n31874), .B(n25360), .Z(n31876) );
  XOR U33162 ( .A(n31878), .B(n31879), .Z(n25360) );
  AND U33163 ( .A(\modmult_1/xin[1023] ), .B(n31880), .Z(n31879) );
  IV U33164 ( .A(n31878), .Z(n31880) );
  XOR U33165 ( .A(n31881), .B(mreg[897]), .Z(n31878) );
  NAND U33166 ( .A(n31882), .B(mul_pow), .Z(n31881) );
  XOR U33167 ( .A(mreg[897]), .B(creg[897]), .Z(n31882) );
  XOR U33168 ( .A(n31883), .B(n31884), .Z(n31874) );
  ANDN U33169 ( .A(n31885), .B(n25367), .Z(n31884) );
  XOR U33170 ( .A(n31886), .B(\modmult_1/zin[0][895] ), .Z(n25367) );
  IV U33171 ( .A(n31883), .Z(n31886) );
  XNOR U33172 ( .A(n31883), .B(n25366), .Z(n31885) );
  XOR U33173 ( .A(n31887), .B(n31888), .Z(n25366) );
  AND U33174 ( .A(\modmult_1/xin[1023] ), .B(n31889), .Z(n31888) );
  IV U33175 ( .A(n31887), .Z(n31889) );
  XOR U33176 ( .A(n31890), .B(mreg[896]), .Z(n31887) );
  NAND U33177 ( .A(n31891), .B(mul_pow), .Z(n31890) );
  XOR U33178 ( .A(mreg[896]), .B(creg[896]), .Z(n31891) );
  XOR U33179 ( .A(n31892), .B(n31893), .Z(n31883) );
  ANDN U33180 ( .A(n31894), .B(n25373), .Z(n31893) );
  XOR U33181 ( .A(n31895), .B(\modmult_1/zin[0][894] ), .Z(n25373) );
  IV U33182 ( .A(n31892), .Z(n31895) );
  XNOR U33183 ( .A(n31892), .B(n25372), .Z(n31894) );
  XOR U33184 ( .A(n31896), .B(n31897), .Z(n25372) );
  AND U33185 ( .A(\modmult_1/xin[1023] ), .B(n31898), .Z(n31897) );
  IV U33186 ( .A(n31896), .Z(n31898) );
  XOR U33187 ( .A(n31899), .B(mreg[895]), .Z(n31896) );
  NAND U33188 ( .A(n31900), .B(mul_pow), .Z(n31899) );
  XOR U33189 ( .A(mreg[895]), .B(creg[895]), .Z(n31900) );
  XOR U33190 ( .A(n31901), .B(n31902), .Z(n31892) );
  ANDN U33191 ( .A(n31903), .B(n25379), .Z(n31902) );
  XOR U33192 ( .A(n31904), .B(\modmult_1/zin[0][893] ), .Z(n25379) );
  IV U33193 ( .A(n31901), .Z(n31904) );
  XNOR U33194 ( .A(n31901), .B(n25378), .Z(n31903) );
  XOR U33195 ( .A(n31905), .B(n31906), .Z(n25378) );
  AND U33196 ( .A(\modmult_1/xin[1023] ), .B(n31907), .Z(n31906) );
  IV U33197 ( .A(n31905), .Z(n31907) );
  XOR U33198 ( .A(n31908), .B(mreg[894]), .Z(n31905) );
  NAND U33199 ( .A(n31909), .B(mul_pow), .Z(n31908) );
  XOR U33200 ( .A(mreg[894]), .B(creg[894]), .Z(n31909) );
  XOR U33201 ( .A(n31910), .B(n31911), .Z(n31901) );
  ANDN U33202 ( .A(n31912), .B(n25385), .Z(n31911) );
  XOR U33203 ( .A(n31913), .B(\modmult_1/zin[0][892] ), .Z(n25385) );
  IV U33204 ( .A(n31910), .Z(n31913) );
  XNOR U33205 ( .A(n31910), .B(n25384), .Z(n31912) );
  XOR U33206 ( .A(n31914), .B(n31915), .Z(n25384) );
  AND U33207 ( .A(\modmult_1/xin[1023] ), .B(n31916), .Z(n31915) );
  IV U33208 ( .A(n31914), .Z(n31916) );
  XOR U33209 ( .A(n31917), .B(mreg[893]), .Z(n31914) );
  NAND U33210 ( .A(n31918), .B(mul_pow), .Z(n31917) );
  XOR U33211 ( .A(mreg[893]), .B(creg[893]), .Z(n31918) );
  XOR U33212 ( .A(n31919), .B(n31920), .Z(n31910) );
  ANDN U33213 ( .A(n31921), .B(n25391), .Z(n31920) );
  XOR U33214 ( .A(n31922), .B(\modmult_1/zin[0][891] ), .Z(n25391) );
  IV U33215 ( .A(n31919), .Z(n31922) );
  XNOR U33216 ( .A(n31919), .B(n25390), .Z(n31921) );
  XOR U33217 ( .A(n31923), .B(n31924), .Z(n25390) );
  AND U33218 ( .A(\modmult_1/xin[1023] ), .B(n31925), .Z(n31924) );
  IV U33219 ( .A(n31923), .Z(n31925) );
  XOR U33220 ( .A(n31926), .B(mreg[892]), .Z(n31923) );
  NAND U33221 ( .A(n31927), .B(mul_pow), .Z(n31926) );
  XOR U33222 ( .A(mreg[892]), .B(creg[892]), .Z(n31927) );
  XOR U33223 ( .A(n31928), .B(n31929), .Z(n31919) );
  ANDN U33224 ( .A(n31930), .B(n25397), .Z(n31929) );
  XOR U33225 ( .A(n31931), .B(\modmult_1/zin[0][890] ), .Z(n25397) );
  IV U33226 ( .A(n31928), .Z(n31931) );
  XNOR U33227 ( .A(n31928), .B(n25396), .Z(n31930) );
  XOR U33228 ( .A(n31932), .B(n31933), .Z(n25396) );
  AND U33229 ( .A(\modmult_1/xin[1023] ), .B(n31934), .Z(n31933) );
  IV U33230 ( .A(n31932), .Z(n31934) );
  XOR U33231 ( .A(n31935), .B(mreg[891]), .Z(n31932) );
  NAND U33232 ( .A(n31936), .B(mul_pow), .Z(n31935) );
  XOR U33233 ( .A(mreg[891]), .B(creg[891]), .Z(n31936) );
  XOR U33234 ( .A(n31937), .B(n31938), .Z(n31928) );
  ANDN U33235 ( .A(n31939), .B(n25403), .Z(n31938) );
  XOR U33236 ( .A(n31940), .B(\modmult_1/zin[0][889] ), .Z(n25403) );
  IV U33237 ( .A(n31937), .Z(n31940) );
  XNOR U33238 ( .A(n31937), .B(n25402), .Z(n31939) );
  XOR U33239 ( .A(n31941), .B(n31942), .Z(n25402) );
  AND U33240 ( .A(\modmult_1/xin[1023] ), .B(n31943), .Z(n31942) );
  IV U33241 ( .A(n31941), .Z(n31943) );
  XOR U33242 ( .A(n31944), .B(mreg[890]), .Z(n31941) );
  NAND U33243 ( .A(n31945), .B(mul_pow), .Z(n31944) );
  XOR U33244 ( .A(mreg[890]), .B(creg[890]), .Z(n31945) );
  XOR U33245 ( .A(n31946), .B(n31947), .Z(n31937) );
  ANDN U33246 ( .A(n31948), .B(n25409), .Z(n31947) );
  XOR U33247 ( .A(n31949), .B(\modmult_1/zin[0][888] ), .Z(n25409) );
  IV U33248 ( .A(n31946), .Z(n31949) );
  XNOR U33249 ( .A(n31946), .B(n25408), .Z(n31948) );
  XOR U33250 ( .A(n31950), .B(n31951), .Z(n25408) );
  AND U33251 ( .A(\modmult_1/xin[1023] ), .B(n31952), .Z(n31951) );
  IV U33252 ( .A(n31950), .Z(n31952) );
  XOR U33253 ( .A(n31953), .B(mreg[889]), .Z(n31950) );
  NAND U33254 ( .A(n31954), .B(mul_pow), .Z(n31953) );
  XOR U33255 ( .A(mreg[889]), .B(creg[889]), .Z(n31954) );
  XOR U33256 ( .A(n31955), .B(n31956), .Z(n31946) );
  ANDN U33257 ( .A(n31957), .B(n25415), .Z(n31956) );
  XOR U33258 ( .A(n31958), .B(\modmult_1/zin[0][887] ), .Z(n25415) );
  IV U33259 ( .A(n31955), .Z(n31958) );
  XNOR U33260 ( .A(n31955), .B(n25414), .Z(n31957) );
  XOR U33261 ( .A(n31959), .B(n31960), .Z(n25414) );
  AND U33262 ( .A(\modmult_1/xin[1023] ), .B(n31961), .Z(n31960) );
  IV U33263 ( .A(n31959), .Z(n31961) );
  XOR U33264 ( .A(n31962), .B(mreg[888]), .Z(n31959) );
  NAND U33265 ( .A(n31963), .B(mul_pow), .Z(n31962) );
  XOR U33266 ( .A(mreg[888]), .B(creg[888]), .Z(n31963) );
  XOR U33267 ( .A(n31964), .B(n31965), .Z(n31955) );
  ANDN U33268 ( .A(n31966), .B(n25421), .Z(n31965) );
  XOR U33269 ( .A(n31967), .B(\modmult_1/zin[0][886] ), .Z(n25421) );
  IV U33270 ( .A(n31964), .Z(n31967) );
  XNOR U33271 ( .A(n31964), .B(n25420), .Z(n31966) );
  XOR U33272 ( .A(n31968), .B(n31969), .Z(n25420) );
  AND U33273 ( .A(\modmult_1/xin[1023] ), .B(n31970), .Z(n31969) );
  IV U33274 ( .A(n31968), .Z(n31970) );
  XOR U33275 ( .A(n31971), .B(mreg[887]), .Z(n31968) );
  NAND U33276 ( .A(n31972), .B(mul_pow), .Z(n31971) );
  XOR U33277 ( .A(mreg[887]), .B(creg[887]), .Z(n31972) );
  XOR U33278 ( .A(n31973), .B(n31974), .Z(n31964) );
  ANDN U33279 ( .A(n31975), .B(n25427), .Z(n31974) );
  XOR U33280 ( .A(n31976), .B(\modmult_1/zin[0][885] ), .Z(n25427) );
  IV U33281 ( .A(n31973), .Z(n31976) );
  XNOR U33282 ( .A(n31973), .B(n25426), .Z(n31975) );
  XOR U33283 ( .A(n31977), .B(n31978), .Z(n25426) );
  AND U33284 ( .A(\modmult_1/xin[1023] ), .B(n31979), .Z(n31978) );
  IV U33285 ( .A(n31977), .Z(n31979) );
  XOR U33286 ( .A(n31980), .B(mreg[886]), .Z(n31977) );
  NAND U33287 ( .A(n31981), .B(mul_pow), .Z(n31980) );
  XOR U33288 ( .A(mreg[886]), .B(creg[886]), .Z(n31981) );
  XOR U33289 ( .A(n31982), .B(n31983), .Z(n31973) );
  ANDN U33290 ( .A(n31984), .B(n25433), .Z(n31983) );
  XOR U33291 ( .A(n31985), .B(\modmult_1/zin[0][884] ), .Z(n25433) );
  IV U33292 ( .A(n31982), .Z(n31985) );
  XNOR U33293 ( .A(n31982), .B(n25432), .Z(n31984) );
  XOR U33294 ( .A(n31986), .B(n31987), .Z(n25432) );
  AND U33295 ( .A(\modmult_1/xin[1023] ), .B(n31988), .Z(n31987) );
  IV U33296 ( .A(n31986), .Z(n31988) );
  XOR U33297 ( .A(n31989), .B(mreg[885]), .Z(n31986) );
  NAND U33298 ( .A(n31990), .B(mul_pow), .Z(n31989) );
  XOR U33299 ( .A(mreg[885]), .B(creg[885]), .Z(n31990) );
  XOR U33300 ( .A(n31991), .B(n31992), .Z(n31982) );
  ANDN U33301 ( .A(n31993), .B(n25439), .Z(n31992) );
  XOR U33302 ( .A(n31994), .B(\modmult_1/zin[0][883] ), .Z(n25439) );
  IV U33303 ( .A(n31991), .Z(n31994) );
  XNOR U33304 ( .A(n31991), .B(n25438), .Z(n31993) );
  XOR U33305 ( .A(n31995), .B(n31996), .Z(n25438) );
  AND U33306 ( .A(\modmult_1/xin[1023] ), .B(n31997), .Z(n31996) );
  IV U33307 ( .A(n31995), .Z(n31997) );
  XOR U33308 ( .A(n31998), .B(mreg[884]), .Z(n31995) );
  NAND U33309 ( .A(n31999), .B(mul_pow), .Z(n31998) );
  XOR U33310 ( .A(mreg[884]), .B(creg[884]), .Z(n31999) );
  XOR U33311 ( .A(n32000), .B(n32001), .Z(n31991) );
  ANDN U33312 ( .A(n32002), .B(n25445), .Z(n32001) );
  XOR U33313 ( .A(n32003), .B(\modmult_1/zin[0][882] ), .Z(n25445) );
  IV U33314 ( .A(n32000), .Z(n32003) );
  XNOR U33315 ( .A(n32000), .B(n25444), .Z(n32002) );
  XOR U33316 ( .A(n32004), .B(n32005), .Z(n25444) );
  AND U33317 ( .A(\modmult_1/xin[1023] ), .B(n32006), .Z(n32005) );
  IV U33318 ( .A(n32004), .Z(n32006) );
  XOR U33319 ( .A(n32007), .B(mreg[883]), .Z(n32004) );
  NAND U33320 ( .A(n32008), .B(mul_pow), .Z(n32007) );
  XOR U33321 ( .A(mreg[883]), .B(creg[883]), .Z(n32008) );
  XOR U33322 ( .A(n32009), .B(n32010), .Z(n32000) );
  ANDN U33323 ( .A(n32011), .B(n25451), .Z(n32010) );
  XOR U33324 ( .A(n32012), .B(\modmult_1/zin[0][881] ), .Z(n25451) );
  IV U33325 ( .A(n32009), .Z(n32012) );
  XNOR U33326 ( .A(n32009), .B(n25450), .Z(n32011) );
  XOR U33327 ( .A(n32013), .B(n32014), .Z(n25450) );
  AND U33328 ( .A(\modmult_1/xin[1023] ), .B(n32015), .Z(n32014) );
  IV U33329 ( .A(n32013), .Z(n32015) );
  XOR U33330 ( .A(n32016), .B(mreg[882]), .Z(n32013) );
  NAND U33331 ( .A(n32017), .B(mul_pow), .Z(n32016) );
  XOR U33332 ( .A(mreg[882]), .B(creg[882]), .Z(n32017) );
  XOR U33333 ( .A(n32018), .B(n32019), .Z(n32009) );
  ANDN U33334 ( .A(n32020), .B(n25457), .Z(n32019) );
  XOR U33335 ( .A(n32021), .B(\modmult_1/zin[0][880] ), .Z(n25457) );
  IV U33336 ( .A(n32018), .Z(n32021) );
  XNOR U33337 ( .A(n32018), .B(n25456), .Z(n32020) );
  XOR U33338 ( .A(n32022), .B(n32023), .Z(n25456) );
  AND U33339 ( .A(\modmult_1/xin[1023] ), .B(n32024), .Z(n32023) );
  IV U33340 ( .A(n32022), .Z(n32024) );
  XOR U33341 ( .A(n32025), .B(mreg[881]), .Z(n32022) );
  NAND U33342 ( .A(n32026), .B(mul_pow), .Z(n32025) );
  XOR U33343 ( .A(mreg[881]), .B(creg[881]), .Z(n32026) );
  XOR U33344 ( .A(n32027), .B(n32028), .Z(n32018) );
  ANDN U33345 ( .A(n32029), .B(n25463), .Z(n32028) );
  XOR U33346 ( .A(n32030), .B(\modmult_1/zin[0][879] ), .Z(n25463) );
  IV U33347 ( .A(n32027), .Z(n32030) );
  XNOR U33348 ( .A(n32027), .B(n25462), .Z(n32029) );
  XOR U33349 ( .A(n32031), .B(n32032), .Z(n25462) );
  AND U33350 ( .A(\modmult_1/xin[1023] ), .B(n32033), .Z(n32032) );
  IV U33351 ( .A(n32031), .Z(n32033) );
  XOR U33352 ( .A(n32034), .B(mreg[880]), .Z(n32031) );
  NAND U33353 ( .A(n32035), .B(mul_pow), .Z(n32034) );
  XOR U33354 ( .A(mreg[880]), .B(creg[880]), .Z(n32035) );
  XOR U33355 ( .A(n32036), .B(n32037), .Z(n32027) );
  ANDN U33356 ( .A(n32038), .B(n25469), .Z(n32037) );
  XOR U33357 ( .A(n32039), .B(\modmult_1/zin[0][878] ), .Z(n25469) );
  IV U33358 ( .A(n32036), .Z(n32039) );
  XNOR U33359 ( .A(n32036), .B(n25468), .Z(n32038) );
  XOR U33360 ( .A(n32040), .B(n32041), .Z(n25468) );
  AND U33361 ( .A(\modmult_1/xin[1023] ), .B(n32042), .Z(n32041) );
  IV U33362 ( .A(n32040), .Z(n32042) );
  XOR U33363 ( .A(n32043), .B(mreg[879]), .Z(n32040) );
  NAND U33364 ( .A(n32044), .B(mul_pow), .Z(n32043) );
  XOR U33365 ( .A(mreg[879]), .B(creg[879]), .Z(n32044) );
  XOR U33366 ( .A(n32045), .B(n32046), .Z(n32036) );
  ANDN U33367 ( .A(n32047), .B(n25475), .Z(n32046) );
  XOR U33368 ( .A(n32048), .B(\modmult_1/zin[0][877] ), .Z(n25475) );
  IV U33369 ( .A(n32045), .Z(n32048) );
  XNOR U33370 ( .A(n32045), .B(n25474), .Z(n32047) );
  XOR U33371 ( .A(n32049), .B(n32050), .Z(n25474) );
  AND U33372 ( .A(\modmult_1/xin[1023] ), .B(n32051), .Z(n32050) );
  IV U33373 ( .A(n32049), .Z(n32051) );
  XOR U33374 ( .A(n32052), .B(mreg[878]), .Z(n32049) );
  NAND U33375 ( .A(n32053), .B(mul_pow), .Z(n32052) );
  XOR U33376 ( .A(mreg[878]), .B(creg[878]), .Z(n32053) );
  XOR U33377 ( .A(n32054), .B(n32055), .Z(n32045) );
  ANDN U33378 ( .A(n32056), .B(n25481), .Z(n32055) );
  XOR U33379 ( .A(n32057), .B(\modmult_1/zin[0][876] ), .Z(n25481) );
  IV U33380 ( .A(n32054), .Z(n32057) );
  XNOR U33381 ( .A(n32054), .B(n25480), .Z(n32056) );
  XOR U33382 ( .A(n32058), .B(n32059), .Z(n25480) );
  AND U33383 ( .A(\modmult_1/xin[1023] ), .B(n32060), .Z(n32059) );
  IV U33384 ( .A(n32058), .Z(n32060) );
  XOR U33385 ( .A(n32061), .B(mreg[877]), .Z(n32058) );
  NAND U33386 ( .A(n32062), .B(mul_pow), .Z(n32061) );
  XOR U33387 ( .A(mreg[877]), .B(creg[877]), .Z(n32062) );
  XOR U33388 ( .A(n32063), .B(n32064), .Z(n32054) );
  ANDN U33389 ( .A(n32065), .B(n25487), .Z(n32064) );
  XOR U33390 ( .A(n32066), .B(\modmult_1/zin[0][875] ), .Z(n25487) );
  IV U33391 ( .A(n32063), .Z(n32066) );
  XNOR U33392 ( .A(n32063), .B(n25486), .Z(n32065) );
  XOR U33393 ( .A(n32067), .B(n32068), .Z(n25486) );
  AND U33394 ( .A(\modmult_1/xin[1023] ), .B(n32069), .Z(n32068) );
  IV U33395 ( .A(n32067), .Z(n32069) );
  XOR U33396 ( .A(n32070), .B(mreg[876]), .Z(n32067) );
  NAND U33397 ( .A(n32071), .B(mul_pow), .Z(n32070) );
  XOR U33398 ( .A(mreg[876]), .B(creg[876]), .Z(n32071) );
  XOR U33399 ( .A(n32072), .B(n32073), .Z(n32063) );
  ANDN U33400 ( .A(n32074), .B(n25493), .Z(n32073) );
  XOR U33401 ( .A(n32075), .B(\modmult_1/zin[0][874] ), .Z(n25493) );
  IV U33402 ( .A(n32072), .Z(n32075) );
  XNOR U33403 ( .A(n32072), .B(n25492), .Z(n32074) );
  XOR U33404 ( .A(n32076), .B(n32077), .Z(n25492) );
  AND U33405 ( .A(\modmult_1/xin[1023] ), .B(n32078), .Z(n32077) );
  IV U33406 ( .A(n32076), .Z(n32078) );
  XOR U33407 ( .A(n32079), .B(mreg[875]), .Z(n32076) );
  NAND U33408 ( .A(n32080), .B(mul_pow), .Z(n32079) );
  XOR U33409 ( .A(mreg[875]), .B(creg[875]), .Z(n32080) );
  XOR U33410 ( .A(n32081), .B(n32082), .Z(n32072) );
  ANDN U33411 ( .A(n32083), .B(n25499), .Z(n32082) );
  XOR U33412 ( .A(n32084), .B(\modmult_1/zin[0][873] ), .Z(n25499) );
  IV U33413 ( .A(n32081), .Z(n32084) );
  XNOR U33414 ( .A(n32081), .B(n25498), .Z(n32083) );
  XOR U33415 ( .A(n32085), .B(n32086), .Z(n25498) );
  AND U33416 ( .A(\modmult_1/xin[1023] ), .B(n32087), .Z(n32086) );
  IV U33417 ( .A(n32085), .Z(n32087) );
  XOR U33418 ( .A(n32088), .B(mreg[874]), .Z(n32085) );
  NAND U33419 ( .A(n32089), .B(mul_pow), .Z(n32088) );
  XOR U33420 ( .A(mreg[874]), .B(creg[874]), .Z(n32089) );
  XOR U33421 ( .A(n32090), .B(n32091), .Z(n32081) );
  ANDN U33422 ( .A(n32092), .B(n25505), .Z(n32091) );
  XOR U33423 ( .A(n32093), .B(\modmult_1/zin[0][872] ), .Z(n25505) );
  IV U33424 ( .A(n32090), .Z(n32093) );
  XNOR U33425 ( .A(n32090), .B(n25504), .Z(n32092) );
  XOR U33426 ( .A(n32094), .B(n32095), .Z(n25504) );
  AND U33427 ( .A(\modmult_1/xin[1023] ), .B(n32096), .Z(n32095) );
  IV U33428 ( .A(n32094), .Z(n32096) );
  XOR U33429 ( .A(n32097), .B(mreg[873]), .Z(n32094) );
  NAND U33430 ( .A(n32098), .B(mul_pow), .Z(n32097) );
  XOR U33431 ( .A(mreg[873]), .B(creg[873]), .Z(n32098) );
  XOR U33432 ( .A(n32099), .B(n32100), .Z(n32090) );
  ANDN U33433 ( .A(n32101), .B(n25511), .Z(n32100) );
  XOR U33434 ( .A(n32102), .B(\modmult_1/zin[0][871] ), .Z(n25511) );
  IV U33435 ( .A(n32099), .Z(n32102) );
  XNOR U33436 ( .A(n32099), .B(n25510), .Z(n32101) );
  XOR U33437 ( .A(n32103), .B(n32104), .Z(n25510) );
  AND U33438 ( .A(\modmult_1/xin[1023] ), .B(n32105), .Z(n32104) );
  IV U33439 ( .A(n32103), .Z(n32105) );
  XOR U33440 ( .A(n32106), .B(mreg[872]), .Z(n32103) );
  NAND U33441 ( .A(n32107), .B(mul_pow), .Z(n32106) );
  XOR U33442 ( .A(mreg[872]), .B(creg[872]), .Z(n32107) );
  XOR U33443 ( .A(n32108), .B(n32109), .Z(n32099) );
  ANDN U33444 ( .A(n32110), .B(n25517), .Z(n32109) );
  XOR U33445 ( .A(n32111), .B(\modmult_1/zin[0][870] ), .Z(n25517) );
  IV U33446 ( .A(n32108), .Z(n32111) );
  XNOR U33447 ( .A(n32108), .B(n25516), .Z(n32110) );
  XOR U33448 ( .A(n32112), .B(n32113), .Z(n25516) );
  AND U33449 ( .A(\modmult_1/xin[1023] ), .B(n32114), .Z(n32113) );
  IV U33450 ( .A(n32112), .Z(n32114) );
  XOR U33451 ( .A(n32115), .B(mreg[871]), .Z(n32112) );
  NAND U33452 ( .A(n32116), .B(mul_pow), .Z(n32115) );
  XOR U33453 ( .A(mreg[871]), .B(creg[871]), .Z(n32116) );
  XOR U33454 ( .A(n32117), .B(n32118), .Z(n32108) );
  ANDN U33455 ( .A(n32119), .B(n25523), .Z(n32118) );
  XOR U33456 ( .A(n32120), .B(\modmult_1/zin[0][869] ), .Z(n25523) );
  IV U33457 ( .A(n32117), .Z(n32120) );
  XNOR U33458 ( .A(n32117), .B(n25522), .Z(n32119) );
  XOR U33459 ( .A(n32121), .B(n32122), .Z(n25522) );
  AND U33460 ( .A(\modmult_1/xin[1023] ), .B(n32123), .Z(n32122) );
  IV U33461 ( .A(n32121), .Z(n32123) );
  XOR U33462 ( .A(n32124), .B(mreg[870]), .Z(n32121) );
  NAND U33463 ( .A(n32125), .B(mul_pow), .Z(n32124) );
  XOR U33464 ( .A(mreg[870]), .B(creg[870]), .Z(n32125) );
  XOR U33465 ( .A(n32126), .B(n32127), .Z(n32117) );
  ANDN U33466 ( .A(n32128), .B(n25529), .Z(n32127) );
  XOR U33467 ( .A(n32129), .B(\modmult_1/zin[0][868] ), .Z(n25529) );
  IV U33468 ( .A(n32126), .Z(n32129) );
  XNOR U33469 ( .A(n32126), .B(n25528), .Z(n32128) );
  XOR U33470 ( .A(n32130), .B(n32131), .Z(n25528) );
  AND U33471 ( .A(\modmult_1/xin[1023] ), .B(n32132), .Z(n32131) );
  IV U33472 ( .A(n32130), .Z(n32132) );
  XOR U33473 ( .A(n32133), .B(mreg[869]), .Z(n32130) );
  NAND U33474 ( .A(n32134), .B(mul_pow), .Z(n32133) );
  XOR U33475 ( .A(mreg[869]), .B(creg[869]), .Z(n32134) );
  XOR U33476 ( .A(n32135), .B(n32136), .Z(n32126) );
  ANDN U33477 ( .A(n32137), .B(n25535), .Z(n32136) );
  XOR U33478 ( .A(n32138), .B(\modmult_1/zin[0][867] ), .Z(n25535) );
  IV U33479 ( .A(n32135), .Z(n32138) );
  XNOR U33480 ( .A(n32135), .B(n25534), .Z(n32137) );
  XOR U33481 ( .A(n32139), .B(n32140), .Z(n25534) );
  AND U33482 ( .A(\modmult_1/xin[1023] ), .B(n32141), .Z(n32140) );
  IV U33483 ( .A(n32139), .Z(n32141) );
  XOR U33484 ( .A(n32142), .B(mreg[868]), .Z(n32139) );
  NAND U33485 ( .A(n32143), .B(mul_pow), .Z(n32142) );
  XOR U33486 ( .A(mreg[868]), .B(creg[868]), .Z(n32143) );
  XOR U33487 ( .A(n32144), .B(n32145), .Z(n32135) );
  ANDN U33488 ( .A(n32146), .B(n25541), .Z(n32145) );
  XOR U33489 ( .A(n32147), .B(\modmult_1/zin[0][866] ), .Z(n25541) );
  IV U33490 ( .A(n32144), .Z(n32147) );
  XNOR U33491 ( .A(n32144), .B(n25540), .Z(n32146) );
  XOR U33492 ( .A(n32148), .B(n32149), .Z(n25540) );
  AND U33493 ( .A(\modmult_1/xin[1023] ), .B(n32150), .Z(n32149) );
  IV U33494 ( .A(n32148), .Z(n32150) );
  XOR U33495 ( .A(n32151), .B(mreg[867]), .Z(n32148) );
  NAND U33496 ( .A(n32152), .B(mul_pow), .Z(n32151) );
  XOR U33497 ( .A(mreg[867]), .B(creg[867]), .Z(n32152) );
  XOR U33498 ( .A(n32153), .B(n32154), .Z(n32144) );
  ANDN U33499 ( .A(n32155), .B(n25547), .Z(n32154) );
  XOR U33500 ( .A(n32156), .B(\modmult_1/zin[0][865] ), .Z(n25547) );
  IV U33501 ( .A(n32153), .Z(n32156) );
  XNOR U33502 ( .A(n32153), .B(n25546), .Z(n32155) );
  XOR U33503 ( .A(n32157), .B(n32158), .Z(n25546) );
  AND U33504 ( .A(\modmult_1/xin[1023] ), .B(n32159), .Z(n32158) );
  IV U33505 ( .A(n32157), .Z(n32159) );
  XOR U33506 ( .A(n32160), .B(mreg[866]), .Z(n32157) );
  NAND U33507 ( .A(n32161), .B(mul_pow), .Z(n32160) );
  XOR U33508 ( .A(mreg[866]), .B(creg[866]), .Z(n32161) );
  XOR U33509 ( .A(n32162), .B(n32163), .Z(n32153) );
  ANDN U33510 ( .A(n32164), .B(n25553), .Z(n32163) );
  XOR U33511 ( .A(n32165), .B(\modmult_1/zin[0][864] ), .Z(n25553) );
  IV U33512 ( .A(n32162), .Z(n32165) );
  XNOR U33513 ( .A(n32162), .B(n25552), .Z(n32164) );
  XOR U33514 ( .A(n32166), .B(n32167), .Z(n25552) );
  AND U33515 ( .A(\modmult_1/xin[1023] ), .B(n32168), .Z(n32167) );
  IV U33516 ( .A(n32166), .Z(n32168) );
  XOR U33517 ( .A(n32169), .B(mreg[865]), .Z(n32166) );
  NAND U33518 ( .A(n32170), .B(mul_pow), .Z(n32169) );
  XOR U33519 ( .A(mreg[865]), .B(creg[865]), .Z(n32170) );
  XOR U33520 ( .A(n32171), .B(n32172), .Z(n32162) );
  ANDN U33521 ( .A(n32173), .B(n25559), .Z(n32172) );
  XOR U33522 ( .A(n32174), .B(\modmult_1/zin[0][863] ), .Z(n25559) );
  IV U33523 ( .A(n32171), .Z(n32174) );
  XNOR U33524 ( .A(n32171), .B(n25558), .Z(n32173) );
  XOR U33525 ( .A(n32175), .B(n32176), .Z(n25558) );
  AND U33526 ( .A(\modmult_1/xin[1023] ), .B(n32177), .Z(n32176) );
  IV U33527 ( .A(n32175), .Z(n32177) );
  XOR U33528 ( .A(n32178), .B(mreg[864]), .Z(n32175) );
  NAND U33529 ( .A(n32179), .B(mul_pow), .Z(n32178) );
  XOR U33530 ( .A(mreg[864]), .B(creg[864]), .Z(n32179) );
  XOR U33531 ( .A(n32180), .B(n32181), .Z(n32171) );
  ANDN U33532 ( .A(n32182), .B(n25565), .Z(n32181) );
  XOR U33533 ( .A(n32183), .B(\modmult_1/zin[0][862] ), .Z(n25565) );
  IV U33534 ( .A(n32180), .Z(n32183) );
  XNOR U33535 ( .A(n32180), .B(n25564), .Z(n32182) );
  XOR U33536 ( .A(n32184), .B(n32185), .Z(n25564) );
  AND U33537 ( .A(\modmult_1/xin[1023] ), .B(n32186), .Z(n32185) );
  IV U33538 ( .A(n32184), .Z(n32186) );
  XOR U33539 ( .A(n32187), .B(mreg[863]), .Z(n32184) );
  NAND U33540 ( .A(n32188), .B(mul_pow), .Z(n32187) );
  XOR U33541 ( .A(mreg[863]), .B(creg[863]), .Z(n32188) );
  XOR U33542 ( .A(n32189), .B(n32190), .Z(n32180) );
  ANDN U33543 ( .A(n32191), .B(n25571), .Z(n32190) );
  XOR U33544 ( .A(n32192), .B(\modmult_1/zin[0][861] ), .Z(n25571) );
  IV U33545 ( .A(n32189), .Z(n32192) );
  XNOR U33546 ( .A(n32189), .B(n25570), .Z(n32191) );
  XOR U33547 ( .A(n32193), .B(n32194), .Z(n25570) );
  AND U33548 ( .A(\modmult_1/xin[1023] ), .B(n32195), .Z(n32194) );
  IV U33549 ( .A(n32193), .Z(n32195) );
  XOR U33550 ( .A(n32196), .B(mreg[862]), .Z(n32193) );
  NAND U33551 ( .A(n32197), .B(mul_pow), .Z(n32196) );
  XOR U33552 ( .A(mreg[862]), .B(creg[862]), .Z(n32197) );
  XOR U33553 ( .A(n32198), .B(n32199), .Z(n32189) );
  ANDN U33554 ( .A(n32200), .B(n25577), .Z(n32199) );
  XOR U33555 ( .A(n32201), .B(\modmult_1/zin[0][860] ), .Z(n25577) );
  IV U33556 ( .A(n32198), .Z(n32201) );
  XNOR U33557 ( .A(n32198), .B(n25576), .Z(n32200) );
  XOR U33558 ( .A(n32202), .B(n32203), .Z(n25576) );
  AND U33559 ( .A(\modmult_1/xin[1023] ), .B(n32204), .Z(n32203) );
  IV U33560 ( .A(n32202), .Z(n32204) );
  XOR U33561 ( .A(n32205), .B(mreg[861]), .Z(n32202) );
  NAND U33562 ( .A(n32206), .B(mul_pow), .Z(n32205) );
  XOR U33563 ( .A(mreg[861]), .B(creg[861]), .Z(n32206) );
  XOR U33564 ( .A(n32207), .B(n32208), .Z(n32198) );
  ANDN U33565 ( .A(n32209), .B(n25583), .Z(n32208) );
  XOR U33566 ( .A(n32210), .B(\modmult_1/zin[0][859] ), .Z(n25583) );
  IV U33567 ( .A(n32207), .Z(n32210) );
  XNOR U33568 ( .A(n32207), .B(n25582), .Z(n32209) );
  XOR U33569 ( .A(n32211), .B(n32212), .Z(n25582) );
  AND U33570 ( .A(\modmult_1/xin[1023] ), .B(n32213), .Z(n32212) );
  IV U33571 ( .A(n32211), .Z(n32213) );
  XOR U33572 ( .A(n32214), .B(mreg[860]), .Z(n32211) );
  NAND U33573 ( .A(n32215), .B(mul_pow), .Z(n32214) );
  XOR U33574 ( .A(mreg[860]), .B(creg[860]), .Z(n32215) );
  XOR U33575 ( .A(n32216), .B(n32217), .Z(n32207) );
  ANDN U33576 ( .A(n32218), .B(n25589), .Z(n32217) );
  XOR U33577 ( .A(n32219), .B(\modmult_1/zin[0][858] ), .Z(n25589) );
  IV U33578 ( .A(n32216), .Z(n32219) );
  XNOR U33579 ( .A(n32216), .B(n25588), .Z(n32218) );
  XOR U33580 ( .A(n32220), .B(n32221), .Z(n25588) );
  AND U33581 ( .A(\modmult_1/xin[1023] ), .B(n32222), .Z(n32221) );
  IV U33582 ( .A(n32220), .Z(n32222) );
  XOR U33583 ( .A(n32223), .B(mreg[859]), .Z(n32220) );
  NAND U33584 ( .A(n32224), .B(mul_pow), .Z(n32223) );
  XOR U33585 ( .A(mreg[859]), .B(creg[859]), .Z(n32224) );
  XOR U33586 ( .A(n32225), .B(n32226), .Z(n32216) );
  ANDN U33587 ( .A(n32227), .B(n25595), .Z(n32226) );
  XOR U33588 ( .A(n32228), .B(\modmult_1/zin[0][857] ), .Z(n25595) );
  IV U33589 ( .A(n32225), .Z(n32228) );
  XNOR U33590 ( .A(n32225), .B(n25594), .Z(n32227) );
  XOR U33591 ( .A(n32229), .B(n32230), .Z(n25594) );
  AND U33592 ( .A(\modmult_1/xin[1023] ), .B(n32231), .Z(n32230) );
  IV U33593 ( .A(n32229), .Z(n32231) );
  XOR U33594 ( .A(n32232), .B(mreg[858]), .Z(n32229) );
  NAND U33595 ( .A(n32233), .B(mul_pow), .Z(n32232) );
  XOR U33596 ( .A(mreg[858]), .B(creg[858]), .Z(n32233) );
  XOR U33597 ( .A(n32234), .B(n32235), .Z(n32225) );
  ANDN U33598 ( .A(n32236), .B(n25601), .Z(n32235) );
  XOR U33599 ( .A(n32237), .B(\modmult_1/zin[0][856] ), .Z(n25601) );
  IV U33600 ( .A(n32234), .Z(n32237) );
  XNOR U33601 ( .A(n32234), .B(n25600), .Z(n32236) );
  XOR U33602 ( .A(n32238), .B(n32239), .Z(n25600) );
  AND U33603 ( .A(\modmult_1/xin[1023] ), .B(n32240), .Z(n32239) );
  IV U33604 ( .A(n32238), .Z(n32240) );
  XOR U33605 ( .A(n32241), .B(mreg[857]), .Z(n32238) );
  NAND U33606 ( .A(n32242), .B(mul_pow), .Z(n32241) );
  XOR U33607 ( .A(mreg[857]), .B(creg[857]), .Z(n32242) );
  XOR U33608 ( .A(n32243), .B(n32244), .Z(n32234) );
  ANDN U33609 ( .A(n32245), .B(n25607), .Z(n32244) );
  XOR U33610 ( .A(n32246), .B(\modmult_1/zin[0][855] ), .Z(n25607) );
  IV U33611 ( .A(n32243), .Z(n32246) );
  XNOR U33612 ( .A(n32243), .B(n25606), .Z(n32245) );
  XOR U33613 ( .A(n32247), .B(n32248), .Z(n25606) );
  AND U33614 ( .A(\modmult_1/xin[1023] ), .B(n32249), .Z(n32248) );
  IV U33615 ( .A(n32247), .Z(n32249) );
  XOR U33616 ( .A(n32250), .B(mreg[856]), .Z(n32247) );
  NAND U33617 ( .A(n32251), .B(mul_pow), .Z(n32250) );
  XOR U33618 ( .A(mreg[856]), .B(creg[856]), .Z(n32251) );
  XOR U33619 ( .A(n32252), .B(n32253), .Z(n32243) );
  ANDN U33620 ( .A(n32254), .B(n25613), .Z(n32253) );
  XOR U33621 ( .A(n32255), .B(\modmult_1/zin[0][854] ), .Z(n25613) );
  IV U33622 ( .A(n32252), .Z(n32255) );
  XNOR U33623 ( .A(n32252), .B(n25612), .Z(n32254) );
  XOR U33624 ( .A(n32256), .B(n32257), .Z(n25612) );
  AND U33625 ( .A(\modmult_1/xin[1023] ), .B(n32258), .Z(n32257) );
  IV U33626 ( .A(n32256), .Z(n32258) );
  XOR U33627 ( .A(n32259), .B(mreg[855]), .Z(n32256) );
  NAND U33628 ( .A(n32260), .B(mul_pow), .Z(n32259) );
  XOR U33629 ( .A(mreg[855]), .B(creg[855]), .Z(n32260) );
  XOR U33630 ( .A(n32261), .B(n32262), .Z(n32252) );
  ANDN U33631 ( .A(n32263), .B(n25619), .Z(n32262) );
  XOR U33632 ( .A(n32264), .B(\modmult_1/zin[0][853] ), .Z(n25619) );
  IV U33633 ( .A(n32261), .Z(n32264) );
  XNOR U33634 ( .A(n32261), .B(n25618), .Z(n32263) );
  XOR U33635 ( .A(n32265), .B(n32266), .Z(n25618) );
  AND U33636 ( .A(\modmult_1/xin[1023] ), .B(n32267), .Z(n32266) );
  IV U33637 ( .A(n32265), .Z(n32267) );
  XOR U33638 ( .A(n32268), .B(mreg[854]), .Z(n32265) );
  NAND U33639 ( .A(n32269), .B(mul_pow), .Z(n32268) );
  XOR U33640 ( .A(mreg[854]), .B(creg[854]), .Z(n32269) );
  XOR U33641 ( .A(n32270), .B(n32271), .Z(n32261) );
  ANDN U33642 ( .A(n32272), .B(n25625), .Z(n32271) );
  XOR U33643 ( .A(n32273), .B(\modmult_1/zin[0][852] ), .Z(n25625) );
  IV U33644 ( .A(n32270), .Z(n32273) );
  XNOR U33645 ( .A(n32270), .B(n25624), .Z(n32272) );
  XOR U33646 ( .A(n32274), .B(n32275), .Z(n25624) );
  AND U33647 ( .A(\modmult_1/xin[1023] ), .B(n32276), .Z(n32275) );
  IV U33648 ( .A(n32274), .Z(n32276) );
  XOR U33649 ( .A(n32277), .B(mreg[853]), .Z(n32274) );
  NAND U33650 ( .A(n32278), .B(mul_pow), .Z(n32277) );
  XOR U33651 ( .A(mreg[853]), .B(creg[853]), .Z(n32278) );
  XOR U33652 ( .A(n32279), .B(n32280), .Z(n32270) );
  ANDN U33653 ( .A(n32281), .B(n25631), .Z(n32280) );
  XOR U33654 ( .A(n32282), .B(\modmult_1/zin[0][851] ), .Z(n25631) );
  IV U33655 ( .A(n32279), .Z(n32282) );
  XNOR U33656 ( .A(n32279), .B(n25630), .Z(n32281) );
  XOR U33657 ( .A(n32283), .B(n32284), .Z(n25630) );
  AND U33658 ( .A(\modmult_1/xin[1023] ), .B(n32285), .Z(n32284) );
  IV U33659 ( .A(n32283), .Z(n32285) );
  XOR U33660 ( .A(n32286), .B(mreg[852]), .Z(n32283) );
  NAND U33661 ( .A(n32287), .B(mul_pow), .Z(n32286) );
  XOR U33662 ( .A(mreg[852]), .B(creg[852]), .Z(n32287) );
  XOR U33663 ( .A(n32288), .B(n32289), .Z(n32279) );
  ANDN U33664 ( .A(n32290), .B(n25637), .Z(n32289) );
  XOR U33665 ( .A(n32291), .B(\modmult_1/zin[0][850] ), .Z(n25637) );
  IV U33666 ( .A(n32288), .Z(n32291) );
  XNOR U33667 ( .A(n32288), .B(n25636), .Z(n32290) );
  XOR U33668 ( .A(n32292), .B(n32293), .Z(n25636) );
  AND U33669 ( .A(\modmult_1/xin[1023] ), .B(n32294), .Z(n32293) );
  IV U33670 ( .A(n32292), .Z(n32294) );
  XOR U33671 ( .A(n32295), .B(mreg[851]), .Z(n32292) );
  NAND U33672 ( .A(n32296), .B(mul_pow), .Z(n32295) );
  XOR U33673 ( .A(mreg[851]), .B(creg[851]), .Z(n32296) );
  XOR U33674 ( .A(n32297), .B(n32298), .Z(n32288) );
  ANDN U33675 ( .A(n32299), .B(n25643), .Z(n32298) );
  XOR U33676 ( .A(n32300), .B(\modmult_1/zin[0][849] ), .Z(n25643) );
  IV U33677 ( .A(n32297), .Z(n32300) );
  XNOR U33678 ( .A(n32297), .B(n25642), .Z(n32299) );
  XOR U33679 ( .A(n32301), .B(n32302), .Z(n25642) );
  AND U33680 ( .A(\modmult_1/xin[1023] ), .B(n32303), .Z(n32302) );
  IV U33681 ( .A(n32301), .Z(n32303) );
  XOR U33682 ( .A(n32304), .B(mreg[850]), .Z(n32301) );
  NAND U33683 ( .A(n32305), .B(mul_pow), .Z(n32304) );
  XOR U33684 ( .A(mreg[850]), .B(creg[850]), .Z(n32305) );
  XOR U33685 ( .A(n32306), .B(n32307), .Z(n32297) );
  ANDN U33686 ( .A(n32308), .B(n25649), .Z(n32307) );
  XOR U33687 ( .A(n32309), .B(\modmult_1/zin[0][848] ), .Z(n25649) );
  IV U33688 ( .A(n32306), .Z(n32309) );
  XNOR U33689 ( .A(n32306), .B(n25648), .Z(n32308) );
  XOR U33690 ( .A(n32310), .B(n32311), .Z(n25648) );
  AND U33691 ( .A(\modmult_1/xin[1023] ), .B(n32312), .Z(n32311) );
  IV U33692 ( .A(n32310), .Z(n32312) );
  XOR U33693 ( .A(n32313), .B(mreg[849]), .Z(n32310) );
  NAND U33694 ( .A(n32314), .B(mul_pow), .Z(n32313) );
  XOR U33695 ( .A(mreg[849]), .B(creg[849]), .Z(n32314) );
  XOR U33696 ( .A(n32315), .B(n32316), .Z(n32306) );
  ANDN U33697 ( .A(n32317), .B(n25655), .Z(n32316) );
  XOR U33698 ( .A(n32318), .B(\modmult_1/zin[0][847] ), .Z(n25655) );
  IV U33699 ( .A(n32315), .Z(n32318) );
  XNOR U33700 ( .A(n32315), .B(n25654), .Z(n32317) );
  XOR U33701 ( .A(n32319), .B(n32320), .Z(n25654) );
  AND U33702 ( .A(\modmult_1/xin[1023] ), .B(n32321), .Z(n32320) );
  IV U33703 ( .A(n32319), .Z(n32321) );
  XOR U33704 ( .A(n32322), .B(mreg[848]), .Z(n32319) );
  NAND U33705 ( .A(n32323), .B(mul_pow), .Z(n32322) );
  XOR U33706 ( .A(mreg[848]), .B(creg[848]), .Z(n32323) );
  XOR U33707 ( .A(n32324), .B(n32325), .Z(n32315) );
  ANDN U33708 ( .A(n32326), .B(n25661), .Z(n32325) );
  XOR U33709 ( .A(n32327), .B(\modmult_1/zin[0][846] ), .Z(n25661) );
  IV U33710 ( .A(n32324), .Z(n32327) );
  XNOR U33711 ( .A(n32324), .B(n25660), .Z(n32326) );
  XOR U33712 ( .A(n32328), .B(n32329), .Z(n25660) );
  AND U33713 ( .A(\modmult_1/xin[1023] ), .B(n32330), .Z(n32329) );
  IV U33714 ( .A(n32328), .Z(n32330) );
  XOR U33715 ( .A(n32331), .B(mreg[847]), .Z(n32328) );
  NAND U33716 ( .A(n32332), .B(mul_pow), .Z(n32331) );
  XOR U33717 ( .A(mreg[847]), .B(creg[847]), .Z(n32332) );
  XOR U33718 ( .A(n32333), .B(n32334), .Z(n32324) );
  ANDN U33719 ( .A(n32335), .B(n25667), .Z(n32334) );
  XOR U33720 ( .A(n32336), .B(\modmult_1/zin[0][845] ), .Z(n25667) );
  IV U33721 ( .A(n32333), .Z(n32336) );
  XNOR U33722 ( .A(n32333), .B(n25666), .Z(n32335) );
  XOR U33723 ( .A(n32337), .B(n32338), .Z(n25666) );
  AND U33724 ( .A(\modmult_1/xin[1023] ), .B(n32339), .Z(n32338) );
  IV U33725 ( .A(n32337), .Z(n32339) );
  XOR U33726 ( .A(n32340), .B(mreg[846]), .Z(n32337) );
  NAND U33727 ( .A(n32341), .B(mul_pow), .Z(n32340) );
  XOR U33728 ( .A(mreg[846]), .B(creg[846]), .Z(n32341) );
  XOR U33729 ( .A(n32342), .B(n32343), .Z(n32333) );
  ANDN U33730 ( .A(n32344), .B(n25673), .Z(n32343) );
  XOR U33731 ( .A(n32345), .B(\modmult_1/zin[0][844] ), .Z(n25673) );
  IV U33732 ( .A(n32342), .Z(n32345) );
  XNOR U33733 ( .A(n32342), .B(n25672), .Z(n32344) );
  XOR U33734 ( .A(n32346), .B(n32347), .Z(n25672) );
  AND U33735 ( .A(\modmult_1/xin[1023] ), .B(n32348), .Z(n32347) );
  IV U33736 ( .A(n32346), .Z(n32348) );
  XOR U33737 ( .A(n32349), .B(mreg[845]), .Z(n32346) );
  NAND U33738 ( .A(n32350), .B(mul_pow), .Z(n32349) );
  XOR U33739 ( .A(mreg[845]), .B(creg[845]), .Z(n32350) );
  XOR U33740 ( .A(n32351), .B(n32352), .Z(n32342) );
  ANDN U33741 ( .A(n32353), .B(n25679), .Z(n32352) );
  XOR U33742 ( .A(n32354), .B(\modmult_1/zin[0][843] ), .Z(n25679) );
  IV U33743 ( .A(n32351), .Z(n32354) );
  XNOR U33744 ( .A(n32351), .B(n25678), .Z(n32353) );
  XOR U33745 ( .A(n32355), .B(n32356), .Z(n25678) );
  AND U33746 ( .A(\modmult_1/xin[1023] ), .B(n32357), .Z(n32356) );
  IV U33747 ( .A(n32355), .Z(n32357) );
  XOR U33748 ( .A(n32358), .B(mreg[844]), .Z(n32355) );
  NAND U33749 ( .A(n32359), .B(mul_pow), .Z(n32358) );
  XOR U33750 ( .A(mreg[844]), .B(creg[844]), .Z(n32359) );
  XOR U33751 ( .A(n32360), .B(n32361), .Z(n32351) );
  ANDN U33752 ( .A(n32362), .B(n25685), .Z(n32361) );
  XOR U33753 ( .A(n32363), .B(\modmult_1/zin[0][842] ), .Z(n25685) );
  IV U33754 ( .A(n32360), .Z(n32363) );
  XNOR U33755 ( .A(n32360), .B(n25684), .Z(n32362) );
  XOR U33756 ( .A(n32364), .B(n32365), .Z(n25684) );
  AND U33757 ( .A(\modmult_1/xin[1023] ), .B(n32366), .Z(n32365) );
  IV U33758 ( .A(n32364), .Z(n32366) );
  XOR U33759 ( .A(n32367), .B(mreg[843]), .Z(n32364) );
  NAND U33760 ( .A(n32368), .B(mul_pow), .Z(n32367) );
  XOR U33761 ( .A(mreg[843]), .B(creg[843]), .Z(n32368) );
  XOR U33762 ( .A(n32369), .B(n32370), .Z(n32360) );
  ANDN U33763 ( .A(n32371), .B(n25691), .Z(n32370) );
  XOR U33764 ( .A(n32372), .B(\modmult_1/zin[0][841] ), .Z(n25691) );
  IV U33765 ( .A(n32369), .Z(n32372) );
  XNOR U33766 ( .A(n32369), .B(n25690), .Z(n32371) );
  XOR U33767 ( .A(n32373), .B(n32374), .Z(n25690) );
  AND U33768 ( .A(\modmult_1/xin[1023] ), .B(n32375), .Z(n32374) );
  IV U33769 ( .A(n32373), .Z(n32375) );
  XOR U33770 ( .A(n32376), .B(mreg[842]), .Z(n32373) );
  NAND U33771 ( .A(n32377), .B(mul_pow), .Z(n32376) );
  XOR U33772 ( .A(mreg[842]), .B(creg[842]), .Z(n32377) );
  XOR U33773 ( .A(n32378), .B(n32379), .Z(n32369) );
  ANDN U33774 ( .A(n32380), .B(n25697), .Z(n32379) );
  XOR U33775 ( .A(n32381), .B(\modmult_1/zin[0][840] ), .Z(n25697) );
  IV U33776 ( .A(n32378), .Z(n32381) );
  XNOR U33777 ( .A(n32378), .B(n25696), .Z(n32380) );
  XOR U33778 ( .A(n32382), .B(n32383), .Z(n25696) );
  AND U33779 ( .A(\modmult_1/xin[1023] ), .B(n32384), .Z(n32383) );
  IV U33780 ( .A(n32382), .Z(n32384) );
  XOR U33781 ( .A(n32385), .B(mreg[841]), .Z(n32382) );
  NAND U33782 ( .A(n32386), .B(mul_pow), .Z(n32385) );
  XOR U33783 ( .A(mreg[841]), .B(creg[841]), .Z(n32386) );
  XOR U33784 ( .A(n32387), .B(n32388), .Z(n32378) );
  ANDN U33785 ( .A(n32389), .B(n25703), .Z(n32388) );
  XOR U33786 ( .A(n32390), .B(\modmult_1/zin[0][839] ), .Z(n25703) );
  IV U33787 ( .A(n32387), .Z(n32390) );
  XNOR U33788 ( .A(n32387), .B(n25702), .Z(n32389) );
  XOR U33789 ( .A(n32391), .B(n32392), .Z(n25702) );
  AND U33790 ( .A(\modmult_1/xin[1023] ), .B(n32393), .Z(n32392) );
  IV U33791 ( .A(n32391), .Z(n32393) );
  XOR U33792 ( .A(n32394), .B(mreg[840]), .Z(n32391) );
  NAND U33793 ( .A(n32395), .B(mul_pow), .Z(n32394) );
  XOR U33794 ( .A(mreg[840]), .B(creg[840]), .Z(n32395) );
  XOR U33795 ( .A(n32396), .B(n32397), .Z(n32387) );
  ANDN U33796 ( .A(n32398), .B(n25709), .Z(n32397) );
  XOR U33797 ( .A(n32399), .B(\modmult_1/zin[0][838] ), .Z(n25709) );
  IV U33798 ( .A(n32396), .Z(n32399) );
  XNOR U33799 ( .A(n32396), .B(n25708), .Z(n32398) );
  XOR U33800 ( .A(n32400), .B(n32401), .Z(n25708) );
  AND U33801 ( .A(\modmult_1/xin[1023] ), .B(n32402), .Z(n32401) );
  IV U33802 ( .A(n32400), .Z(n32402) );
  XOR U33803 ( .A(n32403), .B(mreg[839]), .Z(n32400) );
  NAND U33804 ( .A(n32404), .B(mul_pow), .Z(n32403) );
  XOR U33805 ( .A(mreg[839]), .B(creg[839]), .Z(n32404) );
  XOR U33806 ( .A(n32405), .B(n32406), .Z(n32396) );
  ANDN U33807 ( .A(n32407), .B(n25715), .Z(n32406) );
  XOR U33808 ( .A(n32408), .B(\modmult_1/zin[0][837] ), .Z(n25715) );
  IV U33809 ( .A(n32405), .Z(n32408) );
  XNOR U33810 ( .A(n32405), .B(n25714), .Z(n32407) );
  XOR U33811 ( .A(n32409), .B(n32410), .Z(n25714) );
  AND U33812 ( .A(\modmult_1/xin[1023] ), .B(n32411), .Z(n32410) );
  IV U33813 ( .A(n32409), .Z(n32411) );
  XOR U33814 ( .A(n32412), .B(mreg[838]), .Z(n32409) );
  NAND U33815 ( .A(n32413), .B(mul_pow), .Z(n32412) );
  XOR U33816 ( .A(mreg[838]), .B(creg[838]), .Z(n32413) );
  XOR U33817 ( .A(n32414), .B(n32415), .Z(n32405) );
  ANDN U33818 ( .A(n32416), .B(n25721), .Z(n32415) );
  XOR U33819 ( .A(n32417), .B(\modmult_1/zin[0][836] ), .Z(n25721) );
  IV U33820 ( .A(n32414), .Z(n32417) );
  XNOR U33821 ( .A(n32414), .B(n25720), .Z(n32416) );
  XOR U33822 ( .A(n32418), .B(n32419), .Z(n25720) );
  AND U33823 ( .A(\modmult_1/xin[1023] ), .B(n32420), .Z(n32419) );
  IV U33824 ( .A(n32418), .Z(n32420) );
  XOR U33825 ( .A(n32421), .B(mreg[837]), .Z(n32418) );
  NAND U33826 ( .A(n32422), .B(mul_pow), .Z(n32421) );
  XOR U33827 ( .A(mreg[837]), .B(creg[837]), .Z(n32422) );
  XOR U33828 ( .A(n32423), .B(n32424), .Z(n32414) );
  ANDN U33829 ( .A(n32425), .B(n25727), .Z(n32424) );
  XOR U33830 ( .A(n32426), .B(\modmult_1/zin[0][835] ), .Z(n25727) );
  IV U33831 ( .A(n32423), .Z(n32426) );
  XNOR U33832 ( .A(n32423), .B(n25726), .Z(n32425) );
  XOR U33833 ( .A(n32427), .B(n32428), .Z(n25726) );
  AND U33834 ( .A(\modmult_1/xin[1023] ), .B(n32429), .Z(n32428) );
  IV U33835 ( .A(n32427), .Z(n32429) );
  XOR U33836 ( .A(n32430), .B(mreg[836]), .Z(n32427) );
  NAND U33837 ( .A(n32431), .B(mul_pow), .Z(n32430) );
  XOR U33838 ( .A(mreg[836]), .B(creg[836]), .Z(n32431) );
  XOR U33839 ( .A(n32432), .B(n32433), .Z(n32423) );
  ANDN U33840 ( .A(n32434), .B(n25733), .Z(n32433) );
  XOR U33841 ( .A(n32435), .B(\modmult_1/zin[0][834] ), .Z(n25733) );
  IV U33842 ( .A(n32432), .Z(n32435) );
  XNOR U33843 ( .A(n32432), .B(n25732), .Z(n32434) );
  XOR U33844 ( .A(n32436), .B(n32437), .Z(n25732) );
  AND U33845 ( .A(\modmult_1/xin[1023] ), .B(n32438), .Z(n32437) );
  IV U33846 ( .A(n32436), .Z(n32438) );
  XOR U33847 ( .A(n32439), .B(mreg[835]), .Z(n32436) );
  NAND U33848 ( .A(n32440), .B(mul_pow), .Z(n32439) );
  XOR U33849 ( .A(mreg[835]), .B(creg[835]), .Z(n32440) );
  XOR U33850 ( .A(n32441), .B(n32442), .Z(n32432) );
  ANDN U33851 ( .A(n32443), .B(n25739), .Z(n32442) );
  XOR U33852 ( .A(n32444), .B(\modmult_1/zin[0][833] ), .Z(n25739) );
  IV U33853 ( .A(n32441), .Z(n32444) );
  XNOR U33854 ( .A(n32441), .B(n25738), .Z(n32443) );
  XOR U33855 ( .A(n32445), .B(n32446), .Z(n25738) );
  AND U33856 ( .A(\modmult_1/xin[1023] ), .B(n32447), .Z(n32446) );
  IV U33857 ( .A(n32445), .Z(n32447) );
  XOR U33858 ( .A(n32448), .B(mreg[834]), .Z(n32445) );
  NAND U33859 ( .A(n32449), .B(mul_pow), .Z(n32448) );
  XOR U33860 ( .A(mreg[834]), .B(creg[834]), .Z(n32449) );
  XOR U33861 ( .A(n32450), .B(n32451), .Z(n32441) );
  ANDN U33862 ( .A(n32452), .B(n25745), .Z(n32451) );
  XOR U33863 ( .A(n32453), .B(\modmult_1/zin[0][832] ), .Z(n25745) );
  IV U33864 ( .A(n32450), .Z(n32453) );
  XNOR U33865 ( .A(n32450), .B(n25744), .Z(n32452) );
  XOR U33866 ( .A(n32454), .B(n32455), .Z(n25744) );
  AND U33867 ( .A(\modmult_1/xin[1023] ), .B(n32456), .Z(n32455) );
  IV U33868 ( .A(n32454), .Z(n32456) );
  XOR U33869 ( .A(n32457), .B(mreg[833]), .Z(n32454) );
  NAND U33870 ( .A(n32458), .B(mul_pow), .Z(n32457) );
  XOR U33871 ( .A(mreg[833]), .B(creg[833]), .Z(n32458) );
  XOR U33872 ( .A(n32459), .B(n32460), .Z(n32450) );
  ANDN U33873 ( .A(n32461), .B(n25751), .Z(n32460) );
  XOR U33874 ( .A(n32462), .B(\modmult_1/zin[0][831] ), .Z(n25751) );
  IV U33875 ( .A(n32459), .Z(n32462) );
  XNOR U33876 ( .A(n32459), .B(n25750), .Z(n32461) );
  XOR U33877 ( .A(n32463), .B(n32464), .Z(n25750) );
  AND U33878 ( .A(\modmult_1/xin[1023] ), .B(n32465), .Z(n32464) );
  IV U33879 ( .A(n32463), .Z(n32465) );
  XOR U33880 ( .A(n32466), .B(mreg[832]), .Z(n32463) );
  NAND U33881 ( .A(n32467), .B(mul_pow), .Z(n32466) );
  XOR U33882 ( .A(mreg[832]), .B(creg[832]), .Z(n32467) );
  XOR U33883 ( .A(n32468), .B(n32469), .Z(n32459) );
  ANDN U33884 ( .A(n32470), .B(n25757), .Z(n32469) );
  XOR U33885 ( .A(n32471), .B(\modmult_1/zin[0][830] ), .Z(n25757) );
  IV U33886 ( .A(n32468), .Z(n32471) );
  XNOR U33887 ( .A(n32468), .B(n25756), .Z(n32470) );
  XOR U33888 ( .A(n32472), .B(n32473), .Z(n25756) );
  AND U33889 ( .A(\modmult_1/xin[1023] ), .B(n32474), .Z(n32473) );
  IV U33890 ( .A(n32472), .Z(n32474) );
  XOR U33891 ( .A(n32475), .B(mreg[831]), .Z(n32472) );
  NAND U33892 ( .A(n32476), .B(mul_pow), .Z(n32475) );
  XOR U33893 ( .A(mreg[831]), .B(creg[831]), .Z(n32476) );
  XOR U33894 ( .A(n32477), .B(n32478), .Z(n32468) );
  ANDN U33895 ( .A(n32479), .B(n25763), .Z(n32478) );
  XOR U33896 ( .A(n32480), .B(\modmult_1/zin[0][829] ), .Z(n25763) );
  IV U33897 ( .A(n32477), .Z(n32480) );
  XNOR U33898 ( .A(n32477), .B(n25762), .Z(n32479) );
  XOR U33899 ( .A(n32481), .B(n32482), .Z(n25762) );
  AND U33900 ( .A(\modmult_1/xin[1023] ), .B(n32483), .Z(n32482) );
  IV U33901 ( .A(n32481), .Z(n32483) );
  XOR U33902 ( .A(n32484), .B(mreg[830]), .Z(n32481) );
  NAND U33903 ( .A(n32485), .B(mul_pow), .Z(n32484) );
  XOR U33904 ( .A(mreg[830]), .B(creg[830]), .Z(n32485) );
  XOR U33905 ( .A(n32486), .B(n32487), .Z(n32477) );
  ANDN U33906 ( .A(n32488), .B(n25769), .Z(n32487) );
  XOR U33907 ( .A(n32489), .B(\modmult_1/zin[0][828] ), .Z(n25769) );
  IV U33908 ( .A(n32486), .Z(n32489) );
  XNOR U33909 ( .A(n32486), .B(n25768), .Z(n32488) );
  XOR U33910 ( .A(n32490), .B(n32491), .Z(n25768) );
  AND U33911 ( .A(\modmult_1/xin[1023] ), .B(n32492), .Z(n32491) );
  IV U33912 ( .A(n32490), .Z(n32492) );
  XOR U33913 ( .A(n32493), .B(mreg[829]), .Z(n32490) );
  NAND U33914 ( .A(n32494), .B(mul_pow), .Z(n32493) );
  XOR U33915 ( .A(mreg[829]), .B(creg[829]), .Z(n32494) );
  XOR U33916 ( .A(n32495), .B(n32496), .Z(n32486) );
  ANDN U33917 ( .A(n32497), .B(n25775), .Z(n32496) );
  XOR U33918 ( .A(n32498), .B(\modmult_1/zin[0][827] ), .Z(n25775) );
  IV U33919 ( .A(n32495), .Z(n32498) );
  XNOR U33920 ( .A(n32495), .B(n25774), .Z(n32497) );
  XOR U33921 ( .A(n32499), .B(n32500), .Z(n25774) );
  AND U33922 ( .A(\modmult_1/xin[1023] ), .B(n32501), .Z(n32500) );
  IV U33923 ( .A(n32499), .Z(n32501) );
  XOR U33924 ( .A(n32502), .B(mreg[828]), .Z(n32499) );
  NAND U33925 ( .A(n32503), .B(mul_pow), .Z(n32502) );
  XOR U33926 ( .A(mreg[828]), .B(creg[828]), .Z(n32503) );
  XOR U33927 ( .A(n32504), .B(n32505), .Z(n32495) );
  ANDN U33928 ( .A(n32506), .B(n25781), .Z(n32505) );
  XOR U33929 ( .A(n32507), .B(\modmult_1/zin[0][826] ), .Z(n25781) );
  IV U33930 ( .A(n32504), .Z(n32507) );
  XNOR U33931 ( .A(n32504), .B(n25780), .Z(n32506) );
  XOR U33932 ( .A(n32508), .B(n32509), .Z(n25780) );
  AND U33933 ( .A(\modmult_1/xin[1023] ), .B(n32510), .Z(n32509) );
  IV U33934 ( .A(n32508), .Z(n32510) );
  XOR U33935 ( .A(n32511), .B(mreg[827]), .Z(n32508) );
  NAND U33936 ( .A(n32512), .B(mul_pow), .Z(n32511) );
  XOR U33937 ( .A(mreg[827]), .B(creg[827]), .Z(n32512) );
  XOR U33938 ( .A(n32513), .B(n32514), .Z(n32504) );
  ANDN U33939 ( .A(n32515), .B(n25787), .Z(n32514) );
  XOR U33940 ( .A(n32516), .B(\modmult_1/zin[0][825] ), .Z(n25787) );
  IV U33941 ( .A(n32513), .Z(n32516) );
  XNOR U33942 ( .A(n32513), .B(n25786), .Z(n32515) );
  XOR U33943 ( .A(n32517), .B(n32518), .Z(n25786) );
  AND U33944 ( .A(\modmult_1/xin[1023] ), .B(n32519), .Z(n32518) );
  IV U33945 ( .A(n32517), .Z(n32519) );
  XOR U33946 ( .A(n32520), .B(mreg[826]), .Z(n32517) );
  NAND U33947 ( .A(n32521), .B(mul_pow), .Z(n32520) );
  XOR U33948 ( .A(mreg[826]), .B(creg[826]), .Z(n32521) );
  XOR U33949 ( .A(n32522), .B(n32523), .Z(n32513) );
  ANDN U33950 ( .A(n32524), .B(n25793), .Z(n32523) );
  XOR U33951 ( .A(n32525), .B(\modmult_1/zin[0][824] ), .Z(n25793) );
  IV U33952 ( .A(n32522), .Z(n32525) );
  XNOR U33953 ( .A(n32522), .B(n25792), .Z(n32524) );
  XOR U33954 ( .A(n32526), .B(n32527), .Z(n25792) );
  AND U33955 ( .A(\modmult_1/xin[1023] ), .B(n32528), .Z(n32527) );
  IV U33956 ( .A(n32526), .Z(n32528) );
  XOR U33957 ( .A(n32529), .B(mreg[825]), .Z(n32526) );
  NAND U33958 ( .A(n32530), .B(mul_pow), .Z(n32529) );
  XOR U33959 ( .A(mreg[825]), .B(creg[825]), .Z(n32530) );
  XOR U33960 ( .A(n32531), .B(n32532), .Z(n32522) );
  ANDN U33961 ( .A(n32533), .B(n25799), .Z(n32532) );
  XOR U33962 ( .A(n32534), .B(\modmult_1/zin[0][823] ), .Z(n25799) );
  IV U33963 ( .A(n32531), .Z(n32534) );
  XNOR U33964 ( .A(n32531), .B(n25798), .Z(n32533) );
  XOR U33965 ( .A(n32535), .B(n32536), .Z(n25798) );
  AND U33966 ( .A(\modmult_1/xin[1023] ), .B(n32537), .Z(n32536) );
  IV U33967 ( .A(n32535), .Z(n32537) );
  XOR U33968 ( .A(n32538), .B(mreg[824]), .Z(n32535) );
  NAND U33969 ( .A(n32539), .B(mul_pow), .Z(n32538) );
  XOR U33970 ( .A(mreg[824]), .B(creg[824]), .Z(n32539) );
  XOR U33971 ( .A(n32540), .B(n32541), .Z(n32531) );
  ANDN U33972 ( .A(n32542), .B(n25805), .Z(n32541) );
  XOR U33973 ( .A(n32543), .B(\modmult_1/zin[0][822] ), .Z(n25805) );
  IV U33974 ( .A(n32540), .Z(n32543) );
  XNOR U33975 ( .A(n32540), .B(n25804), .Z(n32542) );
  XOR U33976 ( .A(n32544), .B(n32545), .Z(n25804) );
  AND U33977 ( .A(\modmult_1/xin[1023] ), .B(n32546), .Z(n32545) );
  IV U33978 ( .A(n32544), .Z(n32546) );
  XOR U33979 ( .A(n32547), .B(mreg[823]), .Z(n32544) );
  NAND U33980 ( .A(n32548), .B(mul_pow), .Z(n32547) );
  XOR U33981 ( .A(mreg[823]), .B(creg[823]), .Z(n32548) );
  XOR U33982 ( .A(n32549), .B(n32550), .Z(n32540) );
  ANDN U33983 ( .A(n32551), .B(n25811), .Z(n32550) );
  XOR U33984 ( .A(n32552), .B(\modmult_1/zin[0][821] ), .Z(n25811) );
  IV U33985 ( .A(n32549), .Z(n32552) );
  XNOR U33986 ( .A(n32549), .B(n25810), .Z(n32551) );
  XOR U33987 ( .A(n32553), .B(n32554), .Z(n25810) );
  AND U33988 ( .A(\modmult_1/xin[1023] ), .B(n32555), .Z(n32554) );
  IV U33989 ( .A(n32553), .Z(n32555) );
  XOR U33990 ( .A(n32556), .B(mreg[822]), .Z(n32553) );
  NAND U33991 ( .A(n32557), .B(mul_pow), .Z(n32556) );
  XOR U33992 ( .A(mreg[822]), .B(creg[822]), .Z(n32557) );
  XOR U33993 ( .A(n32558), .B(n32559), .Z(n32549) );
  ANDN U33994 ( .A(n32560), .B(n25817), .Z(n32559) );
  XOR U33995 ( .A(n32561), .B(\modmult_1/zin[0][820] ), .Z(n25817) );
  IV U33996 ( .A(n32558), .Z(n32561) );
  XNOR U33997 ( .A(n32558), .B(n25816), .Z(n32560) );
  XOR U33998 ( .A(n32562), .B(n32563), .Z(n25816) );
  AND U33999 ( .A(\modmult_1/xin[1023] ), .B(n32564), .Z(n32563) );
  IV U34000 ( .A(n32562), .Z(n32564) );
  XOR U34001 ( .A(n32565), .B(mreg[821]), .Z(n32562) );
  NAND U34002 ( .A(n32566), .B(mul_pow), .Z(n32565) );
  XOR U34003 ( .A(mreg[821]), .B(creg[821]), .Z(n32566) );
  XOR U34004 ( .A(n32567), .B(n32568), .Z(n32558) );
  ANDN U34005 ( .A(n32569), .B(n25823), .Z(n32568) );
  XOR U34006 ( .A(n32570), .B(\modmult_1/zin[0][819] ), .Z(n25823) );
  IV U34007 ( .A(n32567), .Z(n32570) );
  XNOR U34008 ( .A(n32567), .B(n25822), .Z(n32569) );
  XOR U34009 ( .A(n32571), .B(n32572), .Z(n25822) );
  AND U34010 ( .A(\modmult_1/xin[1023] ), .B(n32573), .Z(n32572) );
  IV U34011 ( .A(n32571), .Z(n32573) );
  XOR U34012 ( .A(n32574), .B(mreg[820]), .Z(n32571) );
  NAND U34013 ( .A(n32575), .B(mul_pow), .Z(n32574) );
  XOR U34014 ( .A(mreg[820]), .B(creg[820]), .Z(n32575) );
  XOR U34015 ( .A(n32576), .B(n32577), .Z(n32567) );
  ANDN U34016 ( .A(n32578), .B(n25829), .Z(n32577) );
  XOR U34017 ( .A(n32579), .B(\modmult_1/zin[0][818] ), .Z(n25829) );
  IV U34018 ( .A(n32576), .Z(n32579) );
  XNOR U34019 ( .A(n32576), .B(n25828), .Z(n32578) );
  XOR U34020 ( .A(n32580), .B(n32581), .Z(n25828) );
  AND U34021 ( .A(\modmult_1/xin[1023] ), .B(n32582), .Z(n32581) );
  IV U34022 ( .A(n32580), .Z(n32582) );
  XOR U34023 ( .A(n32583), .B(mreg[819]), .Z(n32580) );
  NAND U34024 ( .A(n32584), .B(mul_pow), .Z(n32583) );
  XOR U34025 ( .A(mreg[819]), .B(creg[819]), .Z(n32584) );
  XOR U34026 ( .A(n32585), .B(n32586), .Z(n32576) );
  ANDN U34027 ( .A(n32587), .B(n25835), .Z(n32586) );
  XOR U34028 ( .A(n32588), .B(\modmult_1/zin[0][817] ), .Z(n25835) );
  IV U34029 ( .A(n32585), .Z(n32588) );
  XNOR U34030 ( .A(n32585), .B(n25834), .Z(n32587) );
  XOR U34031 ( .A(n32589), .B(n32590), .Z(n25834) );
  AND U34032 ( .A(\modmult_1/xin[1023] ), .B(n32591), .Z(n32590) );
  IV U34033 ( .A(n32589), .Z(n32591) );
  XOR U34034 ( .A(n32592), .B(mreg[818]), .Z(n32589) );
  NAND U34035 ( .A(n32593), .B(mul_pow), .Z(n32592) );
  XOR U34036 ( .A(mreg[818]), .B(creg[818]), .Z(n32593) );
  XOR U34037 ( .A(n32594), .B(n32595), .Z(n32585) );
  ANDN U34038 ( .A(n32596), .B(n25841), .Z(n32595) );
  XOR U34039 ( .A(n32597), .B(\modmult_1/zin[0][816] ), .Z(n25841) );
  IV U34040 ( .A(n32594), .Z(n32597) );
  XNOR U34041 ( .A(n32594), .B(n25840), .Z(n32596) );
  XOR U34042 ( .A(n32598), .B(n32599), .Z(n25840) );
  AND U34043 ( .A(\modmult_1/xin[1023] ), .B(n32600), .Z(n32599) );
  IV U34044 ( .A(n32598), .Z(n32600) );
  XOR U34045 ( .A(n32601), .B(mreg[817]), .Z(n32598) );
  NAND U34046 ( .A(n32602), .B(mul_pow), .Z(n32601) );
  XOR U34047 ( .A(mreg[817]), .B(creg[817]), .Z(n32602) );
  XOR U34048 ( .A(n32603), .B(n32604), .Z(n32594) );
  ANDN U34049 ( .A(n32605), .B(n25847), .Z(n32604) );
  XOR U34050 ( .A(n32606), .B(\modmult_1/zin[0][815] ), .Z(n25847) );
  IV U34051 ( .A(n32603), .Z(n32606) );
  XNOR U34052 ( .A(n32603), .B(n25846), .Z(n32605) );
  XOR U34053 ( .A(n32607), .B(n32608), .Z(n25846) );
  AND U34054 ( .A(\modmult_1/xin[1023] ), .B(n32609), .Z(n32608) );
  IV U34055 ( .A(n32607), .Z(n32609) );
  XOR U34056 ( .A(n32610), .B(mreg[816]), .Z(n32607) );
  NAND U34057 ( .A(n32611), .B(mul_pow), .Z(n32610) );
  XOR U34058 ( .A(mreg[816]), .B(creg[816]), .Z(n32611) );
  XOR U34059 ( .A(n32612), .B(n32613), .Z(n32603) );
  ANDN U34060 ( .A(n32614), .B(n25853), .Z(n32613) );
  XOR U34061 ( .A(n32615), .B(\modmult_1/zin[0][814] ), .Z(n25853) );
  IV U34062 ( .A(n32612), .Z(n32615) );
  XNOR U34063 ( .A(n32612), .B(n25852), .Z(n32614) );
  XOR U34064 ( .A(n32616), .B(n32617), .Z(n25852) );
  AND U34065 ( .A(\modmult_1/xin[1023] ), .B(n32618), .Z(n32617) );
  IV U34066 ( .A(n32616), .Z(n32618) );
  XOR U34067 ( .A(n32619), .B(mreg[815]), .Z(n32616) );
  NAND U34068 ( .A(n32620), .B(mul_pow), .Z(n32619) );
  XOR U34069 ( .A(mreg[815]), .B(creg[815]), .Z(n32620) );
  XOR U34070 ( .A(n32621), .B(n32622), .Z(n32612) );
  ANDN U34071 ( .A(n32623), .B(n25859), .Z(n32622) );
  XOR U34072 ( .A(n32624), .B(\modmult_1/zin[0][813] ), .Z(n25859) );
  IV U34073 ( .A(n32621), .Z(n32624) );
  XNOR U34074 ( .A(n32621), .B(n25858), .Z(n32623) );
  XOR U34075 ( .A(n32625), .B(n32626), .Z(n25858) );
  AND U34076 ( .A(\modmult_1/xin[1023] ), .B(n32627), .Z(n32626) );
  IV U34077 ( .A(n32625), .Z(n32627) );
  XOR U34078 ( .A(n32628), .B(mreg[814]), .Z(n32625) );
  NAND U34079 ( .A(n32629), .B(mul_pow), .Z(n32628) );
  XOR U34080 ( .A(mreg[814]), .B(creg[814]), .Z(n32629) );
  XOR U34081 ( .A(n32630), .B(n32631), .Z(n32621) );
  ANDN U34082 ( .A(n32632), .B(n25865), .Z(n32631) );
  XOR U34083 ( .A(n32633), .B(\modmult_1/zin[0][812] ), .Z(n25865) );
  IV U34084 ( .A(n32630), .Z(n32633) );
  XNOR U34085 ( .A(n32630), .B(n25864), .Z(n32632) );
  XOR U34086 ( .A(n32634), .B(n32635), .Z(n25864) );
  AND U34087 ( .A(\modmult_1/xin[1023] ), .B(n32636), .Z(n32635) );
  IV U34088 ( .A(n32634), .Z(n32636) );
  XOR U34089 ( .A(n32637), .B(mreg[813]), .Z(n32634) );
  NAND U34090 ( .A(n32638), .B(mul_pow), .Z(n32637) );
  XOR U34091 ( .A(mreg[813]), .B(creg[813]), .Z(n32638) );
  XOR U34092 ( .A(n32639), .B(n32640), .Z(n32630) );
  ANDN U34093 ( .A(n32641), .B(n25871), .Z(n32640) );
  XOR U34094 ( .A(n32642), .B(\modmult_1/zin[0][811] ), .Z(n25871) );
  IV U34095 ( .A(n32639), .Z(n32642) );
  XNOR U34096 ( .A(n32639), .B(n25870), .Z(n32641) );
  XOR U34097 ( .A(n32643), .B(n32644), .Z(n25870) );
  AND U34098 ( .A(\modmult_1/xin[1023] ), .B(n32645), .Z(n32644) );
  IV U34099 ( .A(n32643), .Z(n32645) );
  XOR U34100 ( .A(n32646), .B(mreg[812]), .Z(n32643) );
  NAND U34101 ( .A(n32647), .B(mul_pow), .Z(n32646) );
  XOR U34102 ( .A(mreg[812]), .B(creg[812]), .Z(n32647) );
  XOR U34103 ( .A(n32648), .B(n32649), .Z(n32639) );
  ANDN U34104 ( .A(n32650), .B(n25877), .Z(n32649) );
  XOR U34105 ( .A(n32651), .B(\modmult_1/zin[0][810] ), .Z(n25877) );
  IV U34106 ( .A(n32648), .Z(n32651) );
  XNOR U34107 ( .A(n32648), .B(n25876), .Z(n32650) );
  XOR U34108 ( .A(n32652), .B(n32653), .Z(n25876) );
  AND U34109 ( .A(\modmult_1/xin[1023] ), .B(n32654), .Z(n32653) );
  IV U34110 ( .A(n32652), .Z(n32654) );
  XOR U34111 ( .A(n32655), .B(mreg[811]), .Z(n32652) );
  NAND U34112 ( .A(n32656), .B(mul_pow), .Z(n32655) );
  XOR U34113 ( .A(mreg[811]), .B(creg[811]), .Z(n32656) );
  XOR U34114 ( .A(n32657), .B(n32658), .Z(n32648) );
  ANDN U34115 ( .A(n32659), .B(n25883), .Z(n32658) );
  XOR U34116 ( .A(n32660), .B(\modmult_1/zin[0][809] ), .Z(n25883) );
  IV U34117 ( .A(n32657), .Z(n32660) );
  XNOR U34118 ( .A(n32657), .B(n25882), .Z(n32659) );
  XOR U34119 ( .A(n32661), .B(n32662), .Z(n25882) );
  AND U34120 ( .A(\modmult_1/xin[1023] ), .B(n32663), .Z(n32662) );
  IV U34121 ( .A(n32661), .Z(n32663) );
  XOR U34122 ( .A(n32664), .B(mreg[810]), .Z(n32661) );
  NAND U34123 ( .A(n32665), .B(mul_pow), .Z(n32664) );
  XOR U34124 ( .A(mreg[810]), .B(creg[810]), .Z(n32665) );
  XOR U34125 ( .A(n32666), .B(n32667), .Z(n32657) );
  ANDN U34126 ( .A(n32668), .B(n25889), .Z(n32667) );
  XOR U34127 ( .A(n32669), .B(\modmult_1/zin[0][808] ), .Z(n25889) );
  IV U34128 ( .A(n32666), .Z(n32669) );
  XNOR U34129 ( .A(n32666), .B(n25888), .Z(n32668) );
  XOR U34130 ( .A(n32670), .B(n32671), .Z(n25888) );
  AND U34131 ( .A(\modmult_1/xin[1023] ), .B(n32672), .Z(n32671) );
  IV U34132 ( .A(n32670), .Z(n32672) );
  XOR U34133 ( .A(n32673), .B(mreg[809]), .Z(n32670) );
  NAND U34134 ( .A(n32674), .B(mul_pow), .Z(n32673) );
  XOR U34135 ( .A(mreg[809]), .B(creg[809]), .Z(n32674) );
  XOR U34136 ( .A(n32675), .B(n32676), .Z(n32666) );
  ANDN U34137 ( .A(n32677), .B(n25895), .Z(n32676) );
  XOR U34138 ( .A(n32678), .B(\modmult_1/zin[0][807] ), .Z(n25895) );
  IV U34139 ( .A(n32675), .Z(n32678) );
  XNOR U34140 ( .A(n32675), .B(n25894), .Z(n32677) );
  XOR U34141 ( .A(n32679), .B(n32680), .Z(n25894) );
  AND U34142 ( .A(\modmult_1/xin[1023] ), .B(n32681), .Z(n32680) );
  IV U34143 ( .A(n32679), .Z(n32681) );
  XOR U34144 ( .A(n32682), .B(mreg[808]), .Z(n32679) );
  NAND U34145 ( .A(n32683), .B(mul_pow), .Z(n32682) );
  XOR U34146 ( .A(mreg[808]), .B(creg[808]), .Z(n32683) );
  XOR U34147 ( .A(n32684), .B(n32685), .Z(n32675) );
  ANDN U34148 ( .A(n32686), .B(n25901), .Z(n32685) );
  XOR U34149 ( .A(n32687), .B(\modmult_1/zin[0][806] ), .Z(n25901) );
  IV U34150 ( .A(n32684), .Z(n32687) );
  XNOR U34151 ( .A(n32684), .B(n25900), .Z(n32686) );
  XOR U34152 ( .A(n32688), .B(n32689), .Z(n25900) );
  AND U34153 ( .A(\modmult_1/xin[1023] ), .B(n32690), .Z(n32689) );
  IV U34154 ( .A(n32688), .Z(n32690) );
  XOR U34155 ( .A(n32691), .B(mreg[807]), .Z(n32688) );
  NAND U34156 ( .A(n32692), .B(mul_pow), .Z(n32691) );
  XOR U34157 ( .A(mreg[807]), .B(creg[807]), .Z(n32692) );
  XOR U34158 ( .A(n32693), .B(n32694), .Z(n32684) );
  ANDN U34159 ( .A(n32695), .B(n25907), .Z(n32694) );
  XOR U34160 ( .A(n32696), .B(\modmult_1/zin[0][805] ), .Z(n25907) );
  IV U34161 ( .A(n32693), .Z(n32696) );
  XNOR U34162 ( .A(n32693), .B(n25906), .Z(n32695) );
  XOR U34163 ( .A(n32697), .B(n32698), .Z(n25906) );
  AND U34164 ( .A(\modmult_1/xin[1023] ), .B(n32699), .Z(n32698) );
  IV U34165 ( .A(n32697), .Z(n32699) );
  XOR U34166 ( .A(n32700), .B(mreg[806]), .Z(n32697) );
  NAND U34167 ( .A(n32701), .B(mul_pow), .Z(n32700) );
  XOR U34168 ( .A(mreg[806]), .B(creg[806]), .Z(n32701) );
  XOR U34169 ( .A(n32702), .B(n32703), .Z(n32693) );
  ANDN U34170 ( .A(n32704), .B(n25913), .Z(n32703) );
  XOR U34171 ( .A(n32705), .B(\modmult_1/zin[0][804] ), .Z(n25913) );
  IV U34172 ( .A(n32702), .Z(n32705) );
  XNOR U34173 ( .A(n32702), .B(n25912), .Z(n32704) );
  XOR U34174 ( .A(n32706), .B(n32707), .Z(n25912) );
  AND U34175 ( .A(\modmult_1/xin[1023] ), .B(n32708), .Z(n32707) );
  IV U34176 ( .A(n32706), .Z(n32708) );
  XOR U34177 ( .A(n32709), .B(mreg[805]), .Z(n32706) );
  NAND U34178 ( .A(n32710), .B(mul_pow), .Z(n32709) );
  XOR U34179 ( .A(mreg[805]), .B(creg[805]), .Z(n32710) );
  XOR U34180 ( .A(n32711), .B(n32712), .Z(n32702) );
  ANDN U34181 ( .A(n32713), .B(n25919), .Z(n32712) );
  XOR U34182 ( .A(n32714), .B(\modmult_1/zin[0][803] ), .Z(n25919) );
  IV U34183 ( .A(n32711), .Z(n32714) );
  XNOR U34184 ( .A(n32711), .B(n25918), .Z(n32713) );
  XOR U34185 ( .A(n32715), .B(n32716), .Z(n25918) );
  AND U34186 ( .A(\modmult_1/xin[1023] ), .B(n32717), .Z(n32716) );
  IV U34187 ( .A(n32715), .Z(n32717) );
  XOR U34188 ( .A(n32718), .B(mreg[804]), .Z(n32715) );
  NAND U34189 ( .A(n32719), .B(mul_pow), .Z(n32718) );
  XOR U34190 ( .A(mreg[804]), .B(creg[804]), .Z(n32719) );
  XOR U34191 ( .A(n32720), .B(n32721), .Z(n32711) );
  ANDN U34192 ( .A(n32722), .B(n25925), .Z(n32721) );
  XOR U34193 ( .A(n32723), .B(\modmult_1/zin[0][802] ), .Z(n25925) );
  IV U34194 ( .A(n32720), .Z(n32723) );
  XNOR U34195 ( .A(n32720), .B(n25924), .Z(n32722) );
  XOR U34196 ( .A(n32724), .B(n32725), .Z(n25924) );
  AND U34197 ( .A(\modmult_1/xin[1023] ), .B(n32726), .Z(n32725) );
  IV U34198 ( .A(n32724), .Z(n32726) );
  XOR U34199 ( .A(n32727), .B(mreg[803]), .Z(n32724) );
  NAND U34200 ( .A(n32728), .B(mul_pow), .Z(n32727) );
  XOR U34201 ( .A(mreg[803]), .B(creg[803]), .Z(n32728) );
  XOR U34202 ( .A(n32729), .B(n32730), .Z(n32720) );
  ANDN U34203 ( .A(n32731), .B(n25931), .Z(n32730) );
  XOR U34204 ( .A(n32732), .B(\modmult_1/zin[0][801] ), .Z(n25931) );
  IV U34205 ( .A(n32729), .Z(n32732) );
  XNOR U34206 ( .A(n32729), .B(n25930), .Z(n32731) );
  XOR U34207 ( .A(n32733), .B(n32734), .Z(n25930) );
  AND U34208 ( .A(\modmult_1/xin[1023] ), .B(n32735), .Z(n32734) );
  IV U34209 ( .A(n32733), .Z(n32735) );
  XOR U34210 ( .A(n32736), .B(mreg[802]), .Z(n32733) );
  NAND U34211 ( .A(n32737), .B(mul_pow), .Z(n32736) );
  XOR U34212 ( .A(mreg[802]), .B(creg[802]), .Z(n32737) );
  XOR U34213 ( .A(n32738), .B(n32739), .Z(n32729) );
  ANDN U34214 ( .A(n32740), .B(n25937), .Z(n32739) );
  XOR U34215 ( .A(n32741), .B(\modmult_1/zin[0][800] ), .Z(n25937) );
  IV U34216 ( .A(n32738), .Z(n32741) );
  XNOR U34217 ( .A(n32738), .B(n25936), .Z(n32740) );
  XOR U34218 ( .A(n32742), .B(n32743), .Z(n25936) );
  AND U34219 ( .A(\modmult_1/xin[1023] ), .B(n32744), .Z(n32743) );
  IV U34220 ( .A(n32742), .Z(n32744) );
  XOR U34221 ( .A(n32745), .B(mreg[801]), .Z(n32742) );
  NAND U34222 ( .A(n32746), .B(mul_pow), .Z(n32745) );
  XOR U34223 ( .A(mreg[801]), .B(creg[801]), .Z(n32746) );
  XOR U34224 ( .A(n32747), .B(n32748), .Z(n32738) );
  ANDN U34225 ( .A(n32749), .B(n25943), .Z(n32748) );
  XOR U34226 ( .A(n32750), .B(\modmult_1/zin[0][799] ), .Z(n25943) );
  IV U34227 ( .A(n32747), .Z(n32750) );
  XNOR U34228 ( .A(n32747), .B(n25942), .Z(n32749) );
  XOR U34229 ( .A(n32751), .B(n32752), .Z(n25942) );
  AND U34230 ( .A(\modmult_1/xin[1023] ), .B(n32753), .Z(n32752) );
  IV U34231 ( .A(n32751), .Z(n32753) );
  XOR U34232 ( .A(n32754), .B(mreg[800]), .Z(n32751) );
  NAND U34233 ( .A(n32755), .B(mul_pow), .Z(n32754) );
  XOR U34234 ( .A(mreg[800]), .B(creg[800]), .Z(n32755) );
  XOR U34235 ( .A(n32756), .B(n32757), .Z(n32747) );
  ANDN U34236 ( .A(n32758), .B(n25949), .Z(n32757) );
  XOR U34237 ( .A(n32759), .B(\modmult_1/zin[0][798] ), .Z(n25949) );
  IV U34238 ( .A(n32756), .Z(n32759) );
  XNOR U34239 ( .A(n32756), .B(n25948), .Z(n32758) );
  XOR U34240 ( .A(n32760), .B(n32761), .Z(n25948) );
  AND U34241 ( .A(\modmult_1/xin[1023] ), .B(n32762), .Z(n32761) );
  IV U34242 ( .A(n32760), .Z(n32762) );
  XOR U34243 ( .A(n32763), .B(mreg[799]), .Z(n32760) );
  NAND U34244 ( .A(n32764), .B(mul_pow), .Z(n32763) );
  XOR U34245 ( .A(mreg[799]), .B(creg[799]), .Z(n32764) );
  XOR U34246 ( .A(n32765), .B(n32766), .Z(n32756) );
  ANDN U34247 ( .A(n32767), .B(n25955), .Z(n32766) );
  XOR U34248 ( .A(n32768), .B(\modmult_1/zin[0][797] ), .Z(n25955) );
  IV U34249 ( .A(n32765), .Z(n32768) );
  XNOR U34250 ( .A(n32765), .B(n25954), .Z(n32767) );
  XOR U34251 ( .A(n32769), .B(n32770), .Z(n25954) );
  AND U34252 ( .A(\modmult_1/xin[1023] ), .B(n32771), .Z(n32770) );
  IV U34253 ( .A(n32769), .Z(n32771) );
  XOR U34254 ( .A(n32772), .B(mreg[798]), .Z(n32769) );
  NAND U34255 ( .A(n32773), .B(mul_pow), .Z(n32772) );
  XOR U34256 ( .A(mreg[798]), .B(creg[798]), .Z(n32773) );
  XOR U34257 ( .A(n32774), .B(n32775), .Z(n32765) );
  ANDN U34258 ( .A(n32776), .B(n25961), .Z(n32775) );
  XOR U34259 ( .A(n32777), .B(\modmult_1/zin[0][796] ), .Z(n25961) );
  IV U34260 ( .A(n32774), .Z(n32777) );
  XNOR U34261 ( .A(n32774), .B(n25960), .Z(n32776) );
  XOR U34262 ( .A(n32778), .B(n32779), .Z(n25960) );
  AND U34263 ( .A(\modmult_1/xin[1023] ), .B(n32780), .Z(n32779) );
  IV U34264 ( .A(n32778), .Z(n32780) );
  XOR U34265 ( .A(n32781), .B(mreg[797]), .Z(n32778) );
  NAND U34266 ( .A(n32782), .B(mul_pow), .Z(n32781) );
  XOR U34267 ( .A(mreg[797]), .B(creg[797]), .Z(n32782) );
  XOR U34268 ( .A(n32783), .B(n32784), .Z(n32774) );
  ANDN U34269 ( .A(n32785), .B(n25967), .Z(n32784) );
  XOR U34270 ( .A(n32786), .B(\modmult_1/zin[0][795] ), .Z(n25967) );
  IV U34271 ( .A(n32783), .Z(n32786) );
  XNOR U34272 ( .A(n32783), .B(n25966), .Z(n32785) );
  XOR U34273 ( .A(n32787), .B(n32788), .Z(n25966) );
  AND U34274 ( .A(\modmult_1/xin[1023] ), .B(n32789), .Z(n32788) );
  IV U34275 ( .A(n32787), .Z(n32789) );
  XOR U34276 ( .A(n32790), .B(mreg[796]), .Z(n32787) );
  NAND U34277 ( .A(n32791), .B(mul_pow), .Z(n32790) );
  XOR U34278 ( .A(mreg[796]), .B(creg[796]), .Z(n32791) );
  XOR U34279 ( .A(n32792), .B(n32793), .Z(n32783) );
  ANDN U34280 ( .A(n32794), .B(n25973), .Z(n32793) );
  XOR U34281 ( .A(n32795), .B(\modmult_1/zin[0][794] ), .Z(n25973) );
  IV U34282 ( .A(n32792), .Z(n32795) );
  XNOR U34283 ( .A(n32792), .B(n25972), .Z(n32794) );
  XOR U34284 ( .A(n32796), .B(n32797), .Z(n25972) );
  AND U34285 ( .A(\modmult_1/xin[1023] ), .B(n32798), .Z(n32797) );
  IV U34286 ( .A(n32796), .Z(n32798) );
  XOR U34287 ( .A(n32799), .B(mreg[795]), .Z(n32796) );
  NAND U34288 ( .A(n32800), .B(mul_pow), .Z(n32799) );
  XOR U34289 ( .A(mreg[795]), .B(creg[795]), .Z(n32800) );
  XOR U34290 ( .A(n32801), .B(n32802), .Z(n32792) );
  ANDN U34291 ( .A(n32803), .B(n25979), .Z(n32802) );
  XOR U34292 ( .A(n32804), .B(\modmult_1/zin[0][793] ), .Z(n25979) );
  IV U34293 ( .A(n32801), .Z(n32804) );
  XNOR U34294 ( .A(n32801), .B(n25978), .Z(n32803) );
  XOR U34295 ( .A(n32805), .B(n32806), .Z(n25978) );
  AND U34296 ( .A(\modmult_1/xin[1023] ), .B(n32807), .Z(n32806) );
  IV U34297 ( .A(n32805), .Z(n32807) );
  XOR U34298 ( .A(n32808), .B(mreg[794]), .Z(n32805) );
  NAND U34299 ( .A(n32809), .B(mul_pow), .Z(n32808) );
  XOR U34300 ( .A(mreg[794]), .B(creg[794]), .Z(n32809) );
  XOR U34301 ( .A(n32810), .B(n32811), .Z(n32801) );
  ANDN U34302 ( .A(n32812), .B(n25985), .Z(n32811) );
  XOR U34303 ( .A(n32813), .B(\modmult_1/zin[0][792] ), .Z(n25985) );
  IV U34304 ( .A(n32810), .Z(n32813) );
  XNOR U34305 ( .A(n32810), .B(n25984), .Z(n32812) );
  XOR U34306 ( .A(n32814), .B(n32815), .Z(n25984) );
  AND U34307 ( .A(\modmult_1/xin[1023] ), .B(n32816), .Z(n32815) );
  IV U34308 ( .A(n32814), .Z(n32816) );
  XOR U34309 ( .A(n32817), .B(mreg[793]), .Z(n32814) );
  NAND U34310 ( .A(n32818), .B(mul_pow), .Z(n32817) );
  XOR U34311 ( .A(mreg[793]), .B(creg[793]), .Z(n32818) );
  XOR U34312 ( .A(n32819), .B(n32820), .Z(n32810) );
  ANDN U34313 ( .A(n32821), .B(n25991), .Z(n32820) );
  XOR U34314 ( .A(n32822), .B(\modmult_1/zin[0][791] ), .Z(n25991) );
  IV U34315 ( .A(n32819), .Z(n32822) );
  XNOR U34316 ( .A(n32819), .B(n25990), .Z(n32821) );
  XOR U34317 ( .A(n32823), .B(n32824), .Z(n25990) );
  AND U34318 ( .A(\modmult_1/xin[1023] ), .B(n32825), .Z(n32824) );
  IV U34319 ( .A(n32823), .Z(n32825) );
  XOR U34320 ( .A(n32826), .B(mreg[792]), .Z(n32823) );
  NAND U34321 ( .A(n32827), .B(mul_pow), .Z(n32826) );
  XOR U34322 ( .A(mreg[792]), .B(creg[792]), .Z(n32827) );
  XOR U34323 ( .A(n32828), .B(n32829), .Z(n32819) );
  ANDN U34324 ( .A(n32830), .B(n25997), .Z(n32829) );
  XOR U34325 ( .A(n32831), .B(\modmult_1/zin[0][790] ), .Z(n25997) );
  IV U34326 ( .A(n32828), .Z(n32831) );
  XNOR U34327 ( .A(n32828), .B(n25996), .Z(n32830) );
  XOR U34328 ( .A(n32832), .B(n32833), .Z(n25996) );
  AND U34329 ( .A(\modmult_1/xin[1023] ), .B(n32834), .Z(n32833) );
  IV U34330 ( .A(n32832), .Z(n32834) );
  XOR U34331 ( .A(n32835), .B(mreg[791]), .Z(n32832) );
  NAND U34332 ( .A(n32836), .B(mul_pow), .Z(n32835) );
  XOR U34333 ( .A(mreg[791]), .B(creg[791]), .Z(n32836) );
  XOR U34334 ( .A(n32837), .B(n32838), .Z(n32828) );
  ANDN U34335 ( .A(n32839), .B(n26003), .Z(n32838) );
  XOR U34336 ( .A(n32840), .B(\modmult_1/zin[0][789] ), .Z(n26003) );
  IV U34337 ( .A(n32837), .Z(n32840) );
  XNOR U34338 ( .A(n32837), .B(n26002), .Z(n32839) );
  XOR U34339 ( .A(n32841), .B(n32842), .Z(n26002) );
  AND U34340 ( .A(\modmult_1/xin[1023] ), .B(n32843), .Z(n32842) );
  IV U34341 ( .A(n32841), .Z(n32843) );
  XOR U34342 ( .A(n32844), .B(mreg[790]), .Z(n32841) );
  NAND U34343 ( .A(n32845), .B(mul_pow), .Z(n32844) );
  XOR U34344 ( .A(mreg[790]), .B(creg[790]), .Z(n32845) );
  XOR U34345 ( .A(n32846), .B(n32847), .Z(n32837) );
  ANDN U34346 ( .A(n32848), .B(n26009), .Z(n32847) );
  XOR U34347 ( .A(n32849), .B(\modmult_1/zin[0][788] ), .Z(n26009) );
  IV U34348 ( .A(n32846), .Z(n32849) );
  XNOR U34349 ( .A(n32846), .B(n26008), .Z(n32848) );
  XOR U34350 ( .A(n32850), .B(n32851), .Z(n26008) );
  AND U34351 ( .A(\modmult_1/xin[1023] ), .B(n32852), .Z(n32851) );
  IV U34352 ( .A(n32850), .Z(n32852) );
  XOR U34353 ( .A(n32853), .B(mreg[789]), .Z(n32850) );
  NAND U34354 ( .A(n32854), .B(mul_pow), .Z(n32853) );
  XOR U34355 ( .A(mreg[789]), .B(creg[789]), .Z(n32854) );
  XOR U34356 ( .A(n32855), .B(n32856), .Z(n32846) );
  ANDN U34357 ( .A(n32857), .B(n26015), .Z(n32856) );
  XOR U34358 ( .A(n32858), .B(\modmult_1/zin[0][787] ), .Z(n26015) );
  IV U34359 ( .A(n32855), .Z(n32858) );
  XNOR U34360 ( .A(n32855), .B(n26014), .Z(n32857) );
  XOR U34361 ( .A(n32859), .B(n32860), .Z(n26014) );
  AND U34362 ( .A(\modmult_1/xin[1023] ), .B(n32861), .Z(n32860) );
  IV U34363 ( .A(n32859), .Z(n32861) );
  XOR U34364 ( .A(n32862), .B(mreg[788]), .Z(n32859) );
  NAND U34365 ( .A(n32863), .B(mul_pow), .Z(n32862) );
  XOR U34366 ( .A(mreg[788]), .B(creg[788]), .Z(n32863) );
  XOR U34367 ( .A(n32864), .B(n32865), .Z(n32855) );
  ANDN U34368 ( .A(n32866), .B(n26021), .Z(n32865) );
  XOR U34369 ( .A(n32867), .B(\modmult_1/zin[0][786] ), .Z(n26021) );
  IV U34370 ( .A(n32864), .Z(n32867) );
  XNOR U34371 ( .A(n32864), .B(n26020), .Z(n32866) );
  XOR U34372 ( .A(n32868), .B(n32869), .Z(n26020) );
  AND U34373 ( .A(\modmult_1/xin[1023] ), .B(n32870), .Z(n32869) );
  IV U34374 ( .A(n32868), .Z(n32870) );
  XOR U34375 ( .A(n32871), .B(mreg[787]), .Z(n32868) );
  NAND U34376 ( .A(n32872), .B(mul_pow), .Z(n32871) );
  XOR U34377 ( .A(mreg[787]), .B(creg[787]), .Z(n32872) );
  XOR U34378 ( .A(n32873), .B(n32874), .Z(n32864) );
  ANDN U34379 ( .A(n32875), .B(n26027), .Z(n32874) );
  XOR U34380 ( .A(n32876), .B(\modmult_1/zin[0][785] ), .Z(n26027) );
  IV U34381 ( .A(n32873), .Z(n32876) );
  XNOR U34382 ( .A(n32873), .B(n26026), .Z(n32875) );
  XOR U34383 ( .A(n32877), .B(n32878), .Z(n26026) );
  AND U34384 ( .A(\modmult_1/xin[1023] ), .B(n32879), .Z(n32878) );
  IV U34385 ( .A(n32877), .Z(n32879) );
  XOR U34386 ( .A(n32880), .B(mreg[786]), .Z(n32877) );
  NAND U34387 ( .A(n32881), .B(mul_pow), .Z(n32880) );
  XOR U34388 ( .A(mreg[786]), .B(creg[786]), .Z(n32881) );
  XOR U34389 ( .A(n32882), .B(n32883), .Z(n32873) );
  ANDN U34390 ( .A(n32884), .B(n26033), .Z(n32883) );
  XOR U34391 ( .A(n32885), .B(\modmult_1/zin[0][784] ), .Z(n26033) );
  IV U34392 ( .A(n32882), .Z(n32885) );
  XNOR U34393 ( .A(n32882), .B(n26032), .Z(n32884) );
  XOR U34394 ( .A(n32886), .B(n32887), .Z(n26032) );
  AND U34395 ( .A(\modmult_1/xin[1023] ), .B(n32888), .Z(n32887) );
  IV U34396 ( .A(n32886), .Z(n32888) );
  XOR U34397 ( .A(n32889), .B(mreg[785]), .Z(n32886) );
  NAND U34398 ( .A(n32890), .B(mul_pow), .Z(n32889) );
  XOR U34399 ( .A(mreg[785]), .B(creg[785]), .Z(n32890) );
  XOR U34400 ( .A(n32891), .B(n32892), .Z(n32882) );
  ANDN U34401 ( .A(n32893), .B(n26039), .Z(n32892) );
  XOR U34402 ( .A(n32894), .B(\modmult_1/zin[0][783] ), .Z(n26039) );
  IV U34403 ( .A(n32891), .Z(n32894) );
  XNOR U34404 ( .A(n32891), .B(n26038), .Z(n32893) );
  XOR U34405 ( .A(n32895), .B(n32896), .Z(n26038) );
  AND U34406 ( .A(\modmult_1/xin[1023] ), .B(n32897), .Z(n32896) );
  IV U34407 ( .A(n32895), .Z(n32897) );
  XOR U34408 ( .A(n32898), .B(mreg[784]), .Z(n32895) );
  NAND U34409 ( .A(n32899), .B(mul_pow), .Z(n32898) );
  XOR U34410 ( .A(mreg[784]), .B(creg[784]), .Z(n32899) );
  XOR U34411 ( .A(n32900), .B(n32901), .Z(n32891) );
  ANDN U34412 ( .A(n32902), .B(n26045), .Z(n32901) );
  XOR U34413 ( .A(n32903), .B(\modmult_1/zin[0][782] ), .Z(n26045) );
  IV U34414 ( .A(n32900), .Z(n32903) );
  XNOR U34415 ( .A(n32900), .B(n26044), .Z(n32902) );
  XOR U34416 ( .A(n32904), .B(n32905), .Z(n26044) );
  AND U34417 ( .A(\modmult_1/xin[1023] ), .B(n32906), .Z(n32905) );
  IV U34418 ( .A(n32904), .Z(n32906) );
  XOR U34419 ( .A(n32907), .B(mreg[783]), .Z(n32904) );
  NAND U34420 ( .A(n32908), .B(mul_pow), .Z(n32907) );
  XOR U34421 ( .A(mreg[783]), .B(creg[783]), .Z(n32908) );
  XOR U34422 ( .A(n32909), .B(n32910), .Z(n32900) );
  ANDN U34423 ( .A(n32911), .B(n26051), .Z(n32910) );
  XOR U34424 ( .A(n32912), .B(\modmult_1/zin[0][781] ), .Z(n26051) );
  IV U34425 ( .A(n32909), .Z(n32912) );
  XNOR U34426 ( .A(n32909), .B(n26050), .Z(n32911) );
  XOR U34427 ( .A(n32913), .B(n32914), .Z(n26050) );
  AND U34428 ( .A(\modmult_1/xin[1023] ), .B(n32915), .Z(n32914) );
  IV U34429 ( .A(n32913), .Z(n32915) );
  XOR U34430 ( .A(n32916), .B(mreg[782]), .Z(n32913) );
  NAND U34431 ( .A(n32917), .B(mul_pow), .Z(n32916) );
  XOR U34432 ( .A(mreg[782]), .B(creg[782]), .Z(n32917) );
  XOR U34433 ( .A(n32918), .B(n32919), .Z(n32909) );
  ANDN U34434 ( .A(n32920), .B(n26057), .Z(n32919) );
  XOR U34435 ( .A(n32921), .B(\modmult_1/zin[0][780] ), .Z(n26057) );
  IV U34436 ( .A(n32918), .Z(n32921) );
  XNOR U34437 ( .A(n32918), .B(n26056), .Z(n32920) );
  XOR U34438 ( .A(n32922), .B(n32923), .Z(n26056) );
  AND U34439 ( .A(\modmult_1/xin[1023] ), .B(n32924), .Z(n32923) );
  IV U34440 ( .A(n32922), .Z(n32924) );
  XOR U34441 ( .A(n32925), .B(mreg[781]), .Z(n32922) );
  NAND U34442 ( .A(n32926), .B(mul_pow), .Z(n32925) );
  XOR U34443 ( .A(mreg[781]), .B(creg[781]), .Z(n32926) );
  XOR U34444 ( .A(n32927), .B(n32928), .Z(n32918) );
  ANDN U34445 ( .A(n32929), .B(n26063), .Z(n32928) );
  XOR U34446 ( .A(n32930), .B(\modmult_1/zin[0][779] ), .Z(n26063) );
  IV U34447 ( .A(n32927), .Z(n32930) );
  XNOR U34448 ( .A(n32927), .B(n26062), .Z(n32929) );
  XOR U34449 ( .A(n32931), .B(n32932), .Z(n26062) );
  AND U34450 ( .A(\modmult_1/xin[1023] ), .B(n32933), .Z(n32932) );
  IV U34451 ( .A(n32931), .Z(n32933) );
  XOR U34452 ( .A(n32934), .B(mreg[780]), .Z(n32931) );
  NAND U34453 ( .A(n32935), .B(mul_pow), .Z(n32934) );
  XOR U34454 ( .A(mreg[780]), .B(creg[780]), .Z(n32935) );
  XOR U34455 ( .A(n32936), .B(n32937), .Z(n32927) );
  ANDN U34456 ( .A(n32938), .B(n26069), .Z(n32937) );
  XOR U34457 ( .A(n32939), .B(\modmult_1/zin[0][778] ), .Z(n26069) );
  IV U34458 ( .A(n32936), .Z(n32939) );
  XNOR U34459 ( .A(n32936), .B(n26068), .Z(n32938) );
  XOR U34460 ( .A(n32940), .B(n32941), .Z(n26068) );
  AND U34461 ( .A(\modmult_1/xin[1023] ), .B(n32942), .Z(n32941) );
  IV U34462 ( .A(n32940), .Z(n32942) );
  XOR U34463 ( .A(n32943), .B(mreg[779]), .Z(n32940) );
  NAND U34464 ( .A(n32944), .B(mul_pow), .Z(n32943) );
  XOR U34465 ( .A(mreg[779]), .B(creg[779]), .Z(n32944) );
  XOR U34466 ( .A(n32945), .B(n32946), .Z(n32936) );
  ANDN U34467 ( .A(n32947), .B(n26075), .Z(n32946) );
  XOR U34468 ( .A(n32948), .B(\modmult_1/zin[0][777] ), .Z(n26075) );
  IV U34469 ( .A(n32945), .Z(n32948) );
  XNOR U34470 ( .A(n32945), .B(n26074), .Z(n32947) );
  XOR U34471 ( .A(n32949), .B(n32950), .Z(n26074) );
  AND U34472 ( .A(\modmult_1/xin[1023] ), .B(n32951), .Z(n32950) );
  IV U34473 ( .A(n32949), .Z(n32951) );
  XOR U34474 ( .A(n32952), .B(mreg[778]), .Z(n32949) );
  NAND U34475 ( .A(n32953), .B(mul_pow), .Z(n32952) );
  XOR U34476 ( .A(mreg[778]), .B(creg[778]), .Z(n32953) );
  XOR U34477 ( .A(n32954), .B(n32955), .Z(n32945) );
  ANDN U34478 ( .A(n32956), .B(n26081), .Z(n32955) );
  XOR U34479 ( .A(n32957), .B(\modmult_1/zin[0][776] ), .Z(n26081) );
  IV U34480 ( .A(n32954), .Z(n32957) );
  XNOR U34481 ( .A(n32954), .B(n26080), .Z(n32956) );
  XOR U34482 ( .A(n32958), .B(n32959), .Z(n26080) );
  AND U34483 ( .A(\modmult_1/xin[1023] ), .B(n32960), .Z(n32959) );
  IV U34484 ( .A(n32958), .Z(n32960) );
  XOR U34485 ( .A(n32961), .B(mreg[777]), .Z(n32958) );
  NAND U34486 ( .A(n32962), .B(mul_pow), .Z(n32961) );
  XOR U34487 ( .A(mreg[777]), .B(creg[777]), .Z(n32962) );
  XOR U34488 ( .A(n32963), .B(n32964), .Z(n32954) );
  ANDN U34489 ( .A(n32965), .B(n26087), .Z(n32964) );
  XOR U34490 ( .A(n32966), .B(\modmult_1/zin[0][775] ), .Z(n26087) );
  IV U34491 ( .A(n32963), .Z(n32966) );
  XNOR U34492 ( .A(n32963), .B(n26086), .Z(n32965) );
  XOR U34493 ( .A(n32967), .B(n32968), .Z(n26086) );
  AND U34494 ( .A(\modmult_1/xin[1023] ), .B(n32969), .Z(n32968) );
  IV U34495 ( .A(n32967), .Z(n32969) );
  XOR U34496 ( .A(n32970), .B(mreg[776]), .Z(n32967) );
  NAND U34497 ( .A(n32971), .B(mul_pow), .Z(n32970) );
  XOR U34498 ( .A(mreg[776]), .B(creg[776]), .Z(n32971) );
  XOR U34499 ( .A(n32972), .B(n32973), .Z(n32963) );
  ANDN U34500 ( .A(n32974), .B(n26093), .Z(n32973) );
  XOR U34501 ( .A(n32975), .B(\modmult_1/zin[0][774] ), .Z(n26093) );
  IV U34502 ( .A(n32972), .Z(n32975) );
  XNOR U34503 ( .A(n32972), .B(n26092), .Z(n32974) );
  XOR U34504 ( .A(n32976), .B(n32977), .Z(n26092) );
  AND U34505 ( .A(\modmult_1/xin[1023] ), .B(n32978), .Z(n32977) );
  IV U34506 ( .A(n32976), .Z(n32978) );
  XOR U34507 ( .A(n32979), .B(mreg[775]), .Z(n32976) );
  NAND U34508 ( .A(n32980), .B(mul_pow), .Z(n32979) );
  XOR U34509 ( .A(mreg[775]), .B(creg[775]), .Z(n32980) );
  XOR U34510 ( .A(n32981), .B(n32982), .Z(n32972) );
  ANDN U34511 ( .A(n32983), .B(n26099), .Z(n32982) );
  XOR U34512 ( .A(n32984), .B(\modmult_1/zin[0][773] ), .Z(n26099) );
  IV U34513 ( .A(n32981), .Z(n32984) );
  XNOR U34514 ( .A(n32981), .B(n26098), .Z(n32983) );
  XOR U34515 ( .A(n32985), .B(n32986), .Z(n26098) );
  AND U34516 ( .A(\modmult_1/xin[1023] ), .B(n32987), .Z(n32986) );
  IV U34517 ( .A(n32985), .Z(n32987) );
  XOR U34518 ( .A(n32988), .B(mreg[774]), .Z(n32985) );
  NAND U34519 ( .A(n32989), .B(mul_pow), .Z(n32988) );
  XOR U34520 ( .A(mreg[774]), .B(creg[774]), .Z(n32989) );
  XOR U34521 ( .A(n32990), .B(n32991), .Z(n32981) );
  ANDN U34522 ( .A(n32992), .B(n26105), .Z(n32991) );
  XOR U34523 ( .A(n32993), .B(\modmult_1/zin[0][772] ), .Z(n26105) );
  IV U34524 ( .A(n32990), .Z(n32993) );
  XNOR U34525 ( .A(n32990), .B(n26104), .Z(n32992) );
  XOR U34526 ( .A(n32994), .B(n32995), .Z(n26104) );
  AND U34527 ( .A(\modmult_1/xin[1023] ), .B(n32996), .Z(n32995) );
  IV U34528 ( .A(n32994), .Z(n32996) );
  XOR U34529 ( .A(n32997), .B(mreg[773]), .Z(n32994) );
  NAND U34530 ( .A(n32998), .B(mul_pow), .Z(n32997) );
  XOR U34531 ( .A(mreg[773]), .B(creg[773]), .Z(n32998) );
  XOR U34532 ( .A(n32999), .B(n33000), .Z(n32990) );
  ANDN U34533 ( .A(n33001), .B(n26111), .Z(n33000) );
  XOR U34534 ( .A(n33002), .B(\modmult_1/zin[0][771] ), .Z(n26111) );
  IV U34535 ( .A(n32999), .Z(n33002) );
  XNOR U34536 ( .A(n32999), .B(n26110), .Z(n33001) );
  XOR U34537 ( .A(n33003), .B(n33004), .Z(n26110) );
  AND U34538 ( .A(\modmult_1/xin[1023] ), .B(n33005), .Z(n33004) );
  IV U34539 ( .A(n33003), .Z(n33005) );
  XOR U34540 ( .A(n33006), .B(mreg[772]), .Z(n33003) );
  NAND U34541 ( .A(n33007), .B(mul_pow), .Z(n33006) );
  XOR U34542 ( .A(mreg[772]), .B(creg[772]), .Z(n33007) );
  XOR U34543 ( .A(n33008), .B(n33009), .Z(n32999) );
  ANDN U34544 ( .A(n33010), .B(n26117), .Z(n33009) );
  XOR U34545 ( .A(n33011), .B(\modmult_1/zin[0][770] ), .Z(n26117) );
  IV U34546 ( .A(n33008), .Z(n33011) );
  XNOR U34547 ( .A(n33008), .B(n26116), .Z(n33010) );
  XOR U34548 ( .A(n33012), .B(n33013), .Z(n26116) );
  AND U34549 ( .A(\modmult_1/xin[1023] ), .B(n33014), .Z(n33013) );
  IV U34550 ( .A(n33012), .Z(n33014) );
  XOR U34551 ( .A(n33015), .B(mreg[771]), .Z(n33012) );
  NAND U34552 ( .A(n33016), .B(mul_pow), .Z(n33015) );
  XOR U34553 ( .A(mreg[771]), .B(creg[771]), .Z(n33016) );
  XOR U34554 ( .A(n33017), .B(n33018), .Z(n33008) );
  ANDN U34555 ( .A(n33019), .B(n26123), .Z(n33018) );
  XOR U34556 ( .A(n33020), .B(\modmult_1/zin[0][769] ), .Z(n26123) );
  IV U34557 ( .A(n33017), .Z(n33020) );
  XNOR U34558 ( .A(n33017), .B(n26122), .Z(n33019) );
  XOR U34559 ( .A(n33021), .B(n33022), .Z(n26122) );
  AND U34560 ( .A(\modmult_1/xin[1023] ), .B(n33023), .Z(n33022) );
  IV U34561 ( .A(n33021), .Z(n33023) );
  XOR U34562 ( .A(n33024), .B(mreg[770]), .Z(n33021) );
  NAND U34563 ( .A(n33025), .B(mul_pow), .Z(n33024) );
  XOR U34564 ( .A(mreg[770]), .B(creg[770]), .Z(n33025) );
  XOR U34565 ( .A(n33026), .B(n33027), .Z(n33017) );
  ANDN U34566 ( .A(n33028), .B(n26129), .Z(n33027) );
  XOR U34567 ( .A(n33029), .B(\modmult_1/zin[0][768] ), .Z(n26129) );
  IV U34568 ( .A(n33026), .Z(n33029) );
  XNOR U34569 ( .A(n33026), .B(n26128), .Z(n33028) );
  XOR U34570 ( .A(n33030), .B(n33031), .Z(n26128) );
  AND U34571 ( .A(\modmult_1/xin[1023] ), .B(n33032), .Z(n33031) );
  IV U34572 ( .A(n33030), .Z(n33032) );
  XOR U34573 ( .A(n33033), .B(mreg[769]), .Z(n33030) );
  NAND U34574 ( .A(n33034), .B(mul_pow), .Z(n33033) );
  XOR U34575 ( .A(mreg[769]), .B(creg[769]), .Z(n33034) );
  XOR U34576 ( .A(n33035), .B(n33036), .Z(n33026) );
  ANDN U34577 ( .A(n33037), .B(n26135), .Z(n33036) );
  XOR U34578 ( .A(n33038), .B(\modmult_1/zin[0][767] ), .Z(n26135) );
  IV U34579 ( .A(n33035), .Z(n33038) );
  XNOR U34580 ( .A(n33035), .B(n26134), .Z(n33037) );
  XOR U34581 ( .A(n33039), .B(n33040), .Z(n26134) );
  AND U34582 ( .A(\modmult_1/xin[1023] ), .B(n33041), .Z(n33040) );
  IV U34583 ( .A(n33039), .Z(n33041) );
  XOR U34584 ( .A(n33042), .B(mreg[768]), .Z(n33039) );
  NAND U34585 ( .A(n33043), .B(mul_pow), .Z(n33042) );
  XOR U34586 ( .A(mreg[768]), .B(creg[768]), .Z(n33043) );
  XOR U34587 ( .A(n33044), .B(n33045), .Z(n33035) );
  ANDN U34588 ( .A(n33046), .B(n26141), .Z(n33045) );
  XOR U34589 ( .A(n33047), .B(\modmult_1/zin[0][766] ), .Z(n26141) );
  IV U34590 ( .A(n33044), .Z(n33047) );
  XNOR U34591 ( .A(n33044), .B(n26140), .Z(n33046) );
  XOR U34592 ( .A(n33048), .B(n33049), .Z(n26140) );
  AND U34593 ( .A(\modmult_1/xin[1023] ), .B(n33050), .Z(n33049) );
  IV U34594 ( .A(n33048), .Z(n33050) );
  XOR U34595 ( .A(n33051), .B(mreg[767]), .Z(n33048) );
  NAND U34596 ( .A(n33052), .B(mul_pow), .Z(n33051) );
  XOR U34597 ( .A(mreg[767]), .B(creg[767]), .Z(n33052) );
  XOR U34598 ( .A(n33053), .B(n33054), .Z(n33044) );
  ANDN U34599 ( .A(n33055), .B(n26147), .Z(n33054) );
  XOR U34600 ( .A(n33056), .B(\modmult_1/zin[0][765] ), .Z(n26147) );
  IV U34601 ( .A(n33053), .Z(n33056) );
  XNOR U34602 ( .A(n33053), .B(n26146), .Z(n33055) );
  XOR U34603 ( .A(n33057), .B(n33058), .Z(n26146) );
  AND U34604 ( .A(\modmult_1/xin[1023] ), .B(n33059), .Z(n33058) );
  IV U34605 ( .A(n33057), .Z(n33059) );
  XOR U34606 ( .A(n33060), .B(mreg[766]), .Z(n33057) );
  NAND U34607 ( .A(n33061), .B(mul_pow), .Z(n33060) );
  XOR U34608 ( .A(mreg[766]), .B(creg[766]), .Z(n33061) );
  XOR U34609 ( .A(n33062), .B(n33063), .Z(n33053) );
  ANDN U34610 ( .A(n33064), .B(n26153), .Z(n33063) );
  XOR U34611 ( .A(n33065), .B(\modmult_1/zin[0][764] ), .Z(n26153) );
  IV U34612 ( .A(n33062), .Z(n33065) );
  XNOR U34613 ( .A(n33062), .B(n26152), .Z(n33064) );
  XOR U34614 ( .A(n33066), .B(n33067), .Z(n26152) );
  AND U34615 ( .A(\modmult_1/xin[1023] ), .B(n33068), .Z(n33067) );
  IV U34616 ( .A(n33066), .Z(n33068) );
  XOR U34617 ( .A(n33069), .B(mreg[765]), .Z(n33066) );
  NAND U34618 ( .A(n33070), .B(mul_pow), .Z(n33069) );
  XOR U34619 ( .A(mreg[765]), .B(creg[765]), .Z(n33070) );
  XOR U34620 ( .A(n33071), .B(n33072), .Z(n33062) );
  ANDN U34621 ( .A(n33073), .B(n26159), .Z(n33072) );
  XOR U34622 ( .A(n33074), .B(\modmult_1/zin[0][763] ), .Z(n26159) );
  IV U34623 ( .A(n33071), .Z(n33074) );
  XNOR U34624 ( .A(n33071), .B(n26158), .Z(n33073) );
  XOR U34625 ( .A(n33075), .B(n33076), .Z(n26158) );
  AND U34626 ( .A(\modmult_1/xin[1023] ), .B(n33077), .Z(n33076) );
  IV U34627 ( .A(n33075), .Z(n33077) );
  XOR U34628 ( .A(n33078), .B(mreg[764]), .Z(n33075) );
  NAND U34629 ( .A(n33079), .B(mul_pow), .Z(n33078) );
  XOR U34630 ( .A(mreg[764]), .B(creg[764]), .Z(n33079) );
  XOR U34631 ( .A(n33080), .B(n33081), .Z(n33071) );
  ANDN U34632 ( .A(n33082), .B(n26165), .Z(n33081) );
  XOR U34633 ( .A(n33083), .B(\modmult_1/zin[0][762] ), .Z(n26165) );
  IV U34634 ( .A(n33080), .Z(n33083) );
  XNOR U34635 ( .A(n33080), .B(n26164), .Z(n33082) );
  XOR U34636 ( .A(n33084), .B(n33085), .Z(n26164) );
  AND U34637 ( .A(\modmult_1/xin[1023] ), .B(n33086), .Z(n33085) );
  IV U34638 ( .A(n33084), .Z(n33086) );
  XOR U34639 ( .A(n33087), .B(mreg[763]), .Z(n33084) );
  NAND U34640 ( .A(n33088), .B(mul_pow), .Z(n33087) );
  XOR U34641 ( .A(mreg[763]), .B(creg[763]), .Z(n33088) );
  XOR U34642 ( .A(n33089), .B(n33090), .Z(n33080) );
  ANDN U34643 ( .A(n33091), .B(n26171), .Z(n33090) );
  XOR U34644 ( .A(n33092), .B(\modmult_1/zin[0][761] ), .Z(n26171) );
  IV U34645 ( .A(n33089), .Z(n33092) );
  XNOR U34646 ( .A(n33089), .B(n26170), .Z(n33091) );
  XOR U34647 ( .A(n33093), .B(n33094), .Z(n26170) );
  AND U34648 ( .A(\modmult_1/xin[1023] ), .B(n33095), .Z(n33094) );
  IV U34649 ( .A(n33093), .Z(n33095) );
  XOR U34650 ( .A(n33096), .B(mreg[762]), .Z(n33093) );
  NAND U34651 ( .A(n33097), .B(mul_pow), .Z(n33096) );
  XOR U34652 ( .A(mreg[762]), .B(creg[762]), .Z(n33097) );
  XOR U34653 ( .A(n33098), .B(n33099), .Z(n33089) );
  ANDN U34654 ( .A(n33100), .B(n26177), .Z(n33099) );
  XOR U34655 ( .A(n33101), .B(\modmult_1/zin[0][760] ), .Z(n26177) );
  IV U34656 ( .A(n33098), .Z(n33101) );
  XNOR U34657 ( .A(n33098), .B(n26176), .Z(n33100) );
  XOR U34658 ( .A(n33102), .B(n33103), .Z(n26176) );
  AND U34659 ( .A(\modmult_1/xin[1023] ), .B(n33104), .Z(n33103) );
  IV U34660 ( .A(n33102), .Z(n33104) );
  XOR U34661 ( .A(n33105), .B(mreg[761]), .Z(n33102) );
  NAND U34662 ( .A(n33106), .B(mul_pow), .Z(n33105) );
  XOR U34663 ( .A(mreg[761]), .B(creg[761]), .Z(n33106) );
  XOR U34664 ( .A(n33107), .B(n33108), .Z(n33098) );
  ANDN U34665 ( .A(n33109), .B(n26183), .Z(n33108) );
  XOR U34666 ( .A(n33110), .B(\modmult_1/zin[0][759] ), .Z(n26183) );
  IV U34667 ( .A(n33107), .Z(n33110) );
  XNOR U34668 ( .A(n33107), .B(n26182), .Z(n33109) );
  XOR U34669 ( .A(n33111), .B(n33112), .Z(n26182) );
  AND U34670 ( .A(\modmult_1/xin[1023] ), .B(n33113), .Z(n33112) );
  IV U34671 ( .A(n33111), .Z(n33113) );
  XOR U34672 ( .A(n33114), .B(mreg[760]), .Z(n33111) );
  NAND U34673 ( .A(n33115), .B(mul_pow), .Z(n33114) );
  XOR U34674 ( .A(mreg[760]), .B(creg[760]), .Z(n33115) );
  XOR U34675 ( .A(n33116), .B(n33117), .Z(n33107) );
  ANDN U34676 ( .A(n33118), .B(n26189), .Z(n33117) );
  XOR U34677 ( .A(n33119), .B(\modmult_1/zin[0][758] ), .Z(n26189) );
  IV U34678 ( .A(n33116), .Z(n33119) );
  XNOR U34679 ( .A(n33116), .B(n26188), .Z(n33118) );
  XOR U34680 ( .A(n33120), .B(n33121), .Z(n26188) );
  AND U34681 ( .A(\modmult_1/xin[1023] ), .B(n33122), .Z(n33121) );
  IV U34682 ( .A(n33120), .Z(n33122) );
  XOR U34683 ( .A(n33123), .B(mreg[759]), .Z(n33120) );
  NAND U34684 ( .A(n33124), .B(mul_pow), .Z(n33123) );
  XOR U34685 ( .A(mreg[759]), .B(creg[759]), .Z(n33124) );
  XOR U34686 ( .A(n33125), .B(n33126), .Z(n33116) );
  ANDN U34687 ( .A(n33127), .B(n26195), .Z(n33126) );
  XOR U34688 ( .A(n33128), .B(\modmult_1/zin[0][757] ), .Z(n26195) );
  IV U34689 ( .A(n33125), .Z(n33128) );
  XNOR U34690 ( .A(n33125), .B(n26194), .Z(n33127) );
  XOR U34691 ( .A(n33129), .B(n33130), .Z(n26194) );
  AND U34692 ( .A(\modmult_1/xin[1023] ), .B(n33131), .Z(n33130) );
  IV U34693 ( .A(n33129), .Z(n33131) );
  XOR U34694 ( .A(n33132), .B(mreg[758]), .Z(n33129) );
  NAND U34695 ( .A(n33133), .B(mul_pow), .Z(n33132) );
  XOR U34696 ( .A(mreg[758]), .B(creg[758]), .Z(n33133) );
  XOR U34697 ( .A(n33134), .B(n33135), .Z(n33125) );
  ANDN U34698 ( .A(n33136), .B(n26201), .Z(n33135) );
  XOR U34699 ( .A(n33137), .B(\modmult_1/zin[0][756] ), .Z(n26201) );
  IV U34700 ( .A(n33134), .Z(n33137) );
  XNOR U34701 ( .A(n33134), .B(n26200), .Z(n33136) );
  XOR U34702 ( .A(n33138), .B(n33139), .Z(n26200) );
  AND U34703 ( .A(\modmult_1/xin[1023] ), .B(n33140), .Z(n33139) );
  IV U34704 ( .A(n33138), .Z(n33140) );
  XOR U34705 ( .A(n33141), .B(mreg[757]), .Z(n33138) );
  NAND U34706 ( .A(n33142), .B(mul_pow), .Z(n33141) );
  XOR U34707 ( .A(mreg[757]), .B(creg[757]), .Z(n33142) );
  XOR U34708 ( .A(n33143), .B(n33144), .Z(n33134) );
  ANDN U34709 ( .A(n33145), .B(n26207), .Z(n33144) );
  XOR U34710 ( .A(n33146), .B(\modmult_1/zin[0][755] ), .Z(n26207) );
  IV U34711 ( .A(n33143), .Z(n33146) );
  XNOR U34712 ( .A(n33143), .B(n26206), .Z(n33145) );
  XOR U34713 ( .A(n33147), .B(n33148), .Z(n26206) );
  AND U34714 ( .A(\modmult_1/xin[1023] ), .B(n33149), .Z(n33148) );
  IV U34715 ( .A(n33147), .Z(n33149) );
  XOR U34716 ( .A(n33150), .B(mreg[756]), .Z(n33147) );
  NAND U34717 ( .A(n33151), .B(mul_pow), .Z(n33150) );
  XOR U34718 ( .A(mreg[756]), .B(creg[756]), .Z(n33151) );
  XOR U34719 ( .A(n33152), .B(n33153), .Z(n33143) );
  ANDN U34720 ( .A(n33154), .B(n26213), .Z(n33153) );
  XOR U34721 ( .A(n33155), .B(\modmult_1/zin[0][754] ), .Z(n26213) );
  IV U34722 ( .A(n33152), .Z(n33155) );
  XNOR U34723 ( .A(n33152), .B(n26212), .Z(n33154) );
  XOR U34724 ( .A(n33156), .B(n33157), .Z(n26212) );
  AND U34725 ( .A(\modmult_1/xin[1023] ), .B(n33158), .Z(n33157) );
  IV U34726 ( .A(n33156), .Z(n33158) );
  XOR U34727 ( .A(n33159), .B(mreg[755]), .Z(n33156) );
  NAND U34728 ( .A(n33160), .B(mul_pow), .Z(n33159) );
  XOR U34729 ( .A(mreg[755]), .B(creg[755]), .Z(n33160) );
  XOR U34730 ( .A(n33161), .B(n33162), .Z(n33152) );
  ANDN U34731 ( .A(n33163), .B(n26219), .Z(n33162) );
  XOR U34732 ( .A(n33164), .B(\modmult_1/zin[0][753] ), .Z(n26219) );
  IV U34733 ( .A(n33161), .Z(n33164) );
  XNOR U34734 ( .A(n33161), .B(n26218), .Z(n33163) );
  XOR U34735 ( .A(n33165), .B(n33166), .Z(n26218) );
  AND U34736 ( .A(\modmult_1/xin[1023] ), .B(n33167), .Z(n33166) );
  IV U34737 ( .A(n33165), .Z(n33167) );
  XOR U34738 ( .A(n33168), .B(mreg[754]), .Z(n33165) );
  NAND U34739 ( .A(n33169), .B(mul_pow), .Z(n33168) );
  XOR U34740 ( .A(mreg[754]), .B(creg[754]), .Z(n33169) );
  XOR U34741 ( .A(n33170), .B(n33171), .Z(n33161) );
  ANDN U34742 ( .A(n33172), .B(n26225), .Z(n33171) );
  XOR U34743 ( .A(n33173), .B(\modmult_1/zin[0][752] ), .Z(n26225) );
  IV U34744 ( .A(n33170), .Z(n33173) );
  XNOR U34745 ( .A(n33170), .B(n26224), .Z(n33172) );
  XOR U34746 ( .A(n33174), .B(n33175), .Z(n26224) );
  AND U34747 ( .A(\modmult_1/xin[1023] ), .B(n33176), .Z(n33175) );
  IV U34748 ( .A(n33174), .Z(n33176) );
  XOR U34749 ( .A(n33177), .B(mreg[753]), .Z(n33174) );
  NAND U34750 ( .A(n33178), .B(mul_pow), .Z(n33177) );
  XOR U34751 ( .A(mreg[753]), .B(creg[753]), .Z(n33178) );
  XOR U34752 ( .A(n33179), .B(n33180), .Z(n33170) );
  ANDN U34753 ( .A(n33181), .B(n26231), .Z(n33180) );
  XOR U34754 ( .A(n33182), .B(\modmult_1/zin[0][751] ), .Z(n26231) );
  IV U34755 ( .A(n33179), .Z(n33182) );
  XNOR U34756 ( .A(n33179), .B(n26230), .Z(n33181) );
  XOR U34757 ( .A(n33183), .B(n33184), .Z(n26230) );
  AND U34758 ( .A(\modmult_1/xin[1023] ), .B(n33185), .Z(n33184) );
  IV U34759 ( .A(n33183), .Z(n33185) );
  XOR U34760 ( .A(n33186), .B(mreg[752]), .Z(n33183) );
  NAND U34761 ( .A(n33187), .B(mul_pow), .Z(n33186) );
  XOR U34762 ( .A(mreg[752]), .B(creg[752]), .Z(n33187) );
  XOR U34763 ( .A(n33188), .B(n33189), .Z(n33179) );
  ANDN U34764 ( .A(n33190), .B(n26237), .Z(n33189) );
  XOR U34765 ( .A(n33191), .B(\modmult_1/zin[0][750] ), .Z(n26237) );
  IV U34766 ( .A(n33188), .Z(n33191) );
  XNOR U34767 ( .A(n33188), .B(n26236), .Z(n33190) );
  XOR U34768 ( .A(n33192), .B(n33193), .Z(n26236) );
  AND U34769 ( .A(\modmult_1/xin[1023] ), .B(n33194), .Z(n33193) );
  IV U34770 ( .A(n33192), .Z(n33194) );
  XOR U34771 ( .A(n33195), .B(mreg[751]), .Z(n33192) );
  NAND U34772 ( .A(n33196), .B(mul_pow), .Z(n33195) );
  XOR U34773 ( .A(mreg[751]), .B(creg[751]), .Z(n33196) );
  XOR U34774 ( .A(n33197), .B(n33198), .Z(n33188) );
  ANDN U34775 ( .A(n33199), .B(n26243), .Z(n33198) );
  XOR U34776 ( .A(n33200), .B(\modmult_1/zin[0][749] ), .Z(n26243) );
  IV U34777 ( .A(n33197), .Z(n33200) );
  XNOR U34778 ( .A(n33197), .B(n26242), .Z(n33199) );
  XOR U34779 ( .A(n33201), .B(n33202), .Z(n26242) );
  AND U34780 ( .A(\modmult_1/xin[1023] ), .B(n33203), .Z(n33202) );
  IV U34781 ( .A(n33201), .Z(n33203) );
  XOR U34782 ( .A(n33204), .B(mreg[750]), .Z(n33201) );
  NAND U34783 ( .A(n33205), .B(mul_pow), .Z(n33204) );
  XOR U34784 ( .A(mreg[750]), .B(creg[750]), .Z(n33205) );
  XOR U34785 ( .A(n33206), .B(n33207), .Z(n33197) );
  ANDN U34786 ( .A(n33208), .B(n26249), .Z(n33207) );
  XOR U34787 ( .A(n33209), .B(\modmult_1/zin[0][748] ), .Z(n26249) );
  IV U34788 ( .A(n33206), .Z(n33209) );
  XNOR U34789 ( .A(n33206), .B(n26248), .Z(n33208) );
  XOR U34790 ( .A(n33210), .B(n33211), .Z(n26248) );
  AND U34791 ( .A(\modmult_1/xin[1023] ), .B(n33212), .Z(n33211) );
  IV U34792 ( .A(n33210), .Z(n33212) );
  XOR U34793 ( .A(n33213), .B(mreg[749]), .Z(n33210) );
  NAND U34794 ( .A(n33214), .B(mul_pow), .Z(n33213) );
  XOR U34795 ( .A(mreg[749]), .B(creg[749]), .Z(n33214) );
  XOR U34796 ( .A(n33215), .B(n33216), .Z(n33206) );
  ANDN U34797 ( .A(n33217), .B(n26255), .Z(n33216) );
  XOR U34798 ( .A(n33218), .B(\modmult_1/zin[0][747] ), .Z(n26255) );
  IV U34799 ( .A(n33215), .Z(n33218) );
  XNOR U34800 ( .A(n33215), .B(n26254), .Z(n33217) );
  XOR U34801 ( .A(n33219), .B(n33220), .Z(n26254) );
  AND U34802 ( .A(\modmult_1/xin[1023] ), .B(n33221), .Z(n33220) );
  IV U34803 ( .A(n33219), .Z(n33221) );
  XOR U34804 ( .A(n33222), .B(mreg[748]), .Z(n33219) );
  NAND U34805 ( .A(n33223), .B(mul_pow), .Z(n33222) );
  XOR U34806 ( .A(mreg[748]), .B(creg[748]), .Z(n33223) );
  XOR U34807 ( .A(n33224), .B(n33225), .Z(n33215) );
  ANDN U34808 ( .A(n33226), .B(n26261), .Z(n33225) );
  XOR U34809 ( .A(n33227), .B(\modmult_1/zin[0][746] ), .Z(n26261) );
  IV U34810 ( .A(n33224), .Z(n33227) );
  XNOR U34811 ( .A(n33224), .B(n26260), .Z(n33226) );
  XOR U34812 ( .A(n33228), .B(n33229), .Z(n26260) );
  AND U34813 ( .A(\modmult_1/xin[1023] ), .B(n33230), .Z(n33229) );
  IV U34814 ( .A(n33228), .Z(n33230) );
  XOR U34815 ( .A(n33231), .B(mreg[747]), .Z(n33228) );
  NAND U34816 ( .A(n33232), .B(mul_pow), .Z(n33231) );
  XOR U34817 ( .A(mreg[747]), .B(creg[747]), .Z(n33232) );
  XOR U34818 ( .A(n33233), .B(n33234), .Z(n33224) );
  ANDN U34819 ( .A(n33235), .B(n26267), .Z(n33234) );
  XOR U34820 ( .A(n33236), .B(\modmult_1/zin[0][745] ), .Z(n26267) );
  IV U34821 ( .A(n33233), .Z(n33236) );
  XNOR U34822 ( .A(n33233), .B(n26266), .Z(n33235) );
  XOR U34823 ( .A(n33237), .B(n33238), .Z(n26266) );
  AND U34824 ( .A(\modmult_1/xin[1023] ), .B(n33239), .Z(n33238) );
  IV U34825 ( .A(n33237), .Z(n33239) );
  XOR U34826 ( .A(n33240), .B(mreg[746]), .Z(n33237) );
  NAND U34827 ( .A(n33241), .B(mul_pow), .Z(n33240) );
  XOR U34828 ( .A(mreg[746]), .B(creg[746]), .Z(n33241) );
  XOR U34829 ( .A(n33242), .B(n33243), .Z(n33233) );
  ANDN U34830 ( .A(n33244), .B(n26273), .Z(n33243) );
  XOR U34831 ( .A(n33245), .B(\modmult_1/zin[0][744] ), .Z(n26273) );
  IV U34832 ( .A(n33242), .Z(n33245) );
  XNOR U34833 ( .A(n33242), .B(n26272), .Z(n33244) );
  XOR U34834 ( .A(n33246), .B(n33247), .Z(n26272) );
  AND U34835 ( .A(\modmult_1/xin[1023] ), .B(n33248), .Z(n33247) );
  IV U34836 ( .A(n33246), .Z(n33248) );
  XOR U34837 ( .A(n33249), .B(mreg[745]), .Z(n33246) );
  NAND U34838 ( .A(n33250), .B(mul_pow), .Z(n33249) );
  XOR U34839 ( .A(mreg[745]), .B(creg[745]), .Z(n33250) );
  XOR U34840 ( .A(n33251), .B(n33252), .Z(n33242) );
  ANDN U34841 ( .A(n33253), .B(n26279), .Z(n33252) );
  XOR U34842 ( .A(n33254), .B(\modmult_1/zin[0][743] ), .Z(n26279) );
  IV U34843 ( .A(n33251), .Z(n33254) );
  XNOR U34844 ( .A(n33251), .B(n26278), .Z(n33253) );
  XOR U34845 ( .A(n33255), .B(n33256), .Z(n26278) );
  AND U34846 ( .A(\modmult_1/xin[1023] ), .B(n33257), .Z(n33256) );
  IV U34847 ( .A(n33255), .Z(n33257) );
  XOR U34848 ( .A(n33258), .B(mreg[744]), .Z(n33255) );
  NAND U34849 ( .A(n33259), .B(mul_pow), .Z(n33258) );
  XOR U34850 ( .A(mreg[744]), .B(creg[744]), .Z(n33259) );
  XOR U34851 ( .A(n33260), .B(n33261), .Z(n33251) );
  ANDN U34852 ( .A(n33262), .B(n26285), .Z(n33261) );
  XOR U34853 ( .A(n33263), .B(\modmult_1/zin[0][742] ), .Z(n26285) );
  IV U34854 ( .A(n33260), .Z(n33263) );
  XNOR U34855 ( .A(n33260), .B(n26284), .Z(n33262) );
  XOR U34856 ( .A(n33264), .B(n33265), .Z(n26284) );
  AND U34857 ( .A(\modmult_1/xin[1023] ), .B(n33266), .Z(n33265) );
  IV U34858 ( .A(n33264), .Z(n33266) );
  XOR U34859 ( .A(n33267), .B(mreg[743]), .Z(n33264) );
  NAND U34860 ( .A(n33268), .B(mul_pow), .Z(n33267) );
  XOR U34861 ( .A(mreg[743]), .B(creg[743]), .Z(n33268) );
  XOR U34862 ( .A(n33269), .B(n33270), .Z(n33260) );
  ANDN U34863 ( .A(n33271), .B(n26291), .Z(n33270) );
  XOR U34864 ( .A(n33272), .B(\modmult_1/zin[0][741] ), .Z(n26291) );
  IV U34865 ( .A(n33269), .Z(n33272) );
  XNOR U34866 ( .A(n33269), .B(n26290), .Z(n33271) );
  XOR U34867 ( .A(n33273), .B(n33274), .Z(n26290) );
  AND U34868 ( .A(\modmult_1/xin[1023] ), .B(n33275), .Z(n33274) );
  IV U34869 ( .A(n33273), .Z(n33275) );
  XOR U34870 ( .A(n33276), .B(mreg[742]), .Z(n33273) );
  NAND U34871 ( .A(n33277), .B(mul_pow), .Z(n33276) );
  XOR U34872 ( .A(mreg[742]), .B(creg[742]), .Z(n33277) );
  XOR U34873 ( .A(n33278), .B(n33279), .Z(n33269) );
  ANDN U34874 ( .A(n33280), .B(n26297), .Z(n33279) );
  XOR U34875 ( .A(n33281), .B(\modmult_1/zin[0][740] ), .Z(n26297) );
  IV U34876 ( .A(n33278), .Z(n33281) );
  XNOR U34877 ( .A(n33278), .B(n26296), .Z(n33280) );
  XOR U34878 ( .A(n33282), .B(n33283), .Z(n26296) );
  AND U34879 ( .A(\modmult_1/xin[1023] ), .B(n33284), .Z(n33283) );
  IV U34880 ( .A(n33282), .Z(n33284) );
  XOR U34881 ( .A(n33285), .B(mreg[741]), .Z(n33282) );
  NAND U34882 ( .A(n33286), .B(mul_pow), .Z(n33285) );
  XOR U34883 ( .A(mreg[741]), .B(creg[741]), .Z(n33286) );
  XOR U34884 ( .A(n33287), .B(n33288), .Z(n33278) );
  ANDN U34885 ( .A(n33289), .B(n26303), .Z(n33288) );
  XOR U34886 ( .A(n33290), .B(\modmult_1/zin[0][739] ), .Z(n26303) );
  IV U34887 ( .A(n33287), .Z(n33290) );
  XNOR U34888 ( .A(n33287), .B(n26302), .Z(n33289) );
  XOR U34889 ( .A(n33291), .B(n33292), .Z(n26302) );
  AND U34890 ( .A(\modmult_1/xin[1023] ), .B(n33293), .Z(n33292) );
  IV U34891 ( .A(n33291), .Z(n33293) );
  XOR U34892 ( .A(n33294), .B(mreg[740]), .Z(n33291) );
  NAND U34893 ( .A(n33295), .B(mul_pow), .Z(n33294) );
  XOR U34894 ( .A(mreg[740]), .B(creg[740]), .Z(n33295) );
  XOR U34895 ( .A(n33296), .B(n33297), .Z(n33287) );
  ANDN U34896 ( .A(n33298), .B(n26309), .Z(n33297) );
  XOR U34897 ( .A(n33299), .B(\modmult_1/zin[0][738] ), .Z(n26309) );
  IV U34898 ( .A(n33296), .Z(n33299) );
  XNOR U34899 ( .A(n33296), .B(n26308), .Z(n33298) );
  XOR U34900 ( .A(n33300), .B(n33301), .Z(n26308) );
  AND U34901 ( .A(\modmult_1/xin[1023] ), .B(n33302), .Z(n33301) );
  IV U34902 ( .A(n33300), .Z(n33302) );
  XOR U34903 ( .A(n33303), .B(mreg[739]), .Z(n33300) );
  NAND U34904 ( .A(n33304), .B(mul_pow), .Z(n33303) );
  XOR U34905 ( .A(mreg[739]), .B(creg[739]), .Z(n33304) );
  XOR U34906 ( .A(n33305), .B(n33306), .Z(n33296) );
  ANDN U34907 ( .A(n33307), .B(n26315), .Z(n33306) );
  XOR U34908 ( .A(n33308), .B(\modmult_1/zin[0][737] ), .Z(n26315) );
  IV U34909 ( .A(n33305), .Z(n33308) );
  XNOR U34910 ( .A(n33305), .B(n26314), .Z(n33307) );
  XOR U34911 ( .A(n33309), .B(n33310), .Z(n26314) );
  AND U34912 ( .A(\modmult_1/xin[1023] ), .B(n33311), .Z(n33310) );
  IV U34913 ( .A(n33309), .Z(n33311) );
  XOR U34914 ( .A(n33312), .B(mreg[738]), .Z(n33309) );
  NAND U34915 ( .A(n33313), .B(mul_pow), .Z(n33312) );
  XOR U34916 ( .A(mreg[738]), .B(creg[738]), .Z(n33313) );
  XOR U34917 ( .A(n33314), .B(n33315), .Z(n33305) );
  ANDN U34918 ( .A(n33316), .B(n26321), .Z(n33315) );
  XOR U34919 ( .A(n33317), .B(\modmult_1/zin[0][736] ), .Z(n26321) );
  IV U34920 ( .A(n33314), .Z(n33317) );
  XNOR U34921 ( .A(n33314), .B(n26320), .Z(n33316) );
  XOR U34922 ( .A(n33318), .B(n33319), .Z(n26320) );
  AND U34923 ( .A(\modmult_1/xin[1023] ), .B(n33320), .Z(n33319) );
  IV U34924 ( .A(n33318), .Z(n33320) );
  XOR U34925 ( .A(n33321), .B(mreg[737]), .Z(n33318) );
  NAND U34926 ( .A(n33322), .B(mul_pow), .Z(n33321) );
  XOR U34927 ( .A(mreg[737]), .B(creg[737]), .Z(n33322) );
  XOR U34928 ( .A(n33323), .B(n33324), .Z(n33314) );
  ANDN U34929 ( .A(n33325), .B(n26327), .Z(n33324) );
  XOR U34930 ( .A(n33326), .B(\modmult_1/zin[0][735] ), .Z(n26327) );
  IV U34931 ( .A(n33323), .Z(n33326) );
  XNOR U34932 ( .A(n33323), .B(n26326), .Z(n33325) );
  XOR U34933 ( .A(n33327), .B(n33328), .Z(n26326) );
  AND U34934 ( .A(\modmult_1/xin[1023] ), .B(n33329), .Z(n33328) );
  IV U34935 ( .A(n33327), .Z(n33329) );
  XOR U34936 ( .A(n33330), .B(mreg[736]), .Z(n33327) );
  NAND U34937 ( .A(n33331), .B(mul_pow), .Z(n33330) );
  XOR U34938 ( .A(mreg[736]), .B(creg[736]), .Z(n33331) );
  XOR U34939 ( .A(n33332), .B(n33333), .Z(n33323) );
  ANDN U34940 ( .A(n33334), .B(n26333), .Z(n33333) );
  XOR U34941 ( .A(n33335), .B(\modmult_1/zin[0][734] ), .Z(n26333) );
  IV U34942 ( .A(n33332), .Z(n33335) );
  XNOR U34943 ( .A(n33332), .B(n26332), .Z(n33334) );
  XOR U34944 ( .A(n33336), .B(n33337), .Z(n26332) );
  AND U34945 ( .A(\modmult_1/xin[1023] ), .B(n33338), .Z(n33337) );
  IV U34946 ( .A(n33336), .Z(n33338) );
  XOR U34947 ( .A(n33339), .B(mreg[735]), .Z(n33336) );
  NAND U34948 ( .A(n33340), .B(mul_pow), .Z(n33339) );
  XOR U34949 ( .A(mreg[735]), .B(creg[735]), .Z(n33340) );
  XOR U34950 ( .A(n33341), .B(n33342), .Z(n33332) );
  ANDN U34951 ( .A(n33343), .B(n26339), .Z(n33342) );
  XOR U34952 ( .A(n33344), .B(\modmult_1/zin[0][733] ), .Z(n26339) );
  IV U34953 ( .A(n33341), .Z(n33344) );
  XNOR U34954 ( .A(n33341), .B(n26338), .Z(n33343) );
  XOR U34955 ( .A(n33345), .B(n33346), .Z(n26338) );
  AND U34956 ( .A(\modmult_1/xin[1023] ), .B(n33347), .Z(n33346) );
  IV U34957 ( .A(n33345), .Z(n33347) );
  XOR U34958 ( .A(n33348), .B(mreg[734]), .Z(n33345) );
  NAND U34959 ( .A(n33349), .B(mul_pow), .Z(n33348) );
  XOR U34960 ( .A(mreg[734]), .B(creg[734]), .Z(n33349) );
  XOR U34961 ( .A(n33350), .B(n33351), .Z(n33341) );
  ANDN U34962 ( .A(n33352), .B(n26345), .Z(n33351) );
  XOR U34963 ( .A(n33353), .B(\modmult_1/zin[0][732] ), .Z(n26345) );
  IV U34964 ( .A(n33350), .Z(n33353) );
  XNOR U34965 ( .A(n33350), .B(n26344), .Z(n33352) );
  XOR U34966 ( .A(n33354), .B(n33355), .Z(n26344) );
  AND U34967 ( .A(\modmult_1/xin[1023] ), .B(n33356), .Z(n33355) );
  IV U34968 ( .A(n33354), .Z(n33356) );
  XOR U34969 ( .A(n33357), .B(mreg[733]), .Z(n33354) );
  NAND U34970 ( .A(n33358), .B(mul_pow), .Z(n33357) );
  XOR U34971 ( .A(mreg[733]), .B(creg[733]), .Z(n33358) );
  XOR U34972 ( .A(n33359), .B(n33360), .Z(n33350) );
  ANDN U34973 ( .A(n33361), .B(n26351), .Z(n33360) );
  XOR U34974 ( .A(n33362), .B(\modmult_1/zin[0][731] ), .Z(n26351) );
  IV U34975 ( .A(n33359), .Z(n33362) );
  XNOR U34976 ( .A(n33359), .B(n26350), .Z(n33361) );
  XOR U34977 ( .A(n33363), .B(n33364), .Z(n26350) );
  AND U34978 ( .A(\modmult_1/xin[1023] ), .B(n33365), .Z(n33364) );
  IV U34979 ( .A(n33363), .Z(n33365) );
  XOR U34980 ( .A(n33366), .B(mreg[732]), .Z(n33363) );
  NAND U34981 ( .A(n33367), .B(mul_pow), .Z(n33366) );
  XOR U34982 ( .A(mreg[732]), .B(creg[732]), .Z(n33367) );
  XOR U34983 ( .A(n33368), .B(n33369), .Z(n33359) );
  ANDN U34984 ( .A(n33370), .B(n26357), .Z(n33369) );
  XOR U34985 ( .A(n33371), .B(\modmult_1/zin[0][730] ), .Z(n26357) );
  IV U34986 ( .A(n33368), .Z(n33371) );
  XNOR U34987 ( .A(n33368), .B(n26356), .Z(n33370) );
  XOR U34988 ( .A(n33372), .B(n33373), .Z(n26356) );
  AND U34989 ( .A(\modmult_1/xin[1023] ), .B(n33374), .Z(n33373) );
  IV U34990 ( .A(n33372), .Z(n33374) );
  XOR U34991 ( .A(n33375), .B(mreg[731]), .Z(n33372) );
  NAND U34992 ( .A(n33376), .B(mul_pow), .Z(n33375) );
  XOR U34993 ( .A(mreg[731]), .B(creg[731]), .Z(n33376) );
  XOR U34994 ( .A(n33377), .B(n33378), .Z(n33368) );
  ANDN U34995 ( .A(n33379), .B(n26363), .Z(n33378) );
  XOR U34996 ( .A(n33380), .B(\modmult_1/zin[0][729] ), .Z(n26363) );
  IV U34997 ( .A(n33377), .Z(n33380) );
  XNOR U34998 ( .A(n33377), .B(n26362), .Z(n33379) );
  XOR U34999 ( .A(n33381), .B(n33382), .Z(n26362) );
  AND U35000 ( .A(\modmult_1/xin[1023] ), .B(n33383), .Z(n33382) );
  IV U35001 ( .A(n33381), .Z(n33383) );
  XOR U35002 ( .A(n33384), .B(mreg[730]), .Z(n33381) );
  NAND U35003 ( .A(n33385), .B(mul_pow), .Z(n33384) );
  XOR U35004 ( .A(mreg[730]), .B(creg[730]), .Z(n33385) );
  XOR U35005 ( .A(n33386), .B(n33387), .Z(n33377) );
  ANDN U35006 ( .A(n33388), .B(n26369), .Z(n33387) );
  XOR U35007 ( .A(n33389), .B(\modmult_1/zin[0][728] ), .Z(n26369) );
  IV U35008 ( .A(n33386), .Z(n33389) );
  XNOR U35009 ( .A(n33386), .B(n26368), .Z(n33388) );
  XOR U35010 ( .A(n33390), .B(n33391), .Z(n26368) );
  AND U35011 ( .A(\modmult_1/xin[1023] ), .B(n33392), .Z(n33391) );
  IV U35012 ( .A(n33390), .Z(n33392) );
  XOR U35013 ( .A(n33393), .B(mreg[729]), .Z(n33390) );
  NAND U35014 ( .A(n33394), .B(mul_pow), .Z(n33393) );
  XOR U35015 ( .A(mreg[729]), .B(creg[729]), .Z(n33394) );
  XOR U35016 ( .A(n33395), .B(n33396), .Z(n33386) );
  ANDN U35017 ( .A(n33397), .B(n26375), .Z(n33396) );
  XOR U35018 ( .A(n33398), .B(\modmult_1/zin[0][727] ), .Z(n26375) );
  IV U35019 ( .A(n33395), .Z(n33398) );
  XNOR U35020 ( .A(n33395), .B(n26374), .Z(n33397) );
  XOR U35021 ( .A(n33399), .B(n33400), .Z(n26374) );
  AND U35022 ( .A(\modmult_1/xin[1023] ), .B(n33401), .Z(n33400) );
  IV U35023 ( .A(n33399), .Z(n33401) );
  XOR U35024 ( .A(n33402), .B(mreg[728]), .Z(n33399) );
  NAND U35025 ( .A(n33403), .B(mul_pow), .Z(n33402) );
  XOR U35026 ( .A(mreg[728]), .B(creg[728]), .Z(n33403) );
  XOR U35027 ( .A(n33404), .B(n33405), .Z(n33395) );
  ANDN U35028 ( .A(n33406), .B(n26381), .Z(n33405) );
  XOR U35029 ( .A(n33407), .B(\modmult_1/zin[0][726] ), .Z(n26381) );
  IV U35030 ( .A(n33404), .Z(n33407) );
  XNOR U35031 ( .A(n33404), .B(n26380), .Z(n33406) );
  XOR U35032 ( .A(n33408), .B(n33409), .Z(n26380) );
  AND U35033 ( .A(\modmult_1/xin[1023] ), .B(n33410), .Z(n33409) );
  IV U35034 ( .A(n33408), .Z(n33410) );
  XOR U35035 ( .A(n33411), .B(mreg[727]), .Z(n33408) );
  NAND U35036 ( .A(n33412), .B(mul_pow), .Z(n33411) );
  XOR U35037 ( .A(mreg[727]), .B(creg[727]), .Z(n33412) );
  XOR U35038 ( .A(n33413), .B(n33414), .Z(n33404) );
  ANDN U35039 ( .A(n33415), .B(n26387), .Z(n33414) );
  XOR U35040 ( .A(n33416), .B(\modmult_1/zin[0][725] ), .Z(n26387) );
  IV U35041 ( .A(n33413), .Z(n33416) );
  XNOR U35042 ( .A(n33413), .B(n26386), .Z(n33415) );
  XOR U35043 ( .A(n33417), .B(n33418), .Z(n26386) );
  AND U35044 ( .A(\modmult_1/xin[1023] ), .B(n33419), .Z(n33418) );
  IV U35045 ( .A(n33417), .Z(n33419) );
  XOR U35046 ( .A(n33420), .B(mreg[726]), .Z(n33417) );
  NAND U35047 ( .A(n33421), .B(mul_pow), .Z(n33420) );
  XOR U35048 ( .A(mreg[726]), .B(creg[726]), .Z(n33421) );
  XOR U35049 ( .A(n33422), .B(n33423), .Z(n33413) );
  ANDN U35050 ( .A(n33424), .B(n26393), .Z(n33423) );
  XOR U35051 ( .A(n33425), .B(\modmult_1/zin[0][724] ), .Z(n26393) );
  IV U35052 ( .A(n33422), .Z(n33425) );
  XNOR U35053 ( .A(n33422), .B(n26392), .Z(n33424) );
  XOR U35054 ( .A(n33426), .B(n33427), .Z(n26392) );
  AND U35055 ( .A(\modmult_1/xin[1023] ), .B(n33428), .Z(n33427) );
  IV U35056 ( .A(n33426), .Z(n33428) );
  XOR U35057 ( .A(n33429), .B(mreg[725]), .Z(n33426) );
  NAND U35058 ( .A(n33430), .B(mul_pow), .Z(n33429) );
  XOR U35059 ( .A(mreg[725]), .B(creg[725]), .Z(n33430) );
  XOR U35060 ( .A(n33431), .B(n33432), .Z(n33422) );
  ANDN U35061 ( .A(n33433), .B(n26399), .Z(n33432) );
  XOR U35062 ( .A(n33434), .B(\modmult_1/zin[0][723] ), .Z(n26399) );
  IV U35063 ( .A(n33431), .Z(n33434) );
  XNOR U35064 ( .A(n33431), .B(n26398), .Z(n33433) );
  XOR U35065 ( .A(n33435), .B(n33436), .Z(n26398) );
  AND U35066 ( .A(\modmult_1/xin[1023] ), .B(n33437), .Z(n33436) );
  IV U35067 ( .A(n33435), .Z(n33437) );
  XOR U35068 ( .A(n33438), .B(mreg[724]), .Z(n33435) );
  NAND U35069 ( .A(n33439), .B(mul_pow), .Z(n33438) );
  XOR U35070 ( .A(mreg[724]), .B(creg[724]), .Z(n33439) );
  XOR U35071 ( .A(n33440), .B(n33441), .Z(n33431) );
  ANDN U35072 ( .A(n33442), .B(n26405), .Z(n33441) );
  XOR U35073 ( .A(n33443), .B(\modmult_1/zin[0][722] ), .Z(n26405) );
  IV U35074 ( .A(n33440), .Z(n33443) );
  XNOR U35075 ( .A(n33440), .B(n26404), .Z(n33442) );
  XOR U35076 ( .A(n33444), .B(n33445), .Z(n26404) );
  AND U35077 ( .A(\modmult_1/xin[1023] ), .B(n33446), .Z(n33445) );
  IV U35078 ( .A(n33444), .Z(n33446) );
  XOR U35079 ( .A(n33447), .B(mreg[723]), .Z(n33444) );
  NAND U35080 ( .A(n33448), .B(mul_pow), .Z(n33447) );
  XOR U35081 ( .A(mreg[723]), .B(creg[723]), .Z(n33448) );
  XOR U35082 ( .A(n33449), .B(n33450), .Z(n33440) );
  ANDN U35083 ( .A(n33451), .B(n26411), .Z(n33450) );
  XOR U35084 ( .A(n33452), .B(\modmult_1/zin[0][721] ), .Z(n26411) );
  IV U35085 ( .A(n33449), .Z(n33452) );
  XNOR U35086 ( .A(n33449), .B(n26410), .Z(n33451) );
  XOR U35087 ( .A(n33453), .B(n33454), .Z(n26410) );
  AND U35088 ( .A(\modmult_1/xin[1023] ), .B(n33455), .Z(n33454) );
  IV U35089 ( .A(n33453), .Z(n33455) );
  XOR U35090 ( .A(n33456), .B(mreg[722]), .Z(n33453) );
  NAND U35091 ( .A(n33457), .B(mul_pow), .Z(n33456) );
  XOR U35092 ( .A(mreg[722]), .B(creg[722]), .Z(n33457) );
  XOR U35093 ( .A(n33458), .B(n33459), .Z(n33449) );
  ANDN U35094 ( .A(n33460), .B(n26417), .Z(n33459) );
  XOR U35095 ( .A(n33461), .B(\modmult_1/zin[0][720] ), .Z(n26417) );
  IV U35096 ( .A(n33458), .Z(n33461) );
  XNOR U35097 ( .A(n33458), .B(n26416), .Z(n33460) );
  XOR U35098 ( .A(n33462), .B(n33463), .Z(n26416) );
  AND U35099 ( .A(\modmult_1/xin[1023] ), .B(n33464), .Z(n33463) );
  IV U35100 ( .A(n33462), .Z(n33464) );
  XOR U35101 ( .A(n33465), .B(mreg[721]), .Z(n33462) );
  NAND U35102 ( .A(n33466), .B(mul_pow), .Z(n33465) );
  XOR U35103 ( .A(mreg[721]), .B(creg[721]), .Z(n33466) );
  XOR U35104 ( .A(n33467), .B(n33468), .Z(n33458) );
  ANDN U35105 ( .A(n33469), .B(n26423), .Z(n33468) );
  XOR U35106 ( .A(n33470), .B(\modmult_1/zin[0][719] ), .Z(n26423) );
  IV U35107 ( .A(n33467), .Z(n33470) );
  XNOR U35108 ( .A(n33467), .B(n26422), .Z(n33469) );
  XOR U35109 ( .A(n33471), .B(n33472), .Z(n26422) );
  AND U35110 ( .A(\modmult_1/xin[1023] ), .B(n33473), .Z(n33472) );
  IV U35111 ( .A(n33471), .Z(n33473) );
  XOR U35112 ( .A(n33474), .B(mreg[720]), .Z(n33471) );
  NAND U35113 ( .A(n33475), .B(mul_pow), .Z(n33474) );
  XOR U35114 ( .A(mreg[720]), .B(creg[720]), .Z(n33475) );
  XOR U35115 ( .A(n33476), .B(n33477), .Z(n33467) );
  ANDN U35116 ( .A(n33478), .B(n26429), .Z(n33477) );
  XOR U35117 ( .A(n33479), .B(\modmult_1/zin[0][718] ), .Z(n26429) );
  IV U35118 ( .A(n33476), .Z(n33479) );
  XNOR U35119 ( .A(n33476), .B(n26428), .Z(n33478) );
  XOR U35120 ( .A(n33480), .B(n33481), .Z(n26428) );
  AND U35121 ( .A(\modmult_1/xin[1023] ), .B(n33482), .Z(n33481) );
  IV U35122 ( .A(n33480), .Z(n33482) );
  XOR U35123 ( .A(n33483), .B(mreg[719]), .Z(n33480) );
  NAND U35124 ( .A(n33484), .B(mul_pow), .Z(n33483) );
  XOR U35125 ( .A(mreg[719]), .B(creg[719]), .Z(n33484) );
  XOR U35126 ( .A(n33485), .B(n33486), .Z(n33476) );
  ANDN U35127 ( .A(n33487), .B(n26435), .Z(n33486) );
  XOR U35128 ( .A(n33488), .B(\modmult_1/zin[0][717] ), .Z(n26435) );
  IV U35129 ( .A(n33485), .Z(n33488) );
  XNOR U35130 ( .A(n33485), .B(n26434), .Z(n33487) );
  XOR U35131 ( .A(n33489), .B(n33490), .Z(n26434) );
  AND U35132 ( .A(\modmult_1/xin[1023] ), .B(n33491), .Z(n33490) );
  IV U35133 ( .A(n33489), .Z(n33491) );
  XOR U35134 ( .A(n33492), .B(mreg[718]), .Z(n33489) );
  NAND U35135 ( .A(n33493), .B(mul_pow), .Z(n33492) );
  XOR U35136 ( .A(mreg[718]), .B(creg[718]), .Z(n33493) );
  XOR U35137 ( .A(n33494), .B(n33495), .Z(n33485) );
  ANDN U35138 ( .A(n33496), .B(n26441), .Z(n33495) );
  XOR U35139 ( .A(n33497), .B(\modmult_1/zin[0][716] ), .Z(n26441) );
  IV U35140 ( .A(n33494), .Z(n33497) );
  XNOR U35141 ( .A(n33494), .B(n26440), .Z(n33496) );
  XOR U35142 ( .A(n33498), .B(n33499), .Z(n26440) );
  AND U35143 ( .A(\modmult_1/xin[1023] ), .B(n33500), .Z(n33499) );
  IV U35144 ( .A(n33498), .Z(n33500) );
  XOR U35145 ( .A(n33501), .B(mreg[717]), .Z(n33498) );
  NAND U35146 ( .A(n33502), .B(mul_pow), .Z(n33501) );
  XOR U35147 ( .A(mreg[717]), .B(creg[717]), .Z(n33502) );
  XOR U35148 ( .A(n33503), .B(n33504), .Z(n33494) );
  ANDN U35149 ( .A(n33505), .B(n26447), .Z(n33504) );
  XOR U35150 ( .A(n33506), .B(\modmult_1/zin[0][715] ), .Z(n26447) );
  IV U35151 ( .A(n33503), .Z(n33506) );
  XNOR U35152 ( .A(n33503), .B(n26446), .Z(n33505) );
  XOR U35153 ( .A(n33507), .B(n33508), .Z(n26446) );
  AND U35154 ( .A(\modmult_1/xin[1023] ), .B(n33509), .Z(n33508) );
  IV U35155 ( .A(n33507), .Z(n33509) );
  XOR U35156 ( .A(n33510), .B(mreg[716]), .Z(n33507) );
  NAND U35157 ( .A(n33511), .B(mul_pow), .Z(n33510) );
  XOR U35158 ( .A(mreg[716]), .B(creg[716]), .Z(n33511) );
  XOR U35159 ( .A(n33512), .B(n33513), .Z(n33503) );
  ANDN U35160 ( .A(n33514), .B(n26453), .Z(n33513) );
  XOR U35161 ( .A(n33515), .B(\modmult_1/zin[0][714] ), .Z(n26453) );
  IV U35162 ( .A(n33512), .Z(n33515) );
  XNOR U35163 ( .A(n33512), .B(n26452), .Z(n33514) );
  XOR U35164 ( .A(n33516), .B(n33517), .Z(n26452) );
  AND U35165 ( .A(\modmult_1/xin[1023] ), .B(n33518), .Z(n33517) );
  IV U35166 ( .A(n33516), .Z(n33518) );
  XOR U35167 ( .A(n33519), .B(mreg[715]), .Z(n33516) );
  NAND U35168 ( .A(n33520), .B(mul_pow), .Z(n33519) );
  XOR U35169 ( .A(mreg[715]), .B(creg[715]), .Z(n33520) );
  XOR U35170 ( .A(n33521), .B(n33522), .Z(n33512) );
  ANDN U35171 ( .A(n33523), .B(n26459), .Z(n33522) );
  XOR U35172 ( .A(n33524), .B(\modmult_1/zin[0][713] ), .Z(n26459) );
  IV U35173 ( .A(n33521), .Z(n33524) );
  XNOR U35174 ( .A(n33521), .B(n26458), .Z(n33523) );
  XOR U35175 ( .A(n33525), .B(n33526), .Z(n26458) );
  AND U35176 ( .A(\modmult_1/xin[1023] ), .B(n33527), .Z(n33526) );
  IV U35177 ( .A(n33525), .Z(n33527) );
  XOR U35178 ( .A(n33528), .B(mreg[714]), .Z(n33525) );
  NAND U35179 ( .A(n33529), .B(mul_pow), .Z(n33528) );
  XOR U35180 ( .A(mreg[714]), .B(creg[714]), .Z(n33529) );
  XOR U35181 ( .A(n33530), .B(n33531), .Z(n33521) );
  ANDN U35182 ( .A(n33532), .B(n26465), .Z(n33531) );
  XOR U35183 ( .A(n33533), .B(\modmult_1/zin[0][712] ), .Z(n26465) );
  IV U35184 ( .A(n33530), .Z(n33533) );
  XNOR U35185 ( .A(n33530), .B(n26464), .Z(n33532) );
  XOR U35186 ( .A(n33534), .B(n33535), .Z(n26464) );
  AND U35187 ( .A(\modmult_1/xin[1023] ), .B(n33536), .Z(n33535) );
  IV U35188 ( .A(n33534), .Z(n33536) );
  XOR U35189 ( .A(n33537), .B(mreg[713]), .Z(n33534) );
  NAND U35190 ( .A(n33538), .B(mul_pow), .Z(n33537) );
  XOR U35191 ( .A(mreg[713]), .B(creg[713]), .Z(n33538) );
  XOR U35192 ( .A(n33539), .B(n33540), .Z(n33530) );
  ANDN U35193 ( .A(n33541), .B(n26471), .Z(n33540) );
  XOR U35194 ( .A(n33542), .B(\modmult_1/zin[0][711] ), .Z(n26471) );
  IV U35195 ( .A(n33539), .Z(n33542) );
  XNOR U35196 ( .A(n33539), .B(n26470), .Z(n33541) );
  XOR U35197 ( .A(n33543), .B(n33544), .Z(n26470) );
  AND U35198 ( .A(\modmult_1/xin[1023] ), .B(n33545), .Z(n33544) );
  IV U35199 ( .A(n33543), .Z(n33545) );
  XOR U35200 ( .A(n33546), .B(mreg[712]), .Z(n33543) );
  NAND U35201 ( .A(n33547), .B(mul_pow), .Z(n33546) );
  XOR U35202 ( .A(mreg[712]), .B(creg[712]), .Z(n33547) );
  XOR U35203 ( .A(n33548), .B(n33549), .Z(n33539) );
  ANDN U35204 ( .A(n33550), .B(n26477), .Z(n33549) );
  XOR U35205 ( .A(n33551), .B(\modmult_1/zin[0][710] ), .Z(n26477) );
  IV U35206 ( .A(n33548), .Z(n33551) );
  XNOR U35207 ( .A(n33548), .B(n26476), .Z(n33550) );
  XOR U35208 ( .A(n33552), .B(n33553), .Z(n26476) );
  AND U35209 ( .A(\modmult_1/xin[1023] ), .B(n33554), .Z(n33553) );
  IV U35210 ( .A(n33552), .Z(n33554) );
  XOR U35211 ( .A(n33555), .B(mreg[711]), .Z(n33552) );
  NAND U35212 ( .A(n33556), .B(mul_pow), .Z(n33555) );
  XOR U35213 ( .A(mreg[711]), .B(creg[711]), .Z(n33556) );
  XOR U35214 ( .A(n33557), .B(n33558), .Z(n33548) );
  ANDN U35215 ( .A(n33559), .B(n26483), .Z(n33558) );
  XOR U35216 ( .A(n33560), .B(\modmult_1/zin[0][709] ), .Z(n26483) );
  IV U35217 ( .A(n33557), .Z(n33560) );
  XNOR U35218 ( .A(n33557), .B(n26482), .Z(n33559) );
  XOR U35219 ( .A(n33561), .B(n33562), .Z(n26482) );
  AND U35220 ( .A(\modmult_1/xin[1023] ), .B(n33563), .Z(n33562) );
  IV U35221 ( .A(n33561), .Z(n33563) );
  XOR U35222 ( .A(n33564), .B(mreg[710]), .Z(n33561) );
  NAND U35223 ( .A(n33565), .B(mul_pow), .Z(n33564) );
  XOR U35224 ( .A(mreg[710]), .B(creg[710]), .Z(n33565) );
  XOR U35225 ( .A(n33566), .B(n33567), .Z(n33557) );
  ANDN U35226 ( .A(n33568), .B(n26489), .Z(n33567) );
  XOR U35227 ( .A(n33569), .B(\modmult_1/zin[0][708] ), .Z(n26489) );
  IV U35228 ( .A(n33566), .Z(n33569) );
  XNOR U35229 ( .A(n33566), .B(n26488), .Z(n33568) );
  XOR U35230 ( .A(n33570), .B(n33571), .Z(n26488) );
  AND U35231 ( .A(\modmult_1/xin[1023] ), .B(n33572), .Z(n33571) );
  IV U35232 ( .A(n33570), .Z(n33572) );
  XOR U35233 ( .A(n33573), .B(mreg[709]), .Z(n33570) );
  NAND U35234 ( .A(n33574), .B(mul_pow), .Z(n33573) );
  XOR U35235 ( .A(mreg[709]), .B(creg[709]), .Z(n33574) );
  XOR U35236 ( .A(n33575), .B(n33576), .Z(n33566) );
  ANDN U35237 ( .A(n33577), .B(n26495), .Z(n33576) );
  XOR U35238 ( .A(n33578), .B(\modmult_1/zin[0][707] ), .Z(n26495) );
  IV U35239 ( .A(n33575), .Z(n33578) );
  XNOR U35240 ( .A(n33575), .B(n26494), .Z(n33577) );
  XOR U35241 ( .A(n33579), .B(n33580), .Z(n26494) );
  AND U35242 ( .A(\modmult_1/xin[1023] ), .B(n33581), .Z(n33580) );
  IV U35243 ( .A(n33579), .Z(n33581) );
  XOR U35244 ( .A(n33582), .B(mreg[708]), .Z(n33579) );
  NAND U35245 ( .A(n33583), .B(mul_pow), .Z(n33582) );
  XOR U35246 ( .A(mreg[708]), .B(creg[708]), .Z(n33583) );
  XOR U35247 ( .A(n33584), .B(n33585), .Z(n33575) );
  ANDN U35248 ( .A(n33586), .B(n26501), .Z(n33585) );
  XOR U35249 ( .A(n33587), .B(\modmult_1/zin[0][706] ), .Z(n26501) );
  IV U35250 ( .A(n33584), .Z(n33587) );
  XNOR U35251 ( .A(n33584), .B(n26500), .Z(n33586) );
  XOR U35252 ( .A(n33588), .B(n33589), .Z(n26500) );
  AND U35253 ( .A(\modmult_1/xin[1023] ), .B(n33590), .Z(n33589) );
  IV U35254 ( .A(n33588), .Z(n33590) );
  XOR U35255 ( .A(n33591), .B(mreg[707]), .Z(n33588) );
  NAND U35256 ( .A(n33592), .B(mul_pow), .Z(n33591) );
  XOR U35257 ( .A(mreg[707]), .B(creg[707]), .Z(n33592) );
  XOR U35258 ( .A(n33593), .B(n33594), .Z(n33584) );
  ANDN U35259 ( .A(n33595), .B(n26507), .Z(n33594) );
  XOR U35260 ( .A(n33596), .B(\modmult_1/zin[0][705] ), .Z(n26507) );
  IV U35261 ( .A(n33593), .Z(n33596) );
  XNOR U35262 ( .A(n33593), .B(n26506), .Z(n33595) );
  XOR U35263 ( .A(n33597), .B(n33598), .Z(n26506) );
  AND U35264 ( .A(\modmult_1/xin[1023] ), .B(n33599), .Z(n33598) );
  IV U35265 ( .A(n33597), .Z(n33599) );
  XOR U35266 ( .A(n33600), .B(mreg[706]), .Z(n33597) );
  NAND U35267 ( .A(n33601), .B(mul_pow), .Z(n33600) );
  XOR U35268 ( .A(mreg[706]), .B(creg[706]), .Z(n33601) );
  XOR U35269 ( .A(n33602), .B(n33603), .Z(n33593) );
  ANDN U35270 ( .A(n33604), .B(n26513), .Z(n33603) );
  XOR U35271 ( .A(n33605), .B(\modmult_1/zin[0][704] ), .Z(n26513) );
  IV U35272 ( .A(n33602), .Z(n33605) );
  XNOR U35273 ( .A(n33602), .B(n26512), .Z(n33604) );
  XOR U35274 ( .A(n33606), .B(n33607), .Z(n26512) );
  AND U35275 ( .A(\modmult_1/xin[1023] ), .B(n33608), .Z(n33607) );
  IV U35276 ( .A(n33606), .Z(n33608) );
  XOR U35277 ( .A(n33609), .B(mreg[705]), .Z(n33606) );
  NAND U35278 ( .A(n33610), .B(mul_pow), .Z(n33609) );
  XOR U35279 ( .A(mreg[705]), .B(creg[705]), .Z(n33610) );
  XOR U35280 ( .A(n33611), .B(n33612), .Z(n33602) );
  ANDN U35281 ( .A(n33613), .B(n26519), .Z(n33612) );
  XOR U35282 ( .A(n33614), .B(\modmult_1/zin[0][703] ), .Z(n26519) );
  IV U35283 ( .A(n33611), .Z(n33614) );
  XNOR U35284 ( .A(n33611), .B(n26518), .Z(n33613) );
  XOR U35285 ( .A(n33615), .B(n33616), .Z(n26518) );
  AND U35286 ( .A(\modmult_1/xin[1023] ), .B(n33617), .Z(n33616) );
  IV U35287 ( .A(n33615), .Z(n33617) );
  XOR U35288 ( .A(n33618), .B(mreg[704]), .Z(n33615) );
  NAND U35289 ( .A(n33619), .B(mul_pow), .Z(n33618) );
  XOR U35290 ( .A(mreg[704]), .B(creg[704]), .Z(n33619) );
  XOR U35291 ( .A(n33620), .B(n33621), .Z(n33611) );
  ANDN U35292 ( .A(n33622), .B(n26525), .Z(n33621) );
  XOR U35293 ( .A(n33623), .B(\modmult_1/zin[0][702] ), .Z(n26525) );
  IV U35294 ( .A(n33620), .Z(n33623) );
  XNOR U35295 ( .A(n33620), .B(n26524), .Z(n33622) );
  XOR U35296 ( .A(n33624), .B(n33625), .Z(n26524) );
  AND U35297 ( .A(\modmult_1/xin[1023] ), .B(n33626), .Z(n33625) );
  IV U35298 ( .A(n33624), .Z(n33626) );
  XOR U35299 ( .A(n33627), .B(mreg[703]), .Z(n33624) );
  NAND U35300 ( .A(n33628), .B(mul_pow), .Z(n33627) );
  XOR U35301 ( .A(mreg[703]), .B(creg[703]), .Z(n33628) );
  XOR U35302 ( .A(n33629), .B(n33630), .Z(n33620) );
  ANDN U35303 ( .A(n33631), .B(n26531), .Z(n33630) );
  XOR U35304 ( .A(n33632), .B(\modmult_1/zin[0][701] ), .Z(n26531) );
  IV U35305 ( .A(n33629), .Z(n33632) );
  XNOR U35306 ( .A(n33629), .B(n26530), .Z(n33631) );
  XOR U35307 ( .A(n33633), .B(n33634), .Z(n26530) );
  AND U35308 ( .A(\modmult_1/xin[1023] ), .B(n33635), .Z(n33634) );
  IV U35309 ( .A(n33633), .Z(n33635) );
  XOR U35310 ( .A(n33636), .B(mreg[702]), .Z(n33633) );
  NAND U35311 ( .A(n33637), .B(mul_pow), .Z(n33636) );
  XOR U35312 ( .A(mreg[702]), .B(creg[702]), .Z(n33637) );
  XOR U35313 ( .A(n33638), .B(n33639), .Z(n33629) );
  ANDN U35314 ( .A(n33640), .B(n26537), .Z(n33639) );
  XOR U35315 ( .A(n33641), .B(\modmult_1/zin[0][700] ), .Z(n26537) );
  IV U35316 ( .A(n33638), .Z(n33641) );
  XNOR U35317 ( .A(n33638), .B(n26536), .Z(n33640) );
  XOR U35318 ( .A(n33642), .B(n33643), .Z(n26536) );
  AND U35319 ( .A(\modmult_1/xin[1023] ), .B(n33644), .Z(n33643) );
  IV U35320 ( .A(n33642), .Z(n33644) );
  XOR U35321 ( .A(n33645), .B(mreg[701]), .Z(n33642) );
  NAND U35322 ( .A(n33646), .B(mul_pow), .Z(n33645) );
  XOR U35323 ( .A(mreg[701]), .B(creg[701]), .Z(n33646) );
  XOR U35324 ( .A(n33647), .B(n33648), .Z(n33638) );
  ANDN U35325 ( .A(n33649), .B(n26543), .Z(n33648) );
  XOR U35326 ( .A(n33650), .B(\modmult_1/zin[0][699] ), .Z(n26543) );
  IV U35327 ( .A(n33647), .Z(n33650) );
  XNOR U35328 ( .A(n33647), .B(n26542), .Z(n33649) );
  XOR U35329 ( .A(n33651), .B(n33652), .Z(n26542) );
  AND U35330 ( .A(\modmult_1/xin[1023] ), .B(n33653), .Z(n33652) );
  IV U35331 ( .A(n33651), .Z(n33653) );
  XOR U35332 ( .A(n33654), .B(mreg[700]), .Z(n33651) );
  NAND U35333 ( .A(n33655), .B(mul_pow), .Z(n33654) );
  XOR U35334 ( .A(mreg[700]), .B(creg[700]), .Z(n33655) );
  XOR U35335 ( .A(n33656), .B(n33657), .Z(n33647) );
  ANDN U35336 ( .A(n33658), .B(n26549), .Z(n33657) );
  XOR U35337 ( .A(n33659), .B(\modmult_1/zin[0][698] ), .Z(n26549) );
  IV U35338 ( .A(n33656), .Z(n33659) );
  XNOR U35339 ( .A(n33656), .B(n26548), .Z(n33658) );
  XOR U35340 ( .A(n33660), .B(n33661), .Z(n26548) );
  AND U35341 ( .A(\modmult_1/xin[1023] ), .B(n33662), .Z(n33661) );
  IV U35342 ( .A(n33660), .Z(n33662) );
  XOR U35343 ( .A(n33663), .B(mreg[699]), .Z(n33660) );
  NAND U35344 ( .A(n33664), .B(mul_pow), .Z(n33663) );
  XOR U35345 ( .A(mreg[699]), .B(creg[699]), .Z(n33664) );
  XOR U35346 ( .A(n33665), .B(n33666), .Z(n33656) );
  ANDN U35347 ( .A(n33667), .B(n26555), .Z(n33666) );
  XOR U35348 ( .A(n33668), .B(\modmult_1/zin[0][697] ), .Z(n26555) );
  IV U35349 ( .A(n33665), .Z(n33668) );
  XNOR U35350 ( .A(n33665), .B(n26554), .Z(n33667) );
  XOR U35351 ( .A(n33669), .B(n33670), .Z(n26554) );
  AND U35352 ( .A(\modmult_1/xin[1023] ), .B(n33671), .Z(n33670) );
  IV U35353 ( .A(n33669), .Z(n33671) );
  XOR U35354 ( .A(n33672), .B(mreg[698]), .Z(n33669) );
  NAND U35355 ( .A(n33673), .B(mul_pow), .Z(n33672) );
  XOR U35356 ( .A(mreg[698]), .B(creg[698]), .Z(n33673) );
  XOR U35357 ( .A(n33674), .B(n33675), .Z(n33665) );
  ANDN U35358 ( .A(n33676), .B(n26561), .Z(n33675) );
  XOR U35359 ( .A(n33677), .B(\modmult_1/zin[0][696] ), .Z(n26561) );
  IV U35360 ( .A(n33674), .Z(n33677) );
  XNOR U35361 ( .A(n33674), .B(n26560), .Z(n33676) );
  XOR U35362 ( .A(n33678), .B(n33679), .Z(n26560) );
  AND U35363 ( .A(\modmult_1/xin[1023] ), .B(n33680), .Z(n33679) );
  IV U35364 ( .A(n33678), .Z(n33680) );
  XOR U35365 ( .A(n33681), .B(mreg[697]), .Z(n33678) );
  NAND U35366 ( .A(n33682), .B(mul_pow), .Z(n33681) );
  XOR U35367 ( .A(mreg[697]), .B(creg[697]), .Z(n33682) );
  XOR U35368 ( .A(n33683), .B(n33684), .Z(n33674) );
  ANDN U35369 ( .A(n33685), .B(n26567), .Z(n33684) );
  XOR U35370 ( .A(n33686), .B(\modmult_1/zin[0][695] ), .Z(n26567) );
  IV U35371 ( .A(n33683), .Z(n33686) );
  XNOR U35372 ( .A(n33683), .B(n26566), .Z(n33685) );
  XOR U35373 ( .A(n33687), .B(n33688), .Z(n26566) );
  AND U35374 ( .A(\modmult_1/xin[1023] ), .B(n33689), .Z(n33688) );
  IV U35375 ( .A(n33687), .Z(n33689) );
  XOR U35376 ( .A(n33690), .B(mreg[696]), .Z(n33687) );
  NAND U35377 ( .A(n33691), .B(mul_pow), .Z(n33690) );
  XOR U35378 ( .A(mreg[696]), .B(creg[696]), .Z(n33691) );
  XOR U35379 ( .A(n33692), .B(n33693), .Z(n33683) );
  ANDN U35380 ( .A(n33694), .B(n26573), .Z(n33693) );
  XOR U35381 ( .A(n33695), .B(\modmult_1/zin[0][694] ), .Z(n26573) );
  IV U35382 ( .A(n33692), .Z(n33695) );
  XNOR U35383 ( .A(n33692), .B(n26572), .Z(n33694) );
  XOR U35384 ( .A(n33696), .B(n33697), .Z(n26572) );
  AND U35385 ( .A(\modmult_1/xin[1023] ), .B(n33698), .Z(n33697) );
  IV U35386 ( .A(n33696), .Z(n33698) );
  XOR U35387 ( .A(n33699), .B(mreg[695]), .Z(n33696) );
  NAND U35388 ( .A(n33700), .B(mul_pow), .Z(n33699) );
  XOR U35389 ( .A(mreg[695]), .B(creg[695]), .Z(n33700) );
  XOR U35390 ( .A(n33701), .B(n33702), .Z(n33692) );
  ANDN U35391 ( .A(n33703), .B(n26579), .Z(n33702) );
  XOR U35392 ( .A(n33704), .B(\modmult_1/zin[0][693] ), .Z(n26579) );
  IV U35393 ( .A(n33701), .Z(n33704) );
  XNOR U35394 ( .A(n33701), .B(n26578), .Z(n33703) );
  XOR U35395 ( .A(n33705), .B(n33706), .Z(n26578) );
  AND U35396 ( .A(\modmult_1/xin[1023] ), .B(n33707), .Z(n33706) );
  IV U35397 ( .A(n33705), .Z(n33707) );
  XOR U35398 ( .A(n33708), .B(mreg[694]), .Z(n33705) );
  NAND U35399 ( .A(n33709), .B(mul_pow), .Z(n33708) );
  XOR U35400 ( .A(mreg[694]), .B(creg[694]), .Z(n33709) );
  XOR U35401 ( .A(n33710), .B(n33711), .Z(n33701) );
  ANDN U35402 ( .A(n33712), .B(n26585), .Z(n33711) );
  XOR U35403 ( .A(n33713), .B(\modmult_1/zin[0][692] ), .Z(n26585) );
  IV U35404 ( .A(n33710), .Z(n33713) );
  XNOR U35405 ( .A(n33710), .B(n26584), .Z(n33712) );
  XOR U35406 ( .A(n33714), .B(n33715), .Z(n26584) );
  AND U35407 ( .A(\modmult_1/xin[1023] ), .B(n33716), .Z(n33715) );
  IV U35408 ( .A(n33714), .Z(n33716) );
  XOR U35409 ( .A(n33717), .B(mreg[693]), .Z(n33714) );
  NAND U35410 ( .A(n33718), .B(mul_pow), .Z(n33717) );
  XOR U35411 ( .A(mreg[693]), .B(creg[693]), .Z(n33718) );
  XOR U35412 ( .A(n33719), .B(n33720), .Z(n33710) );
  ANDN U35413 ( .A(n33721), .B(n26591), .Z(n33720) );
  XOR U35414 ( .A(n33722), .B(\modmult_1/zin[0][691] ), .Z(n26591) );
  IV U35415 ( .A(n33719), .Z(n33722) );
  XNOR U35416 ( .A(n33719), .B(n26590), .Z(n33721) );
  XOR U35417 ( .A(n33723), .B(n33724), .Z(n26590) );
  AND U35418 ( .A(\modmult_1/xin[1023] ), .B(n33725), .Z(n33724) );
  IV U35419 ( .A(n33723), .Z(n33725) );
  XOR U35420 ( .A(n33726), .B(mreg[692]), .Z(n33723) );
  NAND U35421 ( .A(n33727), .B(mul_pow), .Z(n33726) );
  XOR U35422 ( .A(mreg[692]), .B(creg[692]), .Z(n33727) );
  XOR U35423 ( .A(n33728), .B(n33729), .Z(n33719) );
  ANDN U35424 ( .A(n33730), .B(n26597), .Z(n33729) );
  XOR U35425 ( .A(n33731), .B(\modmult_1/zin[0][690] ), .Z(n26597) );
  IV U35426 ( .A(n33728), .Z(n33731) );
  XNOR U35427 ( .A(n33728), .B(n26596), .Z(n33730) );
  XOR U35428 ( .A(n33732), .B(n33733), .Z(n26596) );
  AND U35429 ( .A(\modmult_1/xin[1023] ), .B(n33734), .Z(n33733) );
  IV U35430 ( .A(n33732), .Z(n33734) );
  XOR U35431 ( .A(n33735), .B(mreg[691]), .Z(n33732) );
  NAND U35432 ( .A(n33736), .B(mul_pow), .Z(n33735) );
  XOR U35433 ( .A(mreg[691]), .B(creg[691]), .Z(n33736) );
  XOR U35434 ( .A(n33737), .B(n33738), .Z(n33728) );
  ANDN U35435 ( .A(n33739), .B(n26603), .Z(n33738) );
  XOR U35436 ( .A(n33740), .B(\modmult_1/zin[0][689] ), .Z(n26603) );
  IV U35437 ( .A(n33737), .Z(n33740) );
  XNOR U35438 ( .A(n33737), .B(n26602), .Z(n33739) );
  XOR U35439 ( .A(n33741), .B(n33742), .Z(n26602) );
  AND U35440 ( .A(\modmult_1/xin[1023] ), .B(n33743), .Z(n33742) );
  IV U35441 ( .A(n33741), .Z(n33743) );
  XOR U35442 ( .A(n33744), .B(mreg[690]), .Z(n33741) );
  NAND U35443 ( .A(n33745), .B(mul_pow), .Z(n33744) );
  XOR U35444 ( .A(mreg[690]), .B(creg[690]), .Z(n33745) );
  XOR U35445 ( .A(n33746), .B(n33747), .Z(n33737) );
  ANDN U35446 ( .A(n33748), .B(n26609), .Z(n33747) );
  XOR U35447 ( .A(n33749), .B(\modmult_1/zin[0][688] ), .Z(n26609) );
  IV U35448 ( .A(n33746), .Z(n33749) );
  XNOR U35449 ( .A(n33746), .B(n26608), .Z(n33748) );
  XOR U35450 ( .A(n33750), .B(n33751), .Z(n26608) );
  AND U35451 ( .A(\modmult_1/xin[1023] ), .B(n33752), .Z(n33751) );
  IV U35452 ( .A(n33750), .Z(n33752) );
  XOR U35453 ( .A(n33753), .B(mreg[689]), .Z(n33750) );
  NAND U35454 ( .A(n33754), .B(mul_pow), .Z(n33753) );
  XOR U35455 ( .A(mreg[689]), .B(creg[689]), .Z(n33754) );
  XOR U35456 ( .A(n33755), .B(n33756), .Z(n33746) );
  ANDN U35457 ( .A(n33757), .B(n26615), .Z(n33756) );
  XOR U35458 ( .A(n33758), .B(\modmult_1/zin[0][687] ), .Z(n26615) );
  IV U35459 ( .A(n33755), .Z(n33758) );
  XNOR U35460 ( .A(n33755), .B(n26614), .Z(n33757) );
  XOR U35461 ( .A(n33759), .B(n33760), .Z(n26614) );
  AND U35462 ( .A(\modmult_1/xin[1023] ), .B(n33761), .Z(n33760) );
  IV U35463 ( .A(n33759), .Z(n33761) );
  XOR U35464 ( .A(n33762), .B(mreg[688]), .Z(n33759) );
  NAND U35465 ( .A(n33763), .B(mul_pow), .Z(n33762) );
  XOR U35466 ( .A(mreg[688]), .B(creg[688]), .Z(n33763) );
  XOR U35467 ( .A(n33764), .B(n33765), .Z(n33755) );
  ANDN U35468 ( .A(n33766), .B(n26621), .Z(n33765) );
  XOR U35469 ( .A(n33767), .B(\modmult_1/zin[0][686] ), .Z(n26621) );
  IV U35470 ( .A(n33764), .Z(n33767) );
  XNOR U35471 ( .A(n33764), .B(n26620), .Z(n33766) );
  XOR U35472 ( .A(n33768), .B(n33769), .Z(n26620) );
  AND U35473 ( .A(\modmult_1/xin[1023] ), .B(n33770), .Z(n33769) );
  IV U35474 ( .A(n33768), .Z(n33770) );
  XOR U35475 ( .A(n33771), .B(mreg[687]), .Z(n33768) );
  NAND U35476 ( .A(n33772), .B(mul_pow), .Z(n33771) );
  XOR U35477 ( .A(mreg[687]), .B(creg[687]), .Z(n33772) );
  XOR U35478 ( .A(n33773), .B(n33774), .Z(n33764) );
  ANDN U35479 ( .A(n33775), .B(n26627), .Z(n33774) );
  XOR U35480 ( .A(n33776), .B(\modmult_1/zin[0][685] ), .Z(n26627) );
  IV U35481 ( .A(n33773), .Z(n33776) );
  XNOR U35482 ( .A(n33773), .B(n26626), .Z(n33775) );
  XOR U35483 ( .A(n33777), .B(n33778), .Z(n26626) );
  AND U35484 ( .A(\modmult_1/xin[1023] ), .B(n33779), .Z(n33778) );
  IV U35485 ( .A(n33777), .Z(n33779) );
  XOR U35486 ( .A(n33780), .B(mreg[686]), .Z(n33777) );
  NAND U35487 ( .A(n33781), .B(mul_pow), .Z(n33780) );
  XOR U35488 ( .A(mreg[686]), .B(creg[686]), .Z(n33781) );
  XOR U35489 ( .A(n33782), .B(n33783), .Z(n33773) );
  ANDN U35490 ( .A(n33784), .B(n26633), .Z(n33783) );
  XOR U35491 ( .A(n33785), .B(\modmult_1/zin[0][684] ), .Z(n26633) );
  IV U35492 ( .A(n33782), .Z(n33785) );
  XNOR U35493 ( .A(n33782), .B(n26632), .Z(n33784) );
  XOR U35494 ( .A(n33786), .B(n33787), .Z(n26632) );
  AND U35495 ( .A(\modmult_1/xin[1023] ), .B(n33788), .Z(n33787) );
  IV U35496 ( .A(n33786), .Z(n33788) );
  XOR U35497 ( .A(n33789), .B(mreg[685]), .Z(n33786) );
  NAND U35498 ( .A(n33790), .B(mul_pow), .Z(n33789) );
  XOR U35499 ( .A(mreg[685]), .B(creg[685]), .Z(n33790) );
  XOR U35500 ( .A(n33791), .B(n33792), .Z(n33782) );
  ANDN U35501 ( .A(n33793), .B(n26639), .Z(n33792) );
  XOR U35502 ( .A(n33794), .B(\modmult_1/zin[0][683] ), .Z(n26639) );
  IV U35503 ( .A(n33791), .Z(n33794) );
  XNOR U35504 ( .A(n33791), .B(n26638), .Z(n33793) );
  XOR U35505 ( .A(n33795), .B(n33796), .Z(n26638) );
  AND U35506 ( .A(\modmult_1/xin[1023] ), .B(n33797), .Z(n33796) );
  IV U35507 ( .A(n33795), .Z(n33797) );
  XOR U35508 ( .A(n33798), .B(mreg[684]), .Z(n33795) );
  NAND U35509 ( .A(n33799), .B(mul_pow), .Z(n33798) );
  XOR U35510 ( .A(mreg[684]), .B(creg[684]), .Z(n33799) );
  XOR U35511 ( .A(n33800), .B(n33801), .Z(n33791) );
  ANDN U35512 ( .A(n33802), .B(n26645), .Z(n33801) );
  XOR U35513 ( .A(n33803), .B(\modmult_1/zin[0][682] ), .Z(n26645) );
  IV U35514 ( .A(n33800), .Z(n33803) );
  XNOR U35515 ( .A(n33800), .B(n26644), .Z(n33802) );
  XOR U35516 ( .A(n33804), .B(n33805), .Z(n26644) );
  AND U35517 ( .A(\modmult_1/xin[1023] ), .B(n33806), .Z(n33805) );
  IV U35518 ( .A(n33804), .Z(n33806) );
  XOR U35519 ( .A(n33807), .B(mreg[683]), .Z(n33804) );
  NAND U35520 ( .A(n33808), .B(mul_pow), .Z(n33807) );
  XOR U35521 ( .A(mreg[683]), .B(creg[683]), .Z(n33808) );
  XOR U35522 ( .A(n33809), .B(n33810), .Z(n33800) );
  ANDN U35523 ( .A(n33811), .B(n26651), .Z(n33810) );
  XOR U35524 ( .A(n33812), .B(\modmult_1/zin[0][681] ), .Z(n26651) );
  IV U35525 ( .A(n33809), .Z(n33812) );
  XNOR U35526 ( .A(n33809), .B(n26650), .Z(n33811) );
  XOR U35527 ( .A(n33813), .B(n33814), .Z(n26650) );
  AND U35528 ( .A(\modmult_1/xin[1023] ), .B(n33815), .Z(n33814) );
  IV U35529 ( .A(n33813), .Z(n33815) );
  XOR U35530 ( .A(n33816), .B(mreg[682]), .Z(n33813) );
  NAND U35531 ( .A(n33817), .B(mul_pow), .Z(n33816) );
  XOR U35532 ( .A(mreg[682]), .B(creg[682]), .Z(n33817) );
  XOR U35533 ( .A(n33818), .B(n33819), .Z(n33809) );
  ANDN U35534 ( .A(n33820), .B(n26657), .Z(n33819) );
  XOR U35535 ( .A(n33821), .B(\modmult_1/zin[0][680] ), .Z(n26657) );
  IV U35536 ( .A(n33818), .Z(n33821) );
  XNOR U35537 ( .A(n33818), .B(n26656), .Z(n33820) );
  XOR U35538 ( .A(n33822), .B(n33823), .Z(n26656) );
  AND U35539 ( .A(\modmult_1/xin[1023] ), .B(n33824), .Z(n33823) );
  IV U35540 ( .A(n33822), .Z(n33824) );
  XOR U35541 ( .A(n33825), .B(mreg[681]), .Z(n33822) );
  NAND U35542 ( .A(n33826), .B(mul_pow), .Z(n33825) );
  XOR U35543 ( .A(mreg[681]), .B(creg[681]), .Z(n33826) );
  XOR U35544 ( .A(n33827), .B(n33828), .Z(n33818) );
  ANDN U35545 ( .A(n33829), .B(n26663), .Z(n33828) );
  XOR U35546 ( .A(n33830), .B(\modmult_1/zin[0][679] ), .Z(n26663) );
  IV U35547 ( .A(n33827), .Z(n33830) );
  XNOR U35548 ( .A(n33827), .B(n26662), .Z(n33829) );
  XOR U35549 ( .A(n33831), .B(n33832), .Z(n26662) );
  AND U35550 ( .A(\modmult_1/xin[1023] ), .B(n33833), .Z(n33832) );
  IV U35551 ( .A(n33831), .Z(n33833) );
  XOR U35552 ( .A(n33834), .B(mreg[680]), .Z(n33831) );
  NAND U35553 ( .A(n33835), .B(mul_pow), .Z(n33834) );
  XOR U35554 ( .A(mreg[680]), .B(creg[680]), .Z(n33835) );
  XOR U35555 ( .A(n33836), .B(n33837), .Z(n33827) );
  ANDN U35556 ( .A(n33838), .B(n26669), .Z(n33837) );
  XOR U35557 ( .A(n33839), .B(\modmult_1/zin[0][678] ), .Z(n26669) );
  IV U35558 ( .A(n33836), .Z(n33839) );
  XNOR U35559 ( .A(n33836), .B(n26668), .Z(n33838) );
  XOR U35560 ( .A(n33840), .B(n33841), .Z(n26668) );
  AND U35561 ( .A(\modmult_1/xin[1023] ), .B(n33842), .Z(n33841) );
  IV U35562 ( .A(n33840), .Z(n33842) );
  XOR U35563 ( .A(n33843), .B(mreg[679]), .Z(n33840) );
  NAND U35564 ( .A(n33844), .B(mul_pow), .Z(n33843) );
  XOR U35565 ( .A(mreg[679]), .B(creg[679]), .Z(n33844) );
  XOR U35566 ( .A(n33845), .B(n33846), .Z(n33836) );
  ANDN U35567 ( .A(n33847), .B(n26675), .Z(n33846) );
  XOR U35568 ( .A(n33848), .B(\modmult_1/zin[0][677] ), .Z(n26675) );
  IV U35569 ( .A(n33845), .Z(n33848) );
  XNOR U35570 ( .A(n33845), .B(n26674), .Z(n33847) );
  XOR U35571 ( .A(n33849), .B(n33850), .Z(n26674) );
  AND U35572 ( .A(\modmult_1/xin[1023] ), .B(n33851), .Z(n33850) );
  IV U35573 ( .A(n33849), .Z(n33851) );
  XOR U35574 ( .A(n33852), .B(mreg[678]), .Z(n33849) );
  NAND U35575 ( .A(n33853), .B(mul_pow), .Z(n33852) );
  XOR U35576 ( .A(mreg[678]), .B(creg[678]), .Z(n33853) );
  XOR U35577 ( .A(n33854), .B(n33855), .Z(n33845) );
  ANDN U35578 ( .A(n33856), .B(n26681), .Z(n33855) );
  XOR U35579 ( .A(n33857), .B(\modmult_1/zin[0][676] ), .Z(n26681) );
  IV U35580 ( .A(n33854), .Z(n33857) );
  XNOR U35581 ( .A(n33854), .B(n26680), .Z(n33856) );
  XOR U35582 ( .A(n33858), .B(n33859), .Z(n26680) );
  AND U35583 ( .A(\modmult_1/xin[1023] ), .B(n33860), .Z(n33859) );
  IV U35584 ( .A(n33858), .Z(n33860) );
  XOR U35585 ( .A(n33861), .B(mreg[677]), .Z(n33858) );
  NAND U35586 ( .A(n33862), .B(mul_pow), .Z(n33861) );
  XOR U35587 ( .A(mreg[677]), .B(creg[677]), .Z(n33862) );
  XOR U35588 ( .A(n33863), .B(n33864), .Z(n33854) );
  ANDN U35589 ( .A(n33865), .B(n26687), .Z(n33864) );
  XOR U35590 ( .A(n33866), .B(\modmult_1/zin[0][675] ), .Z(n26687) );
  IV U35591 ( .A(n33863), .Z(n33866) );
  XNOR U35592 ( .A(n33863), .B(n26686), .Z(n33865) );
  XOR U35593 ( .A(n33867), .B(n33868), .Z(n26686) );
  AND U35594 ( .A(\modmult_1/xin[1023] ), .B(n33869), .Z(n33868) );
  IV U35595 ( .A(n33867), .Z(n33869) );
  XOR U35596 ( .A(n33870), .B(mreg[676]), .Z(n33867) );
  NAND U35597 ( .A(n33871), .B(mul_pow), .Z(n33870) );
  XOR U35598 ( .A(mreg[676]), .B(creg[676]), .Z(n33871) );
  XOR U35599 ( .A(n33872), .B(n33873), .Z(n33863) );
  ANDN U35600 ( .A(n33874), .B(n26693), .Z(n33873) );
  XOR U35601 ( .A(n33875), .B(\modmult_1/zin[0][674] ), .Z(n26693) );
  IV U35602 ( .A(n33872), .Z(n33875) );
  XNOR U35603 ( .A(n33872), .B(n26692), .Z(n33874) );
  XOR U35604 ( .A(n33876), .B(n33877), .Z(n26692) );
  AND U35605 ( .A(\modmult_1/xin[1023] ), .B(n33878), .Z(n33877) );
  IV U35606 ( .A(n33876), .Z(n33878) );
  XOR U35607 ( .A(n33879), .B(mreg[675]), .Z(n33876) );
  NAND U35608 ( .A(n33880), .B(mul_pow), .Z(n33879) );
  XOR U35609 ( .A(mreg[675]), .B(creg[675]), .Z(n33880) );
  XOR U35610 ( .A(n33881), .B(n33882), .Z(n33872) );
  ANDN U35611 ( .A(n33883), .B(n26699), .Z(n33882) );
  XOR U35612 ( .A(n33884), .B(\modmult_1/zin[0][673] ), .Z(n26699) );
  IV U35613 ( .A(n33881), .Z(n33884) );
  XNOR U35614 ( .A(n33881), .B(n26698), .Z(n33883) );
  XOR U35615 ( .A(n33885), .B(n33886), .Z(n26698) );
  AND U35616 ( .A(\modmult_1/xin[1023] ), .B(n33887), .Z(n33886) );
  IV U35617 ( .A(n33885), .Z(n33887) );
  XOR U35618 ( .A(n33888), .B(mreg[674]), .Z(n33885) );
  NAND U35619 ( .A(n33889), .B(mul_pow), .Z(n33888) );
  XOR U35620 ( .A(mreg[674]), .B(creg[674]), .Z(n33889) );
  XOR U35621 ( .A(n33890), .B(n33891), .Z(n33881) );
  ANDN U35622 ( .A(n33892), .B(n26705), .Z(n33891) );
  XOR U35623 ( .A(n33893), .B(\modmult_1/zin[0][672] ), .Z(n26705) );
  IV U35624 ( .A(n33890), .Z(n33893) );
  XNOR U35625 ( .A(n33890), .B(n26704), .Z(n33892) );
  XOR U35626 ( .A(n33894), .B(n33895), .Z(n26704) );
  AND U35627 ( .A(\modmult_1/xin[1023] ), .B(n33896), .Z(n33895) );
  IV U35628 ( .A(n33894), .Z(n33896) );
  XOR U35629 ( .A(n33897), .B(mreg[673]), .Z(n33894) );
  NAND U35630 ( .A(n33898), .B(mul_pow), .Z(n33897) );
  XOR U35631 ( .A(mreg[673]), .B(creg[673]), .Z(n33898) );
  XOR U35632 ( .A(n33899), .B(n33900), .Z(n33890) );
  ANDN U35633 ( .A(n33901), .B(n26711), .Z(n33900) );
  XOR U35634 ( .A(n33902), .B(\modmult_1/zin[0][671] ), .Z(n26711) );
  IV U35635 ( .A(n33899), .Z(n33902) );
  XNOR U35636 ( .A(n33899), .B(n26710), .Z(n33901) );
  XOR U35637 ( .A(n33903), .B(n33904), .Z(n26710) );
  AND U35638 ( .A(\modmult_1/xin[1023] ), .B(n33905), .Z(n33904) );
  IV U35639 ( .A(n33903), .Z(n33905) );
  XOR U35640 ( .A(n33906), .B(mreg[672]), .Z(n33903) );
  NAND U35641 ( .A(n33907), .B(mul_pow), .Z(n33906) );
  XOR U35642 ( .A(mreg[672]), .B(creg[672]), .Z(n33907) );
  XOR U35643 ( .A(n33908), .B(n33909), .Z(n33899) );
  ANDN U35644 ( .A(n33910), .B(n26717), .Z(n33909) );
  XOR U35645 ( .A(n33911), .B(\modmult_1/zin[0][670] ), .Z(n26717) );
  IV U35646 ( .A(n33908), .Z(n33911) );
  XNOR U35647 ( .A(n33908), .B(n26716), .Z(n33910) );
  XOR U35648 ( .A(n33912), .B(n33913), .Z(n26716) );
  AND U35649 ( .A(\modmult_1/xin[1023] ), .B(n33914), .Z(n33913) );
  IV U35650 ( .A(n33912), .Z(n33914) );
  XOR U35651 ( .A(n33915), .B(mreg[671]), .Z(n33912) );
  NAND U35652 ( .A(n33916), .B(mul_pow), .Z(n33915) );
  XOR U35653 ( .A(mreg[671]), .B(creg[671]), .Z(n33916) );
  XOR U35654 ( .A(n33917), .B(n33918), .Z(n33908) );
  ANDN U35655 ( .A(n33919), .B(n26723), .Z(n33918) );
  XOR U35656 ( .A(n33920), .B(\modmult_1/zin[0][669] ), .Z(n26723) );
  IV U35657 ( .A(n33917), .Z(n33920) );
  XNOR U35658 ( .A(n33917), .B(n26722), .Z(n33919) );
  XOR U35659 ( .A(n33921), .B(n33922), .Z(n26722) );
  AND U35660 ( .A(\modmult_1/xin[1023] ), .B(n33923), .Z(n33922) );
  IV U35661 ( .A(n33921), .Z(n33923) );
  XOR U35662 ( .A(n33924), .B(mreg[670]), .Z(n33921) );
  NAND U35663 ( .A(n33925), .B(mul_pow), .Z(n33924) );
  XOR U35664 ( .A(mreg[670]), .B(creg[670]), .Z(n33925) );
  XOR U35665 ( .A(n33926), .B(n33927), .Z(n33917) );
  ANDN U35666 ( .A(n33928), .B(n26729), .Z(n33927) );
  XOR U35667 ( .A(n33929), .B(\modmult_1/zin[0][668] ), .Z(n26729) );
  IV U35668 ( .A(n33926), .Z(n33929) );
  XNOR U35669 ( .A(n33926), .B(n26728), .Z(n33928) );
  XOR U35670 ( .A(n33930), .B(n33931), .Z(n26728) );
  AND U35671 ( .A(\modmult_1/xin[1023] ), .B(n33932), .Z(n33931) );
  IV U35672 ( .A(n33930), .Z(n33932) );
  XOR U35673 ( .A(n33933), .B(mreg[669]), .Z(n33930) );
  NAND U35674 ( .A(n33934), .B(mul_pow), .Z(n33933) );
  XOR U35675 ( .A(mreg[669]), .B(creg[669]), .Z(n33934) );
  XOR U35676 ( .A(n33935), .B(n33936), .Z(n33926) );
  ANDN U35677 ( .A(n33937), .B(n26735), .Z(n33936) );
  XOR U35678 ( .A(n33938), .B(\modmult_1/zin[0][667] ), .Z(n26735) );
  IV U35679 ( .A(n33935), .Z(n33938) );
  XNOR U35680 ( .A(n33935), .B(n26734), .Z(n33937) );
  XOR U35681 ( .A(n33939), .B(n33940), .Z(n26734) );
  AND U35682 ( .A(\modmult_1/xin[1023] ), .B(n33941), .Z(n33940) );
  IV U35683 ( .A(n33939), .Z(n33941) );
  XOR U35684 ( .A(n33942), .B(mreg[668]), .Z(n33939) );
  NAND U35685 ( .A(n33943), .B(mul_pow), .Z(n33942) );
  XOR U35686 ( .A(mreg[668]), .B(creg[668]), .Z(n33943) );
  XOR U35687 ( .A(n33944), .B(n33945), .Z(n33935) );
  ANDN U35688 ( .A(n33946), .B(n26741), .Z(n33945) );
  XOR U35689 ( .A(n33947), .B(\modmult_1/zin[0][666] ), .Z(n26741) );
  IV U35690 ( .A(n33944), .Z(n33947) );
  XNOR U35691 ( .A(n33944), .B(n26740), .Z(n33946) );
  XOR U35692 ( .A(n33948), .B(n33949), .Z(n26740) );
  AND U35693 ( .A(\modmult_1/xin[1023] ), .B(n33950), .Z(n33949) );
  IV U35694 ( .A(n33948), .Z(n33950) );
  XOR U35695 ( .A(n33951), .B(mreg[667]), .Z(n33948) );
  NAND U35696 ( .A(n33952), .B(mul_pow), .Z(n33951) );
  XOR U35697 ( .A(mreg[667]), .B(creg[667]), .Z(n33952) );
  XOR U35698 ( .A(n33953), .B(n33954), .Z(n33944) );
  ANDN U35699 ( .A(n33955), .B(n26747), .Z(n33954) );
  XOR U35700 ( .A(n33956), .B(\modmult_1/zin[0][665] ), .Z(n26747) );
  IV U35701 ( .A(n33953), .Z(n33956) );
  XNOR U35702 ( .A(n33953), .B(n26746), .Z(n33955) );
  XOR U35703 ( .A(n33957), .B(n33958), .Z(n26746) );
  AND U35704 ( .A(\modmult_1/xin[1023] ), .B(n33959), .Z(n33958) );
  IV U35705 ( .A(n33957), .Z(n33959) );
  XOR U35706 ( .A(n33960), .B(mreg[666]), .Z(n33957) );
  NAND U35707 ( .A(n33961), .B(mul_pow), .Z(n33960) );
  XOR U35708 ( .A(mreg[666]), .B(creg[666]), .Z(n33961) );
  XOR U35709 ( .A(n33962), .B(n33963), .Z(n33953) );
  ANDN U35710 ( .A(n33964), .B(n26753), .Z(n33963) );
  XOR U35711 ( .A(n33965), .B(\modmult_1/zin[0][664] ), .Z(n26753) );
  IV U35712 ( .A(n33962), .Z(n33965) );
  XNOR U35713 ( .A(n33962), .B(n26752), .Z(n33964) );
  XOR U35714 ( .A(n33966), .B(n33967), .Z(n26752) );
  AND U35715 ( .A(\modmult_1/xin[1023] ), .B(n33968), .Z(n33967) );
  IV U35716 ( .A(n33966), .Z(n33968) );
  XOR U35717 ( .A(n33969), .B(mreg[665]), .Z(n33966) );
  NAND U35718 ( .A(n33970), .B(mul_pow), .Z(n33969) );
  XOR U35719 ( .A(mreg[665]), .B(creg[665]), .Z(n33970) );
  XOR U35720 ( .A(n33971), .B(n33972), .Z(n33962) );
  ANDN U35721 ( .A(n33973), .B(n26759), .Z(n33972) );
  XOR U35722 ( .A(n33974), .B(\modmult_1/zin[0][663] ), .Z(n26759) );
  IV U35723 ( .A(n33971), .Z(n33974) );
  XNOR U35724 ( .A(n33971), .B(n26758), .Z(n33973) );
  XOR U35725 ( .A(n33975), .B(n33976), .Z(n26758) );
  AND U35726 ( .A(\modmult_1/xin[1023] ), .B(n33977), .Z(n33976) );
  IV U35727 ( .A(n33975), .Z(n33977) );
  XOR U35728 ( .A(n33978), .B(mreg[664]), .Z(n33975) );
  NAND U35729 ( .A(n33979), .B(mul_pow), .Z(n33978) );
  XOR U35730 ( .A(mreg[664]), .B(creg[664]), .Z(n33979) );
  XOR U35731 ( .A(n33980), .B(n33981), .Z(n33971) );
  ANDN U35732 ( .A(n33982), .B(n26765), .Z(n33981) );
  XOR U35733 ( .A(n33983), .B(\modmult_1/zin[0][662] ), .Z(n26765) );
  IV U35734 ( .A(n33980), .Z(n33983) );
  XNOR U35735 ( .A(n33980), .B(n26764), .Z(n33982) );
  XOR U35736 ( .A(n33984), .B(n33985), .Z(n26764) );
  AND U35737 ( .A(\modmult_1/xin[1023] ), .B(n33986), .Z(n33985) );
  IV U35738 ( .A(n33984), .Z(n33986) );
  XOR U35739 ( .A(n33987), .B(mreg[663]), .Z(n33984) );
  NAND U35740 ( .A(n33988), .B(mul_pow), .Z(n33987) );
  XOR U35741 ( .A(mreg[663]), .B(creg[663]), .Z(n33988) );
  XOR U35742 ( .A(n33989), .B(n33990), .Z(n33980) );
  ANDN U35743 ( .A(n33991), .B(n26771), .Z(n33990) );
  XOR U35744 ( .A(n33992), .B(\modmult_1/zin[0][661] ), .Z(n26771) );
  IV U35745 ( .A(n33989), .Z(n33992) );
  XNOR U35746 ( .A(n33989), .B(n26770), .Z(n33991) );
  XOR U35747 ( .A(n33993), .B(n33994), .Z(n26770) );
  AND U35748 ( .A(\modmult_1/xin[1023] ), .B(n33995), .Z(n33994) );
  IV U35749 ( .A(n33993), .Z(n33995) );
  XOR U35750 ( .A(n33996), .B(mreg[662]), .Z(n33993) );
  NAND U35751 ( .A(n33997), .B(mul_pow), .Z(n33996) );
  XOR U35752 ( .A(mreg[662]), .B(creg[662]), .Z(n33997) );
  XOR U35753 ( .A(n33998), .B(n33999), .Z(n33989) );
  ANDN U35754 ( .A(n34000), .B(n26777), .Z(n33999) );
  XOR U35755 ( .A(n34001), .B(\modmult_1/zin[0][660] ), .Z(n26777) );
  IV U35756 ( .A(n33998), .Z(n34001) );
  XNOR U35757 ( .A(n33998), .B(n26776), .Z(n34000) );
  XOR U35758 ( .A(n34002), .B(n34003), .Z(n26776) );
  AND U35759 ( .A(\modmult_1/xin[1023] ), .B(n34004), .Z(n34003) );
  IV U35760 ( .A(n34002), .Z(n34004) );
  XOR U35761 ( .A(n34005), .B(mreg[661]), .Z(n34002) );
  NAND U35762 ( .A(n34006), .B(mul_pow), .Z(n34005) );
  XOR U35763 ( .A(mreg[661]), .B(creg[661]), .Z(n34006) );
  XOR U35764 ( .A(n34007), .B(n34008), .Z(n33998) );
  ANDN U35765 ( .A(n34009), .B(n26783), .Z(n34008) );
  XOR U35766 ( .A(n34010), .B(\modmult_1/zin[0][659] ), .Z(n26783) );
  IV U35767 ( .A(n34007), .Z(n34010) );
  XNOR U35768 ( .A(n34007), .B(n26782), .Z(n34009) );
  XOR U35769 ( .A(n34011), .B(n34012), .Z(n26782) );
  AND U35770 ( .A(\modmult_1/xin[1023] ), .B(n34013), .Z(n34012) );
  IV U35771 ( .A(n34011), .Z(n34013) );
  XOR U35772 ( .A(n34014), .B(mreg[660]), .Z(n34011) );
  NAND U35773 ( .A(n34015), .B(mul_pow), .Z(n34014) );
  XOR U35774 ( .A(mreg[660]), .B(creg[660]), .Z(n34015) );
  XOR U35775 ( .A(n34016), .B(n34017), .Z(n34007) );
  ANDN U35776 ( .A(n34018), .B(n26789), .Z(n34017) );
  XOR U35777 ( .A(n34019), .B(\modmult_1/zin[0][658] ), .Z(n26789) );
  IV U35778 ( .A(n34016), .Z(n34019) );
  XNOR U35779 ( .A(n34016), .B(n26788), .Z(n34018) );
  XOR U35780 ( .A(n34020), .B(n34021), .Z(n26788) );
  AND U35781 ( .A(\modmult_1/xin[1023] ), .B(n34022), .Z(n34021) );
  IV U35782 ( .A(n34020), .Z(n34022) );
  XOR U35783 ( .A(n34023), .B(mreg[659]), .Z(n34020) );
  NAND U35784 ( .A(n34024), .B(mul_pow), .Z(n34023) );
  XOR U35785 ( .A(mreg[659]), .B(creg[659]), .Z(n34024) );
  XOR U35786 ( .A(n34025), .B(n34026), .Z(n34016) );
  ANDN U35787 ( .A(n34027), .B(n26795), .Z(n34026) );
  XOR U35788 ( .A(n34028), .B(\modmult_1/zin[0][657] ), .Z(n26795) );
  IV U35789 ( .A(n34025), .Z(n34028) );
  XNOR U35790 ( .A(n34025), .B(n26794), .Z(n34027) );
  XOR U35791 ( .A(n34029), .B(n34030), .Z(n26794) );
  AND U35792 ( .A(\modmult_1/xin[1023] ), .B(n34031), .Z(n34030) );
  IV U35793 ( .A(n34029), .Z(n34031) );
  XOR U35794 ( .A(n34032), .B(mreg[658]), .Z(n34029) );
  NAND U35795 ( .A(n34033), .B(mul_pow), .Z(n34032) );
  XOR U35796 ( .A(mreg[658]), .B(creg[658]), .Z(n34033) );
  XOR U35797 ( .A(n34034), .B(n34035), .Z(n34025) );
  ANDN U35798 ( .A(n34036), .B(n26801), .Z(n34035) );
  XOR U35799 ( .A(n34037), .B(\modmult_1/zin[0][656] ), .Z(n26801) );
  IV U35800 ( .A(n34034), .Z(n34037) );
  XNOR U35801 ( .A(n34034), .B(n26800), .Z(n34036) );
  XOR U35802 ( .A(n34038), .B(n34039), .Z(n26800) );
  AND U35803 ( .A(\modmult_1/xin[1023] ), .B(n34040), .Z(n34039) );
  IV U35804 ( .A(n34038), .Z(n34040) );
  XOR U35805 ( .A(n34041), .B(mreg[657]), .Z(n34038) );
  NAND U35806 ( .A(n34042), .B(mul_pow), .Z(n34041) );
  XOR U35807 ( .A(mreg[657]), .B(creg[657]), .Z(n34042) );
  XOR U35808 ( .A(n34043), .B(n34044), .Z(n34034) );
  ANDN U35809 ( .A(n34045), .B(n26807), .Z(n34044) );
  XOR U35810 ( .A(n34046), .B(\modmult_1/zin[0][655] ), .Z(n26807) );
  IV U35811 ( .A(n34043), .Z(n34046) );
  XNOR U35812 ( .A(n34043), .B(n26806), .Z(n34045) );
  XOR U35813 ( .A(n34047), .B(n34048), .Z(n26806) );
  AND U35814 ( .A(\modmult_1/xin[1023] ), .B(n34049), .Z(n34048) );
  IV U35815 ( .A(n34047), .Z(n34049) );
  XOR U35816 ( .A(n34050), .B(mreg[656]), .Z(n34047) );
  NAND U35817 ( .A(n34051), .B(mul_pow), .Z(n34050) );
  XOR U35818 ( .A(mreg[656]), .B(creg[656]), .Z(n34051) );
  XOR U35819 ( .A(n34052), .B(n34053), .Z(n34043) );
  ANDN U35820 ( .A(n34054), .B(n26813), .Z(n34053) );
  XOR U35821 ( .A(n34055), .B(\modmult_1/zin[0][654] ), .Z(n26813) );
  IV U35822 ( .A(n34052), .Z(n34055) );
  XNOR U35823 ( .A(n34052), .B(n26812), .Z(n34054) );
  XOR U35824 ( .A(n34056), .B(n34057), .Z(n26812) );
  AND U35825 ( .A(\modmult_1/xin[1023] ), .B(n34058), .Z(n34057) );
  IV U35826 ( .A(n34056), .Z(n34058) );
  XOR U35827 ( .A(n34059), .B(mreg[655]), .Z(n34056) );
  NAND U35828 ( .A(n34060), .B(mul_pow), .Z(n34059) );
  XOR U35829 ( .A(mreg[655]), .B(creg[655]), .Z(n34060) );
  XOR U35830 ( .A(n34061), .B(n34062), .Z(n34052) );
  ANDN U35831 ( .A(n34063), .B(n26819), .Z(n34062) );
  XOR U35832 ( .A(n34064), .B(\modmult_1/zin[0][653] ), .Z(n26819) );
  IV U35833 ( .A(n34061), .Z(n34064) );
  XNOR U35834 ( .A(n34061), .B(n26818), .Z(n34063) );
  XOR U35835 ( .A(n34065), .B(n34066), .Z(n26818) );
  AND U35836 ( .A(\modmult_1/xin[1023] ), .B(n34067), .Z(n34066) );
  IV U35837 ( .A(n34065), .Z(n34067) );
  XOR U35838 ( .A(n34068), .B(mreg[654]), .Z(n34065) );
  NAND U35839 ( .A(n34069), .B(mul_pow), .Z(n34068) );
  XOR U35840 ( .A(mreg[654]), .B(creg[654]), .Z(n34069) );
  XOR U35841 ( .A(n34070), .B(n34071), .Z(n34061) );
  ANDN U35842 ( .A(n34072), .B(n26825), .Z(n34071) );
  XOR U35843 ( .A(n34073), .B(\modmult_1/zin[0][652] ), .Z(n26825) );
  IV U35844 ( .A(n34070), .Z(n34073) );
  XNOR U35845 ( .A(n34070), .B(n26824), .Z(n34072) );
  XOR U35846 ( .A(n34074), .B(n34075), .Z(n26824) );
  AND U35847 ( .A(\modmult_1/xin[1023] ), .B(n34076), .Z(n34075) );
  IV U35848 ( .A(n34074), .Z(n34076) );
  XOR U35849 ( .A(n34077), .B(mreg[653]), .Z(n34074) );
  NAND U35850 ( .A(n34078), .B(mul_pow), .Z(n34077) );
  XOR U35851 ( .A(mreg[653]), .B(creg[653]), .Z(n34078) );
  XOR U35852 ( .A(n34079), .B(n34080), .Z(n34070) );
  ANDN U35853 ( .A(n34081), .B(n26831), .Z(n34080) );
  XOR U35854 ( .A(n34082), .B(\modmult_1/zin[0][651] ), .Z(n26831) );
  IV U35855 ( .A(n34079), .Z(n34082) );
  XNOR U35856 ( .A(n34079), .B(n26830), .Z(n34081) );
  XOR U35857 ( .A(n34083), .B(n34084), .Z(n26830) );
  AND U35858 ( .A(\modmult_1/xin[1023] ), .B(n34085), .Z(n34084) );
  IV U35859 ( .A(n34083), .Z(n34085) );
  XOR U35860 ( .A(n34086), .B(mreg[652]), .Z(n34083) );
  NAND U35861 ( .A(n34087), .B(mul_pow), .Z(n34086) );
  XOR U35862 ( .A(mreg[652]), .B(creg[652]), .Z(n34087) );
  XOR U35863 ( .A(n34088), .B(n34089), .Z(n34079) );
  ANDN U35864 ( .A(n34090), .B(n26837), .Z(n34089) );
  XOR U35865 ( .A(n34091), .B(\modmult_1/zin[0][650] ), .Z(n26837) );
  IV U35866 ( .A(n34088), .Z(n34091) );
  XNOR U35867 ( .A(n34088), .B(n26836), .Z(n34090) );
  XOR U35868 ( .A(n34092), .B(n34093), .Z(n26836) );
  AND U35869 ( .A(\modmult_1/xin[1023] ), .B(n34094), .Z(n34093) );
  IV U35870 ( .A(n34092), .Z(n34094) );
  XOR U35871 ( .A(n34095), .B(mreg[651]), .Z(n34092) );
  NAND U35872 ( .A(n34096), .B(mul_pow), .Z(n34095) );
  XOR U35873 ( .A(mreg[651]), .B(creg[651]), .Z(n34096) );
  XOR U35874 ( .A(n34097), .B(n34098), .Z(n34088) );
  ANDN U35875 ( .A(n34099), .B(n26843), .Z(n34098) );
  XOR U35876 ( .A(n34100), .B(\modmult_1/zin[0][649] ), .Z(n26843) );
  IV U35877 ( .A(n34097), .Z(n34100) );
  XNOR U35878 ( .A(n34097), .B(n26842), .Z(n34099) );
  XOR U35879 ( .A(n34101), .B(n34102), .Z(n26842) );
  AND U35880 ( .A(\modmult_1/xin[1023] ), .B(n34103), .Z(n34102) );
  IV U35881 ( .A(n34101), .Z(n34103) );
  XOR U35882 ( .A(n34104), .B(mreg[650]), .Z(n34101) );
  NAND U35883 ( .A(n34105), .B(mul_pow), .Z(n34104) );
  XOR U35884 ( .A(mreg[650]), .B(creg[650]), .Z(n34105) );
  XOR U35885 ( .A(n34106), .B(n34107), .Z(n34097) );
  ANDN U35886 ( .A(n34108), .B(n26849), .Z(n34107) );
  XOR U35887 ( .A(n34109), .B(\modmult_1/zin[0][648] ), .Z(n26849) );
  IV U35888 ( .A(n34106), .Z(n34109) );
  XNOR U35889 ( .A(n34106), .B(n26848), .Z(n34108) );
  XOR U35890 ( .A(n34110), .B(n34111), .Z(n26848) );
  AND U35891 ( .A(\modmult_1/xin[1023] ), .B(n34112), .Z(n34111) );
  IV U35892 ( .A(n34110), .Z(n34112) );
  XOR U35893 ( .A(n34113), .B(mreg[649]), .Z(n34110) );
  NAND U35894 ( .A(n34114), .B(mul_pow), .Z(n34113) );
  XOR U35895 ( .A(mreg[649]), .B(creg[649]), .Z(n34114) );
  XOR U35896 ( .A(n34115), .B(n34116), .Z(n34106) );
  ANDN U35897 ( .A(n34117), .B(n26855), .Z(n34116) );
  XOR U35898 ( .A(n34118), .B(\modmult_1/zin[0][647] ), .Z(n26855) );
  IV U35899 ( .A(n34115), .Z(n34118) );
  XNOR U35900 ( .A(n34115), .B(n26854), .Z(n34117) );
  XOR U35901 ( .A(n34119), .B(n34120), .Z(n26854) );
  AND U35902 ( .A(\modmult_1/xin[1023] ), .B(n34121), .Z(n34120) );
  IV U35903 ( .A(n34119), .Z(n34121) );
  XOR U35904 ( .A(n34122), .B(mreg[648]), .Z(n34119) );
  NAND U35905 ( .A(n34123), .B(mul_pow), .Z(n34122) );
  XOR U35906 ( .A(mreg[648]), .B(creg[648]), .Z(n34123) );
  XOR U35907 ( .A(n34124), .B(n34125), .Z(n34115) );
  ANDN U35908 ( .A(n34126), .B(n26861), .Z(n34125) );
  XOR U35909 ( .A(n34127), .B(\modmult_1/zin[0][646] ), .Z(n26861) );
  IV U35910 ( .A(n34124), .Z(n34127) );
  XNOR U35911 ( .A(n34124), .B(n26860), .Z(n34126) );
  XOR U35912 ( .A(n34128), .B(n34129), .Z(n26860) );
  AND U35913 ( .A(\modmult_1/xin[1023] ), .B(n34130), .Z(n34129) );
  IV U35914 ( .A(n34128), .Z(n34130) );
  XOR U35915 ( .A(n34131), .B(mreg[647]), .Z(n34128) );
  NAND U35916 ( .A(n34132), .B(mul_pow), .Z(n34131) );
  XOR U35917 ( .A(mreg[647]), .B(creg[647]), .Z(n34132) );
  XOR U35918 ( .A(n34133), .B(n34134), .Z(n34124) );
  ANDN U35919 ( .A(n34135), .B(n26867), .Z(n34134) );
  XOR U35920 ( .A(n34136), .B(\modmult_1/zin[0][645] ), .Z(n26867) );
  IV U35921 ( .A(n34133), .Z(n34136) );
  XNOR U35922 ( .A(n34133), .B(n26866), .Z(n34135) );
  XOR U35923 ( .A(n34137), .B(n34138), .Z(n26866) );
  AND U35924 ( .A(\modmult_1/xin[1023] ), .B(n34139), .Z(n34138) );
  IV U35925 ( .A(n34137), .Z(n34139) );
  XOR U35926 ( .A(n34140), .B(mreg[646]), .Z(n34137) );
  NAND U35927 ( .A(n34141), .B(mul_pow), .Z(n34140) );
  XOR U35928 ( .A(mreg[646]), .B(creg[646]), .Z(n34141) );
  XOR U35929 ( .A(n34142), .B(n34143), .Z(n34133) );
  ANDN U35930 ( .A(n34144), .B(n26873), .Z(n34143) );
  XOR U35931 ( .A(n34145), .B(\modmult_1/zin[0][644] ), .Z(n26873) );
  IV U35932 ( .A(n34142), .Z(n34145) );
  XNOR U35933 ( .A(n34142), .B(n26872), .Z(n34144) );
  XOR U35934 ( .A(n34146), .B(n34147), .Z(n26872) );
  AND U35935 ( .A(\modmult_1/xin[1023] ), .B(n34148), .Z(n34147) );
  IV U35936 ( .A(n34146), .Z(n34148) );
  XOR U35937 ( .A(n34149), .B(mreg[645]), .Z(n34146) );
  NAND U35938 ( .A(n34150), .B(mul_pow), .Z(n34149) );
  XOR U35939 ( .A(mreg[645]), .B(creg[645]), .Z(n34150) );
  XOR U35940 ( .A(n34151), .B(n34152), .Z(n34142) );
  ANDN U35941 ( .A(n34153), .B(n26879), .Z(n34152) );
  XOR U35942 ( .A(n34154), .B(\modmult_1/zin[0][643] ), .Z(n26879) );
  IV U35943 ( .A(n34151), .Z(n34154) );
  XNOR U35944 ( .A(n34151), .B(n26878), .Z(n34153) );
  XOR U35945 ( .A(n34155), .B(n34156), .Z(n26878) );
  AND U35946 ( .A(\modmult_1/xin[1023] ), .B(n34157), .Z(n34156) );
  IV U35947 ( .A(n34155), .Z(n34157) );
  XOR U35948 ( .A(n34158), .B(mreg[644]), .Z(n34155) );
  NAND U35949 ( .A(n34159), .B(mul_pow), .Z(n34158) );
  XOR U35950 ( .A(mreg[644]), .B(creg[644]), .Z(n34159) );
  XOR U35951 ( .A(n34160), .B(n34161), .Z(n34151) );
  ANDN U35952 ( .A(n34162), .B(n26885), .Z(n34161) );
  XOR U35953 ( .A(n34163), .B(\modmult_1/zin[0][642] ), .Z(n26885) );
  IV U35954 ( .A(n34160), .Z(n34163) );
  XNOR U35955 ( .A(n34160), .B(n26884), .Z(n34162) );
  XOR U35956 ( .A(n34164), .B(n34165), .Z(n26884) );
  AND U35957 ( .A(\modmult_1/xin[1023] ), .B(n34166), .Z(n34165) );
  IV U35958 ( .A(n34164), .Z(n34166) );
  XOR U35959 ( .A(n34167), .B(mreg[643]), .Z(n34164) );
  NAND U35960 ( .A(n34168), .B(mul_pow), .Z(n34167) );
  XOR U35961 ( .A(mreg[643]), .B(creg[643]), .Z(n34168) );
  XOR U35962 ( .A(n34169), .B(n34170), .Z(n34160) );
  ANDN U35963 ( .A(n34171), .B(n26891), .Z(n34170) );
  XOR U35964 ( .A(n34172), .B(\modmult_1/zin[0][641] ), .Z(n26891) );
  IV U35965 ( .A(n34169), .Z(n34172) );
  XNOR U35966 ( .A(n34169), .B(n26890), .Z(n34171) );
  XOR U35967 ( .A(n34173), .B(n34174), .Z(n26890) );
  AND U35968 ( .A(\modmult_1/xin[1023] ), .B(n34175), .Z(n34174) );
  IV U35969 ( .A(n34173), .Z(n34175) );
  XOR U35970 ( .A(n34176), .B(mreg[642]), .Z(n34173) );
  NAND U35971 ( .A(n34177), .B(mul_pow), .Z(n34176) );
  XOR U35972 ( .A(mreg[642]), .B(creg[642]), .Z(n34177) );
  XOR U35973 ( .A(n34178), .B(n34179), .Z(n34169) );
  ANDN U35974 ( .A(n34180), .B(n26897), .Z(n34179) );
  XOR U35975 ( .A(n34181), .B(\modmult_1/zin[0][640] ), .Z(n26897) );
  IV U35976 ( .A(n34178), .Z(n34181) );
  XNOR U35977 ( .A(n34178), .B(n26896), .Z(n34180) );
  XOR U35978 ( .A(n34182), .B(n34183), .Z(n26896) );
  AND U35979 ( .A(\modmult_1/xin[1023] ), .B(n34184), .Z(n34183) );
  IV U35980 ( .A(n34182), .Z(n34184) );
  XOR U35981 ( .A(n34185), .B(mreg[641]), .Z(n34182) );
  NAND U35982 ( .A(n34186), .B(mul_pow), .Z(n34185) );
  XOR U35983 ( .A(mreg[641]), .B(creg[641]), .Z(n34186) );
  XOR U35984 ( .A(n34187), .B(n34188), .Z(n34178) );
  ANDN U35985 ( .A(n34189), .B(n26903), .Z(n34188) );
  XOR U35986 ( .A(n34190), .B(\modmult_1/zin[0][639] ), .Z(n26903) );
  IV U35987 ( .A(n34187), .Z(n34190) );
  XNOR U35988 ( .A(n34187), .B(n26902), .Z(n34189) );
  XOR U35989 ( .A(n34191), .B(n34192), .Z(n26902) );
  AND U35990 ( .A(\modmult_1/xin[1023] ), .B(n34193), .Z(n34192) );
  IV U35991 ( .A(n34191), .Z(n34193) );
  XOR U35992 ( .A(n34194), .B(mreg[640]), .Z(n34191) );
  NAND U35993 ( .A(n34195), .B(mul_pow), .Z(n34194) );
  XOR U35994 ( .A(mreg[640]), .B(creg[640]), .Z(n34195) );
  XOR U35995 ( .A(n34196), .B(n34197), .Z(n34187) );
  ANDN U35996 ( .A(n34198), .B(n26909), .Z(n34197) );
  XOR U35997 ( .A(n34199), .B(\modmult_1/zin[0][638] ), .Z(n26909) );
  IV U35998 ( .A(n34196), .Z(n34199) );
  XNOR U35999 ( .A(n34196), .B(n26908), .Z(n34198) );
  XOR U36000 ( .A(n34200), .B(n34201), .Z(n26908) );
  AND U36001 ( .A(\modmult_1/xin[1023] ), .B(n34202), .Z(n34201) );
  IV U36002 ( .A(n34200), .Z(n34202) );
  XOR U36003 ( .A(n34203), .B(mreg[639]), .Z(n34200) );
  NAND U36004 ( .A(n34204), .B(mul_pow), .Z(n34203) );
  XOR U36005 ( .A(mreg[639]), .B(creg[639]), .Z(n34204) );
  XOR U36006 ( .A(n34205), .B(n34206), .Z(n34196) );
  ANDN U36007 ( .A(n34207), .B(n26915), .Z(n34206) );
  XOR U36008 ( .A(n34208), .B(\modmult_1/zin[0][637] ), .Z(n26915) );
  IV U36009 ( .A(n34205), .Z(n34208) );
  XNOR U36010 ( .A(n34205), .B(n26914), .Z(n34207) );
  XOR U36011 ( .A(n34209), .B(n34210), .Z(n26914) );
  AND U36012 ( .A(\modmult_1/xin[1023] ), .B(n34211), .Z(n34210) );
  IV U36013 ( .A(n34209), .Z(n34211) );
  XOR U36014 ( .A(n34212), .B(mreg[638]), .Z(n34209) );
  NAND U36015 ( .A(n34213), .B(mul_pow), .Z(n34212) );
  XOR U36016 ( .A(mreg[638]), .B(creg[638]), .Z(n34213) );
  XOR U36017 ( .A(n34214), .B(n34215), .Z(n34205) );
  ANDN U36018 ( .A(n34216), .B(n26921), .Z(n34215) );
  XOR U36019 ( .A(n34217), .B(\modmult_1/zin[0][636] ), .Z(n26921) );
  IV U36020 ( .A(n34214), .Z(n34217) );
  XNOR U36021 ( .A(n34214), .B(n26920), .Z(n34216) );
  XOR U36022 ( .A(n34218), .B(n34219), .Z(n26920) );
  AND U36023 ( .A(\modmult_1/xin[1023] ), .B(n34220), .Z(n34219) );
  IV U36024 ( .A(n34218), .Z(n34220) );
  XOR U36025 ( .A(n34221), .B(mreg[637]), .Z(n34218) );
  NAND U36026 ( .A(n34222), .B(mul_pow), .Z(n34221) );
  XOR U36027 ( .A(mreg[637]), .B(creg[637]), .Z(n34222) );
  XOR U36028 ( .A(n34223), .B(n34224), .Z(n34214) );
  ANDN U36029 ( .A(n34225), .B(n26927), .Z(n34224) );
  XOR U36030 ( .A(n34226), .B(\modmult_1/zin[0][635] ), .Z(n26927) );
  IV U36031 ( .A(n34223), .Z(n34226) );
  XNOR U36032 ( .A(n34223), .B(n26926), .Z(n34225) );
  XOR U36033 ( .A(n34227), .B(n34228), .Z(n26926) );
  AND U36034 ( .A(\modmult_1/xin[1023] ), .B(n34229), .Z(n34228) );
  IV U36035 ( .A(n34227), .Z(n34229) );
  XOR U36036 ( .A(n34230), .B(mreg[636]), .Z(n34227) );
  NAND U36037 ( .A(n34231), .B(mul_pow), .Z(n34230) );
  XOR U36038 ( .A(mreg[636]), .B(creg[636]), .Z(n34231) );
  XOR U36039 ( .A(n34232), .B(n34233), .Z(n34223) );
  ANDN U36040 ( .A(n34234), .B(n26933), .Z(n34233) );
  XOR U36041 ( .A(n34235), .B(\modmult_1/zin[0][634] ), .Z(n26933) );
  IV U36042 ( .A(n34232), .Z(n34235) );
  XNOR U36043 ( .A(n34232), .B(n26932), .Z(n34234) );
  XOR U36044 ( .A(n34236), .B(n34237), .Z(n26932) );
  AND U36045 ( .A(\modmult_1/xin[1023] ), .B(n34238), .Z(n34237) );
  IV U36046 ( .A(n34236), .Z(n34238) );
  XOR U36047 ( .A(n34239), .B(mreg[635]), .Z(n34236) );
  NAND U36048 ( .A(n34240), .B(mul_pow), .Z(n34239) );
  XOR U36049 ( .A(mreg[635]), .B(creg[635]), .Z(n34240) );
  XOR U36050 ( .A(n34241), .B(n34242), .Z(n34232) );
  ANDN U36051 ( .A(n34243), .B(n26939), .Z(n34242) );
  XOR U36052 ( .A(n34244), .B(\modmult_1/zin[0][633] ), .Z(n26939) );
  IV U36053 ( .A(n34241), .Z(n34244) );
  XNOR U36054 ( .A(n34241), .B(n26938), .Z(n34243) );
  XOR U36055 ( .A(n34245), .B(n34246), .Z(n26938) );
  AND U36056 ( .A(\modmult_1/xin[1023] ), .B(n34247), .Z(n34246) );
  IV U36057 ( .A(n34245), .Z(n34247) );
  XOR U36058 ( .A(n34248), .B(mreg[634]), .Z(n34245) );
  NAND U36059 ( .A(n34249), .B(mul_pow), .Z(n34248) );
  XOR U36060 ( .A(mreg[634]), .B(creg[634]), .Z(n34249) );
  XOR U36061 ( .A(n34250), .B(n34251), .Z(n34241) );
  ANDN U36062 ( .A(n34252), .B(n26945), .Z(n34251) );
  XOR U36063 ( .A(n34253), .B(\modmult_1/zin[0][632] ), .Z(n26945) );
  IV U36064 ( .A(n34250), .Z(n34253) );
  XNOR U36065 ( .A(n34250), .B(n26944), .Z(n34252) );
  XOR U36066 ( .A(n34254), .B(n34255), .Z(n26944) );
  AND U36067 ( .A(\modmult_1/xin[1023] ), .B(n34256), .Z(n34255) );
  IV U36068 ( .A(n34254), .Z(n34256) );
  XOR U36069 ( .A(n34257), .B(mreg[633]), .Z(n34254) );
  NAND U36070 ( .A(n34258), .B(mul_pow), .Z(n34257) );
  XOR U36071 ( .A(mreg[633]), .B(creg[633]), .Z(n34258) );
  XOR U36072 ( .A(n34259), .B(n34260), .Z(n34250) );
  ANDN U36073 ( .A(n34261), .B(n26951), .Z(n34260) );
  XOR U36074 ( .A(n34262), .B(\modmult_1/zin[0][631] ), .Z(n26951) );
  IV U36075 ( .A(n34259), .Z(n34262) );
  XNOR U36076 ( .A(n34259), .B(n26950), .Z(n34261) );
  XOR U36077 ( .A(n34263), .B(n34264), .Z(n26950) );
  AND U36078 ( .A(\modmult_1/xin[1023] ), .B(n34265), .Z(n34264) );
  IV U36079 ( .A(n34263), .Z(n34265) );
  XOR U36080 ( .A(n34266), .B(mreg[632]), .Z(n34263) );
  NAND U36081 ( .A(n34267), .B(mul_pow), .Z(n34266) );
  XOR U36082 ( .A(mreg[632]), .B(creg[632]), .Z(n34267) );
  XOR U36083 ( .A(n34268), .B(n34269), .Z(n34259) );
  ANDN U36084 ( .A(n34270), .B(n26957), .Z(n34269) );
  XOR U36085 ( .A(n34271), .B(\modmult_1/zin[0][630] ), .Z(n26957) );
  IV U36086 ( .A(n34268), .Z(n34271) );
  XNOR U36087 ( .A(n34268), .B(n26956), .Z(n34270) );
  XOR U36088 ( .A(n34272), .B(n34273), .Z(n26956) );
  AND U36089 ( .A(\modmult_1/xin[1023] ), .B(n34274), .Z(n34273) );
  IV U36090 ( .A(n34272), .Z(n34274) );
  XOR U36091 ( .A(n34275), .B(mreg[631]), .Z(n34272) );
  NAND U36092 ( .A(n34276), .B(mul_pow), .Z(n34275) );
  XOR U36093 ( .A(mreg[631]), .B(creg[631]), .Z(n34276) );
  XOR U36094 ( .A(n34277), .B(n34278), .Z(n34268) );
  ANDN U36095 ( .A(n34279), .B(n26963), .Z(n34278) );
  XOR U36096 ( .A(n34280), .B(\modmult_1/zin[0][629] ), .Z(n26963) );
  IV U36097 ( .A(n34277), .Z(n34280) );
  XNOR U36098 ( .A(n34277), .B(n26962), .Z(n34279) );
  XOR U36099 ( .A(n34281), .B(n34282), .Z(n26962) );
  AND U36100 ( .A(\modmult_1/xin[1023] ), .B(n34283), .Z(n34282) );
  IV U36101 ( .A(n34281), .Z(n34283) );
  XOR U36102 ( .A(n34284), .B(mreg[630]), .Z(n34281) );
  NAND U36103 ( .A(n34285), .B(mul_pow), .Z(n34284) );
  XOR U36104 ( .A(mreg[630]), .B(creg[630]), .Z(n34285) );
  XOR U36105 ( .A(n34286), .B(n34287), .Z(n34277) );
  ANDN U36106 ( .A(n34288), .B(n26969), .Z(n34287) );
  XOR U36107 ( .A(n34289), .B(\modmult_1/zin[0][628] ), .Z(n26969) );
  IV U36108 ( .A(n34286), .Z(n34289) );
  XNOR U36109 ( .A(n34286), .B(n26968), .Z(n34288) );
  XOR U36110 ( .A(n34290), .B(n34291), .Z(n26968) );
  AND U36111 ( .A(\modmult_1/xin[1023] ), .B(n34292), .Z(n34291) );
  IV U36112 ( .A(n34290), .Z(n34292) );
  XOR U36113 ( .A(n34293), .B(mreg[629]), .Z(n34290) );
  NAND U36114 ( .A(n34294), .B(mul_pow), .Z(n34293) );
  XOR U36115 ( .A(mreg[629]), .B(creg[629]), .Z(n34294) );
  XOR U36116 ( .A(n34295), .B(n34296), .Z(n34286) );
  ANDN U36117 ( .A(n34297), .B(n26975), .Z(n34296) );
  XOR U36118 ( .A(n34298), .B(\modmult_1/zin[0][627] ), .Z(n26975) );
  IV U36119 ( .A(n34295), .Z(n34298) );
  XNOR U36120 ( .A(n34295), .B(n26974), .Z(n34297) );
  XOR U36121 ( .A(n34299), .B(n34300), .Z(n26974) );
  AND U36122 ( .A(\modmult_1/xin[1023] ), .B(n34301), .Z(n34300) );
  IV U36123 ( .A(n34299), .Z(n34301) );
  XOR U36124 ( .A(n34302), .B(mreg[628]), .Z(n34299) );
  NAND U36125 ( .A(n34303), .B(mul_pow), .Z(n34302) );
  XOR U36126 ( .A(mreg[628]), .B(creg[628]), .Z(n34303) );
  XOR U36127 ( .A(n34304), .B(n34305), .Z(n34295) );
  ANDN U36128 ( .A(n34306), .B(n26981), .Z(n34305) );
  XOR U36129 ( .A(n34307), .B(\modmult_1/zin[0][626] ), .Z(n26981) );
  IV U36130 ( .A(n34304), .Z(n34307) );
  XNOR U36131 ( .A(n34304), .B(n26980), .Z(n34306) );
  XOR U36132 ( .A(n34308), .B(n34309), .Z(n26980) );
  AND U36133 ( .A(\modmult_1/xin[1023] ), .B(n34310), .Z(n34309) );
  IV U36134 ( .A(n34308), .Z(n34310) );
  XOR U36135 ( .A(n34311), .B(mreg[627]), .Z(n34308) );
  NAND U36136 ( .A(n34312), .B(mul_pow), .Z(n34311) );
  XOR U36137 ( .A(mreg[627]), .B(creg[627]), .Z(n34312) );
  XOR U36138 ( .A(n34313), .B(n34314), .Z(n34304) );
  ANDN U36139 ( .A(n34315), .B(n26987), .Z(n34314) );
  XOR U36140 ( .A(n34316), .B(\modmult_1/zin[0][625] ), .Z(n26987) );
  IV U36141 ( .A(n34313), .Z(n34316) );
  XNOR U36142 ( .A(n34313), .B(n26986), .Z(n34315) );
  XOR U36143 ( .A(n34317), .B(n34318), .Z(n26986) );
  AND U36144 ( .A(\modmult_1/xin[1023] ), .B(n34319), .Z(n34318) );
  IV U36145 ( .A(n34317), .Z(n34319) );
  XOR U36146 ( .A(n34320), .B(mreg[626]), .Z(n34317) );
  NAND U36147 ( .A(n34321), .B(mul_pow), .Z(n34320) );
  XOR U36148 ( .A(mreg[626]), .B(creg[626]), .Z(n34321) );
  XOR U36149 ( .A(n34322), .B(n34323), .Z(n34313) );
  ANDN U36150 ( .A(n34324), .B(n26993), .Z(n34323) );
  XOR U36151 ( .A(n34325), .B(\modmult_1/zin[0][624] ), .Z(n26993) );
  IV U36152 ( .A(n34322), .Z(n34325) );
  XNOR U36153 ( .A(n34322), .B(n26992), .Z(n34324) );
  XOR U36154 ( .A(n34326), .B(n34327), .Z(n26992) );
  AND U36155 ( .A(\modmult_1/xin[1023] ), .B(n34328), .Z(n34327) );
  IV U36156 ( .A(n34326), .Z(n34328) );
  XOR U36157 ( .A(n34329), .B(mreg[625]), .Z(n34326) );
  NAND U36158 ( .A(n34330), .B(mul_pow), .Z(n34329) );
  XOR U36159 ( .A(mreg[625]), .B(creg[625]), .Z(n34330) );
  XOR U36160 ( .A(n34331), .B(n34332), .Z(n34322) );
  ANDN U36161 ( .A(n34333), .B(n26999), .Z(n34332) );
  XOR U36162 ( .A(n34334), .B(\modmult_1/zin[0][623] ), .Z(n26999) );
  IV U36163 ( .A(n34331), .Z(n34334) );
  XNOR U36164 ( .A(n34331), .B(n26998), .Z(n34333) );
  XOR U36165 ( .A(n34335), .B(n34336), .Z(n26998) );
  AND U36166 ( .A(\modmult_1/xin[1023] ), .B(n34337), .Z(n34336) );
  IV U36167 ( .A(n34335), .Z(n34337) );
  XOR U36168 ( .A(n34338), .B(mreg[624]), .Z(n34335) );
  NAND U36169 ( .A(n34339), .B(mul_pow), .Z(n34338) );
  XOR U36170 ( .A(mreg[624]), .B(creg[624]), .Z(n34339) );
  XOR U36171 ( .A(n34340), .B(n34341), .Z(n34331) );
  ANDN U36172 ( .A(n34342), .B(n27005), .Z(n34341) );
  XOR U36173 ( .A(n34343), .B(\modmult_1/zin[0][622] ), .Z(n27005) );
  IV U36174 ( .A(n34340), .Z(n34343) );
  XNOR U36175 ( .A(n34340), .B(n27004), .Z(n34342) );
  XOR U36176 ( .A(n34344), .B(n34345), .Z(n27004) );
  AND U36177 ( .A(\modmult_1/xin[1023] ), .B(n34346), .Z(n34345) );
  IV U36178 ( .A(n34344), .Z(n34346) );
  XOR U36179 ( .A(n34347), .B(mreg[623]), .Z(n34344) );
  NAND U36180 ( .A(n34348), .B(mul_pow), .Z(n34347) );
  XOR U36181 ( .A(mreg[623]), .B(creg[623]), .Z(n34348) );
  XOR U36182 ( .A(n34349), .B(n34350), .Z(n34340) );
  ANDN U36183 ( .A(n34351), .B(n27011), .Z(n34350) );
  XOR U36184 ( .A(n34352), .B(\modmult_1/zin[0][621] ), .Z(n27011) );
  IV U36185 ( .A(n34349), .Z(n34352) );
  XNOR U36186 ( .A(n34349), .B(n27010), .Z(n34351) );
  XOR U36187 ( .A(n34353), .B(n34354), .Z(n27010) );
  AND U36188 ( .A(\modmult_1/xin[1023] ), .B(n34355), .Z(n34354) );
  IV U36189 ( .A(n34353), .Z(n34355) );
  XOR U36190 ( .A(n34356), .B(mreg[622]), .Z(n34353) );
  NAND U36191 ( .A(n34357), .B(mul_pow), .Z(n34356) );
  XOR U36192 ( .A(mreg[622]), .B(creg[622]), .Z(n34357) );
  XOR U36193 ( .A(n34358), .B(n34359), .Z(n34349) );
  ANDN U36194 ( .A(n34360), .B(n27017), .Z(n34359) );
  XOR U36195 ( .A(n34361), .B(\modmult_1/zin[0][620] ), .Z(n27017) );
  IV U36196 ( .A(n34358), .Z(n34361) );
  XNOR U36197 ( .A(n34358), .B(n27016), .Z(n34360) );
  XOR U36198 ( .A(n34362), .B(n34363), .Z(n27016) );
  AND U36199 ( .A(\modmult_1/xin[1023] ), .B(n34364), .Z(n34363) );
  IV U36200 ( .A(n34362), .Z(n34364) );
  XOR U36201 ( .A(n34365), .B(mreg[621]), .Z(n34362) );
  NAND U36202 ( .A(n34366), .B(mul_pow), .Z(n34365) );
  XOR U36203 ( .A(mreg[621]), .B(creg[621]), .Z(n34366) );
  XOR U36204 ( .A(n34367), .B(n34368), .Z(n34358) );
  ANDN U36205 ( .A(n34369), .B(n27023), .Z(n34368) );
  XOR U36206 ( .A(n34370), .B(\modmult_1/zin[0][619] ), .Z(n27023) );
  IV U36207 ( .A(n34367), .Z(n34370) );
  XNOR U36208 ( .A(n34367), .B(n27022), .Z(n34369) );
  XOR U36209 ( .A(n34371), .B(n34372), .Z(n27022) );
  AND U36210 ( .A(\modmult_1/xin[1023] ), .B(n34373), .Z(n34372) );
  IV U36211 ( .A(n34371), .Z(n34373) );
  XOR U36212 ( .A(n34374), .B(mreg[620]), .Z(n34371) );
  NAND U36213 ( .A(n34375), .B(mul_pow), .Z(n34374) );
  XOR U36214 ( .A(mreg[620]), .B(creg[620]), .Z(n34375) );
  XOR U36215 ( .A(n34376), .B(n34377), .Z(n34367) );
  ANDN U36216 ( .A(n34378), .B(n27029), .Z(n34377) );
  XOR U36217 ( .A(n34379), .B(\modmult_1/zin[0][618] ), .Z(n27029) );
  IV U36218 ( .A(n34376), .Z(n34379) );
  XNOR U36219 ( .A(n34376), .B(n27028), .Z(n34378) );
  XOR U36220 ( .A(n34380), .B(n34381), .Z(n27028) );
  AND U36221 ( .A(\modmult_1/xin[1023] ), .B(n34382), .Z(n34381) );
  IV U36222 ( .A(n34380), .Z(n34382) );
  XOR U36223 ( .A(n34383), .B(mreg[619]), .Z(n34380) );
  NAND U36224 ( .A(n34384), .B(mul_pow), .Z(n34383) );
  XOR U36225 ( .A(mreg[619]), .B(creg[619]), .Z(n34384) );
  XOR U36226 ( .A(n34385), .B(n34386), .Z(n34376) );
  ANDN U36227 ( .A(n34387), .B(n27035), .Z(n34386) );
  XOR U36228 ( .A(n34388), .B(\modmult_1/zin[0][617] ), .Z(n27035) );
  IV U36229 ( .A(n34385), .Z(n34388) );
  XNOR U36230 ( .A(n34385), .B(n27034), .Z(n34387) );
  XOR U36231 ( .A(n34389), .B(n34390), .Z(n27034) );
  AND U36232 ( .A(\modmult_1/xin[1023] ), .B(n34391), .Z(n34390) );
  IV U36233 ( .A(n34389), .Z(n34391) );
  XOR U36234 ( .A(n34392), .B(mreg[618]), .Z(n34389) );
  NAND U36235 ( .A(n34393), .B(mul_pow), .Z(n34392) );
  XOR U36236 ( .A(mreg[618]), .B(creg[618]), .Z(n34393) );
  XOR U36237 ( .A(n34394), .B(n34395), .Z(n34385) );
  ANDN U36238 ( .A(n34396), .B(n27041), .Z(n34395) );
  XOR U36239 ( .A(n34397), .B(\modmult_1/zin[0][616] ), .Z(n27041) );
  IV U36240 ( .A(n34394), .Z(n34397) );
  XNOR U36241 ( .A(n34394), .B(n27040), .Z(n34396) );
  XOR U36242 ( .A(n34398), .B(n34399), .Z(n27040) );
  AND U36243 ( .A(\modmult_1/xin[1023] ), .B(n34400), .Z(n34399) );
  IV U36244 ( .A(n34398), .Z(n34400) );
  XOR U36245 ( .A(n34401), .B(mreg[617]), .Z(n34398) );
  NAND U36246 ( .A(n34402), .B(mul_pow), .Z(n34401) );
  XOR U36247 ( .A(mreg[617]), .B(creg[617]), .Z(n34402) );
  XOR U36248 ( .A(n34403), .B(n34404), .Z(n34394) );
  ANDN U36249 ( .A(n34405), .B(n27047), .Z(n34404) );
  XOR U36250 ( .A(n34406), .B(\modmult_1/zin[0][615] ), .Z(n27047) );
  IV U36251 ( .A(n34403), .Z(n34406) );
  XNOR U36252 ( .A(n34403), .B(n27046), .Z(n34405) );
  XOR U36253 ( .A(n34407), .B(n34408), .Z(n27046) );
  AND U36254 ( .A(\modmult_1/xin[1023] ), .B(n34409), .Z(n34408) );
  IV U36255 ( .A(n34407), .Z(n34409) );
  XOR U36256 ( .A(n34410), .B(mreg[616]), .Z(n34407) );
  NAND U36257 ( .A(n34411), .B(mul_pow), .Z(n34410) );
  XOR U36258 ( .A(mreg[616]), .B(creg[616]), .Z(n34411) );
  XOR U36259 ( .A(n34412), .B(n34413), .Z(n34403) );
  ANDN U36260 ( .A(n34414), .B(n27053), .Z(n34413) );
  XOR U36261 ( .A(n34415), .B(\modmult_1/zin[0][614] ), .Z(n27053) );
  IV U36262 ( .A(n34412), .Z(n34415) );
  XNOR U36263 ( .A(n34412), .B(n27052), .Z(n34414) );
  XOR U36264 ( .A(n34416), .B(n34417), .Z(n27052) );
  AND U36265 ( .A(\modmult_1/xin[1023] ), .B(n34418), .Z(n34417) );
  IV U36266 ( .A(n34416), .Z(n34418) );
  XOR U36267 ( .A(n34419), .B(mreg[615]), .Z(n34416) );
  NAND U36268 ( .A(n34420), .B(mul_pow), .Z(n34419) );
  XOR U36269 ( .A(mreg[615]), .B(creg[615]), .Z(n34420) );
  XOR U36270 ( .A(n34421), .B(n34422), .Z(n34412) );
  ANDN U36271 ( .A(n34423), .B(n27059), .Z(n34422) );
  XOR U36272 ( .A(n34424), .B(\modmult_1/zin[0][613] ), .Z(n27059) );
  IV U36273 ( .A(n34421), .Z(n34424) );
  XNOR U36274 ( .A(n34421), .B(n27058), .Z(n34423) );
  XOR U36275 ( .A(n34425), .B(n34426), .Z(n27058) );
  AND U36276 ( .A(\modmult_1/xin[1023] ), .B(n34427), .Z(n34426) );
  IV U36277 ( .A(n34425), .Z(n34427) );
  XOR U36278 ( .A(n34428), .B(mreg[614]), .Z(n34425) );
  NAND U36279 ( .A(n34429), .B(mul_pow), .Z(n34428) );
  XOR U36280 ( .A(mreg[614]), .B(creg[614]), .Z(n34429) );
  XOR U36281 ( .A(n34430), .B(n34431), .Z(n34421) );
  ANDN U36282 ( .A(n34432), .B(n27065), .Z(n34431) );
  XOR U36283 ( .A(n34433), .B(\modmult_1/zin[0][612] ), .Z(n27065) );
  IV U36284 ( .A(n34430), .Z(n34433) );
  XNOR U36285 ( .A(n34430), .B(n27064), .Z(n34432) );
  XOR U36286 ( .A(n34434), .B(n34435), .Z(n27064) );
  AND U36287 ( .A(\modmult_1/xin[1023] ), .B(n34436), .Z(n34435) );
  IV U36288 ( .A(n34434), .Z(n34436) );
  XOR U36289 ( .A(n34437), .B(mreg[613]), .Z(n34434) );
  NAND U36290 ( .A(n34438), .B(mul_pow), .Z(n34437) );
  XOR U36291 ( .A(mreg[613]), .B(creg[613]), .Z(n34438) );
  XOR U36292 ( .A(n34439), .B(n34440), .Z(n34430) );
  ANDN U36293 ( .A(n34441), .B(n27071), .Z(n34440) );
  XOR U36294 ( .A(n34442), .B(\modmult_1/zin[0][611] ), .Z(n27071) );
  IV U36295 ( .A(n34439), .Z(n34442) );
  XNOR U36296 ( .A(n34439), .B(n27070), .Z(n34441) );
  XOR U36297 ( .A(n34443), .B(n34444), .Z(n27070) );
  AND U36298 ( .A(\modmult_1/xin[1023] ), .B(n34445), .Z(n34444) );
  IV U36299 ( .A(n34443), .Z(n34445) );
  XOR U36300 ( .A(n34446), .B(mreg[612]), .Z(n34443) );
  NAND U36301 ( .A(n34447), .B(mul_pow), .Z(n34446) );
  XOR U36302 ( .A(mreg[612]), .B(creg[612]), .Z(n34447) );
  XOR U36303 ( .A(n34448), .B(n34449), .Z(n34439) );
  ANDN U36304 ( .A(n34450), .B(n27077), .Z(n34449) );
  XOR U36305 ( .A(n34451), .B(\modmult_1/zin[0][610] ), .Z(n27077) );
  IV U36306 ( .A(n34448), .Z(n34451) );
  XNOR U36307 ( .A(n34448), .B(n27076), .Z(n34450) );
  XOR U36308 ( .A(n34452), .B(n34453), .Z(n27076) );
  AND U36309 ( .A(\modmult_1/xin[1023] ), .B(n34454), .Z(n34453) );
  IV U36310 ( .A(n34452), .Z(n34454) );
  XOR U36311 ( .A(n34455), .B(mreg[611]), .Z(n34452) );
  NAND U36312 ( .A(n34456), .B(mul_pow), .Z(n34455) );
  XOR U36313 ( .A(mreg[611]), .B(creg[611]), .Z(n34456) );
  XOR U36314 ( .A(n34457), .B(n34458), .Z(n34448) );
  ANDN U36315 ( .A(n34459), .B(n27083), .Z(n34458) );
  XOR U36316 ( .A(n34460), .B(\modmult_1/zin[0][609] ), .Z(n27083) );
  IV U36317 ( .A(n34457), .Z(n34460) );
  XNOR U36318 ( .A(n34457), .B(n27082), .Z(n34459) );
  XOR U36319 ( .A(n34461), .B(n34462), .Z(n27082) );
  AND U36320 ( .A(\modmult_1/xin[1023] ), .B(n34463), .Z(n34462) );
  IV U36321 ( .A(n34461), .Z(n34463) );
  XOR U36322 ( .A(n34464), .B(mreg[610]), .Z(n34461) );
  NAND U36323 ( .A(n34465), .B(mul_pow), .Z(n34464) );
  XOR U36324 ( .A(mreg[610]), .B(creg[610]), .Z(n34465) );
  XOR U36325 ( .A(n34466), .B(n34467), .Z(n34457) );
  ANDN U36326 ( .A(n34468), .B(n27089), .Z(n34467) );
  XOR U36327 ( .A(n34469), .B(\modmult_1/zin[0][608] ), .Z(n27089) );
  IV U36328 ( .A(n34466), .Z(n34469) );
  XNOR U36329 ( .A(n34466), .B(n27088), .Z(n34468) );
  XOR U36330 ( .A(n34470), .B(n34471), .Z(n27088) );
  AND U36331 ( .A(\modmult_1/xin[1023] ), .B(n34472), .Z(n34471) );
  IV U36332 ( .A(n34470), .Z(n34472) );
  XOR U36333 ( .A(n34473), .B(mreg[609]), .Z(n34470) );
  NAND U36334 ( .A(n34474), .B(mul_pow), .Z(n34473) );
  XOR U36335 ( .A(mreg[609]), .B(creg[609]), .Z(n34474) );
  XOR U36336 ( .A(n34475), .B(n34476), .Z(n34466) );
  ANDN U36337 ( .A(n34477), .B(n27095), .Z(n34476) );
  XOR U36338 ( .A(n34478), .B(\modmult_1/zin[0][607] ), .Z(n27095) );
  IV U36339 ( .A(n34475), .Z(n34478) );
  XNOR U36340 ( .A(n34475), .B(n27094), .Z(n34477) );
  XOR U36341 ( .A(n34479), .B(n34480), .Z(n27094) );
  AND U36342 ( .A(\modmult_1/xin[1023] ), .B(n34481), .Z(n34480) );
  IV U36343 ( .A(n34479), .Z(n34481) );
  XOR U36344 ( .A(n34482), .B(mreg[608]), .Z(n34479) );
  NAND U36345 ( .A(n34483), .B(mul_pow), .Z(n34482) );
  XOR U36346 ( .A(mreg[608]), .B(creg[608]), .Z(n34483) );
  XOR U36347 ( .A(n34484), .B(n34485), .Z(n34475) );
  ANDN U36348 ( .A(n34486), .B(n27101), .Z(n34485) );
  XOR U36349 ( .A(n34487), .B(\modmult_1/zin[0][606] ), .Z(n27101) );
  IV U36350 ( .A(n34484), .Z(n34487) );
  XNOR U36351 ( .A(n34484), .B(n27100), .Z(n34486) );
  XOR U36352 ( .A(n34488), .B(n34489), .Z(n27100) );
  AND U36353 ( .A(\modmult_1/xin[1023] ), .B(n34490), .Z(n34489) );
  IV U36354 ( .A(n34488), .Z(n34490) );
  XOR U36355 ( .A(n34491), .B(mreg[607]), .Z(n34488) );
  NAND U36356 ( .A(n34492), .B(mul_pow), .Z(n34491) );
  XOR U36357 ( .A(mreg[607]), .B(creg[607]), .Z(n34492) );
  XOR U36358 ( .A(n34493), .B(n34494), .Z(n34484) );
  ANDN U36359 ( .A(n34495), .B(n27107), .Z(n34494) );
  XOR U36360 ( .A(n34496), .B(\modmult_1/zin[0][605] ), .Z(n27107) );
  IV U36361 ( .A(n34493), .Z(n34496) );
  XNOR U36362 ( .A(n34493), .B(n27106), .Z(n34495) );
  XOR U36363 ( .A(n34497), .B(n34498), .Z(n27106) );
  AND U36364 ( .A(\modmult_1/xin[1023] ), .B(n34499), .Z(n34498) );
  IV U36365 ( .A(n34497), .Z(n34499) );
  XOR U36366 ( .A(n34500), .B(mreg[606]), .Z(n34497) );
  NAND U36367 ( .A(n34501), .B(mul_pow), .Z(n34500) );
  XOR U36368 ( .A(mreg[606]), .B(creg[606]), .Z(n34501) );
  XOR U36369 ( .A(n34502), .B(n34503), .Z(n34493) );
  ANDN U36370 ( .A(n34504), .B(n27113), .Z(n34503) );
  XOR U36371 ( .A(n34505), .B(\modmult_1/zin[0][604] ), .Z(n27113) );
  IV U36372 ( .A(n34502), .Z(n34505) );
  XNOR U36373 ( .A(n34502), .B(n27112), .Z(n34504) );
  XOR U36374 ( .A(n34506), .B(n34507), .Z(n27112) );
  AND U36375 ( .A(\modmult_1/xin[1023] ), .B(n34508), .Z(n34507) );
  IV U36376 ( .A(n34506), .Z(n34508) );
  XOR U36377 ( .A(n34509), .B(mreg[605]), .Z(n34506) );
  NAND U36378 ( .A(n34510), .B(mul_pow), .Z(n34509) );
  XOR U36379 ( .A(mreg[605]), .B(creg[605]), .Z(n34510) );
  XOR U36380 ( .A(n34511), .B(n34512), .Z(n34502) );
  ANDN U36381 ( .A(n34513), .B(n27119), .Z(n34512) );
  XOR U36382 ( .A(n34514), .B(\modmult_1/zin[0][603] ), .Z(n27119) );
  IV U36383 ( .A(n34511), .Z(n34514) );
  XNOR U36384 ( .A(n34511), .B(n27118), .Z(n34513) );
  XOR U36385 ( .A(n34515), .B(n34516), .Z(n27118) );
  AND U36386 ( .A(\modmult_1/xin[1023] ), .B(n34517), .Z(n34516) );
  IV U36387 ( .A(n34515), .Z(n34517) );
  XOR U36388 ( .A(n34518), .B(mreg[604]), .Z(n34515) );
  NAND U36389 ( .A(n34519), .B(mul_pow), .Z(n34518) );
  XOR U36390 ( .A(mreg[604]), .B(creg[604]), .Z(n34519) );
  XOR U36391 ( .A(n34520), .B(n34521), .Z(n34511) );
  ANDN U36392 ( .A(n34522), .B(n27125), .Z(n34521) );
  XOR U36393 ( .A(n34523), .B(\modmult_1/zin[0][602] ), .Z(n27125) );
  IV U36394 ( .A(n34520), .Z(n34523) );
  XNOR U36395 ( .A(n34520), .B(n27124), .Z(n34522) );
  XOR U36396 ( .A(n34524), .B(n34525), .Z(n27124) );
  AND U36397 ( .A(\modmult_1/xin[1023] ), .B(n34526), .Z(n34525) );
  IV U36398 ( .A(n34524), .Z(n34526) );
  XOR U36399 ( .A(n34527), .B(mreg[603]), .Z(n34524) );
  NAND U36400 ( .A(n34528), .B(mul_pow), .Z(n34527) );
  XOR U36401 ( .A(mreg[603]), .B(creg[603]), .Z(n34528) );
  XOR U36402 ( .A(n34529), .B(n34530), .Z(n34520) );
  ANDN U36403 ( .A(n34531), .B(n27131), .Z(n34530) );
  XOR U36404 ( .A(n34532), .B(\modmult_1/zin[0][601] ), .Z(n27131) );
  IV U36405 ( .A(n34529), .Z(n34532) );
  XNOR U36406 ( .A(n34529), .B(n27130), .Z(n34531) );
  XOR U36407 ( .A(n34533), .B(n34534), .Z(n27130) );
  AND U36408 ( .A(\modmult_1/xin[1023] ), .B(n34535), .Z(n34534) );
  IV U36409 ( .A(n34533), .Z(n34535) );
  XOR U36410 ( .A(n34536), .B(mreg[602]), .Z(n34533) );
  NAND U36411 ( .A(n34537), .B(mul_pow), .Z(n34536) );
  XOR U36412 ( .A(mreg[602]), .B(creg[602]), .Z(n34537) );
  XOR U36413 ( .A(n34538), .B(n34539), .Z(n34529) );
  ANDN U36414 ( .A(n34540), .B(n27137), .Z(n34539) );
  XOR U36415 ( .A(n34541), .B(\modmult_1/zin[0][600] ), .Z(n27137) );
  IV U36416 ( .A(n34538), .Z(n34541) );
  XNOR U36417 ( .A(n34538), .B(n27136), .Z(n34540) );
  XOR U36418 ( .A(n34542), .B(n34543), .Z(n27136) );
  AND U36419 ( .A(\modmult_1/xin[1023] ), .B(n34544), .Z(n34543) );
  IV U36420 ( .A(n34542), .Z(n34544) );
  XOR U36421 ( .A(n34545), .B(mreg[601]), .Z(n34542) );
  NAND U36422 ( .A(n34546), .B(mul_pow), .Z(n34545) );
  XOR U36423 ( .A(mreg[601]), .B(creg[601]), .Z(n34546) );
  XOR U36424 ( .A(n34547), .B(n34548), .Z(n34538) );
  ANDN U36425 ( .A(n34549), .B(n27143), .Z(n34548) );
  XOR U36426 ( .A(n34550), .B(\modmult_1/zin[0][599] ), .Z(n27143) );
  IV U36427 ( .A(n34547), .Z(n34550) );
  XNOR U36428 ( .A(n34547), .B(n27142), .Z(n34549) );
  XOR U36429 ( .A(n34551), .B(n34552), .Z(n27142) );
  AND U36430 ( .A(\modmult_1/xin[1023] ), .B(n34553), .Z(n34552) );
  IV U36431 ( .A(n34551), .Z(n34553) );
  XOR U36432 ( .A(n34554), .B(mreg[600]), .Z(n34551) );
  NAND U36433 ( .A(n34555), .B(mul_pow), .Z(n34554) );
  XOR U36434 ( .A(mreg[600]), .B(creg[600]), .Z(n34555) );
  XOR U36435 ( .A(n34556), .B(n34557), .Z(n34547) );
  ANDN U36436 ( .A(n34558), .B(n27149), .Z(n34557) );
  XOR U36437 ( .A(n34559), .B(\modmult_1/zin[0][598] ), .Z(n27149) );
  IV U36438 ( .A(n34556), .Z(n34559) );
  XNOR U36439 ( .A(n34556), .B(n27148), .Z(n34558) );
  XOR U36440 ( .A(n34560), .B(n34561), .Z(n27148) );
  AND U36441 ( .A(\modmult_1/xin[1023] ), .B(n34562), .Z(n34561) );
  IV U36442 ( .A(n34560), .Z(n34562) );
  XOR U36443 ( .A(n34563), .B(mreg[599]), .Z(n34560) );
  NAND U36444 ( .A(n34564), .B(mul_pow), .Z(n34563) );
  XOR U36445 ( .A(mreg[599]), .B(creg[599]), .Z(n34564) );
  XOR U36446 ( .A(n34565), .B(n34566), .Z(n34556) );
  ANDN U36447 ( .A(n34567), .B(n27155), .Z(n34566) );
  XOR U36448 ( .A(n34568), .B(\modmult_1/zin[0][597] ), .Z(n27155) );
  IV U36449 ( .A(n34565), .Z(n34568) );
  XNOR U36450 ( .A(n34565), .B(n27154), .Z(n34567) );
  XOR U36451 ( .A(n34569), .B(n34570), .Z(n27154) );
  AND U36452 ( .A(\modmult_1/xin[1023] ), .B(n34571), .Z(n34570) );
  IV U36453 ( .A(n34569), .Z(n34571) );
  XOR U36454 ( .A(n34572), .B(mreg[598]), .Z(n34569) );
  NAND U36455 ( .A(n34573), .B(mul_pow), .Z(n34572) );
  XOR U36456 ( .A(mreg[598]), .B(creg[598]), .Z(n34573) );
  XOR U36457 ( .A(n34574), .B(n34575), .Z(n34565) );
  ANDN U36458 ( .A(n34576), .B(n27161), .Z(n34575) );
  XOR U36459 ( .A(n34577), .B(\modmult_1/zin[0][596] ), .Z(n27161) );
  IV U36460 ( .A(n34574), .Z(n34577) );
  XNOR U36461 ( .A(n34574), .B(n27160), .Z(n34576) );
  XOR U36462 ( .A(n34578), .B(n34579), .Z(n27160) );
  AND U36463 ( .A(\modmult_1/xin[1023] ), .B(n34580), .Z(n34579) );
  IV U36464 ( .A(n34578), .Z(n34580) );
  XOR U36465 ( .A(n34581), .B(mreg[597]), .Z(n34578) );
  NAND U36466 ( .A(n34582), .B(mul_pow), .Z(n34581) );
  XOR U36467 ( .A(mreg[597]), .B(creg[597]), .Z(n34582) );
  XOR U36468 ( .A(n34583), .B(n34584), .Z(n34574) );
  ANDN U36469 ( .A(n34585), .B(n27167), .Z(n34584) );
  XOR U36470 ( .A(n34586), .B(\modmult_1/zin[0][595] ), .Z(n27167) );
  IV U36471 ( .A(n34583), .Z(n34586) );
  XNOR U36472 ( .A(n34583), .B(n27166), .Z(n34585) );
  XOR U36473 ( .A(n34587), .B(n34588), .Z(n27166) );
  AND U36474 ( .A(\modmult_1/xin[1023] ), .B(n34589), .Z(n34588) );
  IV U36475 ( .A(n34587), .Z(n34589) );
  XOR U36476 ( .A(n34590), .B(mreg[596]), .Z(n34587) );
  NAND U36477 ( .A(n34591), .B(mul_pow), .Z(n34590) );
  XOR U36478 ( .A(mreg[596]), .B(creg[596]), .Z(n34591) );
  XOR U36479 ( .A(n34592), .B(n34593), .Z(n34583) );
  ANDN U36480 ( .A(n34594), .B(n27173), .Z(n34593) );
  XOR U36481 ( .A(n34595), .B(\modmult_1/zin[0][594] ), .Z(n27173) );
  IV U36482 ( .A(n34592), .Z(n34595) );
  XNOR U36483 ( .A(n34592), .B(n27172), .Z(n34594) );
  XOR U36484 ( .A(n34596), .B(n34597), .Z(n27172) );
  AND U36485 ( .A(\modmult_1/xin[1023] ), .B(n34598), .Z(n34597) );
  IV U36486 ( .A(n34596), .Z(n34598) );
  XOR U36487 ( .A(n34599), .B(mreg[595]), .Z(n34596) );
  NAND U36488 ( .A(n34600), .B(mul_pow), .Z(n34599) );
  XOR U36489 ( .A(mreg[595]), .B(creg[595]), .Z(n34600) );
  XOR U36490 ( .A(n34601), .B(n34602), .Z(n34592) );
  ANDN U36491 ( .A(n34603), .B(n27179), .Z(n34602) );
  XOR U36492 ( .A(n34604), .B(\modmult_1/zin[0][593] ), .Z(n27179) );
  IV U36493 ( .A(n34601), .Z(n34604) );
  XNOR U36494 ( .A(n34601), .B(n27178), .Z(n34603) );
  XOR U36495 ( .A(n34605), .B(n34606), .Z(n27178) );
  AND U36496 ( .A(\modmult_1/xin[1023] ), .B(n34607), .Z(n34606) );
  IV U36497 ( .A(n34605), .Z(n34607) );
  XOR U36498 ( .A(n34608), .B(mreg[594]), .Z(n34605) );
  NAND U36499 ( .A(n34609), .B(mul_pow), .Z(n34608) );
  XOR U36500 ( .A(mreg[594]), .B(creg[594]), .Z(n34609) );
  XOR U36501 ( .A(n34610), .B(n34611), .Z(n34601) );
  ANDN U36502 ( .A(n34612), .B(n27185), .Z(n34611) );
  XOR U36503 ( .A(n34613), .B(\modmult_1/zin[0][592] ), .Z(n27185) );
  IV U36504 ( .A(n34610), .Z(n34613) );
  XNOR U36505 ( .A(n34610), .B(n27184), .Z(n34612) );
  XOR U36506 ( .A(n34614), .B(n34615), .Z(n27184) );
  AND U36507 ( .A(\modmult_1/xin[1023] ), .B(n34616), .Z(n34615) );
  IV U36508 ( .A(n34614), .Z(n34616) );
  XOR U36509 ( .A(n34617), .B(mreg[593]), .Z(n34614) );
  NAND U36510 ( .A(n34618), .B(mul_pow), .Z(n34617) );
  XOR U36511 ( .A(mreg[593]), .B(creg[593]), .Z(n34618) );
  XOR U36512 ( .A(n34619), .B(n34620), .Z(n34610) );
  ANDN U36513 ( .A(n34621), .B(n27191), .Z(n34620) );
  XOR U36514 ( .A(n34622), .B(\modmult_1/zin[0][591] ), .Z(n27191) );
  IV U36515 ( .A(n34619), .Z(n34622) );
  XNOR U36516 ( .A(n34619), .B(n27190), .Z(n34621) );
  XOR U36517 ( .A(n34623), .B(n34624), .Z(n27190) );
  AND U36518 ( .A(\modmult_1/xin[1023] ), .B(n34625), .Z(n34624) );
  IV U36519 ( .A(n34623), .Z(n34625) );
  XOR U36520 ( .A(n34626), .B(mreg[592]), .Z(n34623) );
  NAND U36521 ( .A(n34627), .B(mul_pow), .Z(n34626) );
  XOR U36522 ( .A(mreg[592]), .B(creg[592]), .Z(n34627) );
  XOR U36523 ( .A(n34628), .B(n34629), .Z(n34619) );
  ANDN U36524 ( .A(n34630), .B(n27197), .Z(n34629) );
  XOR U36525 ( .A(n34631), .B(\modmult_1/zin[0][590] ), .Z(n27197) );
  IV U36526 ( .A(n34628), .Z(n34631) );
  XNOR U36527 ( .A(n34628), .B(n27196), .Z(n34630) );
  XOR U36528 ( .A(n34632), .B(n34633), .Z(n27196) );
  AND U36529 ( .A(\modmult_1/xin[1023] ), .B(n34634), .Z(n34633) );
  IV U36530 ( .A(n34632), .Z(n34634) );
  XOR U36531 ( .A(n34635), .B(mreg[591]), .Z(n34632) );
  NAND U36532 ( .A(n34636), .B(mul_pow), .Z(n34635) );
  XOR U36533 ( .A(mreg[591]), .B(creg[591]), .Z(n34636) );
  XOR U36534 ( .A(n34637), .B(n34638), .Z(n34628) );
  ANDN U36535 ( .A(n34639), .B(n27203), .Z(n34638) );
  XOR U36536 ( .A(n34640), .B(\modmult_1/zin[0][589] ), .Z(n27203) );
  IV U36537 ( .A(n34637), .Z(n34640) );
  XNOR U36538 ( .A(n34637), .B(n27202), .Z(n34639) );
  XOR U36539 ( .A(n34641), .B(n34642), .Z(n27202) );
  AND U36540 ( .A(\modmult_1/xin[1023] ), .B(n34643), .Z(n34642) );
  IV U36541 ( .A(n34641), .Z(n34643) );
  XOR U36542 ( .A(n34644), .B(mreg[590]), .Z(n34641) );
  NAND U36543 ( .A(n34645), .B(mul_pow), .Z(n34644) );
  XOR U36544 ( .A(mreg[590]), .B(creg[590]), .Z(n34645) );
  XOR U36545 ( .A(n34646), .B(n34647), .Z(n34637) );
  ANDN U36546 ( .A(n34648), .B(n27209), .Z(n34647) );
  XOR U36547 ( .A(n34649), .B(\modmult_1/zin[0][588] ), .Z(n27209) );
  IV U36548 ( .A(n34646), .Z(n34649) );
  XNOR U36549 ( .A(n34646), .B(n27208), .Z(n34648) );
  XOR U36550 ( .A(n34650), .B(n34651), .Z(n27208) );
  AND U36551 ( .A(\modmult_1/xin[1023] ), .B(n34652), .Z(n34651) );
  IV U36552 ( .A(n34650), .Z(n34652) );
  XOR U36553 ( .A(n34653), .B(mreg[589]), .Z(n34650) );
  NAND U36554 ( .A(n34654), .B(mul_pow), .Z(n34653) );
  XOR U36555 ( .A(mreg[589]), .B(creg[589]), .Z(n34654) );
  XOR U36556 ( .A(n34655), .B(n34656), .Z(n34646) );
  ANDN U36557 ( .A(n34657), .B(n27215), .Z(n34656) );
  XOR U36558 ( .A(n34658), .B(\modmult_1/zin[0][587] ), .Z(n27215) );
  IV U36559 ( .A(n34655), .Z(n34658) );
  XNOR U36560 ( .A(n34655), .B(n27214), .Z(n34657) );
  XOR U36561 ( .A(n34659), .B(n34660), .Z(n27214) );
  AND U36562 ( .A(\modmult_1/xin[1023] ), .B(n34661), .Z(n34660) );
  IV U36563 ( .A(n34659), .Z(n34661) );
  XOR U36564 ( .A(n34662), .B(mreg[588]), .Z(n34659) );
  NAND U36565 ( .A(n34663), .B(mul_pow), .Z(n34662) );
  XOR U36566 ( .A(mreg[588]), .B(creg[588]), .Z(n34663) );
  XOR U36567 ( .A(n34664), .B(n34665), .Z(n34655) );
  ANDN U36568 ( .A(n34666), .B(n27221), .Z(n34665) );
  XOR U36569 ( .A(n34667), .B(\modmult_1/zin[0][586] ), .Z(n27221) );
  IV U36570 ( .A(n34664), .Z(n34667) );
  XNOR U36571 ( .A(n34664), .B(n27220), .Z(n34666) );
  XOR U36572 ( .A(n34668), .B(n34669), .Z(n27220) );
  AND U36573 ( .A(\modmult_1/xin[1023] ), .B(n34670), .Z(n34669) );
  IV U36574 ( .A(n34668), .Z(n34670) );
  XOR U36575 ( .A(n34671), .B(mreg[587]), .Z(n34668) );
  NAND U36576 ( .A(n34672), .B(mul_pow), .Z(n34671) );
  XOR U36577 ( .A(mreg[587]), .B(creg[587]), .Z(n34672) );
  XOR U36578 ( .A(n34673), .B(n34674), .Z(n34664) );
  ANDN U36579 ( .A(n34675), .B(n27227), .Z(n34674) );
  XOR U36580 ( .A(n34676), .B(\modmult_1/zin[0][585] ), .Z(n27227) );
  IV U36581 ( .A(n34673), .Z(n34676) );
  XNOR U36582 ( .A(n34673), .B(n27226), .Z(n34675) );
  XOR U36583 ( .A(n34677), .B(n34678), .Z(n27226) );
  AND U36584 ( .A(\modmult_1/xin[1023] ), .B(n34679), .Z(n34678) );
  IV U36585 ( .A(n34677), .Z(n34679) );
  XOR U36586 ( .A(n34680), .B(mreg[586]), .Z(n34677) );
  NAND U36587 ( .A(n34681), .B(mul_pow), .Z(n34680) );
  XOR U36588 ( .A(mreg[586]), .B(creg[586]), .Z(n34681) );
  XOR U36589 ( .A(n34682), .B(n34683), .Z(n34673) );
  ANDN U36590 ( .A(n34684), .B(n27233), .Z(n34683) );
  XOR U36591 ( .A(n34685), .B(\modmult_1/zin[0][584] ), .Z(n27233) );
  IV U36592 ( .A(n34682), .Z(n34685) );
  XNOR U36593 ( .A(n34682), .B(n27232), .Z(n34684) );
  XOR U36594 ( .A(n34686), .B(n34687), .Z(n27232) );
  AND U36595 ( .A(\modmult_1/xin[1023] ), .B(n34688), .Z(n34687) );
  IV U36596 ( .A(n34686), .Z(n34688) );
  XOR U36597 ( .A(n34689), .B(mreg[585]), .Z(n34686) );
  NAND U36598 ( .A(n34690), .B(mul_pow), .Z(n34689) );
  XOR U36599 ( .A(mreg[585]), .B(creg[585]), .Z(n34690) );
  XOR U36600 ( .A(n34691), .B(n34692), .Z(n34682) );
  ANDN U36601 ( .A(n34693), .B(n27239), .Z(n34692) );
  XOR U36602 ( .A(n34694), .B(\modmult_1/zin[0][583] ), .Z(n27239) );
  IV U36603 ( .A(n34691), .Z(n34694) );
  XNOR U36604 ( .A(n34691), .B(n27238), .Z(n34693) );
  XOR U36605 ( .A(n34695), .B(n34696), .Z(n27238) );
  AND U36606 ( .A(\modmult_1/xin[1023] ), .B(n34697), .Z(n34696) );
  IV U36607 ( .A(n34695), .Z(n34697) );
  XOR U36608 ( .A(n34698), .B(mreg[584]), .Z(n34695) );
  NAND U36609 ( .A(n34699), .B(mul_pow), .Z(n34698) );
  XOR U36610 ( .A(mreg[584]), .B(creg[584]), .Z(n34699) );
  XOR U36611 ( .A(n34700), .B(n34701), .Z(n34691) );
  ANDN U36612 ( .A(n34702), .B(n27245), .Z(n34701) );
  XOR U36613 ( .A(n34703), .B(\modmult_1/zin[0][582] ), .Z(n27245) );
  IV U36614 ( .A(n34700), .Z(n34703) );
  XNOR U36615 ( .A(n34700), .B(n27244), .Z(n34702) );
  XOR U36616 ( .A(n34704), .B(n34705), .Z(n27244) );
  AND U36617 ( .A(\modmult_1/xin[1023] ), .B(n34706), .Z(n34705) );
  IV U36618 ( .A(n34704), .Z(n34706) );
  XOR U36619 ( .A(n34707), .B(mreg[583]), .Z(n34704) );
  NAND U36620 ( .A(n34708), .B(mul_pow), .Z(n34707) );
  XOR U36621 ( .A(mreg[583]), .B(creg[583]), .Z(n34708) );
  XOR U36622 ( .A(n34709), .B(n34710), .Z(n34700) );
  ANDN U36623 ( .A(n34711), .B(n27251), .Z(n34710) );
  XOR U36624 ( .A(n34712), .B(\modmult_1/zin[0][581] ), .Z(n27251) );
  IV U36625 ( .A(n34709), .Z(n34712) );
  XNOR U36626 ( .A(n34709), .B(n27250), .Z(n34711) );
  XOR U36627 ( .A(n34713), .B(n34714), .Z(n27250) );
  AND U36628 ( .A(\modmult_1/xin[1023] ), .B(n34715), .Z(n34714) );
  IV U36629 ( .A(n34713), .Z(n34715) );
  XOR U36630 ( .A(n34716), .B(mreg[582]), .Z(n34713) );
  NAND U36631 ( .A(n34717), .B(mul_pow), .Z(n34716) );
  XOR U36632 ( .A(mreg[582]), .B(creg[582]), .Z(n34717) );
  XOR U36633 ( .A(n34718), .B(n34719), .Z(n34709) );
  ANDN U36634 ( .A(n34720), .B(n27257), .Z(n34719) );
  XOR U36635 ( .A(n34721), .B(\modmult_1/zin[0][580] ), .Z(n27257) );
  IV U36636 ( .A(n34718), .Z(n34721) );
  XNOR U36637 ( .A(n34718), .B(n27256), .Z(n34720) );
  XOR U36638 ( .A(n34722), .B(n34723), .Z(n27256) );
  AND U36639 ( .A(\modmult_1/xin[1023] ), .B(n34724), .Z(n34723) );
  IV U36640 ( .A(n34722), .Z(n34724) );
  XOR U36641 ( .A(n34725), .B(mreg[581]), .Z(n34722) );
  NAND U36642 ( .A(n34726), .B(mul_pow), .Z(n34725) );
  XOR U36643 ( .A(mreg[581]), .B(creg[581]), .Z(n34726) );
  XOR U36644 ( .A(n34727), .B(n34728), .Z(n34718) );
  ANDN U36645 ( .A(n34729), .B(n27263), .Z(n34728) );
  XOR U36646 ( .A(n34730), .B(\modmult_1/zin[0][579] ), .Z(n27263) );
  IV U36647 ( .A(n34727), .Z(n34730) );
  XNOR U36648 ( .A(n34727), .B(n27262), .Z(n34729) );
  XOR U36649 ( .A(n34731), .B(n34732), .Z(n27262) );
  AND U36650 ( .A(\modmult_1/xin[1023] ), .B(n34733), .Z(n34732) );
  IV U36651 ( .A(n34731), .Z(n34733) );
  XOR U36652 ( .A(n34734), .B(mreg[580]), .Z(n34731) );
  NAND U36653 ( .A(n34735), .B(mul_pow), .Z(n34734) );
  XOR U36654 ( .A(mreg[580]), .B(creg[580]), .Z(n34735) );
  XOR U36655 ( .A(n34736), .B(n34737), .Z(n34727) );
  ANDN U36656 ( .A(n34738), .B(n27269), .Z(n34737) );
  XOR U36657 ( .A(n34739), .B(\modmult_1/zin[0][578] ), .Z(n27269) );
  IV U36658 ( .A(n34736), .Z(n34739) );
  XNOR U36659 ( .A(n34736), .B(n27268), .Z(n34738) );
  XOR U36660 ( .A(n34740), .B(n34741), .Z(n27268) );
  AND U36661 ( .A(\modmult_1/xin[1023] ), .B(n34742), .Z(n34741) );
  IV U36662 ( .A(n34740), .Z(n34742) );
  XOR U36663 ( .A(n34743), .B(mreg[579]), .Z(n34740) );
  NAND U36664 ( .A(n34744), .B(mul_pow), .Z(n34743) );
  XOR U36665 ( .A(mreg[579]), .B(creg[579]), .Z(n34744) );
  XOR U36666 ( .A(n34745), .B(n34746), .Z(n34736) );
  ANDN U36667 ( .A(n34747), .B(n27275), .Z(n34746) );
  XOR U36668 ( .A(n34748), .B(\modmult_1/zin[0][577] ), .Z(n27275) );
  IV U36669 ( .A(n34745), .Z(n34748) );
  XNOR U36670 ( .A(n34745), .B(n27274), .Z(n34747) );
  XOR U36671 ( .A(n34749), .B(n34750), .Z(n27274) );
  AND U36672 ( .A(\modmult_1/xin[1023] ), .B(n34751), .Z(n34750) );
  IV U36673 ( .A(n34749), .Z(n34751) );
  XOR U36674 ( .A(n34752), .B(mreg[578]), .Z(n34749) );
  NAND U36675 ( .A(n34753), .B(mul_pow), .Z(n34752) );
  XOR U36676 ( .A(mreg[578]), .B(creg[578]), .Z(n34753) );
  XOR U36677 ( .A(n34754), .B(n34755), .Z(n34745) );
  ANDN U36678 ( .A(n34756), .B(n27281), .Z(n34755) );
  XOR U36679 ( .A(n34757), .B(\modmult_1/zin[0][576] ), .Z(n27281) );
  IV U36680 ( .A(n34754), .Z(n34757) );
  XNOR U36681 ( .A(n34754), .B(n27280), .Z(n34756) );
  XOR U36682 ( .A(n34758), .B(n34759), .Z(n27280) );
  AND U36683 ( .A(\modmult_1/xin[1023] ), .B(n34760), .Z(n34759) );
  IV U36684 ( .A(n34758), .Z(n34760) );
  XOR U36685 ( .A(n34761), .B(mreg[577]), .Z(n34758) );
  NAND U36686 ( .A(n34762), .B(mul_pow), .Z(n34761) );
  XOR U36687 ( .A(mreg[577]), .B(creg[577]), .Z(n34762) );
  XOR U36688 ( .A(n34763), .B(n34764), .Z(n34754) );
  ANDN U36689 ( .A(n34765), .B(n27287), .Z(n34764) );
  XOR U36690 ( .A(n34766), .B(\modmult_1/zin[0][575] ), .Z(n27287) );
  IV U36691 ( .A(n34763), .Z(n34766) );
  XNOR U36692 ( .A(n34763), .B(n27286), .Z(n34765) );
  XOR U36693 ( .A(n34767), .B(n34768), .Z(n27286) );
  AND U36694 ( .A(\modmult_1/xin[1023] ), .B(n34769), .Z(n34768) );
  IV U36695 ( .A(n34767), .Z(n34769) );
  XOR U36696 ( .A(n34770), .B(mreg[576]), .Z(n34767) );
  NAND U36697 ( .A(n34771), .B(mul_pow), .Z(n34770) );
  XOR U36698 ( .A(mreg[576]), .B(creg[576]), .Z(n34771) );
  XOR U36699 ( .A(n34772), .B(n34773), .Z(n34763) );
  ANDN U36700 ( .A(n34774), .B(n27293), .Z(n34773) );
  XOR U36701 ( .A(n34775), .B(\modmult_1/zin[0][574] ), .Z(n27293) );
  IV U36702 ( .A(n34772), .Z(n34775) );
  XNOR U36703 ( .A(n34772), .B(n27292), .Z(n34774) );
  XOR U36704 ( .A(n34776), .B(n34777), .Z(n27292) );
  AND U36705 ( .A(\modmult_1/xin[1023] ), .B(n34778), .Z(n34777) );
  IV U36706 ( .A(n34776), .Z(n34778) );
  XOR U36707 ( .A(n34779), .B(mreg[575]), .Z(n34776) );
  NAND U36708 ( .A(n34780), .B(mul_pow), .Z(n34779) );
  XOR U36709 ( .A(mreg[575]), .B(creg[575]), .Z(n34780) );
  XOR U36710 ( .A(n34781), .B(n34782), .Z(n34772) );
  ANDN U36711 ( .A(n34783), .B(n27299), .Z(n34782) );
  XOR U36712 ( .A(n34784), .B(\modmult_1/zin[0][573] ), .Z(n27299) );
  IV U36713 ( .A(n34781), .Z(n34784) );
  XNOR U36714 ( .A(n34781), .B(n27298), .Z(n34783) );
  XOR U36715 ( .A(n34785), .B(n34786), .Z(n27298) );
  AND U36716 ( .A(\modmult_1/xin[1023] ), .B(n34787), .Z(n34786) );
  IV U36717 ( .A(n34785), .Z(n34787) );
  XOR U36718 ( .A(n34788), .B(mreg[574]), .Z(n34785) );
  NAND U36719 ( .A(n34789), .B(mul_pow), .Z(n34788) );
  XOR U36720 ( .A(mreg[574]), .B(creg[574]), .Z(n34789) );
  XOR U36721 ( .A(n34790), .B(n34791), .Z(n34781) );
  ANDN U36722 ( .A(n34792), .B(n27305), .Z(n34791) );
  XOR U36723 ( .A(n34793), .B(\modmult_1/zin[0][572] ), .Z(n27305) );
  IV U36724 ( .A(n34790), .Z(n34793) );
  XNOR U36725 ( .A(n34790), .B(n27304), .Z(n34792) );
  XOR U36726 ( .A(n34794), .B(n34795), .Z(n27304) );
  AND U36727 ( .A(\modmult_1/xin[1023] ), .B(n34796), .Z(n34795) );
  IV U36728 ( .A(n34794), .Z(n34796) );
  XOR U36729 ( .A(n34797), .B(mreg[573]), .Z(n34794) );
  NAND U36730 ( .A(n34798), .B(mul_pow), .Z(n34797) );
  XOR U36731 ( .A(mreg[573]), .B(creg[573]), .Z(n34798) );
  XOR U36732 ( .A(n34799), .B(n34800), .Z(n34790) );
  ANDN U36733 ( .A(n34801), .B(n27311), .Z(n34800) );
  XOR U36734 ( .A(n34802), .B(\modmult_1/zin[0][571] ), .Z(n27311) );
  IV U36735 ( .A(n34799), .Z(n34802) );
  XNOR U36736 ( .A(n34799), .B(n27310), .Z(n34801) );
  XOR U36737 ( .A(n34803), .B(n34804), .Z(n27310) );
  AND U36738 ( .A(\modmult_1/xin[1023] ), .B(n34805), .Z(n34804) );
  IV U36739 ( .A(n34803), .Z(n34805) );
  XOR U36740 ( .A(n34806), .B(mreg[572]), .Z(n34803) );
  NAND U36741 ( .A(n34807), .B(mul_pow), .Z(n34806) );
  XOR U36742 ( .A(mreg[572]), .B(creg[572]), .Z(n34807) );
  XOR U36743 ( .A(n34808), .B(n34809), .Z(n34799) );
  ANDN U36744 ( .A(n34810), .B(n27317), .Z(n34809) );
  XOR U36745 ( .A(n34811), .B(\modmult_1/zin[0][570] ), .Z(n27317) );
  IV U36746 ( .A(n34808), .Z(n34811) );
  XNOR U36747 ( .A(n34808), .B(n27316), .Z(n34810) );
  XOR U36748 ( .A(n34812), .B(n34813), .Z(n27316) );
  AND U36749 ( .A(\modmult_1/xin[1023] ), .B(n34814), .Z(n34813) );
  IV U36750 ( .A(n34812), .Z(n34814) );
  XOR U36751 ( .A(n34815), .B(mreg[571]), .Z(n34812) );
  NAND U36752 ( .A(n34816), .B(mul_pow), .Z(n34815) );
  XOR U36753 ( .A(mreg[571]), .B(creg[571]), .Z(n34816) );
  XOR U36754 ( .A(n34817), .B(n34818), .Z(n34808) );
  ANDN U36755 ( .A(n34819), .B(n27323), .Z(n34818) );
  XOR U36756 ( .A(n34820), .B(\modmult_1/zin[0][569] ), .Z(n27323) );
  IV U36757 ( .A(n34817), .Z(n34820) );
  XNOR U36758 ( .A(n34817), .B(n27322), .Z(n34819) );
  XOR U36759 ( .A(n34821), .B(n34822), .Z(n27322) );
  AND U36760 ( .A(\modmult_1/xin[1023] ), .B(n34823), .Z(n34822) );
  IV U36761 ( .A(n34821), .Z(n34823) );
  XOR U36762 ( .A(n34824), .B(mreg[570]), .Z(n34821) );
  NAND U36763 ( .A(n34825), .B(mul_pow), .Z(n34824) );
  XOR U36764 ( .A(mreg[570]), .B(creg[570]), .Z(n34825) );
  XOR U36765 ( .A(n34826), .B(n34827), .Z(n34817) );
  ANDN U36766 ( .A(n34828), .B(n27329), .Z(n34827) );
  XOR U36767 ( .A(n34829), .B(\modmult_1/zin[0][568] ), .Z(n27329) );
  IV U36768 ( .A(n34826), .Z(n34829) );
  XNOR U36769 ( .A(n34826), .B(n27328), .Z(n34828) );
  XOR U36770 ( .A(n34830), .B(n34831), .Z(n27328) );
  AND U36771 ( .A(\modmult_1/xin[1023] ), .B(n34832), .Z(n34831) );
  IV U36772 ( .A(n34830), .Z(n34832) );
  XOR U36773 ( .A(n34833), .B(mreg[569]), .Z(n34830) );
  NAND U36774 ( .A(n34834), .B(mul_pow), .Z(n34833) );
  XOR U36775 ( .A(mreg[569]), .B(creg[569]), .Z(n34834) );
  XOR U36776 ( .A(n34835), .B(n34836), .Z(n34826) );
  ANDN U36777 ( .A(n34837), .B(n27335), .Z(n34836) );
  XOR U36778 ( .A(n34838), .B(\modmult_1/zin[0][567] ), .Z(n27335) );
  IV U36779 ( .A(n34835), .Z(n34838) );
  XNOR U36780 ( .A(n34835), .B(n27334), .Z(n34837) );
  XOR U36781 ( .A(n34839), .B(n34840), .Z(n27334) );
  AND U36782 ( .A(\modmult_1/xin[1023] ), .B(n34841), .Z(n34840) );
  IV U36783 ( .A(n34839), .Z(n34841) );
  XOR U36784 ( .A(n34842), .B(mreg[568]), .Z(n34839) );
  NAND U36785 ( .A(n34843), .B(mul_pow), .Z(n34842) );
  XOR U36786 ( .A(mreg[568]), .B(creg[568]), .Z(n34843) );
  XOR U36787 ( .A(n34844), .B(n34845), .Z(n34835) );
  ANDN U36788 ( .A(n34846), .B(n27341), .Z(n34845) );
  XOR U36789 ( .A(n34847), .B(\modmult_1/zin[0][566] ), .Z(n27341) );
  IV U36790 ( .A(n34844), .Z(n34847) );
  XNOR U36791 ( .A(n34844), .B(n27340), .Z(n34846) );
  XOR U36792 ( .A(n34848), .B(n34849), .Z(n27340) );
  AND U36793 ( .A(\modmult_1/xin[1023] ), .B(n34850), .Z(n34849) );
  IV U36794 ( .A(n34848), .Z(n34850) );
  XOR U36795 ( .A(n34851), .B(mreg[567]), .Z(n34848) );
  NAND U36796 ( .A(n34852), .B(mul_pow), .Z(n34851) );
  XOR U36797 ( .A(mreg[567]), .B(creg[567]), .Z(n34852) );
  XOR U36798 ( .A(n34853), .B(n34854), .Z(n34844) );
  ANDN U36799 ( .A(n34855), .B(n27347), .Z(n34854) );
  XOR U36800 ( .A(n34856), .B(\modmult_1/zin[0][565] ), .Z(n27347) );
  IV U36801 ( .A(n34853), .Z(n34856) );
  XNOR U36802 ( .A(n34853), .B(n27346), .Z(n34855) );
  XOR U36803 ( .A(n34857), .B(n34858), .Z(n27346) );
  AND U36804 ( .A(\modmult_1/xin[1023] ), .B(n34859), .Z(n34858) );
  IV U36805 ( .A(n34857), .Z(n34859) );
  XOR U36806 ( .A(n34860), .B(mreg[566]), .Z(n34857) );
  NAND U36807 ( .A(n34861), .B(mul_pow), .Z(n34860) );
  XOR U36808 ( .A(mreg[566]), .B(creg[566]), .Z(n34861) );
  XOR U36809 ( .A(n34862), .B(n34863), .Z(n34853) );
  ANDN U36810 ( .A(n34864), .B(n27353), .Z(n34863) );
  XOR U36811 ( .A(n34865), .B(\modmult_1/zin[0][564] ), .Z(n27353) );
  IV U36812 ( .A(n34862), .Z(n34865) );
  XNOR U36813 ( .A(n34862), .B(n27352), .Z(n34864) );
  XOR U36814 ( .A(n34866), .B(n34867), .Z(n27352) );
  AND U36815 ( .A(\modmult_1/xin[1023] ), .B(n34868), .Z(n34867) );
  IV U36816 ( .A(n34866), .Z(n34868) );
  XOR U36817 ( .A(n34869), .B(mreg[565]), .Z(n34866) );
  NAND U36818 ( .A(n34870), .B(mul_pow), .Z(n34869) );
  XOR U36819 ( .A(mreg[565]), .B(creg[565]), .Z(n34870) );
  XOR U36820 ( .A(n34871), .B(n34872), .Z(n34862) );
  ANDN U36821 ( .A(n34873), .B(n27359), .Z(n34872) );
  XOR U36822 ( .A(n34874), .B(\modmult_1/zin[0][563] ), .Z(n27359) );
  IV U36823 ( .A(n34871), .Z(n34874) );
  XNOR U36824 ( .A(n34871), .B(n27358), .Z(n34873) );
  XOR U36825 ( .A(n34875), .B(n34876), .Z(n27358) );
  AND U36826 ( .A(\modmult_1/xin[1023] ), .B(n34877), .Z(n34876) );
  IV U36827 ( .A(n34875), .Z(n34877) );
  XOR U36828 ( .A(n34878), .B(mreg[564]), .Z(n34875) );
  NAND U36829 ( .A(n34879), .B(mul_pow), .Z(n34878) );
  XOR U36830 ( .A(mreg[564]), .B(creg[564]), .Z(n34879) );
  XOR U36831 ( .A(n34880), .B(n34881), .Z(n34871) );
  ANDN U36832 ( .A(n34882), .B(n27365), .Z(n34881) );
  XOR U36833 ( .A(n34883), .B(\modmult_1/zin[0][562] ), .Z(n27365) );
  IV U36834 ( .A(n34880), .Z(n34883) );
  XNOR U36835 ( .A(n34880), .B(n27364), .Z(n34882) );
  XOR U36836 ( .A(n34884), .B(n34885), .Z(n27364) );
  AND U36837 ( .A(\modmult_1/xin[1023] ), .B(n34886), .Z(n34885) );
  IV U36838 ( .A(n34884), .Z(n34886) );
  XOR U36839 ( .A(n34887), .B(mreg[563]), .Z(n34884) );
  NAND U36840 ( .A(n34888), .B(mul_pow), .Z(n34887) );
  XOR U36841 ( .A(mreg[563]), .B(creg[563]), .Z(n34888) );
  XOR U36842 ( .A(n34889), .B(n34890), .Z(n34880) );
  ANDN U36843 ( .A(n34891), .B(n27371), .Z(n34890) );
  XOR U36844 ( .A(n34892), .B(\modmult_1/zin[0][561] ), .Z(n27371) );
  IV U36845 ( .A(n34889), .Z(n34892) );
  XNOR U36846 ( .A(n34889), .B(n27370), .Z(n34891) );
  XOR U36847 ( .A(n34893), .B(n34894), .Z(n27370) );
  AND U36848 ( .A(\modmult_1/xin[1023] ), .B(n34895), .Z(n34894) );
  IV U36849 ( .A(n34893), .Z(n34895) );
  XOR U36850 ( .A(n34896), .B(mreg[562]), .Z(n34893) );
  NAND U36851 ( .A(n34897), .B(mul_pow), .Z(n34896) );
  XOR U36852 ( .A(mreg[562]), .B(creg[562]), .Z(n34897) );
  XOR U36853 ( .A(n34898), .B(n34899), .Z(n34889) );
  ANDN U36854 ( .A(n34900), .B(n27377), .Z(n34899) );
  XOR U36855 ( .A(n34901), .B(\modmult_1/zin[0][560] ), .Z(n27377) );
  IV U36856 ( .A(n34898), .Z(n34901) );
  XNOR U36857 ( .A(n34898), .B(n27376), .Z(n34900) );
  XOR U36858 ( .A(n34902), .B(n34903), .Z(n27376) );
  AND U36859 ( .A(\modmult_1/xin[1023] ), .B(n34904), .Z(n34903) );
  IV U36860 ( .A(n34902), .Z(n34904) );
  XOR U36861 ( .A(n34905), .B(mreg[561]), .Z(n34902) );
  NAND U36862 ( .A(n34906), .B(mul_pow), .Z(n34905) );
  XOR U36863 ( .A(mreg[561]), .B(creg[561]), .Z(n34906) );
  XOR U36864 ( .A(n34907), .B(n34908), .Z(n34898) );
  ANDN U36865 ( .A(n34909), .B(n27383), .Z(n34908) );
  XOR U36866 ( .A(n34910), .B(\modmult_1/zin[0][559] ), .Z(n27383) );
  IV U36867 ( .A(n34907), .Z(n34910) );
  XNOR U36868 ( .A(n34907), .B(n27382), .Z(n34909) );
  XOR U36869 ( .A(n34911), .B(n34912), .Z(n27382) );
  AND U36870 ( .A(\modmult_1/xin[1023] ), .B(n34913), .Z(n34912) );
  IV U36871 ( .A(n34911), .Z(n34913) );
  XOR U36872 ( .A(n34914), .B(mreg[560]), .Z(n34911) );
  NAND U36873 ( .A(n34915), .B(mul_pow), .Z(n34914) );
  XOR U36874 ( .A(mreg[560]), .B(creg[560]), .Z(n34915) );
  XOR U36875 ( .A(n34916), .B(n34917), .Z(n34907) );
  ANDN U36876 ( .A(n34918), .B(n27389), .Z(n34917) );
  XOR U36877 ( .A(n34919), .B(\modmult_1/zin[0][558] ), .Z(n27389) );
  IV U36878 ( .A(n34916), .Z(n34919) );
  XNOR U36879 ( .A(n34916), .B(n27388), .Z(n34918) );
  XOR U36880 ( .A(n34920), .B(n34921), .Z(n27388) );
  AND U36881 ( .A(\modmult_1/xin[1023] ), .B(n34922), .Z(n34921) );
  IV U36882 ( .A(n34920), .Z(n34922) );
  XOR U36883 ( .A(n34923), .B(mreg[559]), .Z(n34920) );
  NAND U36884 ( .A(n34924), .B(mul_pow), .Z(n34923) );
  XOR U36885 ( .A(mreg[559]), .B(creg[559]), .Z(n34924) );
  XOR U36886 ( .A(n34925), .B(n34926), .Z(n34916) );
  ANDN U36887 ( .A(n34927), .B(n27395), .Z(n34926) );
  XOR U36888 ( .A(n34928), .B(\modmult_1/zin[0][557] ), .Z(n27395) );
  IV U36889 ( .A(n34925), .Z(n34928) );
  XNOR U36890 ( .A(n34925), .B(n27394), .Z(n34927) );
  XOR U36891 ( .A(n34929), .B(n34930), .Z(n27394) );
  AND U36892 ( .A(\modmult_1/xin[1023] ), .B(n34931), .Z(n34930) );
  IV U36893 ( .A(n34929), .Z(n34931) );
  XOR U36894 ( .A(n34932), .B(mreg[558]), .Z(n34929) );
  NAND U36895 ( .A(n34933), .B(mul_pow), .Z(n34932) );
  XOR U36896 ( .A(mreg[558]), .B(creg[558]), .Z(n34933) );
  XOR U36897 ( .A(n34934), .B(n34935), .Z(n34925) );
  ANDN U36898 ( .A(n34936), .B(n27401), .Z(n34935) );
  XOR U36899 ( .A(n34937), .B(\modmult_1/zin[0][556] ), .Z(n27401) );
  IV U36900 ( .A(n34934), .Z(n34937) );
  XNOR U36901 ( .A(n34934), .B(n27400), .Z(n34936) );
  XOR U36902 ( .A(n34938), .B(n34939), .Z(n27400) );
  AND U36903 ( .A(\modmult_1/xin[1023] ), .B(n34940), .Z(n34939) );
  IV U36904 ( .A(n34938), .Z(n34940) );
  XOR U36905 ( .A(n34941), .B(mreg[557]), .Z(n34938) );
  NAND U36906 ( .A(n34942), .B(mul_pow), .Z(n34941) );
  XOR U36907 ( .A(mreg[557]), .B(creg[557]), .Z(n34942) );
  XOR U36908 ( .A(n34943), .B(n34944), .Z(n34934) );
  ANDN U36909 ( .A(n34945), .B(n27407), .Z(n34944) );
  XOR U36910 ( .A(n34946), .B(\modmult_1/zin[0][555] ), .Z(n27407) );
  IV U36911 ( .A(n34943), .Z(n34946) );
  XNOR U36912 ( .A(n34943), .B(n27406), .Z(n34945) );
  XOR U36913 ( .A(n34947), .B(n34948), .Z(n27406) );
  AND U36914 ( .A(\modmult_1/xin[1023] ), .B(n34949), .Z(n34948) );
  IV U36915 ( .A(n34947), .Z(n34949) );
  XOR U36916 ( .A(n34950), .B(mreg[556]), .Z(n34947) );
  NAND U36917 ( .A(n34951), .B(mul_pow), .Z(n34950) );
  XOR U36918 ( .A(mreg[556]), .B(creg[556]), .Z(n34951) );
  XOR U36919 ( .A(n34952), .B(n34953), .Z(n34943) );
  ANDN U36920 ( .A(n34954), .B(n27413), .Z(n34953) );
  XOR U36921 ( .A(n34955), .B(\modmult_1/zin[0][554] ), .Z(n27413) );
  IV U36922 ( .A(n34952), .Z(n34955) );
  XNOR U36923 ( .A(n34952), .B(n27412), .Z(n34954) );
  XOR U36924 ( .A(n34956), .B(n34957), .Z(n27412) );
  AND U36925 ( .A(\modmult_1/xin[1023] ), .B(n34958), .Z(n34957) );
  IV U36926 ( .A(n34956), .Z(n34958) );
  XOR U36927 ( .A(n34959), .B(mreg[555]), .Z(n34956) );
  NAND U36928 ( .A(n34960), .B(mul_pow), .Z(n34959) );
  XOR U36929 ( .A(mreg[555]), .B(creg[555]), .Z(n34960) );
  XOR U36930 ( .A(n34961), .B(n34962), .Z(n34952) );
  ANDN U36931 ( .A(n34963), .B(n27419), .Z(n34962) );
  XOR U36932 ( .A(n34964), .B(\modmult_1/zin[0][553] ), .Z(n27419) );
  IV U36933 ( .A(n34961), .Z(n34964) );
  XNOR U36934 ( .A(n34961), .B(n27418), .Z(n34963) );
  XOR U36935 ( .A(n34965), .B(n34966), .Z(n27418) );
  AND U36936 ( .A(\modmult_1/xin[1023] ), .B(n34967), .Z(n34966) );
  IV U36937 ( .A(n34965), .Z(n34967) );
  XOR U36938 ( .A(n34968), .B(mreg[554]), .Z(n34965) );
  NAND U36939 ( .A(n34969), .B(mul_pow), .Z(n34968) );
  XOR U36940 ( .A(mreg[554]), .B(creg[554]), .Z(n34969) );
  XOR U36941 ( .A(n34970), .B(n34971), .Z(n34961) );
  ANDN U36942 ( .A(n34972), .B(n27425), .Z(n34971) );
  XOR U36943 ( .A(n34973), .B(\modmult_1/zin[0][552] ), .Z(n27425) );
  IV U36944 ( .A(n34970), .Z(n34973) );
  XNOR U36945 ( .A(n34970), .B(n27424), .Z(n34972) );
  XOR U36946 ( .A(n34974), .B(n34975), .Z(n27424) );
  AND U36947 ( .A(\modmult_1/xin[1023] ), .B(n34976), .Z(n34975) );
  IV U36948 ( .A(n34974), .Z(n34976) );
  XOR U36949 ( .A(n34977), .B(mreg[553]), .Z(n34974) );
  NAND U36950 ( .A(n34978), .B(mul_pow), .Z(n34977) );
  XOR U36951 ( .A(mreg[553]), .B(creg[553]), .Z(n34978) );
  XOR U36952 ( .A(n34979), .B(n34980), .Z(n34970) );
  ANDN U36953 ( .A(n34981), .B(n27431), .Z(n34980) );
  XOR U36954 ( .A(n34982), .B(\modmult_1/zin[0][551] ), .Z(n27431) );
  IV U36955 ( .A(n34979), .Z(n34982) );
  XNOR U36956 ( .A(n34979), .B(n27430), .Z(n34981) );
  XOR U36957 ( .A(n34983), .B(n34984), .Z(n27430) );
  AND U36958 ( .A(\modmult_1/xin[1023] ), .B(n34985), .Z(n34984) );
  IV U36959 ( .A(n34983), .Z(n34985) );
  XOR U36960 ( .A(n34986), .B(mreg[552]), .Z(n34983) );
  NAND U36961 ( .A(n34987), .B(mul_pow), .Z(n34986) );
  XOR U36962 ( .A(mreg[552]), .B(creg[552]), .Z(n34987) );
  XOR U36963 ( .A(n34988), .B(n34989), .Z(n34979) );
  ANDN U36964 ( .A(n34990), .B(n27437), .Z(n34989) );
  XOR U36965 ( .A(n34991), .B(\modmult_1/zin[0][550] ), .Z(n27437) );
  IV U36966 ( .A(n34988), .Z(n34991) );
  XNOR U36967 ( .A(n34988), .B(n27436), .Z(n34990) );
  XOR U36968 ( .A(n34992), .B(n34993), .Z(n27436) );
  AND U36969 ( .A(\modmult_1/xin[1023] ), .B(n34994), .Z(n34993) );
  IV U36970 ( .A(n34992), .Z(n34994) );
  XOR U36971 ( .A(n34995), .B(mreg[551]), .Z(n34992) );
  NAND U36972 ( .A(n34996), .B(mul_pow), .Z(n34995) );
  XOR U36973 ( .A(mreg[551]), .B(creg[551]), .Z(n34996) );
  XOR U36974 ( .A(n34997), .B(n34998), .Z(n34988) );
  ANDN U36975 ( .A(n34999), .B(n27443), .Z(n34998) );
  XOR U36976 ( .A(n35000), .B(\modmult_1/zin[0][549] ), .Z(n27443) );
  IV U36977 ( .A(n34997), .Z(n35000) );
  XNOR U36978 ( .A(n34997), .B(n27442), .Z(n34999) );
  XOR U36979 ( .A(n35001), .B(n35002), .Z(n27442) );
  AND U36980 ( .A(\modmult_1/xin[1023] ), .B(n35003), .Z(n35002) );
  IV U36981 ( .A(n35001), .Z(n35003) );
  XOR U36982 ( .A(n35004), .B(mreg[550]), .Z(n35001) );
  NAND U36983 ( .A(n35005), .B(mul_pow), .Z(n35004) );
  XOR U36984 ( .A(mreg[550]), .B(creg[550]), .Z(n35005) );
  XOR U36985 ( .A(n35006), .B(n35007), .Z(n34997) );
  ANDN U36986 ( .A(n35008), .B(n27449), .Z(n35007) );
  XOR U36987 ( .A(n35009), .B(\modmult_1/zin[0][548] ), .Z(n27449) );
  IV U36988 ( .A(n35006), .Z(n35009) );
  XNOR U36989 ( .A(n35006), .B(n27448), .Z(n35008) );
  XOR U36990 ( .A(n35010), .B(n35011), .Z(n27448) );
  AND U36991 ( .A(\modmult_1/xin[1023] ), .B(n35012), .Z(n35011) );
  IV U36992 ( .A(n35010), .Z(n35012) );
  XOR U36993 ( .A(n35013), .B(mreg[549]), .Z(n35010) );
  NAND U36994 ( .A(n35014), .B(mul_pow), .Z(n35013) );
  XOR U36995 ( .A(mreg[549]), .B(creg[549]), .Z(n35014) );
  XOR U36996 ( .A(n35015), .B(n35016), .Z(n35006) );
  ANDN U36997 ( .A(n35017), .B(n27455), .Z(n35016) );
  XOR U36998 ( .A(n35018), .B(\modmult_1/zin[0][547] ), .Z(n27455) );
  IV U36999 ( .A(n35015), .Z(n35018) );
  XNOR U37000 ( .A(n35015), .B(n27454), .Z(n35017) );
  XOR U37001 ( .A(n35019), .B(n35020), .Z(n27454) );
  AND U37002 ( .A(\modmult_1/xin[1023] ), .B(n35021), .Z(n35020) );
  IV U37003 ( .A(n35019), .Z(n35021) );
  XOR U37004 ( .A(n35022), .B(mreg[548]), .Z(n35019) );
  NAND U37005 ( .A(n35023), .B(mul_pow), .Z(n35022) );
  XOR U37006 ( .A(mreg[548]), .B(creg[548]), .Z(n35023) );
  XOR U37007 ( .A(n35024), .B(n35025), .Z(n35015) );
  ANDN U37008 ( .A(n35026), .B(n27461), .Z(n35025) );
  XOR U37009 ( .A(n35027), .B(\modmult_1/zin[0][546] ), .Z(n27461) );
  IV U37010 ( .A(n35024), .Z(n35027) );
  XNOR U37011 ( .A(n35024), .B(n27460), .Z(n35026) );
  XOR U37012 ( .A(n35028), .B(n35029), .Z(n27460) );
  AND U37013 ( .A(\modmult_1/xin[1023] ), .B(n35030), .Z(n35029) );
  IV U37014 ( .A(n35028), .Z(n35030) );
  XOR U37015 ( .A(n35031), .B(mreg[547]), .Z(n35028) );
  NAND U37016 ( .A(n35032), .B(mul_pow), .Z(n35031) );
  XOR U37017 ( .A(mreg[547]), .B(creg[547]), .Z(n35032) );
  XOR U37018 ( .A(n35033), .B(n35034), .Z(n35024) );
  ANDN U37019 ( .A(n35035), .B(n27467), .Z(n35034) );
  XOR U37020 ( .A(n35036), .B(\modmult_1/zin[0][545] ), .Z(n27467) );
  IV U37021 ( .A(n35033), .Z(n35036) );
  XNOR U37022 ( .A(n35033), .B(n27466), .Z(n35035) );
  XOR U37023 ( .A(n35037), .B(n35038), .Z(n27466) );
  AND U37024 ( .A(\modmult_1/xin[1023] ), .B(n35039), .Z(n35038) );
  IV U37025 ( .A(n35037), .Z(n35039) );
  XOR U37026 ( .A(n35040), .B(mreg[546]), .Z(n35037) );
  NAND U37027 ( .A(n35041), .B(mul_pow), .Z(n35040) );
  XOR U37028 ( .A(mreg[546]), .B(creg[546]), .Z(n35041) );
  XOR U37029 ( .A(n35042), .B(n35043), .Z(n35033) );
  ANDN U37030 ( .A(n35044), .B(n27473), .Z(n35043) );
  XOR U37031 ( .A(n35045), .B(\modmult_1/zin[0][544] ), .Z(n27473) );
  IV U37032 ( .A(n35042), .Z(n35045) );
  XNOR U37033 ( .A(n35042), .B(n27472), .Z(n35044) );
  XOR U37034 ( .A(n35046), .B(n35047), .Z(n27472) );
  AND U37035 ( .A(\modmult_1/xin[1023] ), .B(n35048), .Z(n35047) );
  IV U37036 ( .A(n35046), .Z(n35048) );
  XOR U37037 ( .A(n35049), .B(mreg[545]), .Z(n35046) );
  NAND U37038 ( .A(n35050), .B(mul_pow), .Z(n35049) );
  XOR U37039 ( .A(mreg[545]), .B(creg[545]), .Z(n35050) );
  XOR U37040 ( .A(n35051), .B(n35052), .Z(n35042) );
  ANDN U37041 ( .A(n35053), .B(n27479), .Z(n35052) );
  XOR U37042 ( .A(n35054), .B(\modmult_1/zin[0][543] ), .Z(n27479) );
  IV U37043 ( .A(n35051), .Z(n35054) );
  XNOR U37044 ( .A(n35051), .B(n27478), .Z(n35053) );
  XOR U37045 ( .A(n35055), .B(n35056), .Z(n27478) );
  AND U37046 ( .A(\modmult_1/xin[1023] ), .B(n35057), .Z(n35056) );
  IV U37047 ( .A(n35055), .Z(n35057) );
  XOR U37048 ( .A(n35058), .B(mreg[544]), .Z(n35055) );
  NAND U37049 ( .A(n35059), .B(mul_pow), .Z(n35058) );
  XOR U37050 ( .A(mreg[544]), .B(creg[544]), .Z(n35059) );
  XOR U37051 ( .A(n35060), .B(n35061), .Z(n35051) );
  ANDN U37052 ( .A(n35062), .B(n27485), .Z(n35061) );
  XOR U37053 ( .A(n35063), .B(\modmult_1/zin[0][542] ), .Z(n27485) );
  IV U37054 ( .A(n35060), .Z(n35063) );
  XNOR U37055 ( .A(n35060), .B(n27484), .Z(n35062) );
  XOR U37056 ( .A(n35064), .B(n35065), .Z(n27484) );
  AND U37057 ( .A(\modmult_1/xin[1023] ), .B(n35066), .Z(n35065) );
  IV U37058 ( .A(n35064), .Z(n35066) );
  XOR U37059 ( .A(n35067), .B(mreg[543]), .Z(n35064) );
  NAND U37060 ( .A(n35068), .B(mul_pow), .Z(n35067) );
  XOR U37061 ( .A(mreg[543]), .B(creg[543]), .Z(n35068) );
  XOR U37062 ( .A(n35069), .B(n35070), .Z(n35060) );
  ANDN U37063 ( .A(n35071), .B(n27491), .Z(n35070) );
  XOR U37064 ( .A(n35072), .B(\modmult_1/zin[0][541] ), .Z(n27491) );
  IV U37065 ( .A(n35069), .Z(n35072) );
  XNOR U37066 ( .A(n35069), .B(n27490), .Z(n35071) );
  XOR U37067 ( .A(n35073), .B(n35074), .Z(n27490) );
  AND U37068 ( .A(\modmult_1/xin[1023] ), .B(n35075), .Z(n35074) );
  IV U37069 ( .A(n35073), .Z(n35075) );
  XOR U37070 ( .A(n35076), .B(mreg[542]), .Z(n35073) );
  NAND U37071 ( .A(n35077), .B(mul_pow), .Z(n35076) );
  XOR U37072 ( .A(mreg[542]), .B(creg[542]), .Z(n35077) );
  XOR U37073 ( .A(n35078), .B(n35079), .Z(n35069) );
  ANDN U37074 ( .A(n35080), .B(n27497), .Z(n35079) );
  XOR U37075 ( .A(n35081), .B(\modmult_1/zin[0][540] ), .Z(n27497) );
  IV U37076 ( .A(n35078), .Z(n35081) );
  XNOR U37077 ( .A(n35078), .B(n27496), .Z(n35080) );
  XOR U37078 ( .A(n35082), .B(n35083), .Z(n27496) );
  AND U37079 ( .A(\modmult_1/xin[1023] ), .B(n35084), .Z(n35083) );
  IV U37080 ( .A(n35082), .Z(n35084) );
  XOR U37081 ( .A(n35085), .B(mreg[541]), .Z(n35082) );
  NAND U37082 ( .A(n35086), .B(mul_pow), .Z(n35085) );
  XOR U37083 ( .A(mreg[541]), .B(creg[541]), .Z(n35086) );
  XOR U37084 ( .A(n35087), .B(n35088), .Z(n35078) );
  ANDN U37085 ( .A(n35089), .B(n27503), .Z(n35088) );
  XOR U37086 ( .A(n35090), .B(\modmult_1/zin[0][539] ), .Z(n27503) );
  IV U37087 ( .A(n35087), .Z(n35090) );
  XNOR U37088 ( .A(n35087), .B(n27502), .Z(n35089) );
  XOR U37089 ( .A(n35091), .B(n35092), .Z(n27502) );
  AND U37090 ( .A(\modmult_1/xin[1023] ), .B(n35093), .Z(n35092) );
  IV U37091 ( .A(n35091), .Z(n35093) );
  XOR U37092 ( .A(n35094), .B(mreg[540]), .Z(n35091) );
  NAND U37093 ( .A(n35095), .B(mul_pow), .Z(n35094) );
  XOR U37094 ( .A(mreg[540]), .B(creg[540]), .Z(n35095) );
  XOR U37095 ( .A(n35096), .B(n35097), .Z(n35087) );
  ANDN U37096 ( .A(n35098), .B(n27509), .Z(n35097) );
  XOR U37097 ( .A(n35099), .B(\modmult_1/zin[0][538] ), .Z(n27509) );
  IV U37098 ( .A(n35096), .Z(n35099) );
  XNOR U37099 ( .A(n35096), .B(n27508), .Z(n35098) );
  XOR U37100 ( .A(n35100), .B(n35101), .Z(n27508) );
  AND U37101 ( .A(\modmult_1/xin[1023] ), .B(n35102), .Z(n35101) );
  IV U37102 ( .A(n35100), .Z(n35102) );
  XOR U37103 ( .A(n35103), .B(mreg[539]), .Z(n35100) );
  NAND U37104 ( .A(n35104), .B(mul_pow), .Z(n35103) );
  XOR U37105 ( .A(mreg[539]), .B(creg[539]), .Z(n35104) );
  XOR U37106 ( .A(n35105), .B(n35106), .Z(n35096) );
  ANDN U37107 ( .A(n35107), .B(n27515), .Z(n35106) );
  XOR U37108 ( .A(n35108), .B(\modmult_1/zin[0][537] ), .Z(n27515) );
  IV U37109 ( .A(n35105), .Z(n35108) );
  XNOR U37110 ( .A(n35105), .B(n27514), .Z(n35107) );
  XOR U37111 ( .A(n35109), .B(n35110), .Z(n27514) );
  AND U37112 ( .A(\modmult_1/xin[1023] ), .B(n35111), .Z(n35110) );
  IV U37113 ( .A(n35109), .Z(n35111) );
  XOR U37114 ( .A(n35112), .B(mreg[538]), .Z(n35109) );
  NAND U37115 ( .A(n35113), .B(mul_pow), .Z(n35112) );
  XOR U37116 ( .A(mreg[538]), .B(creg[538]), .Z(n35113) );
  XOR U37117 ( .A(n35114), .B(n35115), .Z(n35105) );
  ANDN U37118 ( .A(n35116), .B(n27521), .Z(n35115) );
  XOR U37119 ( .A(n35117), .B(\modmult_1/zin[0][536] ), .Z(n27521) );
  IV U37120 ( .A(n35114), .Z(n35117) );
  XNOR U37121 ( .A(n35114), .B(n27520), .Z(n35116) );
  XOR U37122 ( .A(n35118), .B(n35119), .Z(n27520) );
  AND U37123 ( .A(\modmult_1/xin[1023] ), .B(n35120), .Z(n35119) );
  IV U37124 ( .A(n35118), .Z(n35120) );
  XOR U37125 ( .A(n35121), .B(mreg[537]), .Z(n35118) );
  NAND U37126 ( .A(n35122), .B(mul_pow), .Z(n35121) );
  XOR U37127 ( .A(mreg[537]), .B(creg[537]), .Z(n35122) );
  XOR U37128 ( .A(n35123), .B(n35124), .Z(n35114) );
  ANDN U37129 ( .A(n35125), .B(n27527), .Z(n35124) );
  XOR U37130 ( .A(n35126), .B(\modmult_1/zin[0][535] ), .Z(n27527) );
  IV U37131 ( .A(n35123), .Z(n35126) );
  XNOR U37132 ( .A(n35123), .B(n27526), .Z(n35125) );
  XOR U37133 ( .A(n35127), .B(n35128), .Z(n27526) );
  AND U37134 ( .A(\modmult_1/xin[1023] ), .B(n35129), .Z(n35128) );
  IV U37135 ( .A(n35127), .Z(n35129) );
  XOR U37136 ( .A(n35130), .B(mreg[536]), .Z(n35127) );
  NAND U37137 ( .A(n35131), .B(mul_pow), .Z(n35130) );
  XOR U37138 ( .A(mreg[536]), .B(creg[536]), .Z(n35131) );
  XOR U37139 ( .A(n35132), .B(n35133), .Z(n35123) );
  ANDN U37140 ( .A(n35134), .B(n27533), .Z(n35133) );
  XOR U37141 ( .A(n35135), .B(\modmult_1/zin[0][534] ), .Z(n27533) );
  IV U37142 ( .A(n35132), .Z(n35135) );
  XNOR U37143 ( .A(n35132), .B(n27532), .Z(n35134) );
  XOR U37144 ( .A(n35136), .B(n35137), .Z(n27532) );
  AND U37145 ( .A(\modmult_1/xin[1023] ), .B(n35138), .Z(n35137) );
  IV U37146 ( .A(n35136), .Z(n35138) );
  XOR U37147 ( .A(n35139), .B(mreg[535]), .Z(n35136) );
  NAND U37148 ( .A(n35140), .B(mul_pow), .Z(n35139) );
  XOR U37149 ( .A(mreg[535]), .B(creg[535]), .Z(n35140) );
  XOR U37150 ( .A(n35141), .B(n35142), .Z(n35132) );
  ANDN U37151 ( .A(n35143), .B(n27539), .Z(n35142) );
  XOR U37152 ( .A(n35144), .B(\modmult_1/zin[0][533] ), .Z(n27539) );
  IV U37153 ( .A(n35141), .Z(n35144) );
  XNOR U37154 ( .A(n35141), .B(n27538), .Z(n35143) );
  XOR U37155 ( .A(n35145), .B(n35146), .Z(n27538) );
  AND U37156 ( .A(\modmult_1/xin[1023] ), .B(n35147), .Z(n35146) );
  IV U37157 ( .A(n35145), .Z(n35147) );
  XOR U37158 ( .A(n35148), .B(mreg[534]), .Z(n35145) );
  NAND U37159 ( .A(n35149), .B(mul_pow), .Z(n35148) );
  XOR U37160 ( .A(mreg[534]), .B(creg[534]), .Z(n35149) );
  XOR U37161 ( .A(n35150), .B(n35151), .Z(n35141) );
  ANDN U37162 ( .A(n35152), .B(n27545), .Z(n35151) );
  XOR U37163 ( .A(n35153), .B(\modmult_1/zin[0][532] ), .Z(n27545) );
  IV U37164 ( .A(n35150), .Z(n35153) );
  XNOR U37165 ( .A(n35150), .B(n27544), .Z(n35152) );
  XOR U37166 ( .A(n35154), .B(n35155), .Z(n27544) );
  AND U37167 ( .A(\modmult_1/xin[1023] ), .B(n35156), .Z(n35155) );
  IV U37168 ( .A(n35154), .Z(n35156) );
  XOR U37169 ( .A(n35157), .B(mreg[533]), .Z(n35154) );
  NAND U37170 ( .A(n35158), .B(mul_pow), .Z(n35157) );
  XOR U37171 ( .A(mreg[533]), .B(creg[533]), .Z(n35158) );
  XOR U37172 ( .A(n35159), .B(n35160), .Z(n35150) );
  ANDN U37173 ( .A(n35161), .B(n27551), .Z(n35160) );
  XOR U37174 ( .A(n35162), .B(\modmult_1/zin[0][531] ), .Z(n27551) );
  IV U37175 ( .A(n35159), .Z(n35162) );
  XNOR U37176 ( .A(n35159), .B(n27550), .Z(n35161) );
  XOR U37177 ( .A(n35163), .B(n35164), .Z(n27550) );
  AND U37178 ( .A(\modmult_1/xin[1023] ), .B(n35165), .Z(n35164) );
  IV U37179 ( .A(n35163), .Z(n35165) );
  XOR U37180 ( .A(n35166), .B(mreg[532]), .Z(n35163) );
  NAND U37181 ( .A(n35167), .B(mul_pow), .Z(n35166) );
  XOR U37182 ( .A(mreg[532]), .B(creg[532]), .Z(n35167) );
  XOR U37183 ( .A(n35168), .B(n35169), .Z(n35159) );
  ANDN U37184 ( .A(n35170), .B(n27557), .Z(n35169) );
  XOR U37185 ( .A(n35171), .B(\modmult_1/zin[0][530] ), .Z(n27557) );
  IV U37186 ( .A(n35168), .Z(n35171) );
  XNOR U37187 ( .A(n35168), .B(n27556), .Z(n35170) );
  XOR U37188 ( .A(n35172), .B(n35173), .Z(n27556) );
  AND U37189 ( .A(\modmult_1/xin[1023] ), .B(n35174), .Z(n35173) );
  IV U37190 ( .A(n35172), .Z(n35174) );
  XOR U37191 ( .A(n35175), .B(mreg[531]), .Z(n35172) );
  NAND U37192 ( .A(n35176), .B(mul_pow), .Z(n35175) );
  XOR U37193 ( .A(mreg[531]), .B(creg[531]), .Z(n35176) );
  XOR U37194 ( .A(n35177), .B(n35178), .Z(n35168) );
  ANDN U37195 ( .A(n35179), .B(n27563), .Z(n35178) );
  XOR U37196 ( .A(n35180), .B(\modmult_1/zin[0][529] ), .Z(n27563) );
  IV U37197 ( .A(n35177), .Z(n35180) );
  XNOR U37198 ( .A(n35177), .B(n27562), .Z(n35179) );
  XOR U37199 ( .A(n35181), .B(n35182), .Z(n27562) );
  AND U37200 ( .A(\modmult_1/xin[1023] ), .B(n35183), .Z(n35182) );
  IV U37201 ( .A(n35181), .Z(n35183) );
  XOR U37202 ( .A(n35184), .B(mreg[530]), .Z(n35181) );
  NAND U37203 ( .A(n35185), .B(mul_pow), .Z(n35184) );
  XOR U37204 ( .A(mreg[530]), .B(creg[530]), .Z(n35185) );
  XOR U37205 ( .A(n35186), .B(n35187), .Z(n35177) );
  ANDN U37206 ( .A(n35188), .B(n27569), .Z(n35187) );
  XOR U37207 ( .A(n35189), .B(\modmult_1/zin[0][528] ), .Z(n27569) );
  IV U37208 ( .A(n35186), .Z(n35189) );
  XNOR U37209 ( .A(n35186), .B(n27568), .Z(n35188) );
  XOR U37210 ( .A(n35190), .B(n35191), .Z(n27568) );
  AND U37211 ( .A(\modmult_1/xin[1023] ), .B(n35192), .Z(n35191) );
  IV U37212 ( .A(n35190), .Z(n35192) );
  XOR U37213 ( .A(n35193), .B(mreg[529]), .Z(n35190) );
  NAND U37214 ( .A(n35194), .B(mul_pow), .Z(n35193) );
  XOR U37215 ( .A(mreg[529]), .B(creg[529]), .Z(n35194) );
  XOR U37216 ( .A(n35195), .B(n35196), .Z(n35186) );
  ANDN U37217 ( .A(n35197), .B(n27575), .Z(n35196) );
  XOR U37218 ( .A(n35198), .B(\modmult_1/zin[0][527] ), .Z(n27575) );
  IV U37219 ( .A(n35195), .Z(n35198) );
  XNOR U37220 ( .A(n35195), .B(n27574), .Z(n35197) );
  XOR U37221 ( .A(n35199), .B(n35200), .Z(n27574) );
  AND U37222 ( .A(\modmult_1/xin[1023] ), .B(n35201), .Z(n35200) );
  IV U37223 ( .A(n35199), .Z(n35201) );
  XOR U37224 ( .A(n35202), .B(mreg[528]), .Z(n35199) );
  NAND U37225 ( .A(n35203), .B(mul_pow), .Z(n35202) );
  XOR U37226 ( .A(mreg[528]), .B(creg[528]), .Z(n35203) );
  XOR U37227 ( .A(n35204), .B(n35205), .Z(n35195) );
  ANDN U37228 ( .A(n35206), .B(n27581), .Z(n35205) );
  XOR U37229 ( .A(n35207), .B(\modmult_1/zin[0][526] ), .Z(n27581) );
  IV U37230 ( .A(n35204), .Z(n35207) );
  XNOR U37231 ( .A(n35204), .B(n27580), .Z(n35206) );
  XOR U37232 ( .A(n35208), .B(n35209), .Z(n27580) );
  AND U37233 ( .A(\modmult_1/xin[1023] ), .B(n35210), .Z(n35209) );
  IV U37234 ( .A(n35208), .Z(n35210) );
  XOR U37235 ( .A(n35211), .B(mreg[527]), .Z(n35208) );
  NAND U37236 ( .A(n35212), .B(mul_pow), .Z(n35211) );
  XOR U37237 ( .A(mreg[527]), .B(creg[527]), .Z(n35212) );
  XOR U37238 ( .A(n35213), .B(n35214), .Z(n35204) );
  ANDN U37239 ( .A(n35215), .B(n27587), .Z(n35214) );
  XOR U37240 ( .A(n35216), .B(\modmult_1/zin[0][525] ), .Z(n27587) );
  IV U37241 ( .A(n35213), .Z(n35216) );
  XNOR U37242 ( .A(n35213), .B(n27586), .Z(n35215) );
  XOR U37243 ( .A(n35217), .B(n35218), .Z(n27586) );
  AND U37244 ( .A(\modmult_1/xin[1023] ), .B(n35219), .Z(n35218) );
  IV U37245 ( .A(n35217), .Z(n35219) );
  XOR U37246 ( .A(n35220), .B(mreg[526]), .Z(n35217) );
  NAND U37247 ( .A(n35221), .B(mul_pow), .Z(n35220) );
  XOR U37248 ( .A(mreg[526]), .B(creg[526]), .Z(n35221) );
  XOR U37249 ( .A(n35222), .B(n35223), .Z(n35213) );
  ANDN U37250 ( .A(n35224), .B(n27593), .Z(n35223) );
  XOR U37251 ( .A(n35225), .B(\modmult_1/zin[0][524] ), .Z(n27593) );
  IV U37252 ( .A(n35222), .Z(n35225) );
  XNOR U37253 ( .A(n35222), .B(n27592), .Z(n35224) );
  XOR U37254 ( .A(n35226), .B(n35227), .Z(n27592) );
  AND U37255 ( .A(\modmult_1/xin[1023] ), .B(n35228), .Z(n35227) );
  IV U37256 ( .A(n35226), .Z(n35228) );
  XOR U37257 ( .A(n35229), .B(mreg[525]), .Z(n35226) );
  NAND U37258 ( .A(n35230), .B(mul_pow), .Z(n35229) );
  XOR U37259 ( .A(mreg[525]), .B(creg[525]), .Z(n35230) );
  XOR U37260 ( .A(n35231), .B(n35232), .Z(n35222) );
  ANDN U37261 ( .A(n35233), .B(n27599), .Z(n35232) );
  XOR U37262 ( .A(n35234), .B(\modmult_1/zin[0][523] ), .Z(n27599) );
  IV U37263 ( .A(n35231), .Z(n35234) );
  XNOR U37264 ( .A(n35231), .B(n27598), .Z(n35233) );
  XOR U37265 ( .A(n35235), .B(n35236), .Z(n27598) );
  AND U37266 ( .A(\modmult_1/xin[1023] ), .B(n35237), .Z(n35236) );
  IV U37267 ( .A(n35235), .Z(n35237) );
  XOR U37268 ( .A(n35238), .B(mreg[524]), .Z(n35235) );
  NAND U37269 ( .A(n35239), .B(mul_pow), .Z(n35238) );
  XOR U37270 ( .A(mreg[524]), .B(creg[524]), .Z(n35239) );
  XOR U37271 ( .A(n35240), .B(n35241), .Z(n35231) );
  ANDN U37272 ( .A(n35242), .B(n27605), .Z(n35241) );
  XOR U37273 ( .A(n35243), .B(\modmult_1/zin[0][522] ), .Z(n27605) );
  IV U37274 ( .A(n35240), .Z(n35243) );
  XNOR U37275 ( .A(n35240), .B(n27604), .Z(n35242) );
  XOR U37276 ( .A(n35244), .B(n35245), .Z(n27604) );
  AND U37277 ( .A(\modmult_1/xin[1023] ), .B(n35246), .Z(n35245) );
  IV U37278 ( .A(n35244), .Z(n35246) );
  XOR U37279 ( .A(n35247), .B(mreg[523]), .Z(n35244) );
  NAND U37280 ( .A(n35248), .B(mul_pow), .Z(n35247) );
  XOR U37281 ( .A(mreg[523]), .B(creg[523]), .Z(n35248) );
  XOR U37282 ( .A(n35249), .B(n35250), .Z(n35240) );
  ANDN U37283 ( .A(n35251), .B(n27611), .Z(n35250) );
  XOR U37284 ( .A(n35252), .B(\modmult_1/zin[0][521] ), .Z(n27611) );
  IV U37285 ( .A(n35249), .Z(n35252) );
  XNOR U37286 ( .A(n35249), .B(n27610), .Z(n35251) );
  XOR U37287 ( .A(n35253), .B(n35254), .Z(n27610) );
  AND U37288 ( .A(\modmult_1/xin[1023] ), .B(n35255), .Z(n35254) );
  IV U37289 ( .A(n35253), .Z(n35255) );
  XOR U37290 ( .A(n35256), .B(mreg[522]), .Z(n35253) );
  NAND U37291 ( .A(n35257), .B(mul_pow), .Z(n35256) );
  XOR U37292 ( .A(mreg[522]), .B(creg[522]), .Z(n35257) );
  XOR U37293 ( .A(n35258), .B(n35259), .Z(n35249) );
  ANDN U37294 ( .A(n35260), .B(n27617), .Z(n35259) );
  XOR U37295 ( .A(n35261), .B(\modmult_1/zin[0][520] ), .Z(n27617) );
  IV U37296 ( .A(n35258), .Z(n35261) );
  XNOR U37297 ( .A(n35258), .B(n27616), .Z(n35260) );
  XOR U37298 ( .A(n35262), .B(n35263), .Z(n27616) );
  AND U37299 ( .A(\modmult_1/xin[1023] ), .B(n35264), .Z(n35263) );
  IV U37300 ( .A(n35262), .Z(n35264) );
  XOR U37301 ( .A(n35265), .B(mreg[521]), .Z(n35262) );
  NAND U37302 ( .A(n35266), .B(mul_pow), .Z(n35265) );
  XOR U37303 ( .A(mreg[521]), .B(creg[521]), .Z(n35266) );
  XOR U37304 ( .A(n35267), .B(n35268), .Z(n35258) );
  ANDN U37305 ( .A(n35269), .B(n27623), .Z(n35268) );
  XOR U37306 ( .A(n35270), .B(\modmult_1/zin[0][519] ), .Z(n27623) );
  IV U37307 ( .A(n35267), .Z(n35270) );
  XNOR U37308 ( .A(n35267), .B(n27622), .Z(n35269) );
  XOR U37309 ( .A(n35271), .B(n35272), .Z(n27622) );
  AND U37310 ( .A(\modmult_1/xin[1023] ), .B(n35273), .Z(n35272) );
  IV U37311 ( .A(n35271), .Z(n35273) );
  XOR U37312 ( .A(n35274), .B(mreg[520]), .Z(n35271) );
  NAND U37313 ( .A(n35275), .B(mul_pow), .Z(n35274) );
  XOR U37314 ( .A(mreg[520]), .B(creg[520]), .Z(n35275) );
  XOR U37315 ( .A(n35276), .B(n35277), .Z(n35267) );
  ANDN U37316 ( .A(n35278), .B(n27629), .Z(n35277) );
  XOR U37317 ( .A(n35279), .B(\modmult_1/zin[0][518] ), .Z(n27629) );
  IV U37318 ( .A(n35276), .Z(n35279) );
  XNOR U37319 ( .A(n35276), .B(n27628), .Z(n35278) );
  XOR U37320 ( .A(n35280), .B(n35281), .Z(n27628) );
  AND U37321 ( .A(\modmult_1/xin[1023] ), .B(n35282), .Z(n35281) );
  IV U37322 ( .A(n35280), .Z(n35282) );
  XOR U37323 ( .A(n35283), .B(mreg[519]), .Z(n35280) );
  NAND U37324 ( .A(n35284), .B(mul_pow), .Z(n35283) );
  XOR U37325 ( .A(mreg[519]), .B(creg[519]), .Z(n35284) );
  XOR U37326 ( .A(n35285), .B(n35286), .Z(n35276) );
  ANDN U37327 ( .A(n35287), .B(n27635), .Z(n35286) );
  XOR U37328 ( .A(n35288), .B(\modmult_1/zin[0][517] ), .Z(n27635) );
  IV U37329 ( .A(n35285), .Z(n35288) );
  XNOR U37330 ( .A(n35285), .B(n27634), .Z(n35287) );
  XOR U37331 ( .A(n35289), .B(n35290), .Z(n27634) );
  AND U37332 ( .A(\modmult_1/xin[1023] ), .B(n35291), .Z(n35290) );
  IV U37333 ( .A(n35289), .Z(n35291) );
  XOR U37334 ( .A(n35292), .B(mreg[518]), .Z(n35289) );
  NAND U37335 ( .A(n35293), .B(mul_pow), .Z(n35292) );
  XOR U37336 ( .A(mreg[518]), .B(creg[518]), .Z(n35293) );
  XOR U37337 ( .A(n35294), .B(n35295), .Z(n35285) );
  ANDN U37338 ( .A(n35296), .B(n27641), .Z(n35295) );
  XOR U37339 ( .A(n35297), .B(\modmult_1/zin[0][516] ), .Z(n27641) );
  IV U37340 ( .A(n35294), .Z(n35297) );
  XNOR U37341 ( .A(n35294), .B(n27640), .Z(n35296) );
  XOR U37342 ( .A(n35298), .B(n35299), .Z(n27640) );
  AND U37343 ( .A(\modmult_1/xin[1023] ), .B(n35300), .Z(n35299) );
  IV U37344 ( .A(n35298), .Z(n35300) );
  XOR U37345 ( .A(n35301), .B(mreg[517]), .Z(n35298) );
  NAND U37346 ( .A(n35302), .B(mul_pow), .Z(n35301) );
  XOR U37347 ( .A(mreg[517]), .B(creg[517]), .Z(n35302) );
  XOR U37348 ( .A(n35303), .B(n35304), .Z(n35294) );
  ANDN U37349 ( .A(n35305), .B(n27647), .Z(n35304) );
  XOR U37350 ( .A(n35306), .B(\modmult_1/zin[0][515] ), .Z(n27647) );
  IV U37351 ( .A(n35303), .Z(n35306) );
  XNOR U37352 ( .A(n35303), .B(n27646), .Z(n35305) );
  XOR U37353 ( .A(n35307), .B(n35308), .Z(n27646) );
  AND U37354 ( .A(\modmult_1/xin[1023] ), .B(n35309), .Z(n35308) );
  IV U37355 ( .A(n35307), .Z(n35309) );
  XOR U37356 ( .A(n35310), .B(mreg[516]), .Z(n35307) );
  NAND U37357 ( .A(n35311), .B(mul_pow), .Z(n35310) );
  XOR U37358 ( .A(mreg[516]), .B(creg[516]), .Z(n35311) );
  XOR U37359 ( .A(n35312), .B(n35313), .Z(n35303) );
  ANDN U37360 ( .A(n35314), .B(n27653), .Z(n35313) );
  XOR U37361 ( .A(n35315), .B(\modmult_1/zin[0][514] ), .Z(n27653) );
  IV U37362 ( .A(n35312), .Z(n35315) );
  XNOR U37363 ( .A(n35312), .B(n27652), .Z(n35314) );
  XOR U37364 ( .A(n35316), .B(n35317), .Z(n27652) );
  AND U37365 ( .A(\modmult_1/xin[1023] ), .B(n35318), .Z(n35317) );
  IV U37366 ( .A(n35316), .Z(n35318) );
  XOR U37367 ( .A(n35319), .B(mreg[515]), .Z(n35316) );
  NAND U37368 ( .A(n35320), .B(mul_pow), .Z(n35319) );
  XOR U37369 ( .A(mreg[515]), .B(creg[515]), .Z(n35320) );
  XOR U37370 ( .A(n35321), .B(n35322), .Z(n35312) );
  ANDN U37371 ( .A(n35323), .B(n27659), .Z(n35322) );
  XOR U37372 ( .A(n35324), .B(\modmult_1/zin[0][513] ), .Z(n27659) );
  IV U37373 ( .A(n35321), .Z(n35324) );
  XNOR U37374 ( .A(n35321), .B(n27658), .Z(n35323) );
  XOR U37375 ( .A(n35325), .B(n35326), .Z(n27658) );
  AND U37376 ( .A(\modmult_1/xin[1023] ), .B(n35327), .Z(n35326) );
  IV U37377 ( .A(n35325), .Z(n35327) );
  XOR U37378 ( .A(n35328), .B(mreg[514]), .Z(n35325) );
  NAND U37379 ( .A(n35329), .B(mul_pow), .Z(n35328) );
  XOR U37380 ( .A(mreg[514]), .B(creg[514]), .Z(n35329) );
  XOR U37381 ( .A(n35330), .B(n35331), .Z(n35321) );
  ANDN U37382 ( .A(n35332), .B(n27665), .Z(n35331) );
  XOR U37383 ( .A(n35333), .B(\modmult_1/zin[0][512] ), .Z(n27665) );
  IV U37384 ( .A(n35330), .Z(n35333) );
  XNOR U37385 ( .A(n35330), .B(n27664), .Z(n35332) );
  XOR U37386 ( .A(n35334), .B(n35335), .Z(n27664) );
  AND U37387 ( .A(\modmult_1/xin[1023] ), .B(n35336), .Z(n35335) );
  IV U37388 ( .A(n35334), .Z(n35336) );
  XOR U37389 ( .A(n35337), .B(mreg[513]), .Z(n35334) );
  NAND U37390 ( .A(n35338), .B(mul_pow), .Z(n35337) );
  XOR U37391 ( .A(mreg[513]), .B(creg[513]), .Z(n35338) );
  XOR U37392 ( .A(n35339), .B(n35340), .Z(n35330) );
  ANDN U37393 ( .A(n35341), .B(n27671), .Z(n35340) );
  XOR U37394 ( .A(n35342), .B(\modmult_1/zin[0][511] ), .Z(n27671) );
  IV U37395 ( .A(n35339), .Z(n35342) );
  XNOR U37396 ( .A(n35339), .B(n27670), .Z(n35341) );
  XOR U37397 ( .A(n35343), .B(n35344), .Z(n27670) );
  AND U37398 ( .A(\modmult_1/xin[1023] ), .B(n35345), .Z(n35344) );
  IV U37399 ( .A(n35343), .Z(n35345) );
  XOR U37400 ( .A(n35346), .B(mreg[512]), .Z(n35343) );
  NAND U37401 ( .A(n35347), .B(mul_pow), .Z(n35346) );
  XOR U37402 ( .A(mreg[512]), .B(creg[512]), .Z(n35347) );
  XOR U37403 ( .A(n35348), .B(n35349), .Z(n35339) );
  ANDN U37404 ( .A(n35350), .B(n27677), .Z(n35349) );
  XOR U37405 ( .A(n35351), .B(\modmult_1/zin[0][510] ), .Z(n27677) );
  IV U37406 ( .A(n35348), .Z(n35351) );
  XNOR U37407 ( .A(n35348), .B(n27676), .Z(n35350) );
  XOR U37408 ( .A(n35352), .B(n35353), .Z(n27676) );
  AND U37409 ( .A(\modmult_1/xin[1023] ), .B(n35354), .Z(n35353) );
  IV U37410 ( .A(n35352), .Z(n35354) );
  XOR U37411 ( .A(n35355), .B(mreg[511]), .Z(n35352) );
  NAND U37412 ( .A(n35356), .B(mul_pow), .Z(n35355) );
  XOR U37413 ( .A(mreg[511]), .B(creg[511]), .Z(n35356) );
  XOR U37414 ( .A(n35357), .B(n35358), .Z(n35348) );
  ANDN U37415 ( .A(n35359), .B(n27683), .Z(n35358) );
  XOR U37416 ( .A(n35360), .B(\modmult_1/zin[0][509] ), .Z(n27683) );
  IV U37417 ( .A(n35357), .Z(n35360) );
  XNOR U37418 ( .A(n35357), .B(n27682), .Z(n35359) );
  XOR U37419 ( .A(n35361), .B(n35362), .Z(n27682) );
  AND U37420 ( .A(\modmult_1/xin[1023] ), .B(n35363), .Z(n35362) );
  IV U37421 ( .A(n35361), .Z(n35363) );
  XOR U37422 ( .A(n35364), .B(mreg[510]), .Z(n35361) );
  NAND U37423 ( .A(n35365), .B(mul_pow), .Z(n35364) );
  XOR U37424 ( .A(mreg[510]), .B(creg[510]), .Z(n35365) );
  XOR U37425 ( .A(n35366), .B(n35367), .Z(n35357) );
  ANDN U37426 ( .A(n35368), .B(n27689), .Z(n35367) );
  XOR U37427 ( .A(n35369), .B(\modmult_1/zin[0][508] ), .Z(n27689) );
  IV U37428 ( .A(n35366), .Z(n35369) );
  XNOR U37429 ( .A(n35366), .B(n27688), .Z(n35368) );
  XOR U37430 ( .A(n35370), .B(n35371), .Z(n27688) );
  AND U37431 ( .A(\modmult_1/xin[1023] ), .B(n35372), .Z(n35371) );
  IV U37432 ( .A(n35370), .Z(n35372) );
  XOR U37433 ( .A(n35373), .B(mreg[509]), .Z(n35370) );
  NAND U37434 ( .A(n35374), .B(mul_pow), .Z(n35373) );
  XOR U37435 ( .A(mreg[509]), .B(creg[509]), .Z(n35374) );
  XOR U37436 ( .A(n35375), .B(n35376), .Z(n35366) );
  ANDN U37437 ( .A(n35377), .B(n27695), .Z(n35376) );
  XOR U37438 ( .A(n35378), .B(\modmult_1/zin[0][507] ), .Z(n27695) );
  IV U37439 ( .A(n35375), .Z(n35378) );
  XNOR U37440 ( .A(n35375), .B(n27694), .Z(n35377) );
  XOR U37441 ( .A(n35379), .B(n35380), .Z(n27694) );
  AND U37442 ( .A(\modmult_1/xin[1023] ), .B(n35381), .Z(n35380) );
  IV U37443 ( .A(n35379), .Z(n35381) );
  XOR U37444 ( .A(n35382), .B(mreg[508]), .Z(n35379) );
  NAND U37445 ( .A(n35383), .B(mul_pow), .Z(n35382) );
  XOR U37446 ( .A(mreg[508]), .B(creg[508]), .Z(n35383) );
  XOR U37447 ( .A(n35384), .B(n35385), .Z(n35375) );
  ANDN U37448 ( .A(n35386), .B(n27701), .Z(n35385) );
  XOR U37449 ( .A(n35387), .B(\modmult_1/zin[0][506] ), .Z(n27701) );
  IV U37450 ( .A(n35384), .Z(n35387) );
  XNOR U37451 ( .A(n35384), .B(n27700), .Z(n35386) );
  XOR U37452 ( .A(n35388), .B(n35389), .Z(n27700) );
  AND U37453 ( .A(\modmult_1/xin[1023] ), .B(n35390), .Z(n35389) );
  IV U37454 ( .A(n35388), .Z(n35390) );
  XOR U37455 ( .A(n35391), .B(mreg[507]), .Z(n35388) );
  NAND U37456 ( .A(n35392), .B(mul_pow), .Z(n35391) );
  XOR U37457 ( .A(mreg[507]), .B(creg[507]), .Z(n35392) );
  XOR U37458 ( .A(n35393), .B(n35394), .Z(n35384) );
  ANDN U37459 ( .A(n35395), .B(n27707), .Z(n35394) );
  XOR U37460 ( .A(n35396), .B(\modmult_1/zin[0][505] ), .Z(n27707) );
  IV U37461 ( .A(n35393), .Z(n35396) );
  XNOR U37462 ( .A(n35393), .B(n27706), .Z(n35395) );
  XOR U37463 ( .A(n35397), .B(n35398), .Z(n27706) );
  AND U37464 ( .A(\modmult_1/xin[1023] ), .B(n35399), .Z(n35398) );
  IV U37465 ( .A(n35397), .Z(n35399) );
  XOR U37466 ( .A(n35400), .B(mreg[506]), .Z(n35397) );
  NAND U37467 ( .A(n35401), .B(mul_pow), .Z(n35400) );
  XOR U37468 ( .A(mreg[506]), .B(creg[506]), .Z(n35401) );
  XOR U37469 ( .A(n35402), .B(n35403), .Z(n35393) );
  ANDN U37470 ( .A(n35404), .B(n27713), .Z(n35403) );
  XOR U37471 ( .A(n35405), .B(\modmult_1/zin[0][504] ), .Z(n27713) );
  IV U37472 ( .A(n35402), .Z(n35405) );
  XNOR U37473 ( .A(n35402), .B(n27712), .Z(n35404) );
  XOR U37474 ( .A(n35406), .B(n35407), .Z(n27712) );
  AND U37475 ( .A(\modmult_1/xin[1023] ), .B(n35408), .Z(n35407) );
  IV U37476 ( .A(n35406), .Z(n35408) );
  XOR U37477 ( .A(n35409), .B(mreg[505]), .Z(n35406) );
  NAND U37478 ( .A(n35410), .B(mul_pow), .Z(n35409) );
  XOR U37479 ( .A(mreg[505]), .B(creg[505]), .Z(n35410) );
  XOR U37480 ( .A(n35411), .B(n35412), .Z(n35402) );
  ANDN U37481 ( .A(n35413), .B(n27719), .Z(n35412) );
  XOR U37482 ( .A(n35414), .B(\modmult_1/zin[0][503] ), .Z(n27719) );
  IV U37483 ( .A(n35411), .Z(n35414) );
  XNOR U37484 ( .A(n35411), .B(n27718), .Z(n35413) );
  XOR U37485 ( .A(n35415), .B(n35416), .Z(n27718) );
  AND U37486 ( .A(\modmult_1/xin[1023] ), .B(n35417), .Z(n35416) );
  IV U37487 ( .A(n35415), .Z(n35417) );
  XOR U37488 ( .A(n35418), .B(mreg[504]), .Z(n35415) );
  NAND U37489 ( .A(n35419), .B(mul_pow), .Z(n35418) );
  XOR U37490 ( .A(mreg[504]), .B(creg[504]), .Z(n35419) );
  XOR U37491 ( .A(n35420), .B(n35421), .Z(n35411) );
  ANDN U37492 ( .A(n35422), .B(n27725), .Z(n35421) );
  XOR U37493 ( .A(n35423), .B(\modmult_1/zin[0][502] ), .Z(n27725) );
  IV U37494 ( .A(n35420), .Z(n35423) );
  XNOR U37495 ( .A(n35420), .B(n27724), .Z(n35422) );
  XOR U37496 ( .A(n35424), .B(n35425), .Z(n27724) );
  AND U37497 ( .A(\modmult_1/xin[1023] ), .B(n35426), .Z(n35425) );
  IV U37498 ( .A(n35424), .Z(n35426) );
  XOR U37499 ( .A(n35427), .B(mreg[503]), .Z(n35424) );
  NAND U37500 ( .A(n35428), .B(mul_pow), .Z(n35427) );
  XOR U37501 ( .A(mreg[503]), .B(creg[503]), .Z(n35428) );
  XOR U37502 ( .A(n35429), .B(n35430), .Z(n35420) );
  ANDN U37503 ( .A(n35431), .B(n27731), .Z(n35430) );
  XOR U37504 ( .A(n35432), .B(\modmult_1/zin[0][501] ), .Z(n27731) );
  IV U37505 ( .A(n35429), .Z(n35432) );
  XNOR U37506 ( .A(n35429), .B(n27730), .Z(n35431) );
  XOR U37507 ( .A(n35433), .B(n35434), .Z(n27730) );
  AND U37508 ( .A(\modmult_1/xin[1023] ), .B(n35435), .Z(n35434) );
  IV U37509 ( .A(n35433), .Z(n35435) );
  XOR U37510 ( .A(n35436), .B(mreg[502]), .Z(n35433) );
  NAND U37511 ( .A(n35437), .B(mul_pow), .Z(n35436) );
  XOR U37512 ( .A(mreg[502]), .B(creg[502]), .Z(n35437) );
  XOR U37513 ( .A(n35438), .B(n35439), .Z(n35429) );
  ANDN U37514 ( .A(n35440), .B(n27737), .Z(n35439) );
  XOR U37515 ( .A(n35441), .B(\modmult_1/zin[0][500] ), .Z(n27737) );
  IV U37516 ( .A(n35438), .Z(n35441) );
  XNOR U37517 ( .A(n35438), .B(n27736), .Z(n35440) );
  XOR U37518 ( .A(n35442), .B(n35443), .Z(n27736) );
  AND U37519 ( .A(\modmult_1/xin[1023] ), .B(n35444), .Z(n35443) );
  IV U37520 ( .A(n35442), .Z(n35444) );
  XOR U37521 ( .A(n35445), .B(mreg[501]), .Z(n35442) );
  NAND U37522 ( .A(n35446), .B(mul_pow), .Z(n35445) );
  XOR U37523 ( .A(mreg[501]), .B(creg[501]), .Z(n35446) );
  XOR U37524 ( .A(n35447), .B(n35448), .Z(n35438) );
  ANDN U37525 ( .A(n35449), .B(n27743), .Z(n35448) );
  XOR U37526 ( .A(n35450), .B(\modmult_1/zin[0][499] ), .Z(n27743) );
  IV U37527 ( .A(n35447), .Z(n35450) );
  XNOR U37528 ( .A(n35447), .B(n27742), .Z(n35449) );
  XOR U37529 ( .A(n35451), .B(n35452), .Z(n27742) );
  AND U37530 ( .A(\modmult_1/xin[1023] ), .B(n35453), .Z(n35452) );
  IV U37531 ( .A(n35451), .Z(n35453) );
  XOR U37532 ( .A(n35454), .B(mreg[500]), .Z(n35451) );
  NAND U37533 ( .A(n35455), .B(mul_pow), .Z(n35454) );
  XOR U37534 ( .A(mreg[500]), .B(creg[500]), .Z(n35455) );
  XOR U37535 ( .A(n35456), .B(n35457), .Z(n35447) );
  ANDN U37536 ( .A(n35458), .B(n27749), .Z(n35457) );
  XOR U37537 ( .A(n35459), .B(\modmult_1/zin[0][498] ), .Z(n27749) );
  IV U37538 ( .A(n35456), .Z(n35459) );
  XNOR U37539 ( .A(n35456), .B(n27748), .Z(n35458) );
  XOR U37540 ( .A(n35460), .B(n35461), .Z(n27748) );
  AND U37541 ( .A(\modmult_1/xin[1023] ), .B(n35462), .Z(n35461) );
  IV U37542 ( .A(n35460), .Z(n35462) );
  XOR U37543 ( .A(n35463), .B(mreg[499]), .Z(n35460) );
  NAND U37544 ( .A(n35464), .B(mul_pow), .Z(n35463) );
  XOR U37545 ( .A(mreg[499]), .B(creg[499]), .Z(n35464) );
  XOR U37546 ( .A(n35465), .B(n35466), .Z(n35456) );
  ANDN U37547 ( .A(n35467), .B(n27755), .Z(n35466) );
  XOR U37548 ( .A(n35468), .B(\modmult_1/zin[0][497] ), .Z(n27755) );
  IV U37549 ( .A(n35465), .Z(n35468) );
  XNOR U37550 ( .A(n35465), .B(n27754), .Z(n35467) );
  XOR U37551 ( .A(n35469), .B(n35470), .Z(n27754) );
  AND U37552 ( .A(\modmult_1/xin[1023] ), .B(n35471), .Z(n35470) );
  IV U37553 ( .A(n35469), .Z(n35471) );
  XOR U37554 ( .A(n35472), .B(mreg[498]), .Z(n35469) );
  NAND U37555 ( .A(n35473), .B(mul_pow), .Z(n35472) );
  XOR U37556 ( .A(mreg[498]), .B(creg[498]), .Z(n35473) );
  XOR U37557 ( .A(n35474), .B(n35475), .Z(n35465) );
  ANDN U37558 ( .A(n35476), .B(n27761), .Z(n35475) );
  XOR U37559 ( .A(n35477), .B(\modmult_1/zin[0][496] ), .Z(n27761) );
  IV U37560 ( .A(n35474), .Z(n35477) );
  XNOR U37561 ( .A(n35474), .B(n27760), .Z(n35476) );
  XOR U37562 ( .A(n35478), .B(n35479), .Z(n27760) );
  AND U37563 ( .A(\modmult_1/xin[1023] ), .B(n35480), .Z(n35479) );
  IV U37564 ( .A(n35478), .Z(n35480) );
  XOR U37565 ( .A(n35481), .B(mreg[497]), .Z(n35478) );
  NAND U37566 ( .A(n35482), .B(mul_pow), .Z(n35481) );
  XOR U37567 ( .A(mreg[497]), .B(creg[497]), .Z(n35482) );
  XOR U37568 ( .A(n35483), .B(n35484), .Z(n35474) );
  ANDN U37569 ( .A(n35485), .B(n27767), .Z(n35484) );
  XOR U37570 ( .A(n35486), .B(\modmult_1/zin[0][495] ), .Z(n27767) );
  IV U37571 ( .A(n35483), .Z(n35486) );
  XNOR U37572 ( .A(n35483), .B(n27766), .Z(n35485) );
  XOR U37573 ( .A(n35487), .B(n35488), .Z(n27766) );
  AND U37574 ( .A(\modmult_1/xin[1023] ), .B(n35489), .Z(n35488) );
  IV U37575 ( .A(n35487), .Z(n35489) );
  XOR U37576 ( .A(n35490), .B(mreg[496]), .Z(n35487) );
  NAND U37577 ( .A(n35491), .B(mul_pow), .Z(n35490) );
  XOR U37578 ( .A(mreg[496]), .B(creg[496]), .Z(n35491) );
  XOR U37579 ( .A(n35492), .B(n35493), .Z(n35483) );
  ANDN U37580 ( .A(n35494), .B(n27773), .Z(n35493) );
  XOR U37581 ( .A(n35495), .B(\modmult_1/zin[0][494] ), .Z(n27773) );
  IV U37582 ( .A(n35492), .Z(n35495) );
  XNOR U37583 ( .A(n35492), .B(n27772), .Z(n35494) );
  XOR U37584 ( .A(n35496), .B(n35497), .Z(n27772) );
  AND U37585 ( .A(\modmult_1/xin[1023] ), .B(n35498), .Z(n35497) );
  IV U37586 ( .A(n35496), .Z(n35498) );
  XOR U37587 ( .A(n35499), .B(mreg[495]), .Z(n35496) );
  NAND U37588 ( .A(n35500), .B(mul_pow), .Z(n35499) );
  XOR U37589 ( .A(mreg[495]), .B(creg[495]), .Z(n35500) );
  XOR U37590 ( .A(n35501), .B(n35502), .Z(n35492) );
  ANDN U37591 ( .A(n35503), .B(n27779), .Z(n35502) );
  XOR U37592 ( .A(n35504), .B(\modmult_1/zin[0][493] ), .Z(n27779) );
  IV U37593 ( .A(n35501), .Z(n35504) );
  XNOR U37594 ( .A(n35501), .B(n27778), .Z(n35503) );
  XOR U37595 ( .A(n35505), .B(n35506), .Z(n27778) );
  AND U37596 ( .A(\modmult_1/xin[1023] ), .B(n35507), .Z(n35506) );
  IV U37597 ( .A(n35505), .Z(n35507) );
  XOR U37598 ( .A(n35508), .B(mreg[494]), .Z(n35505) );
  NAND U37599 ( .A(n35509), .B(mul_pow), .Z(n35508) );
  XOR U37600 ( .A(mreg[494]), .B(creg[494]), .Z(n35509) );
  XOR U37601 ( .A(n35510), .B(n35511), .Z(n35501) );
  ANDN U37602 ( .A(n35512), .B(n27785), .Z(n35511) );
  XOR U37603 ( .A(n35513), .B(\modmult_1/zin[0][492] ), .Z(n27785) );
  IV U37604 ( .A(n35510), .Z(n35513) );
  XNOR U37605 ( .A(n35510), .B(n27784), .Z(n35512) );
  XOR U37606 ( .A(n35514), .B(n35515), .Z(n27784) );
  AND U37607 ( .A(\modmult_1/xin[1023] ), .B(n35516), .Z(n35515) );
  IV U37608 ( .A(n35514), .Z(n35516) );
  XOR U37609 ( .A(n35517), .B(mreg[493]), .Z(n35514) );
  NAND U37610 ( .A(n35518), .B(mul_pow), .Z(n35517) );
  XOR U37611 ( .A(mreg[493]), .B(creg[493]), .Z(n35518) );
  XOR U37612 ( .A(n35519), .B(n35520), .Z(n35510) );
  ANDN U37613 ( .A(n35521), .B(n27791), .Z(n35520) );
  XOR U37614 ( .A(n35522), .B(\modmult_1/zin[0][491] ), .Z(n27791) );
  IV U37615 ( .A(n35519), .Z(n35522) );
  XNOR U37616 ( .A(n35519), .B(n27790), .Z(n35521) );
  XOR U37617 ( .A(n35523), .B(n35524), .Z(n27790) );
  AND U37618 ( .A(\modmult_1/xin[1023] ), .B(n35525), .Z(n35524) );
  IV U37619 ( .A(n35523), .Z(n35525) );
  XOR U37620 ( .A(n35526), .B(mreg[492]), .Z(n35523) );
  NAND U37621 ( .A(n35527), .B(mul_pow), .Z(n35526) );
  XOR U37622 ( .A(mreg[492]), .B(creg[492]), .Z(n35527) );
  XOR U37623 ( .A(n35528), .B(n35529), .Z(n35519) );
  ANDN U37624 ( .A(n35530), .B(n27797), .Z(n35529) );
  XOR U37625 ( .A(n35531), .B(\modmult_1/zin[0][490] ), .Z(n27797) );
  IV U37626 ( .A(n35528), .Z(n35531) );
  XNOR U37627 ( .A(n35528), .B(n27796), .Z(n35530) );
  XOR U37628 ( .A(n35532), .B(n35533), .Z(n27796) );
  AND U37629 ( .A(\modmult_1/xin[1023] ), .B(n35534), .Z(n35533) );
  IV U37630 ( .A(n35532), .Z(n35534) );
  XOR U37631 ( .A(n35535), .B(mreg[491]), .Z(n35532) );
  NAND U37632 ( .A(n35536), .B(mul_pow), .Z(n35535) );
  XOR U37633 ( .A(mreg[491]), .B(creg[491]), .Z(n35536) );
  XOR U37634 ( .A(n35537), .B(n35538), .Z(n35528) );
  ANDN U37635 ( .A(n35539), .B(n27803), .Z(n35538) );
  XOR U37636 ( .A(n35540), .B(\modmult_1/zin[0][489] ), .Z(n27803) );
  IV U37637 ( .A(n35537), .Z(n35540) );
  XNOR U37638 ( .A(n35537), .B(n27802), .Z(n35539) );
  XOR U37639 ( .A(n35541), .B(n35542), .Z(n27802) );
  AND U37640 ( .A(\modmult_1/xin[1023] ), .B(n35543), .Z(n35542) );
  IV U37641 ( .A(n35541), .Z(n35543) );
  XOR U37642 ( .A(n35544), .B(mreg[490]), .Z(n35541) );
  NAND U37643 ( .A(n35545), .B(mul_pow), .Z(n35544) );
  XOR U37644 ( .A(mreg[490]), .B(creg[490]), .Z(n35545) );
  XOR U37645 ( .A(n35546), .B(n35547), .Z(n35537) );
  ANDN U37646 ( .A(n35548), .B(n27809), .Z(n35547) );
  XOR U37647 ( .A(n35549), .B(\modmult_1/zin[0][488] ), .Z(n27809) );
  IV U37648 ( .A(n35546), .Z(n35549) );
  XNOR U37649 ( .A(n35546), .B(n27808), .Z(n35548) );
  XOR U37650 ( .A(n35550), .B(n35551), .Z(n27808) );
  AND U37651 ( .A(\modmult_1/xin[1023] ), .B(n35552), .Z(n35551) );
  IV U37652 ( .A(n35550), .Z(n35552) );
  XOR U37653 ( .A(n35553), .B(mreg[489]), .Z(n35550) );
  NAND U37654 ( .A(n35554), .B(mul_pow), .Z(n35553) );
  XOR U37655 ( .A(mreg[489]), .B(creg[489]), .Z(n35554) );
  XOR U37656 ( .A(n35555), .B(n35556), .Z(n35546) );
  ANDN U37657 ( .A(n35557), .B(n27815), .Z(n35556) );
  XOR U37658 ( .A(n35558), .B(\modmult_1/zin[0][487] ), .Z(n27815) );
  IV U37659 ( .A(n35555), .Z(n35558) );
  XNOR U37660 ( .A(n35555), .B(n27814), .Z(n35557) );
  XOR U37661 ( .A(n35559), .B(n35560), .Z(n27814) );
  AND U37662 ( .A(\modmult_1/xin[1023] ), .B(n35561), .Z(n35560) );
  IV U37663 ( .A(n35559), .Z(n35561) );
  XOR U37664 ( .A(n35562), .B(mreg[488]), .Z(n35559) );
  NAND U37665 ( .A(n35563), .B(mul_pow), .Z(n35562) );
  XOR U37666 ( .A(mreg[488]), .B(creg[488]), .Z(n35563) );
  XOR U37667 ( .A(n35564), .B(n35565), .Z(n35555) );
  ANDN U37668 ( .A(n35566), .B(n27821), .Z(n35565) );
  XOR U37669 ( .A(n35567), .B(\modmult_1/zin[0][486] ), .Z(n27821) );
  IV U37670 ( .A(n35564), .Z(n35567) );
  XNOR U37671 ( .A(n35564), .B(n27820), .Z(n35566) );
  XOR U37672 ( .A(n35568), .B(n35569), .Z(n27820) );
  AND U37673 ( .A(\modmult_1/xin[1023] ), .B(n35570), .Z(n35569) );
  IV U37674 ( .A(n35568), .Z(n35570) );
  XOR U37675 ( .A(n35571), .B(mreg[487]), .Z(n35568) );
  NAND U37676 ( .A(n35572), .B(mul_pow), .Z(n35571) );
  XOR U37677 ( .A(mreg[487]), .B(creg[487]), .Z(n35572) );
  XOR U37678 ( .A(n35573), .B(n35574), .Z(n35564) );
  ANDN U37679 ( .A(n35575), .B(n27827), .Z(n35574) );
  XOR U37680 ( .A(n35576), .B(\modmult_1/zin[0][485] ), .Z(n27827) );
  IV U37681 ( .A(n35573), .Z(n35576) );
  XNOR U37682 ( .A(n35573), .B(n27826), .Z(n35575) );
  XOR U37683 ( .A(n35577), .B(n35578), .Z(n27826) );
  AND U37684 ( .A(\modmult_1/xin[1023] ), .B(n35579), .Z(n35578) );
  IV U37685 ( .A(n35577), .Z(n35579) );
  XOR U37686 ( .A(n35580), .B(mreg[486]), .Z(n35577) );
  NAND U37687 ( .A(n35581), .B(mul_pow), .Z(n35580) );
  XOR U37688 ( .A(mreg[486]), .B(creg[486]), .Z(n35581) );
  XOR U37689 ( .A(n35582), .B(n35583), .Z(n35573) );
  ANDN U37690 ( .A(n35584), .B(n27833), .Z(n35583) );
  XOR U37691 ( .A(n35585), .B(\modmult_1/zin[0][484] ), .Z(n27833) );
  IV U37692 ( .A(n35582), .Z(n35585) );
  XNOR U37693 ( .A(n35582), .B(n27832), .Z(n35584) );
  XOR U37694 ( .A(n35586), .B(n35587), .Z(n27832) );
  AND U37695 ( .A(\modmult_1/xin[1023] ), .B(n35588), .Z(n35587) );
  IV U37696 ( .A(n35586), .Z(n35588) );
  XOR U37697 ( .A(n35589), .B(mreg[485]), .Z(n35586) );
  NAND U37698 ( .A(n35590), .B(mul_pow), .Z(n35589) );
  XOR U37699 ( .A(mreg[485]), .B(creg[485]), .Z(n35590) );
  XOR U37700 ( .A(n35591), .B(n35592), .Z(n35582) );
  ANDN U37701 ( .A(n35593), .B(n27839), .Z(n35592) );
  XOR U37702 ( .A(n35594), .B(\modmult_1/zin[0][483] ), .Z(n27839) );
  IV U37703 ( .A(n35591), .Z(n35594) );
  XNOR U37704 ( .A(n35591), .B(n27838), .Z(n35593) );
  XOR U37705 ( .A(n35595), .B(n35596), .Z(n27838) );
  AND U37706 ( .A(\modmult_1/xin[1023] ), .B(n35597), .Z(n35596) );
  IV U37707 ( .A(n35595), .Z(n35597) );
  XOR U37708 ( .A(n35598), .B(mreg[484]), .Z(n35595) );
  NAND U37709 ( .A(n35599), .B(mul_pow), .Z(n35598) );
  XOR U37710 ( .A(mreg[484]), .B(creg[484]), .Z(n35599) );
  XOR U37711 ( .A(n35600), .B(n35601), .Z(n35591) );
  ANDN U37712 ( .A(n35602), .B(n27845), .Z(n35601) );
  XOR U37713 ( .A(n35603), .B(\modmult_1/zin[0][482] ), .Z(n27845) );
  IV U37714 ( .A(n35600), .Z(n35603) );
  XNOR U37715 ( .A(n35600), .B(n27844), .Z(n35602) );
  XOR U37716 ( .A(n35604), .B(n35605), .Z(n27844) );
  AND U37717 ( .A(\modmult_1/xin[1023] ), .B(n35606), .Z(n35605) );
  IV U37718 ( .A(n35604), .Z(n35606) );
  XOR U37719 ( .A(n35607), .B(mreg[483]), .Z(n35604) );
  NAND U37720 ( .A(n35608), .B(mul_pow), .Z(n35607) );
  XOR U37721 ( .A(mreg[483]), .B(creg[483]), .Z(n35608) );
  XOR U37722 ( .A(n35609), .B(n35610), .Z(n35600) );
  ANDN U37723 ( .A(n35611), .B(n27851), .Z(n35610) );
  XOR U37724 ( .A(n35612), .B(\modmult_1/zin[0][481] ), .Z(n27851) );
  IV U37725 ( .A(n35609), .Z(n35612) );
  XNOR U37726 ( .A(n35609), .B(n27850), .Z(n35611) );
  XOR U37727 ( .A(n35613), .B(n35614), .Z(n27850) );
  AND U37728 ( .A(\modmult_1/xin[1023] ), .B(n35615), .Z(n35614) );
  IV U37729 ( .A(n35613), .Z(n35615) );
  XOR U37730 ( .A(n35616), .B(mreg[482]), .Z(n35613) );
  NAND U37731 ( .A(n35617), .B(mul_pow), .Z(n35616) );
  XOR U37732 ( .A(mreg[482]), .B(creg[482]), .Z(n35617) );
  XOR U37733 ( .A(n35618), .B(n35619), .Z(n35609) );
  ANDN U37734 ( .A(n35620), .B(n27857), .Z(n35619) );
  XOR U37735 ( .A(n35621), .B(\modmult_1/zin[0][480] ), .Z(n27857) );
  IV U37736 ( .A(n35618), .Z(n35621) );
  XNOR U37737 ( .A(n35618), .B(n27856), .Z(n35620) );
  XOR U37738 ( .A(n35622), .B(n35623), .Z(n27856) );
  AND U37739 ( .A(\modmult_1/xin[1023] ), .B(n35624), .Z(n35623) );
  IV U37740 ( .A(n35622), .Z(n35624) );
  XOR U37741 ( .A(n35625), .B(mreg[481]), .Z(n35622) );
  NAND U37742 ( .A(n35626), .B(mul_pow), .Z(n35625) );
  XOR U37743 ( .A(mreg[481]), .B(creg[481]), .Z(n35626) );
  XOR U37744 ( .A(n35627), .B(n35628), .Z(n35618) );
  ANDN U37745 ( .A(n35629), .B(n27863), .Z(n35628) );
  XOR U37746 ( .A(n35630), .B(\modmult_1/zin[0][479] ), .Z(n27863) );
  IV U37747 ( .A(n35627), .Z(n35630) );
  XNOR U37748 ( .A(n35627), .B(n27862), .Z(n35629) );
  XOR U37749 ( .A(n35631), .B(n35632), .Z(n27862) );
  AND U37750 ( .A(\modmult_1/xin[1023] ), .B(n35633), .Z(n35632) );
  IV U37751 ( .A(n35631), .Z(n35633) );
  XOR U37752 ( .A(n35634), .B(mreg[480]), .Z(n35631) );
  NAND U37753 ( .A(n35635), .B(mul_pow), .Z(n35634) );
  XOR U37754 ( .A(mreg[480]), .B(creg[480]), .Z(n35635) );
  XOR U37755 ( .A(n35636), .B(n35637), .Z(n35627) );
  ANDN U37756 ( .A(n35638), .B(n27869), .Z(n35637) );
  XOR U37757 ( .A(n35639), .B(\modmult_1/zin[0][478] ), .Z(n27869) );
  IV U37758 ( .A(n35636), .Z(n35639) );
  XNOR U37759 ( .A(n35636), .B(n27868), .Z(n35638) );
  XOR U37760 ( .A(n35640), .B(n35641), .Z(n27868) );
  AND U37761 ( .A(\modmult_1/xin[1023] ), .B(n35642), .Z(n35641) );
  IV U37762 ( .A(n35640), .Z(n35642) );
  XOR U37763 ( .A(n35643), .B(mreg[479]), .Z(n35640) );
  NAND U37764 ( .A(n35644), .B(mul_pow), .Z(n35643) );
  XOR U37765 ( .A(mreg[479]), .B(creg[479]), .Z(n35644) );
  XOR U37766 ( .A(n35645), .B(n35646), .Z(n35636) );
  ANDN U37767 ( .A(n35647), .B(n27875), .Z(n35646) );
  XOR U37768 ( .A(n35648), .B(\modmult_1/zin[0][477] ), .Z(n27875) );
  IV U37769 ( .A(n35645), .Z(n35648) );
  XNOR U37770 ( .A(n35645), .B(n27874), .Z(n35647) );
  XOR U37771 ( .A(n35649), .B(n35650), .Z(n27874) );
  AND U37772 ( .A(\modmult_1/xin[1023] ), .B(n35651), .Z(n35650) );
  IV U37773 ( .A(n35649), .Z(n35651) );
  XOR U37774 ( .A(n35652), .B(mreg[478]), .Z(n35649) );
  NAND U37775 ( .A(n35653), .B(mul_pow), .Z(n35652) );
  XOR U37776 ( .A(mreg[478]), .B(creg[478]), .Z(n35653) );
  XOR U37777 ( .A(n35654), .B(n35655), .Z(n35645) );
  ANDN U37778 ( .A(n35656), .B(n27881), .Z(n35655) );
  XOR U37779 ( .A(n35657), .B(\modmult_1/zin[0][476] ), .Z(n27881) );
  IV U37780 ( .A(n35654), .Z(n35657) );
  XNOR U37781 ( .A(n35654), .B(n27880), .Z(n35656) );
  XOR U37782 ( .A(n35658), .B(n35659), .Z(n27880) );
  AND U37783 ( .A(\modmult_1/xin[1023] ), .B(n35660), .Z(n35659) );
  IV U37784 ( .A(n35658), .Z(n35660) );
  XOR U37785 ( .A(n35661), .B(mreg[477]), .Z(n35658) );
  NAND U37786 ( .A(n35662), .B(mul_pow), .Z(n35661) );
  XOR U37787 ( .A(mreg[477]), .B(creg[477]), .Z(n35662) );
  XOR U37788 ( .A(n35663), .B(n35664), .Z(n35654) );
  ANDN U37789 ( .A(n35665), .B(n27887), .Z(n35664) );
  XOR U37790 ( .A(n35666), .B(\modmult_1/zin[0][475] ), .Z(n27887) );
  IV U37791 ( .A(n35663), .Z(n35666) );
  XNOR U37792 ( .A(n35663), .B(n27886), .Z(n35665) );
  XOR U37793 ( .A(n35667), .B(n35668), .Z(n27886) );
  AND U37794 ( .A(\modmult_1/xin[1023] ), .B(n35669), .Z(n35668) );
  IV U37795 ( .A(n35667), .Z(n35669) );
  XOR U37796 ( .A(n35670), .B(mreg[476]), .Z(n35667) );
  NAND U37797 ( .A(n35671), .B(mul_pow), .Z(n35670) );
  XOR U37798 ( .A(mreg[476]), .B(creg[476]), .Z(n35671) );
  XOR U37799 ( .A(n35672), .B(n35673), .Z(n35663) );
  ANDN U37800 ( .A(n35674), .B(n27893), .Z(n35673) );
  XOR U37801 ( .A(n35675), .B(\modmult_1/zin[0][474] ), .Z(n27893) );
  IV U37802 ( .A(n35672), .Z(n35675) );
  XNOR U37803 ( .A(n35672), .B(n27892), .Z(n35674) );
  XOR U37804 ( .A(n35676), .B(n35677), .Z(n27892) );
  AND U37805 ( .A(\modmult_1/xin[1023] ), .B(n35678), .Z(n35677) );
  IV U37806 ( .A(n35676), .Z(n35678) );
  XOR U37807 ( .A(n35679), .B(mreg[475]), .Z(n35676) );
  NAND U37808 ( .A(n35680), .B(mul_pow), .Z(n35679) );
  XOR U37809 ( .A(mreg[475]), .B(creg[475]), .Z(n35680) );
  XOR U37810 ( .A(n35681), .B(n35682), .Z(n35672) );
  ANDN U37811 ( .A(n35683), .B(n27899), .Z(n35682) );
  XOR U37812 ( .A(n35684), .B(\modmult_1/zin[0][473] ), .Z(n27899) );
  IV U37813 ( .A(n35681), .Z(n35684) );
  XNOR U37814 ( .A(n35681), .B(n27898), .Z(n35683) );
  XOR U37815 ( .A(n35685), .B(n35686), .Z(n27898) );
  AND U37816 ( .A(\modmult_1/xin[1023] ), .B(n35687), .Z(n35686) );
  IV U37817 ( .A(n35685), .Z(n35687) );
  XOR U37818 ( .A(n35688), .B(mreg[474]), .Z(n35685) );
  NAND U37819 ( .A(n35689), .B(mul_pow), .Z(n35688) );
  XOR U37820 ( .A(mreg[474]), .B(creg[474]), .Z(n35689) );
  XOR U37821 ( .A(n35690), .B(n35691), .Z(n35681) );
  ANDN U37822 ( .A(n35692), .B(n27905), .Z(n35691) );
  XOR U37823 ( .A(n35693), .B(\modmult_1/zin[0][472] ), .Z(n27905) );
  IV U37824 ( .A(n35690), .Z(n35693) );
  XNOR U37825 ( .A(n35690), .B(n27904), .Z(n35692) );
  XOR U37826 ( .A(n35694), .B(n35695), .Z(n27904) );
  AND U37827 ( .A(\modmult_1/xin[1023] ), .B(n35696), .Z(n35695) );
  IV U37828 ( .A(n35694), .Z(n35696) );
  XOR U37829 ( .A(n35697), .B(mreg[473]), .Z(n35694) );
  NAND U37830 ( .A(n35698), .B(mul_pow), .Z(n35697) );
  XOR U37831 ( .A(mreg[473]), .B(creg[473]), .Z(n35698) );
  XOR U37832 ( .A(n35699), .B(n35700), .Z(n35690) );
  ANDN U37833 ( .A(n35701), .B(n27911), .Z(n35700) );
  XOR U37834 ( .A(n35702), .B(\modmult_1/zin[0][471] ), .Z(n27911) );
  IV U37835 ( .A(n35699), .Z(n35702) );
  XNOR U37836 ( .A(n35699), .B(n27910), .Z(n35701) );
  XOR U37837 ( .A(n35703), .B(n35704), .Z(n27910) );
  AND U37838 ( .A(\modmult_1/xin[1023] ), .B(n35705), .Z(n35704) );
  IV U37839 ( .A(n35703), .Z(n35705) );
  XOR U37840 ( .A(n35706), .B(mreg[472]), .Z(n35703) );
  NAND U37841 ( .A(n35707), .B(mul_pow), .Z(n35706) );
  XOR U37842 ( .A(mreg[472]), .B(creg[472]), .Z(n35707) );
  XOR U37843 ( .A(n35708), .B(n35709), .Z(n35699) );
  ANDN U37844 ( .A(n35710), .B(n27917), .Z(n35709) );
  XOR U37845 ( .A(n35711), .B(\modmult_1/zin[0][470] ), .Z(n27917) );
  IV U37846 ( .A(n35708), .Z(n35711) );
  XNOR U37847 ( .A(n35708), .B(n27916), .Z(n35710) );
  XOR U37848 ( .A(n35712), .B(n35713), .Z(n27916) );
  AND U37849 ( .A(\modmult_1/xin[1023] ), .B(n35714), .Z(n35713) );
  IV U37850 ( .A(n35712), .Z(n35714) );
  XOR U37851 ( .A(n35715), .B(mreg[471]), .Z(n35712) );
  NAND U37852 ( .A(n35716), .B(mul_pow), .Z(n35715) );
  XOR U37853 ( .A(mreg[471]), .B(creg[471]), .Z(n35716) );
  XOR U37854 ( .A(n35717), .B(n35718), .Z(n35708) );
  ANDN U37855 ( .A(n35719), .B(n27923), .Z(n35718) );
  XOR U37856 ( .A(n35720), .B(\modmult_1/zin[0][469] ), .Z(n27923) );
  IV U37857 ( .A(n35717), .Z(n35720) );
  XNOR U37858 ( .A(n35717), .B(n27922), .Z(n35719) );
  XOR U37859 ( .A(n35721), .B(n35722), .Z(n27922) );
  AND U37860 ( .A(\modmult_1/xin[1023] ), .B(n35723), .Z(n35722) );
  IV U37861 ( .A(n35721), .Z(n35723) );
  XOR U37862 ( .A(n35724), .B(mreg[470]), .Z(n35721) );
  NAND U37863 ( .A(n35725), .B(mul_pow), .Z(n35724) );
  XOR U37864 ( .A(mreg[470]), .B(creg[470]), .Z(n35725) );
  XOR U37865 ( .A(n35726), .B(n35727), .Z(n35717) );
  ANDN U37866 ( .A(n35728), .B(n27929), .Z(n35727) );
  XOR U37867 ( .A(n35729), .B(\modmult_1/zin[0][468] ), .Z(n27929) );
  IV U37868 ( .A(n35726), .Z(n35729) );
  XNOR U37869 ( .A(n35726), .B(n27928), .Z(n35728) );
  XOR U37870 ( .A(n35730), .B(n35731), .Z(n27928) );
  AND U37871 ( .A(\modmult_1/xin[1023] ), .B(n35732), .Z(n35731) );
  IV U37872 ( .A(n35730), .Z(n35732) );
  XOR U37873 ( .A(n35733), .B(mreg[469]), .Z(n35730) );
  NAND U37874 ( .A(n35734), .B(mul_pow), .Z(n35733) );
  XOR U37875 ( .A(mreg[469]), .B(creg[469]), .Z(n35734) );
  XOR U37876 ( .A(n35735), .B(n35736), .Z(n35726) );
  ANDN U37877 ( .A(n35737), .B(n27935), .Z(n35736) );
  XOR U37878 ( .A(n35738), .B(\modmult_1/zin[0][467] ), .Z(n27935) );
  IV U37879 ( .A(n35735), .Z(n35738) );
  XNOR U37880 ( .A(n35735), .B(n27934), .Z(n35737) );
  XOR U37881 ( .A(n35739), .B(n35740), .Z(n27934) );
  AND U37882 ( .A(\modmult_1/xin[1023] ), .B(n35741), .Z(n35740) );
  IV U37883 ( .A(n35739), .Z(n35741) );
  XOR U37884 ( .A(n35742), .B(mreg[468]), .Z(n35739) );
  NAND U37885 ( .A(n35743), .B(mul_pow), .Z(n35742) );
  XOR U37886 ( .A(mreg[468]), .B(creg[468]), .Z(n35743) );
  XOR U37887 ( .A(n35744), .B(n35745), .Z(n35735) );
  ANDN U37888 ( .A(n35746), .B(n27941), .Z(n35745) );
  XOR U37889 ( .A(n35747), .B(\modmult_1/zin[0][466] ), .Z(n27941) );
  IV U37890 ( .A(n35744), .Z(n35747) );
  XNOR U37891 ( .A(n35744), .B(n27940), .Z(n35746) );
  XOR U37892 ( .A(n35748), .B(n35749), .Z(n27940) );
  AND U37893 ( .A(\modmult_1/xin[1023] ), .B(n35750), .Z(n35749) );
  IV U37894 ( .A(n35748), .Z(n35750) );
  XOR U37895 ( .A(n35751), .B(mreg[467]), .Z(n35748) );
  NAND U37896 ( .A(n35752), .B(mul_pow), .Z(n35751) );
  XOR U37897 ( .A(mreg[467]), .B(creg[467]), .Z(n35752) );
  XOR U37898 ( .A(n35753), .B(n35754), .Z(n35744) );
  ANDN U37899 ( .A(n35755), .B(n27947), .Z(n35754) );
  XOR U37900 ( .A(n35756), .B(\modmult_1/zin[0][465] ), .Z(n27947) );
  IV U37901 ( .A(n35753), .Z(n35756) );
  XNOR U37902 ( .A(n35753), .B(n27946), .Z(n35755) );
  XOR U37903 ( .A(n35757), .B(n35758), .Z(n27946) );
  AND U37904 ( .A(\modmult_1/xin[1023] ), .B(n35759), .Z(n35758) );
  IV U37905 ( .A(n35757), .Z(n35759) );
  XOR U37906 ( .A(n35760), .B(mreg[466]), .Z(n35757) );
  NAND U37907 ( .A(n35761), .B(mul_pow), .Z(n35760) );
  XOR U37908 ( .A(mreg[466]), .B(creg[466]), .Z(n35761) );
  XOR U37909 ( .A(n35762), .B(n35763), .Z(n35753) );
  ANDN U37910 ( .A(n35764), .B(n27953), .Z(n35763) );
  XOR U37911 ( .A(n35765), .B(\modmult_1/zin[0][464] ), .Z(n27953) );
  IV U37912 ( .A(n35762), .Z(n35765) );
  XNOR U37913 ( .A(n35762), .B(n27952), .Z(n35764) );
  XOR U37914 ( .A(n35766), .B(n35767), .Z(n27952) );
  AND U37915 ( .A(\modmult_1/xin[1023] ), .B(n35768), .Z(n35767) );
  IV U37916 ( .A(n35766), .Z(n35768) );
  XOR U37917 ( .A(n35769), .B(mreg[465]), .Z(n35766) );
  NAND U37918 ( .A(n35770), .B(mul_pow), .Z(n35769) );
  XOR U37919 ( .A(mreg[465]), .B(creg[465]), .Z(n35770) );
  XOR U37920 ( .A(n35771), .B(n35772), .Z(n35762) );
  ANDN U37921 ( .A(n35773), .B(n27959), .Z(n35772) );
  XOR U37922 ( .A(n35774), .B(\modmult_1/zin[0][463] ), .Z(n27959) );
  IV U37923 ( .A(n35771), .Z(n35774) );
  XNOR U37924 ( .A(n35771), .B(n27958), .Z(n35773) );
  XOR U37925 ( .A(n35775), .B(n35776), .Z(n27958) );
  AND U37926 ( .A(\modmult_1/xin[1023] ), .B(n35777), .Z(n35776) );
  IV U37927 ( .A(n35775), .Z(n35777) );
  XOR U37928 ( .A(n35778), .B(mreg[464]), .Z(n35775) );
  NAND U37929 ( .A(n35779), .B(mul_pow), .Z(n35778) );
  XOR U37930 ( .A(mreg[464]), .B(creg[464]), .Z(n35779) );
  XOR U37931 ( .A(n35780), .B(n35781), .Z(n35771) );
  ANDN U37932 ( .A(n35782), .B(n27965), .Z(n35781) );
  XOR U37933 ( .A(n35783), .B(\modmult_1/zin[0][462] ), .Z(n27965) );
  IV U37934 ( .A(n35780), .Z(n35783) );
  XNOR U37935 ( .A(n35780), .B(n27964), .Z(n35782) );
  XOR U37936 ( .A(n35784), .B(n35785), .Z(n27964) );
  AND U37937 ( .A(\modmult_1/xin[1023] ), .B(n35786), .Z(n35785) );
  IV U37938 ( .A(n35784), .Z(n35786) );
  XOR U37939 ( .A(n35787), .B(mreg[463]), .Z(n35784) );
  NAND U37940 ( .A(n35788), .B(mul_pow), .Z(n35787) );
  XOR U37941 ( .A(mreg[463]), .B(creg[463]), .Z(n35788) );
  XOR U37942 ( .A(n35789), .B(n35790), .Z(n35780) );
  ANDN U37943 ( .A(n35791), .B(n27971), .Z(n35790) );
  XOR U37944 ( .A(n35792), .B(\modmult_1/zin[0][461] ), .Z(n27971) );
  IV U37945 ( .A(n35789), .Z(n35792) );
  XNOR U37946 ( .A(n35789), .B(n27970), .Z(n35791) );
  XOR U37947 ( .A(n35793), .B(n35794), .Z(n27970) );
  AND U37948 ( .A(\modmult_1/xin[1023] ), .B(n35795), .Z(n35794) );
  IV U37949 ( .A(n35793), .Z(n35795) );
  XOR U37950 ( .A(n35796), .B(mreg[462]), .Z(n35793) );
  NAND U37951 ( .A(n35797), .B(mul_pow), .Z(n35796) );
  XOR U37952 ( .A(mreg[462]), .B(creg[462]), .Z(n35797) );
  XOR U37953 ( .A(n35798), .B(n35799), .Z(n35789) );
  ANDN U37954 ( .A(n35800), .B(n27977), .Z(n35799) );
  XOR U37955 ( .A(n35801), .B(\modmult_1/zin[0][460] ), .Z(n27977) );
  IV U37956 ( .A(n35798), .Z(n35801) );
  XNOR U37957 ( .A(n35798), .B(n27976), .Z(n35800) );
  XOR U37958 ( .A(n35802), .B(n35803), .Z(n27976) );
  AND U37959 ( .A(\modmult_1/xin[1023] ), .B(n35804), .Z(n35803) );
  IV U37960 ( .A(n35802), .Z(n35804) );
  XOR U37961 ( .A(n35805), .B(mreg[461]), .Z(n35802) );
  NAND U37962 ( .A(n35806), .B(mul_pow), .Z(n35805) );
  XOR U37963 ( .A(mreg[461]), .B(creg[461]), .Z(n35806) );
  XOR U37964 ( .A(n35807), .B(n35808), .Z(n35798) );
  ANDN U37965 ( .A(n35809), .B(n27983), .Z(n35808) );
  XOR U37966 ( .A(n35810), .B(\modmult_1/zin[0][459] ), .Z(n27983) );
  IV U37967 ( .A(n35807), .Z(n35810) );
  XNOR U37968 ( .A(n35807), .B(n27982), .Z(n35809) );
  XOR U37969 ( .A(n35811), .B(n35812), .Z(n27982) );
  AND U37970 ( .A(\modmult_1/xin[1023] ), .B(n35813), .Z(n35812) );
  IV U37971 ( .A(n35811), .Z(n35813) );
  XOR U37972 ( .A(n35814), .B(mreg[460]), .Z(n35811) );
  NAND U37973 ( .A(n35815), .B(mul_pow), .Z(n35814) );
  XOR U37974 ( .A(mreg[460]), .B(creg[460]), .Z(n35815) );
  XOR U37975 ( .A(n35816), .B(n35817), .Z(n35807) );
  ANDN U37976 ( .A(n35818), .B(n27989), .Z(n35817) );
  XOR U37977 ( .A(n35819), .B(\modmult_1/zin[0][458] ), .Z(n27989) );
  IV U37978 ( .A(n35816), .Z(n35819) );
  XNOR U37979 ( .A(n35816), .B(n27988), .Z(n35818) );
  XOR U37980 ( .A(n35820), .B(n35821), .Z(n27988) );
  AND U37981 ( .A(\modmult_1/xin[1023] ), .B(n35822), .Z(n35821) );
  IV U37982 ( .A(n35820), .Z(n35822) );
  XOR U37983 ( .A(n35823), .B(mreg[459]), .Z(n35820) );
  NAND U37984 ( .A(n35824), .B(mul_pow), .Z(n35823) );
  XOR U37985 ( .A(mreg[459]), .B(creg[459]), .Z(n35824) );
  XOR U37986 ( .A(n35825), .B(n35826), .Z(n35816) );
  ANDN U37987 ( .A(n35827), .B(n27995), .Z(n35826) );
  XOR U37988 ( .A(n35828), .B(\modmult_1/zin[0][457] ), .Z(n27995) );
  IV U37989 ( .A(n35825), .Z(n35828) );
  XNOR U37990 ( .A(n35825), .B(n27994), .Z(n35827) );
  XOR U37991 ( .A(n35829), .B(n35830), .Z(n27994) );
  AND U37992 ( .A(\modmult_1/xin[1023] ), .B(n35831), .Z(n35830) );
  IV U37993 ( .A(n35829), .Z(n35831) );
  XOR U37994 ( .A(n35832), .B(mreg[458]), .Z(n35829) );
  NAND U37995 ( .A(n35833), .B(mul_pow), .Z(n35832) );
  XOR U37996 ( .A(mreg[458]), .B(creg[458]), .Z(n35833) );
  XOR U37997 ( .A(n35834), .B(n35835), .Z(n35825) );
  ANDN U37998 ( .A(n35836), .B(n28001), .Z(n35835) );
  XOR U37999 ( .A(n35837), .B(\modmult_1/zin[0][456] ), .Z(n28001) );
  IV U38000 ( .A(n35834), .Z(n35837) );
  XNOR U38001 ( .A(n35834), .B(n28000), .Z(n35836) );
  XOR U38002 ( .A(n35838), .B(n35839), .Z(n28000) );
  AND U38003 ( .A(\modmult_1/xin[1023] ), .B(n35840), .Z(n35839) );
  IV U38004 ( .A(n35838), .Z(n35840) );
  XOR U38005 ( .A(n35841), .B(mreg[457]), .Z(n35838) );
  NAND U38006 ( .A(n35842), .B(mul_pow), .Z(n35841) );
  XOR U38007 ( .A(mreg[457]), .B(creg[457]), .Z(n35842) );
  XOR U38008 ( .A(n35843), .B(n35844), .Z(n35834) );
  ANDN U38009 ( .A(n35845), .B(n28007), .Z(n35844) );
  XOR U38010 ( .A(n35846), .B(\modmult_1/zin[0][455] ), .Z(n28007) );
  IV U38011 ( .A(n35843), .Z(n35846) );
  XNOR U38012 ( .A(n35843), .B(n28006), .Z(n35845) );
  XOR U38013 ( .A(n35847), .B(n35848), .Z(n28006) );
  AND U38014 ( .A(\modmult_1/xin[1023] ), .B(n35849), .Z(n35848) );
  IV U38015 ( .A(n35847), .Z(n35849) );
  XOR U38016 ( .A(n35850), .B(mreg[456]), .Z(n35847) );
  NAND U38017 ( .A(n35851), .B(mul_pow), .Z(n35850) );
  XOR U38018 ( .A(mreg[456]), .B(creg[456]), .Z(n35851) );
  XOR U38019 ( .A(n35852), .B(n35853), .Z(n35843) );
  ANDN U38020 ( .A(n35854), .B(n28013), .Z(n35853) );
  XOR U38021 ( .A(n35855), .B(\modmult_1/zin[0][454] ), .Z(n28013) );
  IV U38022 ( .A(n35852), .Z(n35855) );
  XNOR U38023 ( .A(n35852), .B(n28012), .Z(n35854) );
  XOR U38024 ( .A(n35856), .B(n35857), .Z(n28012) );
  AND U38025 ( .A(\modmult_1/xin[1023] ), .B(n35858), .Z(n35857) );
  IV U38026 ( .A(n35856), .Z(n35858) );
  XOR U38027 ( .A(n35859), .B(mreg[455]), .Z(n35856) );
  NAND U38028 ( .A(n35860), .B(mul_pow), .Z(n35859) );
  XOR U38029 ( .A(mreg[455]), .B(creg[455]), .Z(n35860) );
  XOR U38030 ( .A(n35861), .B(n35862), .Z(n35852) );
  ANDN U38031 ( .A(n35863), .B(n28019), .Z(n35862) );
  XOR U38032 ( .A(n35864), .B(\modmult_1/zin[0][453] ), .Z(n28019) );
  IV U38033 ( .A(n35861), .Z(n35864) );
  XNOR U38034 ( .A(n35861), .B(n28018), .Z(n35863) );
  XOR U38035 ( .A(n35865), .B(n35866), .Z(n28018) );
  AND U38036 ( .A(\modmult_1/xin[1023] ), .B(n35867), .Z(n35866) );
  IV U38037 ( .A(n35865), .Z(n35867) );
  XOR U38038 ( .A(n35868), .B(mreg[454]), .Z(n35865) );
  NAND U38039 ( .A(n35869), .B(mul_pow), .Z(n35868) );
  XOR U38040 ( .A(mreg[454]), .B(creg[454]), .Z(n35869) );
  XOR U38041 ( .A(n35870), .B(n35871), .Z(n35861) );
  ANDN U38042 ( .A(n35872), .B(n28025), .Z(n35871) );
  XOR U38043 ( .A(n35873), .B(\modmult_1/zin[0][452] ), .Z(n28025) );
  IV U38044 ( .A(n35870), .Z(n35873) );
  XNOR U38045 ( .A(n35870), .B(n28024), .Z(n35872) );
  XOR U38046 ( .A(n35874), .B(n35875), .Z(n28024) );
  AND U38047 ( .A(\modmult_1/xin[1023] ), .B(n35876), .Z(n35875) );
  IV U38048 ( .A(n35874), .Z(n35876) );
  XOR U38049 ( .A(n35877), .B(mreg[453]), .Z(n35874) );
  NAND U38050 ( .A(n35878), .B(mul_pow), .Z(n35877) );
  XOR U38051 ( .A(mreg[453]), .B(creg[453]), .Z(n35878) );
  XOR U38052 ( .A(n35879), .B(n35880), .Z(n35870) );
  ANDN U38053 ( .A(n35881), .B(n28031), .Z(n35880) );
  XOR U38054 ( .A(n35882), .B(\modmult_1/zin[0][451] ), .Z(n28031) );
  IV U38055 ( .A(n35879), .Z(n35882) );
  XNOR U38056 ( .A(n35879), .B(n28030), .Z(n35881) );
  XOR U38057 ( .A(n35883), .B(n35884), .Z(n28030) );
  AND U38058 ( .A(\modmult_1/xin[1023] ), .B(n35885), .Z(n35884) );
  IV U38059 ( .A(n35883), .Z(n35885) );
  XOR U38060 ( .A(n35886), .B(mreg[452]), .Z(n35883) );
  NAND U38061 ( .A(n35887), .B(mul_pow), .Z(n35886) );
  XOR U38062 ( .A(mreg[452]), .B(creg[452]), .Z(n35887) );
  XOR U38063 ( .A(n35888), .B(n35889), .Z(n35879) );
  ANDN U38064 ( .A(n35890), .B(n28037), .Z(n35889) );
  XOR U38065 ( .A(n35891), .B(\modmult_1/zin[0][450] ), .Z(n28037) );
  IV U38066 ( .A(n35888), .Z(n35891) );
  XNOR U38067 ( .A(n35888), .B(n28036), .Z(n35890) );
  XOR U38068 ( .A(n35892), .B(n35893), .Z(n28036) );
  AND U38069 ( .A(\modmult_1/xin[1023] ), .B(n35894), .Z(n35893) );
  IV U38070 ( .A(n35892), .Z(n35894) );
  XOR U38071 ( .A(n35895), .B(mreg[451]), .Z(n35892) );
  NAND U38072 ( .A(n35896), .B(mul_pow), .Z(n35895) );
  XOR U38073 ( .A(mreg[451]), .B(creg[451]), .Z(n35896) );
  XOR U38074 ( .A(n35897), .B(n35898), .Z(n35888) );
  ANDN U38075 ( .A(n35899), .B(n28043), .Z(n35898) );
  XOR U38076 ( .A(n35900), .B(\modmult_1/zin[0][449] ), .Z(n28043) );
  IV U38077 ( .A(n35897), .Z(n35900) );
  XNOR U38078 ( .A(n35897), .B(n28042), .Z(n35899) );
  XOR U38079 ( .A(n35901), .B(n35902), .Z(n28042) );
  AND U38080 ( .A(\modmult_1/xin[1023] ), .B(n35903), .Z(n35902) );
  IV U38081 ( .A(n35901), .Z(n35903) );
  XOR U38082 ( .A(n35904), .B(mreg[450]), .Z(n35901) );
  NAND U38083 ( .A(n35905), .B(mul_pow), .Z(n35904) );
  XOR U38084 ( .A(mreg[450]), .B(creg[450]), .Z(n35905) );
  XOR U38085 ( .A(n35906), .B(n35907), .Z(n35897) );
  ANDN U38086 ( .A(n35908), .B(n28049), .Z(n35907) );
  XOR U38087 ( .A(n35909), .B(\modmult_1/zin[0][448] ), .Z(n28049) );
  IV U38088 ( .A(n35906), .Z(n35909) );
  XNOR U38089 ( .A(n35906), .B(n28048), .Z(n35908) );
  XOR U38090 ( .A(n35910), .B(n35911), .Z(n28048) );
  AND U38091 ( .A(\modmult_1/xin[1023] ), .B(n35912), .Z(n35911) );
  IV U38092 ( .A(n35910), .Z(n35912) );
  XOR U38093 ( .A(n35913), .B(mreg[449]), .Z(n35910) );
  NAND U38094 ( .A(n35914), .B(mul_pow), .Z(n35913) );
  XOR U38095 ( .A(mreg[449]), .B(creg[449]), .Z(n35914) );
  XOR U38096 ( .A(n35915), .B(n35916), .Z(n35906) );
  ANDN U38097 ( .A(n35917), .B(n28055), .Z(n35916) );
  XOR U38098 ( .A(n35918), .B(\modmult_1/zin[0][447] ), .Z(n28055) );
  IV U38099 ( .A(n35915), .Z(n35918) );
  XNOR U38100 ( .A(n35915), .B(n28054), .Z(n35917) );
  XOR U38101 ( .A(n35919), .B(n35920), .Z(n28054) );
  AND U38102 ( .A(\modmult_1/xin[1023] ), .B(n35921), .Z(n35920) );
  IV U38103 ( .A(n35919), .Z(n35921) );
  XOR U38104 ( .A(n35922), .B(mreg[448]), .Z(n35919) );
  NAND U38105 ( .A(n35923), .B(mul_pow), .Z(n35922) );
  XOR U38106 ( .A(mreg[448]), .B(creg[448]), .Z(n35923) );
  XOR U38107 ( .A(n35924), .B(n35925), .Z(n35915) );
  ANDN U38108 ( .A(n35926), .B(n28061), .Z(n35925) );
  XOR U38109 ( .A(n35927), .B(\modmult_1/zin[0][446] ), .Z(n28061) );
  IV U38110 ( .A(n35924), .Z(n35927) );
  XNOR U38111 ( .A(n35924), .B(n28060), .Z(n35926) );
  XOR U38112 ( .A(n35928), .B(n35929), .Z(n28060) );
  AND U38113 ( .A(\modmult_1/xin[1023] ), .B(n35930), .Z(n35929) );
  IV U38114 ( .A(n35928), .Z(n35930) );
  XOR U38115 ( .A(n35931), .B(mreg[447]), .Z(n35928) );
  NAND U38116 ( .A(n35932), .B(mul_pow), .Z(n35931) );
  XOR U38117 ( .A(mreg[447]), .B(creg[447]), .Z(n35932) );
  XOR U38118 ( .A(n35933), .B(n35934), .Z(n35924) );
  ANDN U38119 ( .A(n35935), .B(n28067), .Z(n35934) );
  XOR U38120 ( .A(n35936), .B(\modmult_1/zin[0][445] ), .Z(n28067) );
  IV U38121 ( .A(n35933), .Z(n35936) );
  XNOR U38122 ( .A(n35933), .B(n28066), .Z(n35935) );
  XOR U38123 ( .A(n35937), .B(n35938), .Z(n28066) );
  AND U38124 ( .A(\modmult_1/xin[1023] ), .B(n35939), .Z(n35938) );
  IV U38125 ( .A(n35937), .Z(n35939) );
  XOR U38126 ( .A(n35940), .B(mreg[446]), .Z(n35937) );
  NAND U38127 ( .A(n35941), .B(mul_pow), .Z(n35940) );
  XOR U38128 ( .A(mreg[446]), .B(creg[446]), .Z(n35941) );
  XOR U38129 ( .A(n35942), .B(n35943), .Z(n35933) );
  ANDN U38130 ( .A(n35944), .B(n28073), .Z(n35943) );
  XOR U38131 ( .A(n35945), .B(\modmult_1/zin[0][444] ), .Z(n28073) );
  IV U38132 ( .A(n35942), .Z(n35945) );
  XNOR U38133 ( .A(n35942), .B(n28072), .Z(n35944) );
  XOR U38134 ( .A(n35946), .B(n35947), .Z(n28072) );
  AND U38135 ( .A(\modmult_1/xin[1023] ), .B(n35948), .Z(n35947) );
  IV U38136 ( .A(n35946), .Z(n35948) );
  XOR U38137 ( .A(n35949), .B(mreg[445]), .Z(n35946) );
  NAND U38138 ( .A(n35950), .B(mul_pow), .Z(n35949) );
  XOR U38139 ( .A(mreg[445]), .B(creg[445]), .Z(n35950) );
  XOR U38140 ( .A(n35951), .B(n35952), .Z(n35942) );
  ANDN U38141 ( .A(n35953), .B(n28079), .Z(n35952) );
  XOR U38142 ( .A(n35954), .B(\modmult_1/zin[0][443] ), .Z(n28079) );
  IV U38143 ( .A(n35951), .Z(n35954) );
  XNOR U38144 ( .A(n35951), .B(n28078), .Z(n35953) );
  XOR U38145 ( .A(n35955), .B(n35956), .Z(n28078) );
  AND U38146 ( .A(\modmult_1/xin[1023] ), .B(n35957), .Z(n35956) );
  IV U38147 ( .A(n35955), .Z(n35957) );
  XOR U38148 ( .A(n35958), .B(mreg[444]), .Z(n35955) );
  NAND U38149 ( .A(n35959), .B(mul_pow), .Z(n35958) );
  XOR U38150 ( .A(mreg[444]), .B(creg[444]), .Z(n35959) );
  XOR U38151 ( .A(n35960), .B(n35961), .Z(n35951) );
  ANDN U38152 ( .A(n35962), .B(n28085), .Z(n35961) );
  XOR U38153 ( .A(n35963), .B(\modmult_1/zin[0][442] ), .Z(n28085) );
  IV U38154 ( .A(n35960), .Z(n35963) );
  XNOR U38155 ( .A(n35960), .B(n28084), .Z(n35962) );
  XOR U38156 ( .A(n35964), .B(n35965), .Z(n28084) );
  AND U38157 ( .A(\modmult_1/xin[1023] ), .B(n35966), .Z(n35965) );
  IV U38158 ( .A(n35964), .Z(n35966) );
  XOR U38159 ( .A(n35967), .B(mreg[443]), .Z(n35964) );
  NAND U38160 ( .A(n35968), .B(mul_pow), .Z(n35967) );
  XOR U38161 ( .A(mreg[443]), .B(creg[443]), .Z(n35968) );
  XOR U38162 ( .A(n35969), .B(n35970), .Z(n35960) );
  ANDN U38163 ( .A(n35971), .B(n28091), .Z(n35970) );
  XOR U38164 ( .A(n35972), .B(\modmult_1/zin[0][441] ), .Z(n28091) );
  IV U38165 ( .A(n35969), .Z(n35972) );
  XNOR U38166 ( .A(n35969), .B(n28090), .Z(n35971) );
  XOR U38167 ( .A(n35973), .B(n35974), .Z(n28090) );
  AND U38168 ( .A(\modmult_1/xin[1023] ), .B(n35975), .Z(n35974) );
  IV U38169 ( .A(n35973), .Z(n35975) );
  XOR U38170 ( .A(n35976), .B(mreg[442]), .Z(n35973) );
  NAND U38171 ( .A(n35977), .B(mul_pow), .Z(n35976) );
  XOR U38172 ( .A(mreg[442]), .B(creg[442]), .Z(n35977) );
  XOR U38173 ( .A(n35978), .B(n35979), .Z(n35969) );
  ANDN U38174 ( .A(n35980), .B(n28097), .Z(n35979) );
  XOR U38175 ( .A(n35981), .B(\modmult_1/zin[0][440] ), .Z(n28097) );
  IV U38176 ( .A(n35978), .Z(n35981) );
  XNOR U38177 ( .A(n35978), .B(n28096), .Z(n35980) );
  XOR U38178 ( .A(n35982), .B(n35983), .Z(n28096) );
  AND U38179 ( .A(\modmult_1/xin[1023] ), .B(n35984), .Z(n35983) );
  IV U38180 ( .A(n35982), .Z(n35984) );
  XOR U38181 ( .A(n35985), .B(mreg[441]), .Z(n35982) );
  NAND U38182 ( .A(n35986), .B(mul_pow), .Z(n35985) );
  XOR U38183 ( .A(mreg[441]), .B(creg[441]), .Z(n35986) );
  XOR U38184 ( .A(n35987), .B(n35988), .Z(n35978) );
  ANDN U38185 ( .A(n35989), .B(n28103), .Z(n35988) );
  XOR U38186 ( .A(n35990), .B(\modmult_1/zin[0][439] ), .Z(n28103) );
  IV U38187 ( .A(n35987), .Z(n35990) );
  XNOR U38188 ( .A(n35987), .B(n28102), .Z(n35989) );
  XOR U38189 ( .A(n35991), .B(n35992), .Z(n28102) );
  AND U38190 ( .A(\modmult_1/xin[1023] ), .B(n35993), .Z(n35992) );
  IV U38191 ( .A(n35991), .Z(n35993) );
  XOR U38192 ( .A(n35994), .B(mreg[440]), .Z(n35991) );
  NAND U38193 ( .A(n35995), .B(mul_pow), .Z(n35994) );
  XOR U38194 ( .A(mreg[440]), .B(creg[440]), .Z(n35995) );
  XOR U38195 ( .A(n35996), .B(n35997), .Z(n35987) );
  ANDN U38196 ( .A(n35998), .B(n28109), .Z(n35997) );
  XOR U38197 ( .A(n35999), .B(\modmult_1/zin[0][438] ), .Z(n28109) );
  IV U38198 ( .A(n35996), .Z(n35999) );
  XNOR U38199 ( .A(n35996), .B(n28108), .Z(n35998) );
  XOR U38200 ( .A(n36000), .B(n36001), .Z(n28108) );
  AND U38201 ( .A(\modmult_1/xin[1023] ), .B(n36002), .Z(n36001) );
  IV U38202 ( .A(n36000), .Z(n36002) );
  XOR U38203 ( .A(n36003), .B(mreg[439]), .Z(n36000) );
  NAND U38204 ( .A(n36004), .B(mul_pow), .Z(n36003) );
  XOR U38205 ( .A(mreg[439]), .B(creg[439]), .Z(n36004) );
  XOR U38206 ( .A(n36005), .B(n36006), .Z(n35996) );
  ANDN U38207 ( .A(n36007), .B(n28115), .Z(n36006) );
  XOR U38208 ( .A(n36008), .B(\modmult_1/zin[0][437] ), .Z(n28115) );
  IV U38209 ( .A(n36005), .Z(n36008) );
  XNOR U38210 ( .A(n36005), .B(n28114), .Z(n36007) );
  XOR U38211 ( .A(n36009), .B(n36010), .Z(n28114) );
  AND U38212 ( .A(\modmult_1/xin[1023] ), .B(n36011), .Z(n36010) );
  IV U38213 ( .A(n36009), .Z(n36011) );
  XOR U38214 ( .A(n36012), .B(mreg[438]), .Z(n36009) );
  NAND U38215 ( .A(n36013), .B(mul_pow), .Z(n36012) );
  XOR U38216 ( .A(mreg[438]), .B(creg[438]), .Z(n36013) );
  XOR U38217 ( .A(n36014), .B(n36015), .Z(n36005) );
  ANDN U38218 ( .A(n36016), .B(n28121), .Z(n36015) );
  XOR U38219 ( .A(n36017), .B(\modmult_1/zin[0][436] ), .Z(n28121) );
  IV U38220 ( .A(n36014), .Z(n36017) );
  XNOR U38221 ( .A(n36014), .B(n28120), .Z(n36016) );
  XOR U38222 ( .A(n36018), .B(n36019), .Z(n28120) );
  AND U38223 ( .A(\modmult_1/xin[1023] ), .B(n36020), .Z(n36019) );
  IV U38224 ( .A(n36018), .Z(n36020) );
  XOR U38225 ( .A(n36021), .B(mreg[437]), .Z(n36018) );
  NAND U38226 ( .A(n36022), .B(mul_pow), .Z(n36021) );
  XOR U38227 ( .A(mreg[437]), .B(creg[437]), .Z(n36022) );
  XOR U38228 ( .A(n36023), .B(n36024), .Z(n36014) );
  ANDN U38229 ( .A(n36025), .B(n28127), .Z(n36024) );
  XOR U38230 ( .A(n36026), .B(\modmult_1/zin[0][435] ), .Z(n28127) );
  IV U38231 ( .A(n36023), .Z(n36026) );
  XNOR U38232 ( .A(n36023), .B(n28126), .Z(n36025) );
  XOR U38233 ( .A(n36027), .B(n36028), .Z(n28126) );
  AND U38234 ( .A(\modmult_1/xin[1023] ), .B(n36029), .Z(n36028) );
  IV U38235 ( .A(n36027), .Z(n36029) );
  XOR U38236 ( .A(n36030), .B(mreg[436]), .Z(n36027) );
  NAND U38237 ( .A(n36031), .B(mul_pow), .Z(n36030) );
  XOR U38238 ( .A(mreg[436]), .B(creg[436]), .Z(n36031) );
  XOR U38239 ( .A(n36032), .B(n36033), .Z(n36023) );
  ANDN U38240 ( .A(n36034), .B(n28133), .Z(n36033) );
  XOR U38241 ( .A(n36035), .B(\modmult_1/zin[0][434] ), .Z(n28133) );
  IV U38242 ( .A(n36032), .Z(n36035) );
  XNOR U38243 ( .A(n36032), .B(n28132), .Z(n36034) );
  XOR U38244 ( .A(n36036), .B(n36037), .Z(n28132) );
  AND U38245 ( .A(\modmult_1/xin[1023] ), .B(n36038), .Z(n36037) );
  IV U38246 ( .A(n36036), .Z(n36038) );
  XOR U38247 ( .A(n36039), .B(mreg[435]), .Z(n36036) );
  NAND U38248 ( .A(n36040), .B(mul_pow), .Z(n36039) );
  XOR U38249 ( .A(mreg[435]), .B(creg[435]), .Z(n36040) );
  XOR U38250 ( .A(n36041), .B(n36042), .Z(n36032) );
  ANDN U38251 ( .A(n36043), .B(n28139), .Z(n36042) );
  XOR U38252 ( .A(n36044), .B(\modmult_1/zin[0][433] ), .Z(n28139) );
  IV U38253 ( .A(n36041), .Z(n36044) );
  XNOR U38254 ( .A(n36041), .B(n28138), .Z(n36043) );
  XOR U38255 ( .A(n36045), .B(n36046), .Z(n28138) );
  AND U38256 ( .A(\modmult_1/xin[1023] ), .B(n36047), .Z(n36046) );
  IV U38257 ( .A(n36045), .Z(n36047) );
  XOR U38258 ( .A(n36048), .B(mreg[434]), .Z(n36045) );
  NAND U38259 ( .A(n36049), .B(mul_pow), .Z(n36048) );
  XOR U38260 ( .A(mreg[434]), .B(creg[434]), .Z(n36049) );
  XOR U38261 ( .A(n36050), .B(n36051), .Z(n36041) );
  ANDN U38262 ( .A(n36052), .B(n28145), .Z(n36051) );
  XOR U38263 ( .A(n36053), .B(\modmult_1/zin[0][432] ), .Z(n28145) );
  IV U38264 ( .A(n36050), .Z(n36053) );
  XNOR U38265 ( .A(n36050), .B(n28144), .Z(n36052) );
  XOR U38266 ( .A(n36054), .B(n36055), .Z(n28144) );
  AND U38267 ( .A(\modmult_1/xin[1023] ), .B(n36056), .Z(n36055) );
  IV U38268 ( .A(n36054), .Z(n36056) );
  XOR U38269 ( .A(n36057), .B(mreg[433]), .Z(n36054) );
  NAND U38270 ( .A(n36058), .B(mul_pow), .Z(n36057) );
  XOR U38271 ( .A(mreg[433]), .B(creg[433]), .Z(n36058) );
  XOR U38272 ( .A(n36059), .B(n36060), .Z(n36050) );
  ANDN U38273 ( .A(n36061), .B(n28151), .Z(n36060) );
  XOR U38274 ( .A(n36062), .B(\modmult_1/zin[0][431] ), .Z(n28151) );
  IV U38275 ( .A(n36059), .Z(n36062) );
  XNOR U38276 ( .A(n36059), .B(n28150), .Z(n36061) );
  XOR U38277 ( .A(n36063), .B(n36064), .Z(n28150) );
  AND U38278 ( .A(\modmult_1/xin[1023] ), .B(n36065), .Z(n36064) );
  IV U38279 ( .A(n36063), .Z(n36065) );
  XOR U38280 ( .A(n36066), .B(mreg[432]), .Z(n36063) );
  NAND U38281 ( .A(n36067), .B(mul_pow), .Z(n36066) );
  XOR U38282 ( .A(mreg[432]), .B(creg[432]), .Z(n36067) );
  XOR U38283 ( .A(n36068), .B(n36069), .Z(n36059) );
  ANDN U38284 ( .A(n36070), .B(n28157), .Z(n36069) );
  XOR U38285 ( .A(n36071), .B(\modmult_1/zin[0][430] ), .Z(n28157) );
  IV U38286 ( .A(n36068), .Z(n36071) );
  XNOR U38287 ( .A(n36068), .B(n28156), .Z(n36070) );
  XOR U38288 ( .A(n36072), .B(n36073), .Z(n28156) );
  AND U38289 ( .A(\modmult_1/xin[1023] ), .B(n36074), .Z(n36073) );
  IV U38290 ( .A(n36072), .Z(n36074) );
  XOR U38291 ( .A(n36075), .B(mreg[431]), .Z(n36072) );
  NAND U38292 ( .A(n36076), .B(mul_pow), .Z(n36075) );
  XOR U38293 ( .A(mreg[431]), .B(creg[431]), .Z(n36076) );
  XOR U38294 ( .A(n36077), .B(n36078), .Z(n36068) );
  ANDN U38295 ( .A(n36079), .B(n28163), .Z(n36078) );
  XOR U38296 ( .A(n36080), .B(\modmult_1/zin[0][429] ), .Z(n28163) );
  IV U38297 ( .A(n36077), .Z(n36080) );
  XNOR U38298 ( .A(n36077), .B(n28162), .Z(n36079) );
  XOR U38299 ( .A(n36081), .B(n36082), .Z(n28162) );
  AND U38300 ( .A(\modmult_1/xin[1023] ), .B(n36083), .Z(n36082) );
  IV U38301 ( .A(n36081), .Z(n36083) );
  XOR U38302 ( .A(n36084), .B(mreg[430]), .Z(n36081) );
  NAND U38303 ( .A(n36085), .B(mul_pow), .Z(n36084) );
  XOR U38304 ( .A(mreg[430]), .B(creg[430]), .Z(n36085) );
  XOR U38305 ( .A(n36086), .B(n36087), .Z(n36077) );
  ANDN U38306 ( .A(n36088), .B(n28169), .Z(n36087) );
  XOR U38307 ( .A(n36089), .B(\modmult_1/zin[0][428] ), .Z(n28169) );
  IV U38308 ( .A(n36086), .Z(n36089) );
  XNOR U38309 ( .A(n36086), .B(n28168), .Z(n36088) );
  XOR U38310 ( .A(n36090), .B(n36091), .Z(n28168) );
  AND U38311 ( .A(\modmult_1/xin[1023] ), .B(n36092), .Z(n36091) );
  IV U38312 ( .A(n36090), .Z(n36092) );
  XOR U38313 ( .A(n36093), .B(mreg[429]), .Z(n36090) );
  NAND U38314 ( .A(n36094), .B(mul_pow), .Z(n36093) );
  XOR U38315 ( .A(mreg[429]), .B(creg[429]), .Z(n36094) );
  XOR U38316 ( .A(n36095), .B(n36096), .Z(n36086) );
  ANDN U38317 ( .A(n36097), .B(n28175), .Z(n36096) );
  XOR U38318 ( .A(n36098), .B(\modmult_1/zin[0][427] ), .Z(n28175) );
  IV U38319 ( .A(n36095), .Z(n36098) );
  XNOR U38320 ( .A(n36095), .B(n28174), .Z(n36097) );
  XOR U38321 ( .A(n36099), .B(n36100), .Z(n28174) );
  AND U38322 ( .A(\modmult_1/xin[1023] ), .B(n36101), .Z(n36100) );
  IV U38323 ( .A(n36099), .Z(n36101) );
  XOR U38324 ( .A(n36102), .B(mreg[428]), .Z(n36099) );
  NAND U38325 ( .A(n36103), .B(mul_pow), .Z(n36102) );
  XOR U38326 ( .A(mreg[428]), .B(creg[428]), .Z(n36103) );
  XOR U38327 ( .A(n36104), .B(n36105), .Z(n36095) );
  ANDN U38328 ( .A(n36106), .B(n28181), .Z(n36105) );
  XOR U38329 ( .A(n36107), .B(\modmult_1/zin[0][426] ), .Z(n28181) );
  IV U38330 ( .A(n36104), .Z(n36107) );
  XNOR U38331 ( .A(n36104), .B(n28180), .Z(n36106) );
  XOR U38332 ( .A(n36108), .B(n36109), .Z(n28180) );
  AND U38333 ( .A(\modmult_1/xin[1023] ), .B(n36110), .Z(n36109) );
  IV U38334 ( .A(n36108), .Z(n36110) );
  XOR U38335 ( .A(n36111), .B(mreg[427]), .Z(n36108) );
  NAND U38336 ( .A(n36112), .B(mul_pow), .Z(n36111) );
  XOR U38337 ( .A(mreg[427]), .B(creg[427]), .Z(n36112) );
  XOR U38338 ( .A(n36113), .B(n36114), .Z(n36104) );
  ANDN U38339 ( .A(n36115), .B(n28187), .Z(n36114) );
  XOR U38340 ( .A(n36116), .B(\modmult_1/zin[0][425] ), .Z(n28187) );
  IV U38341 ( .A(n36113), .Z(n36116) );
  XNOR U38342 ( .A(n36113), .B(n28186), .Z(n36115) );
  XOR U38343 ( .A(n36117), .B(n36118), .Z(n28186) );
  AND U38344 ( .A(\modmult_1/xin[1023] ), .B(n36119), .Z(n36118) );
  IV U38345 ( .A(n36117), .Z(n36119) );
  XOR U38346 ( .A(n36120), .B(mreg[426]), .Z(n36117) );
  NAND U38347 ( .A(n36121), .B(mul_pow), .Z(n36120) );
  XOR U38348 ( .A(mreg[426]), .B(creg[426]), .Z(n36121) );
  XOR U38349 ( .A(n36122), .B(n36123), .Z(n36113) );
  ANDN U38350 ( .A(n36124), .B(n28193), .Z(n36123) );
  XOR U38351 ( .A(n36125), .B(\modmult_1/zin[0][424] ), .Z(n28193) );
  IV U38352 ( .A(n36122), .Z(n36125) );
  XNOR U38353 ( .A(n36122), .B(n28192), .Z(n36124) );
  XOR U38354 ( .A(n36126), .B(n36127), .Z(n28192) );
  AND U38355 ( .A(\modmult_1/xin[1023] ), .B(n36128), .Z(n36127) );
  IV U38356 ( .A(n36126), .Z(n36128) );
  XOR U38357 ( .A(n36129), .B(mreg[425]), .Z(n36126) );
  NAND U38358 ( .A(n36130), .B(mul_pow), .Z(n36129) );
  XOR U38359 ( .A(mreg[425]), .B(creg[425]), .Z(n36130) );
  XOR U38360 ( .A(n36131), .B(n36132), .Z(n36122) );
  ANDN U38361 ( .A(n36133), .B(n28199), .Z(n36132) );
  XOR U38362 ( .A(n36134), .B(\modmult_1/zin[0][423] ), .Z(n28199) );
  IV U38363 ( .A(n36131), .Z(n36134) );
  XNOR U38364 ( .A(n36131), .B(n28198), .Z(n36133) );
  XOR U38365 ( .A(n36135), .B(n36136), .Z(n28198) );
  AND U38366 ( .A(\modmult_1/xin[1023] ), .B(n36137), .Z(n36136) );
  IV U38367 ( .A(n36135), .Z(n36137) );
  XOR U38368 ( .A(n36138), .B(mreg[424]), .Z(n36135) );
  NAND U38369 ( .A(n36139), .B(mul_pow), .Z(n36138) );
  XOR U38370 ( .A(mreg[424]), .B(creg[424]), .Z(n36139) );
  XOR U38371 ( .A(n36140), .B(n36141), .Z(n36131) );
  ANDN U38372 ( .A(n36142), .B(n28205), .Z(n36141) );
  XOR U38373 ( .A(n36143), .B(\modmult_1/zin[0][422] ), .Z(n28205) );
  IV U38374 ( .A(n36140), .Z(n36143) );
  XNOR U38375 ( .A(n36140), .B(n28204), .Z(n36142) );
  XOR U38376 ( .A(n36144), .B(n36145), .Z(n28204) );
  AND U38377 ( .A(\modmult_1/xin[1023] ), .B(n36146), .Z(n36145) );
  IV U38378 ( .A(n36144), .Z(n36146) );
  XOR U38379 ( .A(n36147), .B(mreg[423]), .Z(n36144) );
  NAND U38380 ( .A(n36148), .B(mul_pow), .Z(n36147) );
  XOR U38381 ( .A(mreg[423]), .B(creg[423]), .Z(n36148) );
  XOR U38382 ( .A(n36149), .B(n36150), .Z(n36140) );
  ANDN U38383 ( .A(n36151), .B(n28211), .Z(n36150) );
  XOR U38384 ( .A(n36152), .B(\modmult_1/zin[0][421] ), .Z(n28211) );
  IV U38385 ( .A(n36149), .Z(n36152) );
  XNOR U38386 ( .A(n36149), .B(n28210), .Z(n36151) );
  XOR U38387 ( .A(n36153), .B(n36154), .Z(n28210) );
  AND U38388 ( .A(\modmult_1/xin[1023] ), .B(n36155), .Z(n36154) );
  IV U38389 ( .A(n36153), .Z(n36155) );
  XOR U38390 ( .A(n36156), .B(mreg[422]), .Z(n36153) );
  NAND U38391 ( .A(n36157), .B(mul_pow), .Z(n36156) );
  XOR U38392 ( .A(mreg[422]), .B(creg[422]), .Z(n36157) );
  XOR U38393 ( .A(n36158), .B(n36159), .Z(n36149) );
  ANDN U38394 ( .A(n36160), .B(n28217), .Z(n36159) );
  XOR U38395 ( .A(n36161), .B(\modmult_1/zin[0][420] ), .Z(n28217) );
  IV U38396 ( .A(n36158), .Z(n36161) );
  XNOR U38397 ( .A(n36158), .B(n28216), .Z(n36160) );
  XOR U38398 ( .A(n36162), .B(n36163), .Z(n28216) );
  AND U38399 ( .A(\modmult_1/xin[1023] ), .B(n36164), .Z(n36163) );
  IV U38400 ( .A(n36162), .Z(n36164) );
  XOR U38401 ( .A(n36165), .B(mreg[421]), .Z(n36162) );
  NAND U38402 ( .A(n36166), .B(mul_pow), .Z(n36165) );
  XOR U38403 ( .A(mreg[421]), .B(creg[421]), .Z(n36166) );
  XOR U38404 ( .A(n36167), .B(n36168), .Z(n36158) );
  ANDN U38405 ( .A(n36169), .B(n28223), .Z(n36168) );
  XOR U38406 ( .A(n36170), .B(\modmult_1/zin[0][419] ), .Z(n28223) );
  IV U38407 ( .A(n36167), .Z(n36170) );
  XNOR U38408 ( .A(n36167), .B(n28222), .Z(n36169) );
  XOR U38409 ( .A(n36171), .B(n36172), .Z(n28222) );
  AND U38410 ( .A(\modmult_1/xin[1023] ), .B(n36173), .Z(n36172) );
  IV U38411 ( .A(n36171), .Z(n36173) );
  XOR U38412 ( .A(n36174), .B(mreg[420]), .Z(n36171) );
  NAND U38413 ( .A(n36175), .B(mul_pow), .Z(n36174) );
  XOR U38414 ( .A(mreg[420]), .B(creg[420]), .Z(n36175) );
  XOR U38415 ( .A(n36176), .B(n36177), .Z(n36167) );
  ANDN U38416 ( .A(n36178), .B(n28229), .Z(n36177) );
  XOR U38417 ( .A(n36179), .B(\modmult_1/zin[0][418] ), .Z(n28229) );
  IV U38418 ( .A(n36176), .Z(n36179) );
  XNOR U38419 ( .A(n36176), .B(n28228), .Z(n36178) );
  XOR U38420 ( .A(n36180), .B(n36181), .Z(n28228) );
  AND U38421 ( .A(\modmult_1/xin[1023] ), .B(n36182), .Z(n36181) );
  IV U38422 ( .A(n36180), .Z(n36182) );
  XOR U38423 ( .A(n36183), .B(mreg[419]), .Z(n36180) );
  NAND U38424 ( .A(n36184), .B(mul_pow), .Z(n36183) );
  XOR U38425 ( .A(mreg[419]), .B(creg[419]), .Z(n36184) );
  XOR U38426 ( .A(n36185), .B(n36186), .Z(n36176) );
  ANDN U38427 ( .A(n36187), .B(n28235), .Z(n36186) );
  XOR U38428 ( .A(n36188), .B(\modmult_1/zin[0][417] ), .Z(n28235) );
  IV U38429 ( .A(n36185), .Z(n36188) );
  XNOR U38430 ( .A(n36185), .B(n28234), .Z(n36187) );
  XOR U38431 ( .A(n36189), .B(n36190), .Z(n28234) );
  AND U38432 ( .A(\modmult_1/xin[1023] ), .B(n36191), .Z(n36190) );
  IV U38433 ( .A(n36189), .Z(n36191) );
  XOR U38434 ( .A(n36192), .B(mreg[418]), .Z(n36189) );
  NAND U38435 ( .A(n36193), .B(mul_pow), .Z(n36192) );
  XOR U38436 ( .A(mreg[418]), .B(creg[418]), .Z(n36193) );
  XOR U38437 ( .A(n36194), .B(n36195), .Z(n36185) );
  ANDN U38438 ( .A(n36196), .B(n28241), .Z(n36195) );
  XOR U38439 ( .A(n36197), .B(\modmult_1/zin[0][416] ), .Z(n28241) );
  IV U38440 ( .A(n36194), .Z(n36197) );
  XNOR U38441 ( .A(n36194), .B(n28240), .Z(n36196) );
  XOR U38442 ( .A(n36198), .B(n36199), .Z(n28240) );
  AND U38443 ( .A(\modmult_1/xin[1023] ), .B(n36200), .Z(n36199) );
  IV U38444 ( .A(n36198), .Z(n36200) );
  XOR U38445 ( .A(n36201), .B(mreg[417]), .Z(n36198) );
  NAND U38446 ( .A(n36202), .B(mul_pow), .Z(n36201) );
  XOR U38447 ( .A(mreg[417]), .B(creg[417]), .Z(n36202) );
  XOR U38448 ( .A(n36203), .B(n36204), .Z(n36194) );
  ANDN U38449 ( .A(n36205), .B(n28247), .Z(n36204) );
  XOR U38450 ( .A(n36206), .B(\modmult_1/zin[0][415] ), .Z(n28247) );
  IV U38451 ( .A(n36203), .Z(n36206) );
  XNOR U38452 ( .A(n36203), .B(n28246), .Z(n36205) );
  XOR U38453 ( .A(n36207), .B(n36208), .Z(n28246) );
  AND U38454 ( .A(\modmult_1/xin[1023] ), .B(n36209), .Z(n36208) );
  IV U38455 ( .A(n36207), .Z(n36209) );
  XOR U38456 ( .A(n36210), .B(mreg[416]), .Z(n36207) );
  NAND U38457 ( .A(n36211), .B(mul_pow), .Z(n36210) );
  XOR U38458 ( .A(mreg[416]), .B(creg[416]), .Z(n36211) );
  XOR U38459 ( .A(n36212), .B(n36213), .Z(n36203) );
  ANDN U38460 ( .A(n36214), .B(n28253), .Z(n36213) );
  XOR U38461 ( .A(n36215), .B(\modmult_1/zin[0][414] ), .Z(n28253) );
  IV U38462 ( .A(n36212), .Z(n36215) );
  XNOR U38463 ( .A(n36212), .B(n28252), .Z(n36214) );
  XOR U38464 ( .A(n36216), .B(n36217), .Z(n28252) );
  AND U38465 ( .A(\modmult_1/xin[1023] ), .B(n36218), .Z(n36217) );
  IV U38466 ( .A(n36216), .Z(n36218) );
  XOR U38467 ( .A(n36219), .B(mreg[415]), .Z(n36216) );
  NAND U38468 ( .A(n36220), .B(mul_pow), .Z(n36219) );
  XOR U38469 ( .A(mreg[415]), .B(creg[415]), .Z(n36220) );
  XOR U38470 ( .A(n36221), .B(n36222), .Z(n36212) );
  ANDN U38471 ( .A(n36223), .B(n28259), .Z(n36222) );
  XOR U38472 ( .A(n36224), .B(\modmult_1/zin[0][413] ), .Z(n28259) );
  IV U38473 ( .A(n36221), .Z(n36224) );
  XNOR U38474 ( .A(n36221), .B(n28258), .Z(n36223) );
  XOR U38475 ( .A(n36225), .B(n36226), .Z(n28258) );
  AND U38476 ( .A(\modmult_1/xin[1023] ), .B(n36227), .Z(n36226) );
  IV U38477 ( .A(n36225), .Z(n36227) );
  XOR U38478 ( .A(n36228), .B(mreg[414]), .Z(n36225) );
  NAND U38479 ( .A(n36229), .B(mul_pow), .Z(n36228) );
  XOR U38480 ( .A(mreg[414]), .B(creg[414]), .Z(n36229) );
  XOR U38481 ( .A(n36230), .B(n36231), .Z(n36221) );
  ANDN U38482 ( .A(n36232), .B(n28265), .Z(n36231) );
  XOR U38483 ( .A(n36233), .B(\modmult_1/zin[0][412] ), .Z(n28265) );
  IV U38484 ( .A(n36230), .Z(n36233) );
  XNOR U38485 ( .A(n36230), .B(n28264), .Z(n36232) );
  XOR U38486 ( .A(n36234), .B(n36235), .Z(n28264) );
  AND U38487 ( .A(\modmult_1/xin[1023] ), .B(n36236), .Z(n36235) );
  IV U38488 ( .A(n36234), .Z(n36236) );
  XOR U38489 ( .A(n36237), .B(mreg[413]), .Z(n36234) );
  NAND U38490 ( .A(n36238), .B(mul_pow), .Z(n36237) );
  XOR U38491 ( .A(mreg[413]), .B(creg[413]), .Z(n36238) );
  XOR U38492 ( .A(n36239), .B(n36240), .Z(n36230) );
  ANDN U38493 ( .A(n36241), .B(n28271), .Z(n36240) );
  XOR U38494 ( .A(n36242), .B(\modmult_1/zin[0][411] ), .Z(n28271) );
  IV U38495 ( .A(n36239), .Z(n36242) );
  XNOR U38496 ( .A(n36239), .B(n28270), .Z(n36241) );
  XOR U38497 ( .A(n36243), .B(n36244), .Z(n28270) );
  AND U38498 ( .A(\modmult_1/xin[1023] ), .B(n36245), .Z(n36244) );
  IV U38499 ( .A(n36243), .Z(n36245) );
  XOR U38500 ( .A(n36246), .B(mreg[412]), .Z(n36243) );
  NAND U38501 ( .A(n36247), .B(mul_pow), .Z(n36246) );
  XOR U38502 ( .A(mreg[412]), .B(creg[412]), .Z(n36247) );
  XOR U38503 ( .A(n36248), .B(n36249), .Z(n36239) );
  ANDN U38504 ( .A(n36250), .B(n28277), .Z(n36249) );
  XOR U38505 ( .A(n36251), .B(\modmult_1/zin[0][410] ), .Z(n28277) );
  IV U38506 ( .A(n36248), .Z(n36251) );
  XNOR U38507 ( .A(n36248), .B(n28276), .Z(n36250) );
  XOR U38508 ( .A(n36252), .B(n36253), .Z(n28276) );
  AND U38509 ( .A(\modmult_1/xin[1023] ), .B(n36254), .Z(n36253) );
  IV U38510 ( .A(n36252), .Z(n36254) );
  XOR U38511 ( .A(n36255), .B(mreg[411]), .Z(n36252) );
  NAND U38512 ( .A(n36256), .B(mul_pow), .Z(n36255) );
  XOR U38513 ( .A(mreg[411]), .B(creg[411]), .Z(n36256) );
  XOR U38514 ( .A(n36257), .B(n36258), .Z(n36248) );
  ANDN U38515 ( .A(n36259), .B(n28283), .Z(n36258) );
  XOR U38516 ( .A(n36260), .B(\modmult_1/zin[0][409] ), .Z(n28283) );
  IV U38517 ( .A(n36257), .Z(n36260) );
  XNOR U38518 ( .A(n36257), .B(n28282), .Z(n36259) );
  XOR U38519 ( .A(n36261), .B(n36262), .Z(n28282) );
  AND U38520 ( .A(\modmult_1/xin[1023] ), .B(n36263), .Z(n36262) );
  IV U38521 ( .A(n36261), .Z(n36263) );
  XOR U38522 ( .A(n36264), .B(mreg[410]), .Z(n36261) );
  NAND U38523 ( .A(n36265), .B(mul_pow), .Z(n36264) );
  XOR U38524 ( .A(mreg[410]), .B(creg[410]), .Z(n36265) );
  XOR U38525 ( .A(n36266), .B(n36267), .Z(n36257) );
  ANDN U38526 ( .A(n36268), .B(n28289), .Z(n36267) );
  XOR U38527 ( .A(n36269), .B(\modmult_1/zin[0][408] ), .Z(n28289) );
  IV U38528 ( .A(n36266), .Z(n36269) );
  XNOR U38529 ( .A(n36266), .B(n28288), .Z(n36268) );
  XOR U38530 ( .A(n36270), .B(n36271), .Z(n28288) );
  AND U38531 ( .A(\modmult_1/xin[1023] ), .B(n36272), .Z(n36271) );
  IV U38532 ( .A(n36270), .Z(n36272) );
  XOR U38533 ( .A(n36273), .B(mreg[409]), .Z(n36270) );
  NAND U38534 ( .A(n36274), .B(mul_pow), .Z(n36273) );
  XOR U38535 ( .A(mreg[409]), .B(creg[409]), .Z(n36274) );
  XOR U38536 ( .A(n36275), .B(n36276), .Z(n36266) );
  ANDN U38537 ( .A(n36277), .B(n28295), .Z(n36276) );
  XOR U38538 ( .A(n36278), .B(\modmult_1/zin[0][407] ), .Z(n28295) );
  IV U38539 ( .A(n36275), .Z(n36278) );
  XNOR U38540 ( .A(n36275), .B(n28294), .Z(n36277) );
  XOR U38541 ( .A(n36279), .B(n36280), .Z(n28294) );
  AND U38542 ( .A(\modmult_1/xin[1023] ), .B(n36281), .Z(n36280) );
  IV U38543 ( .A(n36279), .Z(n36281) );
  XOR U38544 ( .A(n36282), .B(mreg[408]), .Z(n36279) );
  NAND U38545 ( .A(n36283), .B(mul_pow), .Z(n36282) );
  XOR U38546 ( .A(mreg[408]), .B(creg[408]), .Z(n36283) );
  XOR U38547 ( .A(n36284), .B(n36285), .Z(n36275) );
  ANDN U38548 ( .A(n36286), .B(n28301), .Z(n36285) );
  XOR U38549 ( .A(n36287), .B(\modmult_1/zin[0][406] ), .Z(n28301) );
  IV U38550 ( .A(n36284), .Z(n36287) );
  XNOR U38551 ( .A(n36284), .B(n28300), .Z(n36286) );
  XOR U38552 ( .A(n36288), .B(n36289), .Z(n28300) );
  AND U38553 ( .A(\modmult_1/xin[1023] ), .B(n36290), .Z(n36289) );
  IV U38554 ( .A(n36288), .Z(n36290) );
  XOR U38555 ( .A(n36291), .B(mreg[407]), .Z(n36288) );
  NAND U38556 ( .A(n36292), .B(mul_pow), .Z(n36291) );
  XOR U38557 ( .A(mreg[407]), .B(creg[407]), .Z(n36292) );
  XOR U38558 ( .A(n36293), .B(n36294), .Z(n36284) );
  ANDN U38559 ( .A(n36295), .B(n28307), .Z(n36294) );
  XOR U38560 ( .A(n36296), .B(\modmult_1/zin[0][405] ), .Z(n28307) );
  IV U38561 ( .A(n36293), .Z(n36296) );
  XNOR U38562 ( .A(n36293), .B(n28306), .Z(n36295) );
  XOR U38563 ( .A(n36297), .B(n36298), .Z(n28306) );
  AND U38564 ( .A(\modmult_1/xin[1023] ), .B(n36299), .Z(n36298) );
  IV U38565 ( .A(n36297), .Z(n36299) );
  XOR U38566 ( .A(n36300), .B(mreg[406]), .Z(n36297) );
  NAND U38567 ( .A(n36301), .B(mul_pow), .Z(n36300) );
  XOR U38568 ( .A(mreg[406]), .B(creg[406]), .Z(n36301) );
  XOR U38569 ( .A(n36302), .B(n36303), .Z(n36293) );
  ANDN U38570 ( .A(n36304), .B(n28313), .Z(n36303) );
  XOR U38571 ( .A(n36305), .B(\modmult_1/zin[0][404] ), .Z(n28313) );
  IV U38572 ( .A(n36302), .Z(n36305) );
  XNOR U38573 ( .A(n36302), .B(n28312), .Z(n36304) );
  XOR U38574 ( .A(n36306), .B(n36307), .Z(n28312) );
  AND U38575 ( .A(\modmult_1/xin[1023] ), .B(n36308), .Z(n36307) );
  IV U38576 ( .A(n36306), .Z(n36308) );
  XOR U38577 ( .A(n36309), .B(mreg[405]), .Z(n36306) );
  NAND U38578 ( .A(n36310), .B(mul_pow), .Z(n36309) );
  XOR U38579 ( .A(mreg[405]), .B(creg[405]), .Z(n36310) );
  XOR U38580 ( .A(n36311), .B(n36312), .Z(n36302) );
  ANDN U38581 ( .A(n36313), .B(n28319), .Z(n36312) );
  XOR U38582 ( .A(n36314), .B(\modmult_1/zin[0][403] ), .Z(n28319) );
  IV U38583 ( .A(n36311), .Z(n36314) );
  XNOR U38584 ( .A(n36311), .B(n28318), .Z(n36313) );
  XOR U38585 ( .A(n36315), .B(n36316), .Z(n28318) );
  AND U38586 ( .A(\modmult_1/xin[1023] ), .B(n36317), .Z(n36316) );
  IV U38587 ( .A(n36315), .Z(n36317) );
  XOR U38588 ( .A(n36318), .B(mreg[404]), .Z(n36315) );
  NAND U38589 ( .A(n36319), .B(mul_pow), .Z(n36318) );
  XOR U38590 ( .A(mreg[404]), .B(creg[404]), .Z(n36319) );
  XOR U38591 ( .A(n36320), .B(n36321), .Z(n36311) );
  ANDN U38592 ( .A(n36322), .B(n28325), .Z(n36321) );
  XOR U38593 ( .A(n36323), .B(\modmult_1/zin[0][402] ), .Z(n28325) );
  IV U38594 ( .A(n36320), .Z(n36323) );
  XNOR U38595 ( .A(n36320), .B(n28324), .Z(n36322) );
  XOR U38596 ( .A(n36324), .B(n36325), .Z(n28324) );
  AND U38597 ( .A(\modmult_1/xin[1023] ), .B(n36326), .Z(n36325) );
  IV U38598 ( .A(n36324), .Z(n36326) );
  XOR U38599 ( .A(n36327), .B(mreg[403]), .Z(n36324) );
  NAND U38600 ( .A(n36328), .B(mul_pow), .Z(n36327) );
  XOR U38601 ( .A(mreg[403]), .B(creg[403]), .Z(n36328) );
  XOR U38602 ( .A(n36329), .B(n36330), .Z(n36320) );
  ANDN U38603 ( .A(n36331), .B(n28331), .Z(n36330) );
  XOR U38604 ( .A(n36332), .B(\modmult_1/zin[0][401] ), .Z(n28331) );
  IV U38605 ( .A(n36329), .Z(n36332) );
  XNOR U38606 ( .A(n36329), .B(n28330), .Z(n36331) );
  XOR U38607 ( .A(n36333), .B(n36334), .Z(n28330) );
  AND U38608 ( .A(\modmult_1/xin[1023] ), .B(n36335), .Z(n36334) );
  IV U38609 ( .A(n36333), .Z(n36335) );
  XOR U38610 ( .A(n36336), .B(mreg[402]), .Z(n36333) );
  NAND U38611 ( .A(n36337), .B(mul_pow), .Z(n36336) );
  XOR U38612 ( .A(mreg[402]), .B(creg[402]), .Z(n36337) );
  XOR U38613 ( .A(n36338), .B(n36339), .Z(n36329) );
  ANDN U38614 ( .A(n36340), .B(n28337), .Z(n36339) );
  XOR U38615 ( .A(n36341), .B(\modmult_1/zin[0][400] ), .Z(n28337) );
  IV U38616 ( .A(n36338), .Z(n36341) );
  XNOR U38617 ( .A(n36338), .B(n28336), .Z(n36340) );
  XOR U38618 ( .A(n36342), .B(n36343), .Z(n28336) );
  AND U38619 ( .A(\modmult_1/xin[1023] ), .B(n36344), .Z(n36343) );
  IV U38620 ( .A(n36342), .Z(n36344) );
  XOR U38621 ( .A(n36345), .B(mreg[401]), .Z(n36342) );
  NAND U38622 ( .A(n36346), .B(mul_pow), .Z(n36345) );
  XOR U38623 ( .A(mreg[401]), .B(creg[401]), .Z(n36346) );
  XOR U38624 ( .A(n36347), .B(n36348), .Z(n36338) );
  ANDN U38625 ( .A(n36349), .B(n28343), .Z(n36348) );
  XOR U38626 ( .A(n36350), .B(\modmult_1/zin[0][399] ), .Z(n28343) );
  IV U38627 ( .A(n36347), .Z(n36350) );
  XNOR U38628 ( .A(n36347), .B(n28342), .Z(n36349) );
  XOR U38629 ( .A(n36351), .B(n36352), .Z(n28342) );
  AND U38630 ( .A(\modmult_1/xin[1023] ), .B(n36353), .Z(n36352) );
  IV U38631 ( .A(n36351), .Z(n36353) );
  XOR U38632 ( .A(n36354), .B(mreg[400]), .Z(n36351) );
  NAND U38633 ( .A(n36355), .B(mul_pow), .Z(n36354) );
  XOR U38634 ( .A(mreg[400]), .B(creg[400]), .Z(n36355) );
  XOR U38635 ( .A(n36356), .B(n36357), .Z(n36347) );
  ANDN U38636 ( .A(n36358), .B(n28349), .Z(n36357) );
  XOR U38637 ( .A(n36359), .B(\modmult_1/zin[0][398] ), .Z(n28349) );
  IV U38638 ( .A(n36356), .Z(n36359) );
  XNOR U38639 ( .A(n36356), .B(n28348), .Z(n36358) );
  XOR U38640 ( .A(n36360), .B(n36361), .Z(n28348) );
  AND U38641 ( .A(\modmult_1/xin[1023] ), .B(n36362), .Z(n36361) );
  IV U38642 ( .A(n36360), .Z(n36362) );
  XOR U38643 ( .A(n36363), .B(mreg[399]), .Z(n36360) );
  NAND U38644 ( .A(n36364), .B(mul_pow), .Z(n36363) );
  XOR U38645 ( .A(mreg[399]), .B(creg[399]), .Z(n36364) );
  XOR U38646 ( .A(n36365), .B(n36366), .Z(n36356) );
  ANDN U38647 ( .A(n36367), .B(n28355), .Z(n36366) );
  XOR U38648 ( .A(n36368), .B(\modmult_1/zin[0][397] ), .Z(n28355) );
  IV U38649 ( .A(n36365), .Z(n36368) );
  XNOR U38650 ( .A(n36365), .B(n28354), .Z(n36367) );
  XOR U38651 ( .A(n36369), .B(n36370), .Z(n28354) );
  AND U38652 ( .A(\modmult_1/xin[1023] ), .B(n36371), .Z(n36370) );
  IV U38653 ( .A(n36369), .Z(n36371) );
  XOR U38654 ( .A(n36372), .B(mreg[398]), .Z(n36369) );
  NAND U38655 ( .A(n36373), .B(mul_pow), .Z(n36372) );
  XOR U38656 ( .A(mreg[398]), .B(creg[398]), .Z(n36373) );
  XOR U38657 ( .A(n36374), .B(n36375), .Z(n36365) );
  ANDN U38658 ( .A(n36376), .B(n28361), .Z(n36375) );
  XOR U38659 ( .A(n36377), .B(\modmult_1/zin[0][396] ), .Z(n28361) );
  IV U38660 ( .A(n36374), .Z(n36377) );
  XNOR U38661 ( .A(n36374), .B(n28360), .Z(n36376) );
  XOR U38662 ( .A(n36378), .B(n36379), .Z(n28360) );
  AND U38663 ( .A(\modmult_1/xin[1023] ), .B(n36380), .Z(n36379) );
  IV U38664 ( .A(n36378), .Z(n36380) );
  XOR U38665 ( .A(n36381), .B(mreg[397]), .Z(n36378) );
  NAND U38666 ( .A(n36382), .B(mul_pow), .Z(n36381) );
  XOR U38667 ( .A(mreg[397]), .B(creg[397]), .Z(n36382) );
  XOR U38668 ( .A(n36383), .B(n36384), .Z(n36374) );
  ANDN U38669 ( .A(n36385), .B(n28367), .Z(n36384) );
  XOR U38670 ( .A(n36386), .B(\modmult_1/zin[0][395] ), .Z(n28367) );
  IV U38671 ( .A(n36383), .Z(n36386) );
  XNOR U38672 ( .A(n36383), .B(n28366), .Z(n36385) );
  XOR U38673 ( .A(n36387), .B(n36388), .Z(n28366) );
  AND U38674 ( .A(\modmult_1/xin[1023] ), .B(n36389), .Z(n36388) );
  IV U38675 ( .A(n36387), .Z(n36389) );
  XOR U38676 ( .A(n36390), .B(mreg[396]), .Z(n36387) );
  NAND U38677 ( .A(n36391), .B(mul_pow), .Z(n36390) );
  XOR U38678 ( .A(mreg[396]), .B(creg[396]), .Z(n36391) );
  XOR U38679 ( .A(n36392), .B(n36393), .Z(n36383) );
  ANDN U38680 ( .A(n36394), .B(n28373), .Z(n36393) );
  XOR U38681 ( .A(n36395), .B(\modmult_1/zin[0][394] ), .Z(n28373) );
  IV U38682 ( .A(n36392), .Z(n36395) );
  XNOR U38683 ( .A(n36392), .B(n28372), .Z(n36394) );
  XOR U38684 ( .A(n36396), .B(n36397), .Z(n28372) );
  AND U38685 ( .A(\modmult_1/xin[1023] ), .B(n36398), .Z(n36397) );
  IV U38686 ( .A(n36396), .Z(n36398) );
  XOR U38687 ( .A(n36399), .B(mreg[395]), .Z(n36396) );
  NAND U38688 ( .A(n36400), .B(mul_pow), .Z(n36399) );
  XOR U38689 ( .A(mreg[395]), .B(creg[395]), .Z(n36400) );
  XOR U38690 ( .A(n36401), .B(n36402), .Z(n36392) );
  ANDN U38691 ( .A(n36403), .B(n28379), .Z(n36402) );
  XOR U38692 ( .A(n36404), .B(\modmult_1/zin[0][393] ), .Z(n28379) );
  IV U38693 ( .A(n36401), .Z(n36404) );
  XNOR U38694 ( .A(n36401), .B(n28378), .Z(n36403) );
  XOR U38695 ( .A(n36405), .B(n36406), .Z(n28378) );
  AND U38696 ( .A(\modmult_1/xin[1023] ), .B(n36407), .Z(n36406) );
  IV U38697 ( .A(n36405), .Z(n36407) );
  XOR U38698 ( .A(n36408), .B(mreg[394]), .Z(n36405) );
  NAND U38699 ( .A(n36409), .B(mul_pow), .Z(n36408) );
  XOR U38700 ( .A(mreg[394]), .B(creg[394]), .Z(n36409) );
  XOR U38701 ( .A(n36410), .B(n36411), .Z(n36401) );
  ANDN U38702 ( .A(n36412), .B(n28385), .Z(n36411) );
  XOR U38703 ( .A(n36413), .B(\modmult_1/zin[0][392] ), .Z(n28385) );
  IV U38704 ( .A(n36410), .Z(n36413) );
  XNOR U38705 ( .A(n36410), .B(n28384), .Z(n36412) );
  XOR U38706 ( .A(n36414), .B(n36415), .Z(n28384) );
  AND U38707 ( .A(\modmult_1/xin[1023] ), .B(n36416), .Z(n36415) );
  IV U38708 ( .A(n36414), .Z(n36416) );
  XOR U38709 ( .A(n36417), .B(mreg[393]), .Z(n36414) );
  NAND U38710 ( .A(n36418), .B(mul_pow), .Z(n36417) );
  XOR U38711 ( .A(mreg[393]), .B(creg[393]), .Z(n36418) );
  XOR U38712 ( .A(n36419), .B(n36420), .Z(n36410) );
  ANDN U38713 ( .A(n36421), .B(n28391), .Z(n36420) );
  XOR U38714 ( .A(n36422), .B(\modmult_1/zin[0][391] ), .Z(n28391) );
  IV U38715 ( .A(n36419), .Z(n36422) );
  XNOR U38716 ( .A(n36419), .B(n28390), .Z(n36421) );
  XOR U38717 ( .A(n36423), .B(n36424), .Z(n28390) );
  AND U38718 ( .A(\modmult_1/xin[1023] ), .B(n36425), .Z(n36424) );
  IV U38719 ( .A(n36423), .Z(n36425) );
  XOR U38720 ( .A(n36426), .B(mreg[392]), .Z(n36423) );
  NAND U38721 ( .A(n36427), .B(mul_pow), .Z(n36426) );
  XOR U38722 ( .A(mreg[392]), .B(creg[392]), .Z(n36427) );
  XOR U38723 ( .A(n36428), .B(n36429), .Z(n36419) );
  ANDN U38724 ( .A(n36430), .B(n28397), .Z(n36429) );
  XOR U38725 ( .A(n36431), .B(\modmult_1/zin[0][390] ), .Z(n28397) );
  IV U38726 ( .A(n36428), .Z(n36431) );
  XNOR U38727 ( .A(n36428), .B(n28396), .Z(n36430) );
  XOR U38728 ( .A(n36432), .B(n36433), .Z(n28396) );
  AND U38729 ( .A(\modmult_1/xin[1023] ), .B(n36434), .Z(n36433) );
  IV U38730 ( .A(n36432), .Z(n36434) );
  XOR U38731 ( .A(n36435), .B(mreg[391]), .Z(n36432) );
  NAND U38732 ( .A(n36436), .B(mul_pow), .Z(n36435) );
  XOR U38733 ( .A(mreg[391]), .B(creg[391]), .Z(n36436) );
  XOR U38734 ( .A(n36437), .B(n36438), .Z(n36428) );
  ANDN U38735 ( .A(n36439), .B(n28403), .Z(n36438) );
  XOR U38736 ( .A(n36440), .B(\modmult_1/zin[0][389] ), .Z(n28403) );
  IV U38737 ( .A(n36437), .Z(n36440) );
  XNOR U38738 ( .A(n36437), .B(n28402), .Z(n36439) );
  XOR U38739 ( .A(n36441), .B(n36442), .Z(n28402) );
  AND U38740 ( .A(\modmult_1/xin[1023] ), .B(n36443), .Z(n36442) );
  IV U38741 ( .A(n36441), .Z(n36443) );
  XOR U38742 ( .A(n36444), .B(mreg[390]), .Z(n36441) );
  NAND U38743 ( .A(n36445), .B(mul_pow), .Z(n36444) );
  XOR U38744 ( .A(mreg[390]), .B(creg[390]), .Z(n36445) );
  XOR U38745 ( .A(n36446), .B(n36447), .Z(n36437) );
  ANDN U38746 ( .A(n36448), .B(n28409), .Z(n36447) );
  XOR U38747 ( .A(n36449), .B(\modmult_1/zin[0][388] ), .Z(n28409) );
  IV U38748 ( .A(n36446), .Z(n36449) );
  XNOR U38749 ( .A(n36446), .B(n28408), .Z(n36448) );
  XOR U38750 ( .A(n36450), .B(n36451), .Z(n28408) );
  AND U38751 ( .A(\modmult_1/xin[1023] ), .B(n36452), .Z(n36451) );
  IV U38752 ( .A(n36450), .Z(n36452) );
  XOR U38753 ( .A(n36453), .B(mreg[389]), .Z(n36450) );
  NAND U38754 ( .A(n36454), .B(mul_pow), .Z(n36453) );
  XOR U38755 ( .A(mreg[389]), .B(creg[389]), .Z(n36454) );
  XOR U38756 ( .A(n36455), .B(n36456), .Z(n36446) );
  ANDN U38757 ( .A(n36457), .B(n28415), .Z(n36456) );
  XOR U38758 ( .A(n36458), .B(\modmult_1/zin[0][387] ), .Z(n28415) );
  IV U38759 ( .A(n36455), .Z(n36458) );
  XNOR U38760 ( .A(n36455), .B(n28414), .Z(n36457) );
  XOR U38761 ( .A(n36459), .B(n36460), .Z(n28414) );
  AND U38762 ( .A(\modmult_1/xin[1023] ), .B(n36461), .Z(n36460) );
  IV U38763 ( .A(n36459), .Z(n36461) );
  XOR U38764 ( .A(n36462), .B(mreg[388]), .Z(n36459) );
  NAND U38765 ( .A(n36463), .B(mul_pow), .Z(n36462) );
  XOR U38766 ( .A(mreg[388]), .B(creg[388]), .Z(n36463) );
  XOR U38767 ( .A(n36464), .B(n36465), .Z(n36455) );
  ANDN U38768 ( .A(n36466), .B(n28421), .Z(n36465) );
  XOR U38769 ( .A(n36467), .B(\modmult_1/zin[0][386] ), .Z(n28421) );
  IV U38770 ( .A(n36464), .Z(n36467) );
  XNOR U38771 ( .A(n36464), .B(n28420), .Z(n36466) );
  XOR U38772 ( .A(n36468), .B(n36469), .Z(n28420) );
  AND U38773 ( .A(\modmult_1/xin[1023] ), .B(n36470), .Z(n36469) );
  IV U38774 ( .A(n36468), .Z(n36470) );
  XOR U38775 ( .A(n36471), .B(mreg[387]), .Z(n36468) );
  NAND U38776 ( .A(n36472), .B(mul_pow), .Z(n36471) );
  XOR U38777 ( .A(mreg[387]), .B(creg[387]), .Z(n36472) );
  XOR U38778 ( .A(n36473), .B(n36474), .Z(n36464) );
  ANDN U38779 ( .A(n36475), .B(n28427), .Z(n36474) );
  XOR U38780 ( .A(n36476), .B(\modmult_1/zin[0][385] ), .Z(n28427) );
  IV U38781 ( .A(n36473), .Z(n36476) );
  XNOR U38782 ( .A(n36473), .B(n28426), .Z(n36475) );
  XOR U38783 ( .A(n36477), .B(n36478), .Z(n28426) );
  AND U38784 ( .A(\modmult_1/xin[1023] ), .B(n36479), .Z(n36478) );
  IV U38785 ( .A(n36477), .Z(n36479) );
  XOR U38786 ( .A(n36480), .B(mreg[386]), .Z(n36477) );
  NAND U38787 ( .A(n36481), .B(mul_pow), .Z(n36480) );
  XOR U38788 ( .A(mreg[386]), .B(creg[386]), .Z(n36481) );
  XOR U38789 ( .A(n36482), .B(n36483), .Z(n36473) );
  ANDN U38790 ( .A(n36484), .B(n28433), .Z(n36483) );
  XOR U38791 ( .A(n36485), .B(\modmult_1/zin[0][384] ), .Z(n28433) );
  IV U38792 ( .A(n36482), .Z(n36485) );
  XNOR U38793 ( .A(n36482), .B(n28432), .Z(n36484) );
  XOR U38794 ( .A(n36486), .B(n36487), .Z(n28432) );
  AND U38795 ( .A(\modmult_1/xin[1023] ), .B(n36488), .Z(n36487) );
  IV U38796 ( .A(n36486), .Z(n36488) );
  XOR U38797 ( .A(n36489), .B(mreg[385]), .Z(n36486) );
  NAND U38798 ( .A(n36490), .B(mul_pow), .Z(n36489) );
  XOR U38799 ( .A(mreg[385]), .B(creg[385]), .Z(n36490) );
  XOR U38800 ( .A(n36491), .B(n36492), .Z(n36482) );
  ANDN U38801 ( .A(n36493), .B(n28439), .Z(n36492) );
  XOR U38802 ( .A(n36494), .B(\modmult_1/zin[0][383] ), .Z(n28439) );
  IV U38803 ( .A(n36491), .Z(n36494) );
  XNOR U38804 ( .A(n36491), .B(n28438), .Z(n36493) );
  XOR U38805 ( .A(n36495), .B(n36496), .Z(n28438) );
  AND U38806 ( .A(\modmult_1/xin[1023] ), .B(n36497), .Z(n36496) );
  IV U38807 ( .A(n36495), .Z(n36497) );
  XOR U38808 ( .A(n36498), .B(mreg[384]), .Z(n36495) );
  NAND U38809 ( .A(n36499), .B(mul_pow), .Z(n36498) );
  XOR U38810 ( .A(mreg[384]), .B(creg[384]), .Z(n36499) );
  XOR U38811 ( .A(n36500), .B(n36501), .Z(n36491) );
  ANDN U38812 ( .A(n36502), .B(n28445), .Z(n36501) );
  XOR U38813 ( .A(n36503), .B(\modmult_1/zin[0][382] ), .Z(n28445) );
  IV U38814 ( .A(n36500), .Z(n36503) );
  XNOR U38815 ( .A(n36500), .B(n28444), .Z(n36502) );
  XOR U38816 ( .A(n36504), .B(n36505), .Z(n28444) );
  AND U38817 ( .A(\modmult_1/xin[1023] ), .B(n36506), .Z(n36505) );
  IV U38818 ( .A(n36504), .Z(n36506) );
  XOR U38819 ( .A(n36507), .B(mreg[383]), .Z(n36504) );
  NAND U38820 ( .A(n36508), .B(mul_pow), .Z(n36507) );
  XOR U38821 ( .A(mreg[383]), .B(creg[383]), .Z(n36508) );
  XOR U38822 ( .A(n36509), .B(n36510), .Z(n36500) );
  ANDN U38823 ( .A(n36511), .B(n28451), .Z(n36510) );
  XOR U38824 ( .A(n36512), .B(\modmult_1/zin[0][381] ), .Z(n28451) );
  IV U38825 ( .A(n36509), .Z(n36512) );
  XNOR U38826 ( .A(n36509), .B(n28450), .Z(n36511) );
  XOR U38827 ( .A(n36513), .B(n36514), .Z(n28450) );
  AND U38828 ( .A(\modmult_1/xin[1023] ), .B(n36515), .Z(n36514) );
  IV U38829 ( .A(n36513), .Z(n36515) );
  XOR U38830 ( .A(n36516), .B(mreg[382]), .Z(n36513) );
  NAND U38831 ( .A(n36517), .B(mul_pow), .Z(n36516) );
  XOR U38832 ( .A(mreg[382]), .B(creg[382]), .Z(n36517) );
  XOR U38833 ( .A(n36518), .B(n36519), .Z(n36509) );
  ANDN U38834 ( .A(n36520), .B(n28457), .Z(n36519) );
  XOR U38835 ( .A(n36521), .B(\modmult_1/zin[0][380] ), .Z(n28457) );
  IV U38836 ( .A(n36518), .Z(n36521) );
  XNOR U38837 ( .A(n36518), .B(n28456), .Z(n36520) );
  XOR U38838 ( .A(n36522), .B(n36523), .Z(n28456) );
  AND U38839 ( .A(\modmult_1/xin[1023] ), .B(n36524), .Z(n36523) );
  IV U38840 ( .A(n36522), .Z(n36524) );
  XOR U38841 ( .A(n36525), .B(mreg[381]), .Z(n36522) );
  NAND U38842 ( .A(n36526), .B(mul_pow), .Z(n36525) );
  XOR U38843 ( .A(mreg[381]), .B(creg[381]), .Z(n36526) );
  XOR U38844 ( .A(n36527), .B(n36528), .Z(n36518) );
  ANDN U38845 ( .A(n36529), .B(n28463), .Z(n36528) );
  XOR U38846 ( .A(n36530), .B(\modmult_1/zin[0][379] ), .Z(n28463) );
  IV U38847 ( .A(n36527), .Z(n36530) );
  XNOR U38848 ( .A(n36527), .B(n28462), .Z(n36529) );
  XOR U38849 ( .A(n36531), .B(n36532), .Z(n28462) );
  AND U38850 ( .A(\modmult_1/xin[1023] ), .B(n36533), .Z(n36532) );
  IV U38851 ( .A(n36531), .Z(n36533) );
  XOR U38852 ( .A(n36534), .B(mreg[380]), .Z(n36531) );
  NAND U38853 ( .A(n36535), .B(mul_pow), .Z(n36534) );
  XOR U38854 ( .A(mreg[380]), .B(creg[380]), .Z(n36535) );
  XOR U38855 ( .A(n36536), .B(n36537), .Z(n36527) );
  ANDN U38856 ( .A(n36538), .B(n28469), .Z(n36537) );
  XOR U38857 ( .A(n36539), .B(\modmult_1/zin[0][378] ), .Z(n28469) );
  IV U38858 ( .A(n36536), .Z(n36539) );
  XNOR U38859 ( .A(n36536), .B(n28468), .Z(n36538) );
  XOR U38860 ( .A(n36540), .B(n36541), .Z(n28468) );
  AND U38861 ( .A(\modmult_1/xin[1023] ), .B(n36542), .Z(n36541) );
  IV U38862 ( .A(n36540), .Z(n36542) );
  XOR U38863 ( .A(n36543), .B(mreg[379]), .Z(n36540) );
  NAND U38864 ( .A(n36544), .B(mul_pow), .Z(n36543) );
  XOR U38865 ( .A(mreg[379]), .B(creg[379]), .Z(n36544) );
  XOR U38866 ( .A(n36545), .B(n36546), .Z(n36536) );
  ANDN U38867 ( .A(n36547), .B(n28475), .Z(n36546) );
  XOR U38868 ( .A(n36548), .B(\modmult_1/zin[0][377] ), .Z(n28475) );
  IV U38869 ( .A(n36545), .Z(n36548) );
  XNOR U38870 ( .A(n36545), .B(n28474), .Z(n36547) );
  XOR U38871 ( .A(n36549), .B(n36550), .Z(n28474) );
  AND U38872 ( .A(\modmult_1/xin[1023] ), .B(n36551), .Z(n36550) );
  IV U38873 ( .A(n36549), .Z(n36551) );
  XOR U38874 ( .A(n36552), .B(mreg[378]), .Z(n36549) );
  NAND U38875 ( .A(n36553), .B(mul_pow), .Z(n36552) );
  XOR U38876 ( .A(mreg[378]), .B(creg[378]), .Z(n36553) );
  XOR U38877 ( .A(n36554), .B(n36555), .Z(n36545) );
  ANDN U38878 ( .A(n36556), .B(n28481), .Z(n36555) );
  XOR U38879 ( .A(n36557), .B(\modmult_1/zin[0][376] ), .Z(n28481) );
  IV U38880 ( .A(n36554), .Z(n36557) );
  XNOR U38881 ( .A(n36554), .B(n28480), .Z(n36556) );
  XOR U38882 ( .A(n36558), .B(n36559), .Z(n28480) );
  AND U38883 ( .A(\modmult_1/xin[1023] ), .B(n36560), .Z(n36559) );
  IV U38884 ( .A(n36558), .Z(n36560) );
  XOR U38885 ( .A(n36561), .B(mreg[377]), .Z(n36558) );
  NAND U38886 ( .A(n36562), .B(mul_pow), .Z(n36561) );
  XOR U38887 ( .A(mreg[377]), .B(creg[377]), .Z(n36562) );
  XOR U38888 ( .A(n36563), .B(n36564), .Z(n36554) );
  ANDN U38889 ( .A(n36565), .B(n28487), .Z(n36564) );
  XOR U38890 ( .A(n36566), .B(\modmult_1/zin[0][375] ), .Z(n28487) );
  IV U38891 ( .A(n36563), .Z(n36566) );
  XNOR U38892 ( .A(n36563), .B(n28486), .Z(n36565) );
  XOR U38893 ( .A(n36567), .B(n36568), .Z(n28486) );
  AND U38894 ( .A(\modmult_1/xin[1023] ), .B(n36569), .Z(n36568) );
  IV U38895 ( .A(n36567), .Z(n36569) );
  XOR U38896 ( .A(n36570), .B(mreg[376]), .Z(n36567) );
  NAND U38897 ( .A(n36571), .B(mul_pow), .Z(n36570) );
  XOR U38898 ( .A(mreg[376]), .B(creg[376]), .Z(n36571) );
  XOR U38899 ( .A(n36572), .B(n36573), .Z(n36563) );
  ANDN U38900 ( .A(n36574), .B(n28493), .Z(n36573) );
  XOR U38901 ( .A(n36575), .B(\modmult_1/zin[0][374] ), .Z(n28493) );
  IV U38902 ( .A(n36572), .Z(n36575) );
  XNOR U38903 ( .A(n36572), .B(n28492), .Z(n36574) );
  XOR U38904 ( .A(n36576), .B(n36577), .Z(n28492) );
  AND U38905 ( .A(\modmult_1/xin[1023] ), .B(n36578), .Z(n36577) );
  IV U38906 ( .A(n36576), .Z(n36578) );
  XOR U38907 ( .A(n36579), .B(mreg[375]), .Z(n36576) );
  NAND U38908 ( .A(n36580), .B(mul_pow), .Z(n36579) );
  XOR U38909 ( .A(mreg[375]), .B(creg[375]), .Z(n36580) );
  XOR U38910 ( .A(n36581), .B(n36582), .Z(n36572) );
  ANDN U38911 ( .A(n36583), .B(n28499), .Z(n36582) );
  XOR U38912 ( .A(n36584), .B(\modmult_1/zin[0][373] ), .Z(n28499) );
  IV U38913 ( .A(n36581), .Z(n36584) );
  XNOR U38914 ( .A(n36581), .B(n28498), .Z(n36583) );
  XOR U38915 ( .A(n36585), .B(n36586), .Z(n28498) );
  AND U38916 ( .A(\modmult_1/xin[1023] ), .B(n36587), .Z(n36586) );
  IV U38917 ( .A(n36585), .Z(n36587) );
  XOR U38918 ( .A(n36588), .B(mreg[374]), .Z(n36585) );
  NAND U38919 ( .A(n36589), .B(mul_pow), .Z(n36588) );
  XOR U38920 ( .A(mreg[374]), .B(creg[374]), .Z(n36589) );
  XOR U38921 ( .A(n36590), .B(n36591), .Z(n36581) );
  ANDN U38922 ( .A(n36592), .B(n28505), .Z(n36591) );
  XOR U38923 ( .A(n36593), .B(\modmult_1/zin[0][372] ), .Z(n28505) );
  IV U38924 ( .A(n36590), .Z(n36593) );
  XNOR U38925 ( .A(n36590), .B(n28504), .Z(n36592) );
  XOR U38926 ( .A(n36594), .B(n36595), .Z(n28504) );
  AND U38927 ( .A(\modmult_1/xin[1023] ), .B(n36596), .Z(n36595) );
  IV U38928 ( .A(n36594), .Z(n36596) );
  XOR U38929 ( .A(n36597), .B(mreg[373]), .Z(n36594) );
  NAND U38930 ( .A(n36598), .B(mul_pow), .Z(n36597) );
  XOR U38931 ( .A(mreg[373]), .B(creg[373]), .Z(n36598) );
  XOR U38932 ( .A(n36599), .B(n36600), .Z(n36590) );
  ANDN U38933 ( .A(n36601), .B(n28511), .Z(n36600) );
  XOR U38934 ( .A(n36602), .B(\modmult_1/zin[0][371] ), .Z(n28511) );
  IV U38935 ( .A(n36599), .Z(n36602) );
  XNOR U38936 ( .A(n36599), .B(n28510), .Z(n36601) );
  XOR U38937 ( .A(n36603), .B(n36604), .Z(n28510) );
  AND U38938 ( .A(\modmult_1/xin[1023] ), .B(n36605), .Z(n36604) );
  IV U38939 ( .A(n36603), .Z(n36605) );
  XOR U38940 ( .A(n36606), .B(mreg[372]), .Z(n36603) );
  NAND U38941 ( .A(n36607), .B(mul_pow), .Z(n36606) );
  XOR U38942 ( .A(mreg[372]), .B(creg[372]), .Z(n36607) );
  XOR U38943 ( .A(n36608), .B(n36609), .Z(n36599) );
  ANDN U38944 ( .A(n36610), .B(n28517), .Z(n36609) );
  XOR U38945 ( .A(n36611), .B(\modmult_1/zin[0][370] ), .Z(n28517) );
  IV U38946 ( .A(n36608), .Z(n36611) );
  XNOR U38947 ( .A(n36608), .B(n28516), .Z(n36610) );
  XOR U38948 ( .A(n36612), .B(n36613), .Z(n28516) );
  AND U38949 ( .A(\modmult_1/xin[1023] ), .B(n36614), .Z(n36613) );
  IV U38950 ( .A(n36612), .Z(n36614) );
  XOR U38951 ( .A(n36615), .B(mreg[371]), .Z(n36612) );
  NAND U38952 ( .A(n36616), .B(mul_pow), .Z(n36615) );
  XOR U38953 ( .A(mreg[371]), .B(creg[371]), .Z(n36616) );
  XOR U38954 ( .A(n36617), .B(n36618), .Z(n36608) );
  ANDN U38955 ( .A(n36619), .B(n28523), .Z(n36618) );
  XOR U38956 ( .A(n36620), .B(\modmult_1/zin[0][369] ), .Z(n28523) );
  IV U38957 ( .A(n36617), .Z(n36620) );
  XNOR U38958 ( .A(n36617), .B(n28522), .Z(n36619) );
  XOR U38959 ( .A(n36621), .B(n36622), .Z(n28522) );
  AND U38960 ( .A(\modmult_1/xin[1023] ), .B(n36623), .Z(n36622) );
  IV U38961 ( .A(n36621), .Z(n36623) );
  XOR U38962 ( .A(n36624), .B(mreg[370]), .Z(n36621) );
  NAND U38963 ( .A(n36625), .B(mul_pow), .Z(n36624) );
  XOR U38964 ( .A(mreg[370]), .B(creg[370]), .Z(n36625) );
  XOR U38965 ( .A(n36626), .B(n36627), .Z(n36617) );
  ANDN U38966 ( .A(n36628), .B(n28529), .Z(n36627) );
  XOR U38967 ( .A(n36629), .B(\modmult_1/zin[0][368] ), .Z(n28529) );
  IV U38968 ( .A(n36626), .Z(n36629) );
  XNOR U38969 ( .A(n36626), .B(n28528), .Z(n36628) );
  XOR U38970 ( .A(n36630), .B(n36631), .Z(n28528) );
  AND U38971 ( .A(\modmult_1/xin[1023] ), .B(n36632), .Z(n36631) );
  IV U38972 ( .A(n36630), .Z(n36632) );
  XOR U38973 ( .A(n36633), .B(mreg[369]), .Z(n36630) );
  NAND U38974 ( .A(n36634), .B(mul_pow), .Z(n36633) );
  XOR U38975 ( .A(mreg[369]), .B(creg[369]), .Z(n36634) );
  XOR U38976 ( .A(n36635), .B(n36636), .Z(n36626) );
  ANDN U38977 ( .A(n36637), .B(n28535), .Z(n36636) );
  XOR U38978 ( .A(n36638), .B(\modmult_1/zin[0][367] ), .Z(n28535) );
  IV U38979 ( .A(n36635), .Z(n36638) );
  XNOR U38980 ( .A(n36635), .B(n28534), .Z(n36637) );
  XOR U38981 ( .A(n36639), .B(n36640), .Z(n28534) );
  AND U38982 ( .A(\modmult_1/xin[1023] ), .B(n36641), .Z(n36640) );
  IV U38983 ( .A(n36639), .Z(n36641) );
  XOR U38984 ( .A(n36642), .B(mreg[368]), .Z(n36639) );
  NAND U38985 ( .A(n36643), .B(mul_pow), .Z(n36642) );
  XOR U38986 ( .A(mreg[368]), .B(creg[368]), .Z(n36643) );
  XOR U38987 ( .A(n36644), .B(n36645), .Z(n36635) );
  ANDN U38988 ( .A(n36646), .B(n28541), .Z(n36645) );
  XOR U38989 ( .A(n36647), .B(\modmult_1/zin[0][366] ), .Z(n28541) );
  IV U38990 ( .A(n36644), .Z(n36647) );
  XNOR U38991 ( .A(n36644), .B(n28540), .Z(n36646) );
  XOR U38992 ( .A(n36648), .B(n36649), .Z(n28540) );
  AND U38993 ( .A(\modmult_1/xin[1023] ), .B(n36650), .Z(n36649) );
  IV U38994 ( .A(n36648), .Z(n36650) );
  XOR U38995 ( .A(n36651), .B(mreg[367]), .Z(n36648) );
  NAND U38996 ( .A(n36652), .B(mul_pow), .Z(n36651) );
  XOR U38997 ( .A(mreg[367]), .B(creg[367]), .Z(n36652) );
  XOR U38998 ( .A(n36653), .B(n36654), .Z(n36644) );
  ANDN U38999 ( .A(n36655), .B(n28547), .Z(n36654) );
  XOR U39000 ( .A(n36656), .B(\modmult_1/zin[0][365] ), .Z(n28547) );
  IV U39001 ( .A(n36653), .Z(n36656) );
  XNOR U39002 ( .A(n36653), .B(n28546), .Z(n36655) );
  XOR U39003 ( .A(n36657), .B(n36658), .Z(n28546) );
  AND U39004 ( .A(\modmult_1/xin[1023] ), .B(n36659), .Z(n36658) );
  IV U39005 ( .A(n36657), .Z(n36659) );
  XOR U39006 ( .A(n36660), .B(mreg[366]), .Z(n36657) );
  NAND U39007 ( .A(n36661), .B(mul_pow), .Z(n36660) );
  XOR U39008 ( .A(mreg[366]), .B(creg[366]), .Z(n36661) );
  XOR U39009 ( .A(n36662), .B(n36663), .Z(n36653) );
  ANDN U39010 ( .A(n36664), .B(n28553), .Z(n36663) );
  XOR U39011 ( .A(n36665), .B(\modmult_1/zin[0][364] ), .Z(n28553) );
  IV U39012 ( .A(n36662), .Z(n36665) );
  XNOR U39013 ( .A(n36662), .B(n28552), .Z(n36664) );
  XOR U39014 ( .A(n36666), .B(n36667), .Z(n28552) );
  AND U39015 ( .A(\modmult_1/xin[1023] ), .B(n36668), .Z(n36667) );
  IV U39016 ( .A(n36666), .Z(n36668) );
  XOR U39017 ( .A(n36669), .B(mreg[365]), .Z(n36666) );
  NAND U39018 ( .A(n36670), .B(mul_pow), .Z(n36669) );
  XOR U39019 ( .A(mreg[365]), .B(creg[365]), .Z(n36670) );
  XOR U39020 ( .A(n36671), .B(n36672), .Z(n36662) );
  ANDN U39021 ( .A(n36673), .B(n28559), .Z(n36672) );
  XOR U39022 ( .A(n36674), .B(\modmult_1/zin[0][363] ), .Z(n28559) );
  IV U39023 ( .A(n36671), .Z(n36674) );
  XNOR U39024 ( .A(n36671), .B(n28558), .Z(n36673) );
  XOR U39025 ( .A(n36675), .B(n36676), .Z(n28558) );
  AND U39026 ( .A(\modmult_1/xin[1023] ), .B(n36677), .Z(n36676) );
  IV U39027 ( .A(n36675), .Z(n36677) );
  XOR U39028 ( .A(n36678), .B(mreg[364]), .Z(n36675) );
  NAND U39029 ( .A(n36679), .B(mul_pow), .Z(n36678) );
  XOR U39030 ( .A(mreg[364]), .B(creg[364]), .Z(n36679) );
  XOR U39031 ( .A(n36680), .B(n36681), .Z(n36671) );
  ANDN U39032 ( .A(n36682), .B(n28565), .Z(n36681) );
  XOR U39033 ( .A(n36683), .B(\modmult_1/zin[0][362] ), .Z(n28565) );
  IV U39034 ( .A(n36680), .Z(n36683) );
  XNOR U39035 ( .A(n36680), .B(n28564), .Z(n36682) );
  XOR U39036 ( .A(n36684), .B(n36685), .Z(n28564) );
  AND U39037 ( .A(\modmult_1/xin[1023] ), .B(n36686), .Z(n36685) );
  IV U39038 ( .A(n36684), .Z(n36686) );
  XOR U39039 ( .A(n36687), .B(mreg[363]), .Z(n36684) );
  NAND U39040 ( .A(n36688), .B(mul_pow), .Z(n36687) );
  XOR U39041 ( .A(mreg[363]), .B(creg[363]), .Z(n36688) );
  XOR U39042 ( .A(n36689), .B(n36690), .Z(n36680) );
  ANDN U39043 ( .A(n36691), .B(n28571), .Z(n36690) );
  XOR U39044 ( .A(n36692), .B(\modmult_1/zin[0][361] ), .Z(n28571) );
  IV U39045 ( .A(n36689), .Z(n36692) );
  XNOR U39046 ( .A(n36689), .B(n28570), .Z(n36691) );
  XOR U39047 ( .A(n36693), .B(n36694), .Z(n28570) );
  AND U39048 ( .A(\modmult_1/xin[1023] ), .B(n36695), .Z(n36694) );
  IV U39049 ( .A(n36693), .Z(n36695) );
  XOR U39050 ( .A(n36696), .B(mreg[362]), .Z(n36693) );
  NAND U39051 ( .A(n36697), .B(mul_pow), .Z(n36696) );
  XOR U39052 ( .A(mreg[362]), .B(creg[362]), .Z(n36697) );
  XOR U39053 ( .A(n36698), .B(n36699), .Z(n36689) );
  ANDN U39054 ( .A(n36700), .B(n28577), .Z(n36699) );
  XOR U39055 ( .A(n36701), .B(\modmult_1/zin[0][360] ), .Z(n28577) );
  IV U39056 ( .A(n36698), .Z(n36701) );
  XNOR U39057 ( .A(n36698), .B(n28576), .Z(n36700) );
  XOR U39058 ( .A(n36702), .B(n36703), .Z(n28576) );
  AND U39059 ( .A(\modmult_1/xin[1023] ), .B(n36704), .Z(n36703) );
  IV U39060 ( .A(n36702), .Z(n36704) );
  XOR U39061 ( .A(n36705), .B(mreg[361]), .Z(n36702) );
  NAND U39062 ( .A(n36706), .B(mul_pow), .Z(n36705) );
  XOR U39063 ( .A(mreg[361]), .B(creg[361]), .Z(n36706) );
  XOR U39064 ( .A(n36707), .B(n36708), .Z(n36698) );
  ANDN U39065 ( .A(n36709), .B(n28583), .Z(n36708) );
  XOR U39066 ( .A(n36710), .B(\modmult_1/zin[0][359] ), .Z(n28583) );
  IV U39067 ( .A(n36707), .Z(n36710) );
  XNOR U39068 ( .A(n36707), .B(n28582), .Z(n36709) );
  XOR U39069 ( .A(n36711), .B(n36712), .Z(n28582) );
  AND U39070 ( .A(\modmult_1/xin[1023] ), .B(n36713), .Z(n36712) );
  IV U39071 ( .A(n36711), .Z(n36713) );
  XOR U39072 ( .A(n36714), .B(mreg[360]), .Z(n36711) );
  NAND U39073 ( .A(n36715), .B(mul_pow), .Z(n36714) );
  XOR U39074 ( .A(mreg[360]), .B(creg[360]), .Z(n36715) );
  XOR U39075 ( .A(n36716), .B(n36717), .Z(n36707) );
  ANDN U39076 ( .A(n36718), .B(n28589), .Z(n36717) );
  XOR U39077 ( .A(n36719), .B(\modmult_1/zin[0][358] ), .Z(n28589) );
  IV U39078 ( .A(n36716), .Z(n36719) );
  XNOR U39079 ( .A(n36716), .B(n28588), .Z(n36718) );
  XOR U39080 ( .A(n36720), .B(n36721), .Z(n28588) );
  AND U39081 ( .A(\modmult_1/xin[1023] ), .B(n36722), .Z(n36721) );
  IV U39082 ( .A(n36720), .Z(n36722) );
  XOR U39083 ( .A(n36723), .B(mreg[359]), .Z(n36720) );
  NAND U39084 ( .A(n36724), .B(mul_pow), .Z(n36723) );
  XOR U39085 ( .A(mreg[359]), .B(creg[359]), .Z(n36724) );
  XOR U39086 ( .A(n36725), .B(n36726), .Z(n36716) );
  ANDN U39087 ( .A(n36727), .B(n28595), .Z(n36726) );
  XOR U39088 ( .A(n36728), .B(\modmult_1/zin[0][357] ), .Z(n28595) );
  IV U39089 ( .A(n36725), .Z(n36728) );
  XNOR U39090 ( .A(n36725), .B(n28594), .Z(n36727) );
  XOR U39091 ( .A(n36729), .B(n36730), .Z(n28594) );
  AND U39092 ( .A(\modmult_1/xin[1023] ), .B(n36731), .Z(n36730) );
  IV U39093 ( .A(n36729), .Z(n36731) );
  XOR U39094 ( .A(n36732), .B(mreg[358]), .Z(n36729) );
  NAND U39095 ( .A(n36733), .B(mul_pow), .Z(n36732) );
  XOR U39096 ( .A(mreg[358]), .B(creg[358]), .Z(n36733) );
  XOR U39097 ( .A(n36734), .B(n36735), .Z(n36725) );
  ANDN U39098 ( .A(n36736), .B(n28601), .Z(n36735) );
  XOR U39099 ( .A(n36737), .B(\modmult_1/zin[0][356] ), .Z(n28601) );
  IV U39100 ( .A(n36734), .Z(n36737) );
  XNOR U39101 ( .A(n36734), .B(n28600), .Z(n36736) );
  XOR U39102 ( .A(n36738), .B(n36739), .Z(n28600) );
  AND U39103 ( .A(\modmult_1/xin[1023] ), .B(n36740), .Z(n36739) );
  IV U39104 ( .A(n36738), .Z(n36740) );
  XOR U39105 ( .A(n36741), .B(mreg[357]), .Z(n36738) );
  NAND U39106 ( .A(n36742), .B(mul_pow), .Z(n36741) );
  XOR U39107 ( .A(mreg[357]), .B(creg[357]), .Z(n36742) );
  XOR U39108 ( .A(n36743), .B(n36744), .Z(n36734) );
  ANDN U39109 ( .A(n36745), .B(n28607), .Z(n36744) );
  XOR U39110 ( .A(n36746), .B(\modmult_1/zin[0][355] ), .Z(n28607) );
  IV U39111 ( .A(n36743), .Z(n36746) );
  XNOR U39112 ( .A(n36743), .B(n28606), .Z(n36745) );
  XOR U39113 ( .A(n36747), .B(n36748), .Z(n28606) );
  AND U39114 ( .A(\modmult_1/xin[1023] ), .B(n36749), .Z(n36748) );
  IV U39115 ( .A(n36747), .Z(n36749) );
  XOR U39116 ( .A(n36750), .B(mreg[356]), .Z(n36747) );
  NAND U39117 ( .A(n36751), .B(mul_pow), .Z(n36750) );
  XOR U39118 ( .A(mreg[356]), .B(creg[356]), .Z(n36751) );
  XOR U39119 ( .A(n36752), .B(n36753), .Z(n36743) );
  ANDN U39120 ( .A(n36754), .B(n28613), .Z(n36753) );
  XOR U39121 ( .A(n36755), .B(\modmult_1/zin[0][354] ), .Z(n28613) );
  IV U39122 ( .A(n36752), .Z(n36755) );
  XNOR U39123 ( .A(n36752), .B(n28612), .Z(n36754) );
  XOR U39124 ( .A(n36756), .B(n36757), .Z(n28612) );
  AND U39125 ( .A(\modmult_1/xin[1023] ), .B(n36758), .Z(n36757) );
  IV U39126 ( .A(n36756), .Z(n36758) );
  XOR U39127 ( .A(n36759), .B(mreg[355]), .Z(n36756) );
  NAND U39128 ( .A(n36760), .B(mul_pow), .Z(n36759) );
  XOR U39129 ( .A(mreg[355]), .B(creg[355]), .Z(n36760) );
  XOR U39130 ( .A(n36761), .B(n36762), .Z(n36752) );
  ANDN U39131 ( .A(n36763), .B(n28619), .Z(n36762) );
  XOR U39132 ( .A(n36764), .B(\modmult_1/zin[0][353] ), .Z(n28619) );
  IV U39133 ( .A(n36761), .Z(n36764) );
  XNOR U39134 ( .A(n36761), .B(n28618), .Z(n36763) );
  XOR U39135 ( .A(n36765), .B(n36766), .Z(n28618) );
  AND U39136 ( .A(\modmult_1/xin[1023] ), .B(n36767), .Z(n36766) );
  IV U39137 ( .A(n36765), .Z(n36767) );
  XOR U39138 ( .A(n36768), .B(mreg[354]), .Z(n36765) );
  NAND U39139 ( .A(n36769), .B(mul_pow), .Z(n36768) );
  XOR U39140 ( .A(mreg[354]), .B(creg[354]), .Z(n36769) );
  XOR U39141 ( .A(n36770), .B(n36771), .Z(n36761) );
  ANDN U39142 ( .A(n36772), .B(n28625), .Z(n36771) );
  XOR U39143 ( .A(n36773), .B(\modmult_1/zin[0][352] ), .Z(n28625) );
  IV U39144 ( .A(n36770), .Z(n36773) );
  XNOR U39145 ( .A(n36770), .B(n28624), .Z(n36772) );
  XOR U39146 ( .A(n36774), .B(n36775), .Z(n28624) );
  AND U39147 ( .A(\modmult_1/xin[1023] ), .B(n36776), .Z(n36775) );
  IV U39148 ( .A(n36774), .Z(n36776) );
  XOR U39149 ( .A(n36777), .B(mreg[353]), .Z(n36774) );
  NAND U39150 ( .A(n36778), .B(mul_pow), .Z(n36777) );
  XOR U39151 ( .A(mreg[353]), .B(creg[353]), .Z(n36778) );
  XOR U39152 ( .A(n36779), .B(n36780), .Z(n36770) );
  ANDN U39153 ( .A(n36781), .B(n28631), .Z(n36780) );
  XOR U39154 ( .A(n36782), .B(\modmult_1/zin[0][351] ), .Z(n28631) );
  IV U39155 ( .A(n36779), .Z(n36782) );
  XNOR U39156 ( .A(n36779), .B(n28630), .Z(n36781) );
  XOR U39157 ( .A(n36783), .B(n36784), .Z(n28630) );
  AND U39158 ( .A(\modmult_1/xin[1023] ), .B(n36785), .Z(n36784) );
  IV U39159 ( .A(n36783), .Z(n36785) );
  XOR U39160 ( .A(n36786), .B(mreg[352]), .Z(n36783) );
  NAND U39161 ( .A(n36787), .B(mul_pow), .Z(n36786) );
  XOR U39162 ( .A(mreg[352]), .B(creg[352]), .Z(n36787) );
  XOR U39163 ( .A(n36788), .B(n36789), .Z(n36779) );
  ANDN U39164 ( .A(n36790), .B(n28637), .Z(n36789) );
  XOR U39165 ( .A(n36791), .B(\modmult_1/zin[0][350] ), .Z(n28637) );
  IV U39166 ( .A(n36788), .Z(n36791) );
  XNOR U39167 ( .A(n36788), .B(n28636), .Z(n36790) );
  XOR U39168 ( .A(n36792), .B(n36793), .Z(n28636) );
  AND U39169 ( .A(\modmult_1/xin[1023] ), .B(n36794), .Z(n36793) );
  IV U39170 ( .A(n36792), .Z(n36794) );
  XOR U39171 ( .A(n36795), .B(mreg[351]), .Z(n36792) );
  NAND U39172 ( .A(n36796), .B(mul_pow), .Z(n36795) );
  XOR U39173 ( .A(mreg[351]), .B(creg[351]), .Z(n36796) );
  XOR U39174 ( .A(n36797), .B(n36798), .Z(n36788) );
  ANDN U39175 ( .A(n36799), .B(n28643), .Z(n36798) );
  XOR U39176 ( .A(n36800), .B(\modmult_1/zin[0][349] ), .Z(n28643) );
  IV U39177 ( .A(n36797), .Z(n36800) );
  XNOR U39178 ( .A(n36797), .B(n28642), .Z(n36799) );
  XOR U39179 ( .A(n36801), .B(n36802), .Z(n28642) );
  AND U39180 ( .A(\modmult_1/xin[1023] ), .B(n36803), .Z(n36802) );
  IV U39181 ( .A(n36801), .Z(n36803) );
  XOR U39182 ( .A(n36804), .B(mreg[350]), .Z(n36801) );
  NAND U39183 ( .A(n36805), .B(mul_pow), .Z(n36804) );
  XOR U39184 ( .A(mreg[350]), .B(creg[350]), .Z(n36805) );
  XOR U39185 ( .A(n36806), .B(n36807), .Z(n36797) );
  ANDN U39186 ( .A(n36808), .B(n28649), .Z(n36807) );
  XOR U39187 ( .A(n36809), .B(\modmult_1/zin[0][348] ), .Z(n28649) );
  IV U39188 ( .A(n36806), .Z(n36809) );
  XNOR U39189 ( .A(n36806), .B(n28648), .Z(n36808) );
  XOR U39190 ( .A(n36810), .B(n36811), .Z(n28648) );
  AND U39191 ( .A(\modmult_1/xin[1023] ), .B(n36812), .Z(n36811) );
  IV U39192 ( .A(n36810), .Z(n36812) );
  XOR U39193 ( .A(n36813), .B(mreg[349]), .Z(n36810) );
  NAND U39194 ( .A(n36814), .B(mul_pow), .Z(n36813) );
  XOR U39195 ( .A(mreg[349]), .B(creg[349]), .Z(n36814) );
  XOR U39196 ( .A(n36815), .B(n36816), .Z(n36806) );
  ANDN U39197 ( .A(n36817), .B(n28655), .Z(n36816) );
  XOR U39198 ( .A(n36818), .B(\modmult_1/zin[0][347] ), .Z(n28655) );
  IV U39199 ( .A(n36815), .Z(n36818) );
  XNOR U39200 ( .A(n36815), .B(n28654), .Z(n36817) );
  XOR U39201 ( .A(n36819), .B(n36820), .Z(n28654) );
  AND U39202 ( .A(\modmult_1/xin[1023] ), .B(n36821), .Z(n36820) );
  IV U39203 ( .A(n36819), .Z(n36821) );
  XOR U39204 ( .A(n36822), .B(mreg[348]), .Z(n36819) );
  NAND U39205 ( .A(n36823), .B(mul_pow), .Z(n36822) );
  XOR U39206 ( .A(mreg[348]), .B(creg[348]), .Z(n36823) );
  XOR U39207 ( .A(n36824), .B(n36825), .Z(n36815) );
  ANDN U39208 ( .A(n36826), .B(n28661), .Z(n36825) );
  XOR U39209 ( .A(n36827), .B(\modmult_1/zin[0][346] ), .Z(n28661) );
  IV U39210 ( .A(n36824), .Z(n36827) );
  XNOR U39211 ( .A(n36824), .B(n28660), .Z(n36826) );
  XOR U39212 ( .A(n36828), .B(n36829), .Z(n28660) );
  AND U39213 ( .A(\modmult_1/xin[1023] ), .B(n36830), .Z(n36829) );
  IV U39214 ( .A(n36828), .Z(n36830) );
  XOR U39215 ( .A(n36831), .B(mreg[347]), .Z(n36828) );
  NAND U39216 ( .A(n36832), .B(mul_pow), .Z(n36831) );
  XOR U39217 ( .A(mreg[347]), .B(creg[347]), .Z(n36832) );
  XOR U39218 ( .A(n36833), .B(n36834), .Z(n36824) );
  ANDN U39219 ( .A(n36835), .B(n28667), .Z(n36834) );
  XOR U39220 ( .A(n36836), .B(\modmult_1/zin[0][345] ), .Z(n28667) );
  IV U39221 ( .A(n36833), .Z(n36836) );
  XNOR U39222 ( .A(n36833), .B(n28666), .Z(n36835) );
  XOR U39223 ( .A(n36837), .B(n36838), .Z(n28666) );
  AND U39224 ( .A(\modmult_1/xin[1023] ), .B(n36839), .Z(n36838) );
  IV U39225 ( .A(n36837), .Z(n36839) );
  XOR U39226 ( .A(n36840), .B(mreg[346]), .Z(n36837) );
  NAND U39227 ( .A(n36841), .B(mul_pow), .Z(n36840) );
  XOR U39228 ( .A(mreg[346]), .B(creg[346]), .Z(n36841) );
  XOR U39229 ( .A(n36842), .B(n36843), .Z(n36833) );
  ANDN U39230 ( .A(n36844), .B(n28673), .Z(n36843) );
  XOR U39231 ( .A(n36845), .B(\modmult_1/zin[0][344] ), .Z(n28673) );
  IV U39232 ( .A(n36842), .Z(n36845) );
  XNOR U39233 ( .A(n36842), .B(n28672), .Z(n36844) );
  XOR U39234 ( .A(n36846), .B(n36847), .Z(n28672) );
  AND U39235 ( .A(\modmult_1/xin[1023] ), .B(n36848), .Z(n36847) );
  IV U39236 ( .A(n36846), .Z(n36848) );
  XOR U39237 ( .A(n36849), .B(mreg[345]), .Z(n36846) );
  NAND U39238 ( .A(n36850), .B(mul_pow), .Z(n36849) );
  XOR U39239 ( .A(mreg[345]), .B(creg[345]), .Z(n36850) );
  XOR U39240 ( .A(n36851), .B(n36852), .Z(n36842) );
  ANDN U39241 ( .A(n36853), .B(n28679), .Z(n36852) );
  XOR U39242 ( .A(n36854), .B(\modmult_1/zin[0][343] ), .Z(n28679) );
  IV U39243 ( .A(n36851), .Z(n36854) );
  XNOR U39244 ( .A(n36851), .B(n28678), .Z(n36853) );
  XOR U39245 ( .A(n36855), .B(n36856), .Z(n28678) );
  AND U39246 ( .A(\modmult_1/xin[1023] ), .B(n36857), .Z(n36856) );
  IV U39247 ( .A(n36855), .Z(n36857) );
  XOR U39248 ( .A(n36858), .B(mreg[344]), .Z(n36855) );
  NAND U39249 ( .A(n36859), .B(mul_pow), .Z(n36858) );
  XOR U39250 ( .A(mreg[344]), .B(creg[344]), .Z(n36859) );
  XOR U39251 ( .A(n36860), .B(n36861), .Z(n36851) );
  ANDN U39252 ( .A(n36862), .B(n28685), .Z(n36861) );
  XOR U39253 ( .A(n36863), .B(\modmult_1/zin[0][342] ), .Z(n28685) );
  IV U39254 ( .A(n36860), .Z(n36863) );
  XNOR U39255 ( .A(n36860), .B(n28684), .Z(n36862) );
  XOR U39256 ( .A(n36864), .B(n36865), .Z(n28684) );
  AND U39257 ( .A(\modmult_1/xin[1023] ), .B(n36866), .Z(n36865) );
  IV U39258 ( .A(n36864), .Z(n36866) );
  XOR U39259 ( .A(n36867), .B(mreg[343]), .Z(n36864) );
  NAND U39260 ( .A(n36868), .B(mul_pow), .Z(n36867) );
  XOR U39261 ( .A(mreg[343]), .B(creg[343]), .Z(n36868) );
  XOR U39262 ( .A(n36869), .B(n36870), .Z(n36860) );
  ANDN U39263 ( .A(n36871), .B(n28691), .Z(n36870) );
  XOR U39264 ( .A(n36872), .B(\modmult_1/zin[0][341] ), .Z(n28691) );
  IV U39265 ( .A(n36869), .Z(n36872) );
  XNOR U39266 ( .A(n36869), .B(n28690), .Z(n36871) );
  XOR U39267 ( .A(n36873), .B(n36874), .Z(n28690) );
  AND U39268 ( .A(\modmult_1/xin[1023] ), .B(n36875), .Z(n36874) );
  IV U39269 ( .A(n36873), .Z(n36875) );
  XOR U39270 ( .A(n36876), .B(mreg[342]), .Z(n36873) );
  NAND U39271 ( .A(n36877), .B(mul_pow), .Z(n36876) );
  XOR U39272 ( .A(mreg[342]), .B(creg[342]), .Z(n36877) );
  XOR U39273 ( .A(n36878), .B(n36879), .Z(n36869) );
  ANDN U39274 ( .A(n36880), .B(n28697), .Z(n36879) );
  XOR U39275 ( .A(n36881), .B(\modmult_1/zin[0][340] ), .Z(n28697) );
  IV U39276 ( .A(n36878), .Z(n36881) );
  XNOR U39277 ( .A(n36878), .B(n28696), .Z(n36880) );
  XOR U39278 ( .A(n36882), .B(n36883), .Z(n28696) );
  AND U39279 ( .A(\modmult_1/xin[1023] ), .B(n36884), .Z(n36883) );
  IV U39280 ( .A(n36882), .Z(n36884) );
  XOR U39281 ( .A(n36885), .B(mreg[341]), .Z(n36882) );
  NAND U39282 ( .A(n36886), .B(mul_pow), .Z(n36885) );
  XOR U39283 ( .A(mreg[341]), .B(creg[341]), .Z(n36886) );
  XOR U39284 ( .A(n36887), .B(n36888), .Z(n36878) );
  ANDN U39285 ( .A(n36889), .B(n28703), .Z(n36888) );
  XOR U39286 ( .A(n36890), .B(\modmult_1/zin[0][339] ), .Z(n28703) );
  IV U39287 ( .A(n36887), .Z(n36890) );
  XNOR U39288 ( .A(n36887), .B(n28702), .Z(n36889) );
  XOR U39289 ( .A(n36891), .B(n36892), .Z(n28702) );
  AND U39290 ( .A(\modmult_1/xin[1023] ), .B(n36893), .Z(n36892) );
  IV U39291 ( .A(n36891), .Z(n36893) );
  XOR U39292 ( .A(n36894), .B(mreg[340]), .Z(n36891) );
  NAND U39293 ( .A(n36895), .B(mul_pow), .Z(n36894) );
  XOR U39294 ( .A(mreg[340]), .B(creg[340]), .Z(n36895) );
  XOR U39295 ( .A(n36896), .B(n36897), .Z(n36887) );
  ANDN U39296 ( .A(n36898), .B(n28709), .Z(n36897) );
  XOR U39297 ( .A(n36899), .B(\modmult_1/zin[0][338] ), .Z(n28709) );
  IV U39298 ( .A(n36896), .Z(n36899) );
  XNOR U39299 ( .A(n36896), .B(n28708), .Z(n36898) );
  XOR U39300 ( .A(n36900), .B(n36901), .Z(n28708) );
  AND U39301 ( .A(\modmult_1/xin[1023] ), .B(n36902), .Z(n36901) );
  IV U39302 ( .A(n36900), .Z(n36902) );
  XOR U39303 ( .A(n36903), .B(mreg[339]), .Z(n36900) );
  NAND U39304 ( .A(n36904), .B(mul_pow), .Z(n36903) );
  XOR U39305 ( .A(mreg[339]), .B(creg[339]), .Z(n36904) );
  XOR U39306 ( .A(n36905), .B(n36906), .Z(n36896) );
  ANDN U39307 ( .A(n36907), .B(n28715), .Z(n36906) );
  XOR U39308 ( .A(n36908), .B(\modmult_1/zin[0][337] ), .Z(n28715) );
  IV U39309 ( .A(n36905), .Z(n36908) );
  XNOR U39310 ( .A(n36905), .B(n28714), .Z(n36907) );
  XOR U39311 ( .A(n36909), .B(n36910), .Z(n28714) );
  AND U39312 ( .A(\modmult_1/xin[1023] ), .B(n36911), .Z(n36910) );
  IV U39313 ( .A(n36909), .Z(n36911) );
  XOR U39314 ( .A(n36912), .B(mreg[338]), .Z(n36909) );
  NAND U39315 ( .A(n36913), .B(mul_pow), .Z(n36912) );
  XOR U39316 ( .A(mreg[338]), .B(creg[338]), .Z(n36913) );
  XOR U39317 ( .A(n36914), .B(n36915), .Z(n36905) );
  ANDN U39318 ( .A(n36916), .B(n28721), .Z(n36915) );
  XOR U39319 ( .A(n36917), .B(\modmult_1/zin[0][336] ), .Z(n28721) );
  IV U39320 ( .A(n36914), .Z(n36917) );
  XNOR U39321 ( .A(n36914), .B(n28720), .Z(n36916) );
  XOR U39322 ( .A(n36918), .B(n36919), .Z(n28720) );
  AND U39323 ( .A(\modmult_1/xin[1023] ), .B(n36920), .Z(n36919) );
  IV U39324 ( .A(n36918), .Z(n36920) );
  XOR U39325 ( .A(n36921), .B(mreg[337]), .Z(n36918) );
  NAND U39326 ( .A(n36922), .B(mul_pow), .Z(n36921) );
  XOR U39327 ( .A(mreg[337]), .B(creg[337]), .Z(n36922) );
  XOR U39328 ( .A(n36923), .B(n36924), .Z(n36914) );
  ANDN U39329 ( .A(n36925), .B(n28727), .Z(n36924) );
  XOR U39330 ( .A(n36926), .B(\modmult_1/zin[0][335] ), .Z(n28727) );
  IV U39331 ( .A(n36923), .Z(n36926) );
  XNOR U39332 ( .A(n36923), .B(n28726), .Z(n36925) );
  XOR U39333 ( .A(n36927), .B(n36928), .Z(n28726) );
  AND U39334 ( .A(\modmult_1/xin[1023] ), .B(n36929), .Z(n36928) );
  IV U39335 ( .A(n36927), .Z(n36929) );
  XOR U39336 ( .A(n36930), .B(mreg[336]), .Z(n36927) );
  NAND U39337 ( .A(n36931), .B(mul_pow), .Z(n36930) );
  XOR U39338 ( .A(mreg[336]), .B(creg[336]), .Z(n36931) );
  XOR U39339 ( .A(n36932), .B(n36933), .Z(n36923) );
  ANDN U39340 ( .A(n36934), .B(n28733), .Z(n36933) );
  XOR U39341 ( .A(n36935), .B(\modmult_1/zin[0][334] ), .Z(n28733) );
  IV U39342 ( .A(n36932), .Z(n36935) );
  XNOR U39343 ( .A(n36932), .B(n28732), .Z(n36934) );
  XOR U39344 ( .A(n36936), .B(n36937), .Z(n28732) );
  AND U39345 ( .A(\modmult_1/xin[1023] ), .B(n36938), .Z(n36937) );
  IV U39346 ( .A(n36936), .Z(n36938) );
  XOR U39347 ( .A(n36939), .B(mreg[335]), .Z(n36936) );
  NAND U39348 ( .A(n36940), .B(mul_pow), .Z(n36939) );
  XOR U39349 ( .A(mreg[335]), .B(creg[335]), .Z(n36940) );
  XOR U39350 ( .A(n36941), .B(n36942), .Z(n36932) );
  ANDN U39351 ( .A(n36943), .B(n28739), .Z(n36942) );
  XOR U39352 ( .A(n36944), .B(\modmult_1/zin[0][333] ), .Z(n28739) );
  IV U39353 ( .A(n36941), .Z(n36944) );
  XNOR U39354 ( .A(n36941), .B(n28738), .Z(n36943) );
  XOR U39355 ( .A(n36945), .B(n36946), .Z(n28738) );
  AND U39356 ( .A(\modmult_1/xin[1023] ), .B(n36947), .Z(n36946) );
  IV U39357 ( .A(n36945), .Z(n36947) );
  XOR U39358 ( .A(n36948), .B(mreg[334]), .Z(n36945) );
  NAND U39359 ( .A(n36949), .B(mul_pow), .Z(n36948) );
  XOR U39360 ( .A(mreg[334]), .B(creg[334]), .Z(n36949) );
  XOR U39361 ( .A(n36950), .B(n36951), .Z(n36941) );
  ANDN U39362 ( .A(n36952), .B(n28745), .Z(n36951) );
  XOR U39363 ( .A(n36953), .B(\modmult_1/zin[0][332] ), .Z(n28745) );
  IV U39364 ( .A(n36950), .Z(n36953) );
  XNOR U39365 ( .A(n36950), .B(n28744), .Z(n36952) );
  XOR U39366 ( .A(n36954), .B(n36955), .Z(n28744) );
  AND U39367 ( .A(\modmult_1/xin[1023] ), .B(n36956), .Z(n36955) );
  IV U39368 ( .A(n36954), .Z(n36956) );
  XOR U39369 ( .A(n36957), .B(mreg[333]), .Z(n36954) );
  NAND U39370 ( .A(n36958), .B(mul_pow), .Z(n36957) );
  XOR U39371 ( .A(mreg[333]), .B(creg[333]), .Z(n36958) );
  XOR U39372 ( .A(n36959), .B(n36960), .Z(n36950) );
  ANDN U39373 ( .A(n36961), .B(n28751), .Z(n36960) );
  XOR U39374 ( .A(n36962), .B(\modmult_1/zin[0][331] ), .Z(n28751) );
  IV U39375 ( .A(n36959), .Z(n36962) );
  XNOR U39376 ( .A(n36959), .B(n28750), .Z(n36961) );
  XOR U39377 ( .A(n36963), .B(n36964), .Z(n28750) );
  AND U39378 ( .A(\modmult_1/xin[1023] ), .B(n36965), .Z(n36964) );
  IV U39379 ( .A(n36963), .Z(n36965) );
  XOR U39380 ( .A(n36966), .B(mreg[332]), .Z(n36963) );
  NAND U39381 ( .A(n36967), .B(mul_pow), .Z(n36966) );
  XOR U39382 ( .A(mreg[332]), .B(creg[332]), .Z(n36967) );
  XOR U39383 ( .A(n36968), .B(n36969), .Z(n36959) );
  ANDN U39384 ( .A(n36970), .B(n28757), .Z(n36969) );
  XOR U39385 ( .A(n36971), .B(\modmult_1/zin[0][330] ), .Z(n28757) );
  IV U39386 ( .A(n36968), .Z(n36971) );
  XNOR U39387 ( .A(n36968), .B(n28756), .Z(n36970) );
  XOR U39388 ( .A(n36972), .B(n36973), .Z(n28756) );
  AND U39389 ( .A(\modmult_1/xin[1023] ), .B(n36974), .Z(n36973) );
  IV U39390 ( .A(n36972), .Z(n36974) );
  XOR U39391 ( .A(n36975), .B(mreg[331]), .Z(n36972) );
  NAND U39392 ( .A(n36976), .B(mul_pow), .Z(n36975) );
  XOR U39393 ( .A(mreg[331]), .B(creg[331]), .Z(n36976) );
  XOR U39394 ( .A(n36977), .B(n36978), .Z(n36968) );
  ANDN U39395 ( .A(n36979), .B(n28763), .Z(n36978) );
  XOR U39396 ( .A(n36980), .B(\modmult_1/zin[0][329] ), .Z(n28763) );
  IV U39397 ( .A(n36977), .Z(n36980) );
  XNOR U39398 ( .A(n36977), .B(n28762), .Z(n36979) );
  XOR U39399 ( .A(n36981), .B(n36982), .Z(n28762) );
  AND U39400 ( .A(\modmult_1/xin[1023] ), .B(n36983), .Z(n36982) );
  IV U39401 ( .A(n36981), .Z(n36983) );
  XOR U39402 ( .A(n36984), .B(mreg[330]), .Z(n36981) );
  NAND U39403 ( .A(n36985), .B(mul_pow), .Z(n36984) );
  XOR U39404 ( .A(mreg[330]), .B(creg[330]), .Z(n36985) );
  XOR U39405 ( .A(n36986), .B(n36987), .Z(n36977) );
  ANDN U39406 ( .A(n36988), .B(n28769), .Z(n36987) );
  XOR U39407 ( .A(n36989), .B(\modmult_1/zin[0][328] ), .Z(n28769) );
  IV U39408 ( .A(n36986), .Z(n36989) );
  XNOR U39409 ( .A(n36986), .B(n28768), .Z(n36988) );
  XOR U39410 ( .A(n36990), .B(n36991), .Z(n28768) );
  AND U39411 ( .A(\modmult_1/xin[1023] ), .B(n36992), .Z(n36991) );
  IV U39412 ( .A(n36990), .Z(n36992) );
  XOR U39413 ( .A(n36993), .B(mreg[329]), .Z(n36990) );
  NAND U39414 ( .A(n36994), .B(mul_pow), .Z(n36993) );
  XOR U39415 ( .A(mreg[329]), .B(creg[329]), .Z(n36994) );
  XOR U39416 ( .A(n36995), .B(n36996), .Z(n36986) );
  ANDN U39417 ( .A(n36997), .B(n28775), .Z(n36996) );
  XOR U39418 ( .A(n36998), .B(\modmult_1/zin[0][327] ), .Z(n28775) );
  IV U39419 ( .A(n36995), .Z(n36998) );
  XNOR U39420 ( .A(n36995), .B(n28774), .Z(n36997) );
  XOR U39421 ( .A(n36999), .B(n37000), .Z(n28774) );
  AND U39422 ( .A(\modmult_1/xin[1023] ), .B(n37001), .Z(n37000) );
  IV U39423 ( .A(n36999), .Z(n37001) );
  XOR U39424 ( .A(n37002), .B(mreg[328]), .Z(n36999) );
  NAND U39425 ( .A(n37003), .B(mul_pow), .Z(n37002) );
  XOR U39426 ( .A(mreg[328]), .B(creg[328]), .Z(n37003) );
  XOR U39427 ( .A(n37004), .B(n37005), .Z(n36995) );
  ANDN U39428 ( .A(n37006), .B(n28781), .Z(n37005) );
  XOR U39429 ( .A(n37007), .B(\modmult_1/zin[0][326] ), .Z(n28781) );
  IV U39430 ( .A(n37004), .Z(n37007) );
  XNOR U39431 ( .A(n37004), .B(n28780), .Z(n37006) );
  XOR U39432 ( .A(n37008), .B(n37009), .Z(n28780) );
  AND U39433 ( .A(\modmult_1/xin[1023] ), .B(n37010), .Z(n37009) );
  IV U39434 ( .A(n37008), .Z(n37010) );
  XOR U39435 ( .A(n37011), .B(mreg[327]), .Z(n37008) );
  NAND U39436 ( .A(n37012), .B(mul_pow), .Z(n37011) );
  XOR U39437 ( .A(mreg[327]), .B(creg[327]), .Z(n37012) );
  XOR U39438 ( .A(n37013), .B(n37014), .Z(n37004) );
  ANDN U39439 ( .A(n37015), .B(n28787), .Z(n37014) );
  XOR U39440 ( .A(n37016), .B(\modmult_1/zin[0][325] ), .Z(n28787) );
  IV U39441 ( .A(n37013), .Z(n37016) );
  XNOR U39442 ( .A(n37013), .B(n28786), .Z(n37015) );
  XOR U39443 ( .A(n37017), .B(n37018), .Z(n28786) );
  AND U39444 ( .A(\modmult_1/xin[1023] ), .B(n37019), .Z(n37018) );
  IV U39445 ( .A(n37017), .Z(n37019) );
  XOR U39446 ( .A(n37020), .B(mreg[326]), .Z(n37017) );
  NAND U39447 ( .A(n37021), .B(mul_pow), .Z(n37020) );
  XOR U39448 ( .A(mreg[326]), .B(creg[326]), .Z(n37021) );
  XOR U39449 ( .A(n37022), .B(n37023), .Z(n37013) );
  ANDN U39450 ( .A(n37024), .B(n28793), .Z(n37023) );
  XOR U39451 ( .A(n37025), .B(\modmult_1/zin[0][324] ), .Z(n28793) );
  IV U39452 ( .A(n37022), .Z(n37025) );
  XNOR U39453 ( .A(n37022), .B(n28792), .Z(n37024) );
  XOR U39454 ( .A(n37026), .B(n37027), .Z(n28792) );
  AND U39455 ( .A(\modmult_1/xin[1023] ), .B(n37028), .Z(n37027) );
  IV U39456 ( .A(n37026), .Z(n37028) );
  XOR U39457 ( .A(n37029), .B(mreg[325]), .Z(n37026) );
  NAND U39458 ( .A(n37030), .B(mul_pow), .Z(n37029) );
  XOR U39459 ( .A(mreg[325]), .B(creg[325]), .Z(n37030) );
  XOR U39460 ( .A(n37031), .B(n37032), .Z(n37022) );
  ANDN U39461 ( .A(n37033), .B(n28799), .Z(n37032) );
  XOR U39462 ( .A(n37034), .B(\modmult_1/zin[0][323] ), .Z(n28799) );
  IV U39463 ( .A(n37031), .Z(n37034) );
  XNOR U39464 ( .A(n37031), .B(n28798), .Z(n37033) );
  XOR U39465 ( .A(n37035), .B(n37036), .Z(n28798) );
  AND U39466 ( .A(\modmult_1/xin[1023] ), .B(n37037), .Z(n37036) );
  IV U39467 ( .A(n37035), .Z(n37037) );
  XOR U39468 ( .A(n37038), .B(mreg[324]), .Z(n37035) );
  NAND U39469 ( .A(n37039), .B(mul_pow), .Z(n37038) );
  XOR U39470 ( .A(mreg[324]), .B(creg[324]), .Z(n37039) );
  XOR U39471 ( .A(n37040), .B(n37041), .Z(n37031) );
  ANDN U39472 ( .A(n37042), .B(n28805), .Z(n37041) );
  XOR U39473 ( .A(n37043), .B(\modmult_1/zin[0][322] ), .Z(n28805) );
  IV U39474 ( .A(n37040), .Z(n37043) );
  XNOR U39475 ( .A(n37040), .B(n28804), .Z(n37042) );
  XOR U39476 ( .A(n37044), .B(n37045), .Z(n28804) );
  AND U39477 ( .A(\modmult_1/xin[1023] ), .B(n37046), .Z(n37045) );
  IV U39478 ( .A(n37044), .Z(n37046) );
  XOR U39479 ( .A(n37047), .B(mreg[323]), .Z(n37044) );
  NAND U39480 ( .A(n37048), .B(mul_pow), .Z(n37047) );
  XOR U39481 ( .A(mreg[323]), .B(creg[323]), .Z(n37048) );
  XOR U39482 ( .A(n37049), .B(n37050), .Z(n37040) );
  ANDN U39483 ( .A(n37051), .B(n28811), .Z(n37050) );
  XOR U39484 ( .A(n37052), .B(\modmult_1/zin[0][321] ), .Z(n28811) );
  IV U39485 ( .A(n37049), .Z(n37052) );
  XNOR U39486 ( .A(n37049), .B(n28810), .Z(n37051) );
  XOR U39487 ( .A(n37053), .B(n37054), .Z(n28810) );
  AND U39488 ( .A(\modmult_1/xin[1023] ), .B(n37055), .Z(n37054) );
  IV U39489 ( .A(n37053), .Z(n37055) );
  XOR U39490 ( .A(n37056), .B(mreg[322]), .Z(n37053) );
  NAND U39491 ( .A(n37057), .B(mul_pow), .Z(n37056) );
  XOR U39492 ( .A(mreg[322]), .B(creg[322]), .Z(n37057) );
  XOR U39493 ( .A(n37058), .B(n37059), .Z(n37049) );
  ANDN U39494 ( .A(n37060), .B(n28817), .Z(n37059) );
  XOR U39495 ( .A(n37061), .B(\modmult_1/zin[0][320] ), .Z(n28817) );
  IV U39496 ( .A(n37058), .Z(n37061) );
  XNOR U39497 ( .A(n37058), .B(n28816), .Z(n37060) );
  XOR U39498 ( .A(n37062), .B(n37063), .Z(n28816) );
  AND U39499 ( .A(\modmult_1/xin[1023] ), .B(n37064), .Z(n37063) );
  IV U39500 ( .A(n37062), .Z(n37064) );
  XOR U39501 ( .A(n37065), .B(mreg[321]), .Z(n37062) );
  NAND U39502 ( .A(n37066), .B(mul_pow), .Z(n37065) );
  XOR U39503 ( .A(mreg[321]), .B(creg[321]), .Z(n37066) );
  XOR U39504 ( .A(n37067), .B(n37068), .Z(n37058) );
  ANDN U39505 ( .A(n37069), .B(n28823), .Z(n37068) );
  XOR U39506 ( .A(n37070), .B(\modmult_1/zin[0][319] ), .Z(n28823) );
  IV U39507 ( .A(n37067), .Z(n37070) );
  XNOR U39508 ( .A(n37067), .B(n28822), .Z(n37069) );
  XOR U39509 ( .A(n37071), .B(n37072), .Z(n28822) );
  AND U39510 ( .A(\modmult_1/xin[1023] ), .B(n37073), .Z(n37072) );
  IV U39511 ( .A(n37071), .Z(n37073) );
  XOR U39512 ( .A(n37074), .B(mreg[320]), .Z(n37071) );
  NAND U39513 ( .A(n37075), .B(mul_pow), .Z(n37074) );
  XOR U39514 ( .A(mreg[320]), .B(creg[320]), .Z(n37075) );
  XOR U39515 ( .A(n37076), .B(n37077), .Z(n37067) );
  ANDN U39516 ( .A(n37078), .B(n28829), .Z(n37077) );
  XOR U39517 ( .A(n37079), .B(\modmult_1/zin[0][318] ), .Z(n28829) );
  IV U39518 ( .A(n37076), .Z(n37079) );
  XNOR U39519 ( .A(n37076), .B(n28828), .Z(n37078) );
  XOR U39520 ( .A(n37080), .B(n37081), .Z(n28828) );
  AND U39521 ( .A(\modmult_1/xin[1023] ), .B(n37082), .Z(n37081) );
  IV U39522 ( .A(n37080), .Z(n37082) );
  XOR U39523 ( .A(n37083), .B(mreg[319]), .Z(n37080) );
  NAND U39524 ( .A(n37084), .B(mul_pow), .Z(n37083) );
  XOR U39525 ( .A(mreg[319]), .B(creg[319]), .Z(n37084) );
  XOR U39526 ( .A(n37085), .B(n37086), .Z(n37076) );
  ANDN U39527 ( .A(n37087), .B(n28835), .Z(n37086) );
  XOR U39528 ( .A(n37088), .B(\modmult_1/zin[0][317] ), .Z(n28835) );
  IV U39529 ( .A(n37085), .Z(n37088) );
  XNOR U39530 ( .A(n37085), .B(n28834), .Z(n37087) );
  XOR U39531 ( .A(n37089), .B(n37090), .Z(n28834) );
  AND U39532 ( .A(\modmult_1/xin[1023] ), .B(n37091), .Z(n37090) );
  IV U39533 ( .A(n37089), .Z(n37091) );
  XOR U39534 ( .A(n37092), .B(mreg[318]), .Z(n37089) );
  NAND U39535 ( .A(n37093), .B(mul_pow), .Z(n37092) );
  XOR U39536 ( .A(mreg[318]), .B(creg[318]), .Z(n37093) );
  XOR U39537 ( .A(n37094), .B(n37095), .Z(n37085) );
  ANDN U39538 ( .A(n37096), .B(n28841), .Z(n37095) );
  XOR U39539 ( .A(n37097), .B(\modmult_1/zin[0][316] ), .Z(n28841) );
  IV U39540 ( .A(n37094), .Z(n37097) );
  XNOR U39541 ( .A(n37094), .B(n28840), .Z(n37096) );
  XOR U39542 ( .A(n37098), .B(n37099), .Z(n28840) );
  AND U39543 ( .A(\modmult_1/xin[1023] ), .B(n37100), .Z(n37099) );
  IV U39544 ( .A(n37098), .Z(n37100) );
  XOR U39545 ( .A(n37101), .B(mreg[317]), .Z(n37098) );
  NAND U39546 ( .A(n37102), .B(mul_pow), .Z(n37101) );
  XOR U39547 ( .A(mreg[317]), .B(creg[317]), .Z(n37102) );
  XOR U39548 ( .A(n37103), .B(n37104), .Z(n37094) );
  ANDN U39549 ( .A(n37105), .B(n28847), .Z(n37104) );
  XOR U39550 ( .A(n37106), .B(\modmult_1/zin[0][315] ), .Z(n28847) );
  IV U39551 ( .A(n37103), .Z(n37106) );
  XNOR U39552 ( .A(n37103), .B(n28846), .Z(n37105) );
  XOR U39553 ( .A(n37107), .B(n37108), .Z(n28846) );
  AND U39554 ( .A(\modmult_1/xin[1023] ), .B(n37109), .Z(n37108) );
  IV U39555 ( .A(n37107), .Z(n37109) );
  XOR U39556 ( .A(n37110), .B(mreg[316]), .Z(n37107) );
  NAND U39557 ( .A(n37111), .B(mul_pow), .Z(n37110) );
  XOR U39558 ( .A(mreg[316]), .B(creg[316]), .Z(n37111) );
  XOR U39559 ( .A(n37112), .B(n37113), .Z(n37103) );
  ANDN U39560 ( .A(n37114), .B(n28853), .Z(n37113) );
  XOR U39561 ( .A(n37115), .B(\modmult_1/zin[0][314] ), .Z(n28853) );
  IV U39562 ( .A(n37112), .Z(n37115) );
  XNOR U39563 ( .A(n37112), .B(n28852), .Z(n37114) );
  XOR U39564 ( .A(n37116), .B(n37117), .Z(n28852) );
  AND U39565 ( .A(\modmult_1/xin[1023] ), .B(n37118), .Z(n37117) );
  IV U39566 ( .A(n37116), .Z(n37118) );
  XOR U39567 ( .A(n37119), .B(mreg[315]), .Z(n37116) );
  NAND U39568 ( .A(n37120), .B(mul_pow), .Z(n37119) );
  XOR U39569 ( .A(mreg[315]), .B(creg[315]), .Z(n37120) );
  XOR U39570 ( .A(n37121), .B(n37122), .Z(n37112) );
  ANDN U39571 ( .A(n37123), .B(n28859), .Z(n37122) );
  XOR U39572 ( .A(n37124), .B(\modmult_1/zin[0][313] ), .Z(n28859) );
  IV U39573 ( .A(n37121), .Z(n37124) );
  XNOR U39574 ( .A(n37121), .B(n28858), .Z(n37123) );
  XOR U39575 ( .A(n37125), .B(n37126), .Z(n28858) );
  AND U39576 ( .A(\modmult_1/xin[1023] ), .B(n37127), .Z(n37126) );
  IV U39577 ( .A(n37125), .Z(n37127) );
  XOR U39578 ( .A(n37128), .B(mreg[314]), .Z(n37125) );
  NAND U39579 ( .A(n37129), .B(mul_pow), .Z(n37128) );
  XOR U39580 ( .A(mreg[314]), .B(creg[314]), .Z(n37129) );
  XOR U39581 ( .A(n37130), .B(n37131), .Z(n37121) );
  ANDN U39582 ( .A(n37132), .B(n28865), .Z(n37131) );
  XOR U39583 ( .A(n37133), .B(\modmult_1/zin[0][312] ), .Z(n28865) );
  IV U39584 ( .A(n37130), .Z(n37133) );
  XNOR U39585 ( .A(n37130), .B(n28864), .Z(n37132) );
  XOR U39586 ( .A(n37134), .B(n37135), .Z(n28864) );
  AND U39587 ( .A(\modmult_1/xin[1023] ), .B(n37136), .Z(n37135) );
  IV U39588 ( .A(n37134), .Z(n37136) );
  XOR U39589 ( .A(n37137), .B(mreg[313]), .Z(n37134) );
  NAND U39590 ( .A(n37138), .B(mul_pow), .Z(n37137) );
  XOR U39591 ( .A(mreg[313]), .B(creg[313]), .Z(n37138) );
  XOR U39592 ( .A(n37139), .B(n37140), .Z(n37130) );
  ANDN U39593 ( .A(n37141), .B(n28871), .Z(n37140) );
  XOR U39594 ( .A(n37142), .B(\modmult_1/zin[0][311] ), .Z(n28871) );
  IV U39595 ( .A(n37139), .Z(n37142) );
  XNOR U39596 ( .A(n37139), .B(n28870), .Z(n37141) );
  XOR U39597 ( .A(n37143), .B(n37144), .Z(n28870) );
  AND U39598 ( .A(\modmult_1/xin[1023] ), .B(n37145), .Z(n37144) );
  IV U39599 ( .A(n37143), .Z(n37145) );
  XOR U39600 ( .A(n37146), .B(mreg[312]), .Z(n37143) );
  NAND U39601 ( .A(n37147), .B(mul_pow), .Z(n37146) );
  XOR U39602 ( .A(mreg[312]), .B(creg[312]), .Z(n37147) );
  XOR U39603 ( .A(n37148), .B(n37149), .Z(n37139) );
  ANDN U39604 ( .A(n37150), .B(n28877), .Z(n37149) );
  XOR U39605 ( .A(n37151), .B(\modmult_1/zin[0][310] ), .Z(n28877) );
  IV U39606 ( .A(n37148), .Z(n37151) );
  XNOR U39607 ( .A(n37148), .B(n28876), .Z(n37150) );
  XOR U39608 ( .A(n37152), .B(n37153), .Z(n28876) );
  AND U39609 ( .A(\modmult_1/xin[1023] ), .B(n37154), .Z(n37153) );
  IV U39610 ( .A(n37152), .Z(n37154) );
  XOR U39611 ( .A(n37155), .B(mreg[311]), .Z(n37152) );
  NAND U39612 ( .A(n37156), .B(mul_pow), .Z(n37155) );
  XOR U39613 ( .A(mreg[311]), .B(creg[311]), .Z(n37156) );
  XOR U39614 ( .A(n37157), .B(n37158), .Z(n37148) );
  ANDN U39615 ( .A(n37159), .B(n28883), .Z(n37158) );
  XOR U39616 ( .A(n37160), .B(\modmult_1/zin[0][309] ), .Z(n28883) );
  IV U39617 ( .A(n37157), .Z(n37160) );
  XNOR U39618 ( .A(n37157), .B(n28882), .Z(n37159) );
  XOR U39619 ( .A(n37161), .B(n37162), .Z(n28882) );
  AND U39620 ( .A(\modmult_1/xin[1023] ), .B(n37163), .Z(n37162) );
  IV U39621 ( .A(n37161), .Z(n37163) );
  XOR U39622 ( .A(n37164), .B(mreg[310]), .Z(n37161) );
  NAND U39623 ( .A(n37165), .B(mul_pow), .Z(n37164) );
  XOR U39624 ( .A(mreg[310]), .B(creg[310]), .Z(n37165) );
  XOR U39625 ( .A(n37166), .B(n37167), .Z(n37157) );
  ANDN U39626 ( .A(n37168), .B(n28889), .Z(n37167) );
  XOR U39627 ( .A(n37169), .B(\modmult_1/zin[0][308] ), .Z(n28889) );
  IV U39628 ( .A(n37166), .Z(n37169) );
  XNOR U39629 ( .A(n37166), .B(n28888), .Z(n37168) );
  XOR U39630 ( .A(n37170), .B(n37171), .Z(n28888) );
  AND U39631 ( .A(\modmult_1/xin[1023] ), .B(n37172), .Z(n37171) );
  IV U39632 ( .A(n37170), .Z(n37172) );
  XOR U39633 ( .A(n37173), .B(mreg[309]), .Z(n37170) );
  NAND U39634 ( .A(n37174), .B(mul_pow), .Z(n37173) );
  XOR U39635 ( .A(mreg[309]), .B(creg[309]), .Z(n37174) );
  XOR U39636 ( .A(n37175), .B(n37176), .Z(n37166) );
  ANDN U39637 ( .A(n37177), .B(n28895), .Z(n37176) );
  XOR U39638 ( .A(n37178), .B(\modmult_1/zin[0][307] ), .Z(n28895) );
  IV U39639 ( .A(n37175), .Z(n37178) );
  XNOR U39640 ( .A(n37175), .B(n28894), .Z(n37177) );
  XOR U39641 ( .A(n37179), .B(n37180), .Z(n28894) );
  AND U39642 ( .A(\modmult_1/xin[1023] ), .B(n37181), .Z(n37180) );
  IV U39643 ( .A(n37179), .Z(n37181) );
  XOR U39644 ( .A(n37182), .B(mreg[308]), .Z(n37179) );
  NAND U39645 ( .A(n37183), .B(mul_pow), .Z(n37182) );
  XOR U39646 ( .A(mreg[308]), .B(creg[308]), .Z(n37183) );
  XOR U39647 ( .A(n37184), .B(n37185), .Z(n37175) );
  ANDN U39648 ( .A(n37186), .B(n28901), .Z(n37185) );
  XOR U39649 ( .A(n37187), .B(\modmult_1/zin[0][306] ), .Z(n28901) );
  IV U39650 ( .A(n37184), .Z(n37187) );
  XNOR U39651 ( .A(n37184), .B(n28900), .Z(n37186) );
  XOR U39652 ( .A(n37188), .B(n37189), .Z(n28900) );
  AND U39653 ( .A(\modmult_1/xin[1023] ), .B(n37190), .Z(n37189) );
  IV U39654 ( .A(n37188), .Z(n37190) );
  XOR U39655 ( .A(n37191), .B(mreg[307]), .Z(n37188) );
  NAND U39656 ( .A(n37192), .B(mul_pow), .Z(n37191) );
  XOR U39657 ( .A(mreg[307]), .B(creg[307]), .Z(n37192) );
  XOR U39658 ( .A(n37193), .B(n37194), .Z(n37184) );
  ANDN U39659 ( .A(n37195), .B(n28907), .Z(n37194) );
  XOR U39660 ( .A(n37196), .B(\modmult_1/zin[0][305] ), .Z(n28907) );
  IV U39661 ( .A(n37193), .Z(n37196) );
  XNOR U39662 ( .A(n37193), .B(n28906), .Z(n37195) );
  XOR U39663 ( .A(n37197), .B(n37198), .Z(n28906) );
  AND U39664 ( .A(\modmult_1/xin[1023] ), .B(n37199), .Z(n37198) );
  IV U39665 ( .A(n37197), .Z(n37199) );
  XOR U39666 ( .A(n37200), .B(mreg[306]), .Z(n37197) );
  NAND U39667 ( .A(n37201), .B(mul_pow), .Z(n37200) );
  XOR U39668 ( .A(mreg[306]), .B(creg[306]), .Z(n37201) );
  XOR U39669 ( .A(n37202), .B(n37203), .Z(n37193) );
  ANDN U39670 ( .A(n37204), .B(n28913), .Z(n37203) );
  XOR U39671 ( .A(n37205), .B(\modmult_1/zin[0][304] ), .Z(n28913) );
  IV U39672 ( .A(n37202), .Z(n37205) );
  XNOR U39673 ( .A(n37202), .B(n28912), .Z(n37204) );
  XOR U39674 ( .A(n37206), .B(n37207), .Z(n28912) );
  AND U39675 ( .A(\modmult_1/xin[1023] ), .B(n37208), .Z(n37207) );
  IV U39676 ( .A(n37206), .Z(n37208) );
  XOR U39677 ( .A(n37209), .B(mreg[305]), .Z(n37206) );
  NAND U39678 ( .A(n37210), .B(mul_pow), .Z(n37209) );
  XOR U39679 ( .A(mreg[305]), .B(creg[305]), .Z(n37210) );
  XOR U39680 ( .A(n37211), .B(n37212), .Z(n37202) );
  ANDN U39681 ( .A(n37213), .B(n28919), .Z(n37212) );
  XOR U39682 ( .A(n37214), .B(\modmult_1/zin[0][303] ), .Z(n28919) );
  IV U39683 ( .A(n37211), .Z(n37214) );
  XNOR U39684 ( .A(n37211), .B(n28918), .Z(n37213) );
  XOR U39685 ( .A(n37215), .B(n37216), .Z(n28918) );
  AND U39686 ( .A(\modmult_1/xin[1023] ), .B(n37217), .Z(n37216) );
  IV U39687 ( .A(n37215), .Z(n37217) );
  XOR U39688 ( .A(n37218), .B(mreg[304]), .Z(n37215) );
  NAND U39689 ( .A(n37219), .B(mul_pow), .Z(n37218) );
  XOR U39690 ( .A(mreg[304]), .B(creg[304]), .Z(n37219) );
  XOR U39691 ( .A(n37220), .B(n37221), .Z(n37211) );
  ANDN U39692 ( .A(n37222), .B(n28925), .Z(n37221) );
  XOR U39693 ( .A(n37223), .B(\modmult_1/zin[0][302] ), .Z(n28925) );
  IV U39694 ( .A(n37220), .Z(n37223) );
  XNOR U39695 ( .A(n37220), .B(n28924), .Z(n37222) );
  XOR U39696 ( .A(n37224), .B(n37225), .Z(n28924) );
  AND U39697 ( .A(\modmult_1/xin[1023] ), .B(n37226), .Z(n37225) );
  IV U39698 ( .A(n37224), .Z(n37226) );
  XOR U39699 ( .A(n37227), .B(mreg[303]), .Z(n37224) );
  NAND U39700 ( .A(n37228), .B(mul_pow), .Z(n37227) );
  XOR U39701 ( .A(mreg[303]), .B(creg[303]), .Z(n37228) );
  XOR U39702 ( .A(n37229), .B(n37230), .Z(n37220) );
  ANDN U39703 ( .A(n37231), .B(n28931), .Z(n37230) );
  XOR U39704 ( .A(n37232), .B(\modmult_1/zin[0][301] ), .Z(n28931) );
  IV U39705 ( .A(n37229), .Z(n37232) );
  XNOR U39706 ( .A(n37229), .B(n28930), .Z(n37231) );
  XOR U39707 ( .A(n37233), .B(n37234), .Z(n28930) );
  AND U39708 ( .A(\modmult_1/xin[1023] ), .B(n37235), .Z(n37234) );
  IV U39709 ( .A(n37233), .Z(n37235) );
  XOR U39710 ( .A(n37236), .B(mreg[302]), .Z(n37233) );
  NAND U39711 ( .A(n37237), .B(mul_pow), .Z(n37236) );
  XOR U39712 ( .A(mreg[302]), .B(creg[302]), .Z(n37237) );
  XOR U39713 ( .A(n37238), .B(n37239), .Z(n37229) );
  ANDN U39714 ( .A(n37240), .B(n28937), .Z(n37239) );
  XOR U39715 ( .A(n37241), .B(\modmult_1/zin[0][300] ), .Z(n28937) );
  IV U39716 ( .A(n37238), .Z(n37241) );
  XNOR U39717 ( .A(n37238), .B(n28936), .Z(n37240) );
  XOR U39718 ( .A(n37242), .B(n37243), .Z(n28936) );
  AND U39719 ( .A(\modmult_1/xin[1023] ), .B(n37244), .Z(n37243) );
  IV U39720 ( .A(n37242), .Z(n37244) );
  XOR U39721 ( .A(n37245), .B(mreg[301]), .Z(n37242) );
  NAND U39722 ( .A(n37246), .B(mul_pow), .Z(n37245) );
  XOR U39723 ( .A(mreg[301]), .B(creg[301]), .Z(n37246) );
  XOR U39724 ( .A(n37247), .B(n37248), .Z(n37238) );
  ANDN U39725 ( .A(n37249), .B(n28943), .Z(n37248) );
  XOR U39726 ( .A(n37250), .B(\modmult_1/zin[0][299] ), .Z(n28943) );
  IV U39727 ( .A(n37247), .Z(n37250) );
  XNOR U39728 ( .A(n37247), .B(n28942), .Z(n37249) );
  XOR U39729 ( .A(n37251), .B(n37252), .Z(n28942) );
  AND U39730 ( .A(\modmult_1/xin[1023] ), .B(n37253), .Z(n37252) );
  IV U39731 ( .A(n37251), .Z(n37253) );
  XOR U39732 ( .A(n37254), .B(mreg[300]), .Z(n37251) );
  NAND U39733 ( .A(n37255), .B(mul_pow), .Z(n37254) );
  XOR U39734 ( .A(mreg[300]), .B(creg[300]), .Z(n37255) );
  XOR U39735 ( .A(n37256), .B(n37257), .Z(n37247) );
  ANDN U39736 ( .A(n37258), .B(n28949), .Z(n37257) );
  XOR U39737 ( .A(n37259), .B(\modmult_1/zin[0][298] ), .Z(n28949) );
  IV U39738 ( .A(n37256), .Z(n37259) );
  XNOR U39739 ( .A(n37256), .B(n28948), .Z(n37258) );
  XOR U39740 ( .A(n37260), .B(n37261), .Z(n28948) );
  AND U39741 ( .A(\modmult_1/xin[1023] ), .B(n37262), .Z(n37261) );
  IV U39742 ( .A(n37260), .Z(n37262) );
  XOR U39743 ( .A(n37263), .B(mreg[299]), .Z(n37260) );
  NAND U39744 ( .A(n37264), .B(mul_pow), .Z(n37263) );
  XOR U39745 ( .A(mreg[299]), .B(creg[299]), .Z(n37264) );
  XOR U39746 ( .A(n37265), .B(n37266), .Z(n37256) );
  ANDN U39747 ( .A(n37267), .B(n28955), .Z(n37266) );
  XOR U39748 ( .A(n37268), .B(\modmult_1/zin[0][297] ), .Z(n28955) );
  IV U39749 ( .A(n37265), .Z(n37268) );
  XNOR U39750 ( .A(n37265), .B(n28954), .Z(n37267) );
  XOR U39751 ( .A(n37269), .B(n37270), .Z(n28954) );
  AND U39752 ( .A(\modmult_1/xin[1023] ), .B(n37271), .Z(n37270) );
  IV U39753 ( .A(n37269), .Z(n37271) );
  XOR U39754 ( .A(n37272), .B(mreg[298]), .Z(n37269) );
  NAND U39755 ( .A(n37273), .B(mul_pow), .Z(n37272) );
  XOR U39756 ( .A(mreg[298]), .B(creg[298]), .Z(n37273) );
  XOR U39757 ( .A(n37274), .B(n37275), .Z(n37265) );
  ANDN U39758 ( .A(n37276), .B(n28961), .Z(n37275) );
  XOR U39759 ( .A(n37277), .B(\modmult_1/zin[0][296] ), .Z(n28961) );
  IV U39760 ( .A(n37274), .Z(n37277) );
  XNOR U39761 ( .A(n37274), .B(n28960), .Z(n37276) );
  XOR U39762 ( .A(n37278), .B(n37279), .Z(n28960) );
  AND U39763 ( .A(\modmult_1/xin[1023] ), .B(n37280), .Z(n37279) );
  IV U39764 ( .A(n37278), .Z(n37280) );
  XOR U39765 ( .A(n37281), .B(mreg[297]), .Z(n37278) );
  NAND U39766 ( .A(n37282), .B(mul_pow), .Z(n37281) );
  XOR U39767 ( .A(mreg[297]), .B(creg[297]), .Z(n37282) );
  XOR U39768 ( .A(n37283), .B(n37284), .Z(n37274) );
  ANDN U39769 ( .A(n37285), .B(n28967), .Z(n37284) );
  XOR U39770 ( .A(n37286), .B(\modmult_1/zin[0][295] ), .Z(n28967) );
  IV U39771 ( .A(n37283), .Z(n37286) );
  XNOR U39772 ( .A(n37283), .B(n28966), .Z(n37285) );
  XOR U39773 ( .A(n37287), .B(n37288), .Z(n28966) );
  AND U39774 ( .A(\modmult_1/xin[1023] ), .B(n37289), .Z(n37288) );
  IV U39775 ( .A(n37287), .Z(n37289) );
  XOR U39776 ( .A(n37290), .B(mreg[296]), .Z(n37287) );
  NAND U39777 ( .A(n37291), .B(mul_pow), .Z(n37290) );
  XOR U39778 ( .A(mreg[296]), .B(creg[296]), .Z(n37291) );
  XOR U39779 ( .A(n37292), .B(n37293), .Z(n37283) );
  ANDN U39780 ( .A(n37294), .B(n28973), .Z(n37293) );
  XOR U39781 ( .A(n37295), .B(\modmult_1/zin[0][294] ), .Z(n28973) );
  IV U39782 ( .A(n37292), .Z(n37295) );
  XNOR U39783 ( .A(n37292), .B(n28972), .Z(n37294) );
  XOR U39784 ( .A(n37296), .B(n37297), .Z(n28972) );
  AND U39785 ( .A(\modmult_1/xin[1023] ), .B(n37298), .Z(n37297) );
  IV U39786 ( .A(n37296), .Z(n37298) );
  XOR U39787 ( .A(n37299), .B(mreg[295]), .Z(n37296) );
  NAND U39788 ( .A(n37300), .B(mul_pow), .Z(n37299) );
  XOR U39789 ( .A(mreg[295]), .B(creg[295]), .Z(n37300) );
  XOR U39790 ( .A(n37301), .B(n37302), .Z(n37292) );
  ANDN U39791 ( .A(n37303), .B(n28979), .Z(n37302) );
  XOR U39792 ( .A(n37304), .B(\modmult_1/zin[0][293] ), .Z(n28979) );
  IV U39793 ( .A(n37301), .Z(n37304) );
  XNOR U39794 ( .A(n37301), .B(n28978), .Z(n37303) );
  XOR U39795 ( .A(n37305), .B(n37306), .Z(n28978) );
  AND U39796 ( .A(\modmult_1/xin[1023] ), .B(n37307), .Z(n37306) );
  IV U39797 ( .A(n37305), .Z(n37307) );
  XOR U39798 ( .A(n37308), .B(mreg[294]), .Z(n37305) );
  NAND U39799 ( .A(n37309), .B(mul_pow), .Z(n37308) );
  XOR U39800 ( .A(mreg[294]), .B(creg[294]), .Z(n37309) );
  XOR U39801 ( .A(n37310), .B(n37311), .Z(n37301) );
  ANDN U39802 ( .A(n37312), .B(n28985), .Z(n37311) );
  XOR U39803 ( .A(n37313), .B(\modmult_1/zin[0][292] ), .Z(n28985) );
  IV U39804 ( .A(n37310), .Z(n37313) );
  XNOR U39805 ( .A(n37310), .B(n28984), .Z(n37312) );
  XOR U39806 ( .A(n37314), .B(n37315), .Z(n28984) );
  AND U39807 ( .A(\modmult_1/xin[1023] ), .B(n37316), .Z(n37315) );
  IV U39808 ( .A(n37314), .Z(n37316) );
  XOR U39809 ( .A(n37317), .B(mreg[293]), .Z(n37314) );
  NAND U39810 ( .A(n37318), .B(mul_pow), .Z(n37317) );
  XOR U39811 ( .A(mreg[293]), .B(creg[293]), .Z(n37318) );
  XOR U39812 ( .A(n37319), .B(n37320), .Z(n37310) );
  ANDN U39813 ( .A(n37321), .B(n28991), .Z(n37320) );
  XOR U39814 ( .A(n37322), .B(\modmult_1/zin[0][291] ), .Z(n28991) );
  IV U39815 ( .A(n37319), .Z(n37322) );
  XNOR U39816 ( .A(n37319), .B(n28990), .Z(n37321) );
  XOR U39817 ( .A(n37323), .B(n37324), .Z(n28990) );
  AND U39818 ( .A(\modmult_1/xin[1023] ), .B(n37325), .Z(n37324) );
  IV U39819 ( .A(n37323), .Z(n37325) );
  XOR U39820 ( .A(n37326), .B(mreg[292]), .Z(n37323) );
  NAND U39821 ( .A(n37327), .B(mul_pow), .Z(n37326) );
  XOR U39822 ( .A(mreg[292]), .B(creg[292]), .Z(n37327) );
  XOR U39823 ( .A(n37328), .B(n37329), .Z(n37319) );
  ANDN U39824 ( .A(n37330), .B(n28997), .Z(n37329) );
  XOR U39825 ( .A(n37331), .B(\modmult_1/zin[0][290] ), .Z(n28997) );
  IV U39826 ( .A(n37328), .Z(n37331) );
  XNOR U39827 ( .A(n37328), .B(n28996), .Z(n37330) );
  XOR U39828 ( .A(n37332), .B(n37333), .Z(n28996) );
  AND U39829 ( .A(\modmult_1/xin[1023] ), .B(n37334), .Z(n37333) );
  IV U39830 ( .A(n37332), .Z(n37334) );
  XOR U39831 ( .A(n37335), .B(mreg[291]), .Z(n37332) );
  NAND U39832 ( .A(n37336), .B(mul_pow), .Z(n37335) );
  XOR U39833 ( .A(mreg[291]), .B(creg[291]), .Z(n37336) );
  XOR U39834 ( .A(n37337), .B(n37338), .Z(n37328) );
  ANDN U39835 ( .A(n37339), .B(n29003), .Z(n37338) );
  XOR U39836 ( .A(n37340), .B(\modmult_1/zin[0][289] ), .Z(n29003) );
  IV U39837 ( .A(n37337), .Z(n37340) );
  XNOR U39838 ( .A(n37337), .B(n29002), .Z(n37339) );
  XOR U39839 ( .A(n37341), .B(n37342), .Z(n29002) );
  AND U39840 ( .A(\modmult_1/xin[1023] ), .B(n37343), .Z(n37342) );
  IV U39841 ( .A(n37341), .Z(n37343) );
  XOR U39842 ( .A(n37344), .B(mreg[290]), .Z(n37341) );
  NAND U39843 ( .A(n37345), .B(mul_pow), .Z(n37344) );
  XOR U39844 ( .A(mreg[290]), .B(creg[290]), .Z(n37345) );
  XOR U39845 ( .A(n37346), .B(n37347), .Z(n37337) );
  ANDN U39846 ( .A(n37348), .B(n29009), .Z(n37347) );
  XOR U39847 ( .A(n37349), .B(\modmult_1/zin[0][288] ), .Z(n29009) );
  IV U39848 ( .A(n37346), .Z(n37349) );
  XNOR U39849 ( .A(n37346), .B(n29008), .Z(n37348) );
  XOR U39850 ( .A(n37350), .B(n37351), .Z(n29008) );
  AND U39851 ( .A(\modmult_1/xin[1023] ), .B(n37352), .Z(n37351) );
  IV U39852 ( .A(n37350), .Z(n37352) );
  XOR U39853 ( .A(n37353), .B(mreg[289]), .Z(n37350) );
  NAND U39854 ( .A(n37354), .B(mul_pow), .Z(n37353) );
  XOR U39855 ( .A(mreg[289]), .B(creg[289]), .Z(n37354) );
  XOR U39856 ( .A(n37355), .B(n37356), .Z(n37346) );
  ANDN U39857 ( .A(n37357), .B(n29015), .Z(n37356) );
  XOR U39858 ( .A(n37358), .B(\modmult_1/zin[0][287] ), .Z(n29015) );
  IV U39859 ( .A(n37355), .Z(n37358) );
  XNOR U39860 ( .A(n37355), .B(n29014), .Z(n37357) );
  XOR U39861 ( .A(n37359), .B(n37360), .Z(n29014) );
  AND U39862 ( .A(\modmult_1/xin[1023] ), .B(n37361), .Z(n37360) );
  IV U39863 ( .A(n37359), .Z(n37361) );
  XOR U39864 ( .A(n37362), .B(mreg[288]), .Z(n37359) );
  NAND U39865 ( .A(n37363), .B(mul_pow), .Z(n37362) );
  XOR U39866 ( .A(mreg[288]), .B(creg[288]), .Z(n37363) );
  XOR U39867 ( .A(n37364), .B(n37365), .Z(n37355) );
  ANDN U39868 ( .A(n37366), .B(n29021), .Z(n37365) );
  XOR U39869 ( .A(n37367), .B(\modmult_1/zin[0][286] ), .Z(n29021) );
  IV U39870 ( .A(n37364), .Z(n37367) );
  XNOR U39871 ( .A(n37364), .B(n29020), .Z(n37366) );
  XOR U39872 ( .A(n37368), .B(n37369), .Z(n29020) );
  AND U39873 ( .A(\modmult_1/xin[1023] ), .B(n37370), .Z(n37369) );
  IV U39874 ( .A(n37368), .Z(n37370) );
  XOR U39875 ( .A(n37371), .B(mreg[287]), .Z(n37368) );
  NAND U39876 ( .A(n37372), .B(mul_pow), .Z(n37371) );
  XOR U39877 ( .A(mreg[287]), .B(creg[287]), .Z(n37372) );
  XOR U39878 ( .A(n37373), .B(n37374), .Z(n37364) );
  ANDN U39879 ( .A(n37375), .B(n29027), .Z(n37374) );
  XOR U39880 ( .A(n37376), .B(\modmult_1/zin[0][285] ), .Z(n29027) );
  IV U39881 ( .A(n37373), .Z(n37376) );
  XNOR U39882 ( .A(n37373), .B(n29026), .Z(n37375) );
  XOR U39883 ( .A(n37377), .B(n37378), .Z(n29026) );
  AND U39884 ( .A(\modmult_1/xin[1023] ), .B(n37379), .Z(n37378) );
  IV U39885 ( .A(n37377), .Z(n37379) );
  XOR U39886 ( .A(n37380), .B(mreg[286]), .Z(n37377) );
  NAND U39887 ( .A(n37381), .B(mul_pow), .Z(n37380) );
  XOR U39888 ( .A(mreg[286]), .B(creg[286]), .Z(n37381) );
  XOR U39889 ( .A(n37382), .B(n37383), .Z(n37373) );
  ANDN U39890 ( .A(n37384), .B(n29033), .Z(n37383) );
  XOR U39891 ( .A(n37385), .B(\modmult_1/zin[0][284] ), .Z(n29033) );
  IV U39892 ( .A(n37382), .Z(n37385) );
  XNOR U39893 ( .A(n37382), .B(n29032), .Z(n37384) );
  XOR U39894 ( .A(n37386), .B(n37387), .Z(n29032) );
  AND U39895 ( .A(\modmult_1/xin[1023] ), .B(n37388), .Z(n37387) );
  IV U39896 ( .A(n37386), .Z(n37388) );
  XOR U39897 ( .A(n37389), .B(mreg[285]), .Z(n37386) );
  NAND U39898 ( .A(n37390), .B(mul_pow), .Z(n37389) );
  XOR U39899 ( .A(mreg[285]), .B(creg[285]), .Z(n37390) );
  XOR U39900 ( .A(n37391), .B(n37392), .Z(n37382) );
  ANDN U39901 ( .A(n37393), .B(n29039), .Z(n37392) );
  XOR U39902 ( .A(n37394), .B(\modmult_1/zin[0][283] ), .Z(n29039) );
  IV U39903 ( .A(n37391), .Z(n37394) );
  XNOR U39904 ( .A(n37391), .B(n29038), .Z(n37393) );
  XOR U39905 ( .A(n37395), .B(n37396), .Z(n29038) );
  AND U39906 ( .A(\modmult_1/xin[1023] ), .B(n37397), .Z(n37396) );
  IV U39907 ( .A(n37395), .Z(n37397) );
  XOR U39908 ( .A(n37398), .B(mreg[284]), .Z(n37395) );
  NAND U39909 ( .A(n37399), .B(mul_pow), .Z(n37398) );
  XOR U39910 ( .A(mreg[284]), .B(creg[284]), .Z(n37399) );
  XOR U39911 ( .A(n37400), .B(n37401), .Z(n37391) );
  ANDN U39912 ( .A(n37402), .B(n29045), .Z(n37401) );
  XOR U39913 ( .A(n37403), .B(\modmult_1/zin[0][282] ), .Z(n29045) );
  IV U39914 ( .A(n37400), .Z(n37403) );
  XNOR U39915 ( .A(n37400), .B(n29044), .Z(n37402) );
  XOR U39916 ( .A(n37404), .B(n37405), .Z(n29044) );
  AND U39917 ( .A(\modmult_1/xin[1023] ), .B(n37406), .Z(n37405) );
  IV U39918 ( .A(n37404), .Z(n37406) );
  XOR U39919 ( .A(n37407), .B(mreg[283]), .Z(n37404) );
  NAND U39920 ( .A(n37408), .B(mul_pow), .Z(n37407) );
  XOR U39921 ( .A(mreg[283]), .B(creg[283]), .Z(n37408) );
  XOR U39922 ( .A(n37409), .B(n37410), .Z(n37400) );
  ANDN U39923 ( .A(n37411), .B(n29051), .Z(n37410) );
  XOR U39924 ( .A(n37412), .B(\modmult_1/zin[0][281] ), .Z(n29051) );
  IV U39925 ( .A(n37409), .Z(n37412) );
  XNOR U39926 ( .A(n37409), .B(n29050), .Z(n37411) );
  XOR U39927 ( .A(n37413), .B(n37414), .Z(n29050) );
  AND U39928 ( .A(\modmult_1/xin[1023] ), .B(n37415), .Z(n37414) );
  IV U39929 ( .A(n37413), .Z(n37415) );
  XOR U39930 ( .A(n37416), .B(mreg[282]), .Z(n37413) );
  NAND U39931 ( .A(n37417), .B(mul_pow), .Z(n37416) );
  XOR U39932 ( .A(mreg[282]), .B(creg[282]), .Z(n37417) );
  XOR U39933 ( .A(n37418), .B(n37419), .Z(n37409) );
  ANDN U39934 ( .A(n37420), .B(n29057), .Z(n37419) );
  XOR U39935 ( .A(n37421), .B(\modmult_1/zin[0][280] ), .Z(n29057) );
  IV U39936 ( .A(n37418), .Z(n37421) );
  XNOR U39937 ( .A(n37418), .B(n29056), .Z(n37420) );
  XOR U39938 ( .A(n37422), .B(n37423), .Z(n29056) );
  AND U39939 ( .A(\modmult_1/xin[1023] ), .B(n37424), .Z(n37423) );
  IV U39940 ( .A(n37422), .Z(n37424) );
  XOR U39941 ( .A(n37425), .B(mreg[281]), .Z(n37422) );
  NAND U39942 ( .A(n37426), .B(mul_pow), .Z(n37425) );
  XOR U39943 ( .A(mreg[281]), .B(creg[281]), .Z(n37426) );
  XOR U39944 ( .A(n37427), .B(n37428), .Z(n37418) );
  ANDN U39945 ( .A(n37429), .B(n29063), .Z(n37428) );
  XOR U39946 ( .A(n37430), .B(\modmult_1/zin[0][279] ), .Z(n29063) );
  IV U39947 ( .A(n37427), .Z(n37430) );
  XNOR U39948 ( .A(n37427), .B(n29062), .Z(n37429) );
  XOR U39949 ( .A(n37431), .B(n37432), .Z(n29062) );
  AND U39950 ( .A(\modmult_1/xin[1023] ), .B(n37433), .Z(n37432) );
  IV U39951 ( .A(n37431), .Z(n37433) );
  XOR U39952 ( .A(n37434), .B(mreg[280]), .Z(n37431) );
  NAND U39953 ( .A(n37435), .B(mul_pow), .Z(n37434) );
  XOR U39954 ( .A(mreg[280]), .B(creg[280]), .Z(n37435) );
  XOR U39955 ( .A(n37436), .B(n37437), .Z(n37427) );
  ANDN U39956 ( .A(n37438), .B(n29069), .Z(n37437) );
  XOR U39957 ( .A(n37439), .B(\modmult_1/zin[0][278] ), .Z(n29069) );
  IV U39958 ( .A(n37436), .Z(n37439) );
  XNOR U39959 ( .A(n37436), .B(n29068), .Z(n37438) );
  XOR U39960 ( .A(n37440), .B(n37441), .Z(n29068) );
  AND U39961 ( .A(\modmult_1/xin[1023] ), .B(n37442), .Z(n37441) );
  IV U39962 ( .A(n37440), .Z(n37442) );
  XOR U39963 ( .A(n37443), .B(mreg[279]), .Z(n37440) );
  NAND U39964 ( .A(n37444), .B(mul_pow), .Z(n37443) );
  XOR U39965 ( .A(mreg[279]), .B(creg[279]), .Z(n37444) );
  XOR U39966 ( .A(n37445), .B(n37446), .Z(n37436) );
  ANDN U39967 ( .A(n37447), .B(n29075), .Z(n37446) );
  XOR U39968 ( .A(n37448), .B(\modmult_1/zin[0][277] ), .Z(n29075) );
  IV U39969 ( .A(n37445), .Z(n37448) );
  XNOR U39970 ( .A(n37445), .B(n29074), .Z(n37447) );
  XOR U39971 ( .A(n37449), .B(n37450), .Z(n29074) );
  AND U39972 ( .A(\modmult_1/xin[1023] ), .B(n37451), .Z(n37450) );
  IV U39973 ( .A(n37449), .Z(n37451) );
  XOR U39974 ( .A(n37452), .B(mreg[278]), .Z(n37449) );
  NAND U39975 ( .A(n37453), .B(mul_pow), .Z(n37452) );
  XOR U39976 ( .A(mreg[278]), .B(creg[278]), .Z(n37453) );
  XOR U39977 ( .A(n37454), .B(n37455), .Z(n37445) );
  ANDN U39978 ( .A(n37456), .B(n29081), .Z(n37455) );
  XOR U39979 ( .A(n37457), .B(\modmult_1/zin[0][276] ), .Z(n29081) );
  IV U39980 ( .A(n37454), .Z(n37457) );
  XNOR U39981 ( .A(n37454), .B(n29080), .Z(n37456) );
  XOR U39982 ( .A(n37458), .B(n37459), .Z(n29080) );
  AND U39983 ( .A(\modmult_1/xin[1023] ), .B(n37460), .Z(n37459) );
  IV U39984 ( .A(n37458), .Z(n37460) );
  XOR U39985 ( .A(n37461), .B(mreg[277]), .Z(n37458) );
  NAND U39986 ( .A(n37462), .B(mul_pow), .Z(n37461) );
  XOR U39987 ( .A(mreg[277]), .B(creg[277]), .Z(n37462) );
  XOR U39988 ( .A(n37463), .B(n37464), .Z(n37454) );
  ANDN U39989 ( .A(n37465), .B(n29087), .Z(n37464) );
  XOR U39990 ( .A(n37466), .B(\modmult_1/zin[0][275] ), .Z(n29087) );
  IV U39991 ( .A(n37463), .Z(n37466) );
  XNOR U39992 ( .A(n37463), .B(n29086), .Z(n37465) );
  XOR U39993 ( .A(n37467), .B(n37468), .Z(n29086) );
  AND U39994 ( .A(\modmult_1/xin[1023] ), .B(n37469), .Z(n37468) );
  IV U39995 ( .A(n37467), .Z(n37469) );
  XOR U39996 ( .A(n37470), .B(mreg[276]), .Z(n37467) );
  NAND U39997 ( .A(n37471), .B(mul_pow), .Z(n37470) );
  XOR U39998 ( .A(mreg[276]), .B(creg[276]), .Z(n37471) );
  XOR U39999 ( .A(n37472), .B(n37473), .Z(n37463) );
  ANDN U40000 ( .A(n37474), .B(n29093), .Z(n37473) );
  XOR U40001 ( .A(n37475), .B(\modmult_1/zin[0][274] ), .Z(n29093) );
  IV U40002 ( .A(n37472), .Z(n37475) );
  XNOR U40003 ( .A(n37472), .B(n29092), .Z(n37474) );
  XOR U40004 ( .A(n37476), .B(n37477), .Z(n29092) );
  AND U40005 ( .A(\modmult_1/xin[1023] ), .B(n37478), .Z(n37477) );
  IV U40006 ( .A(n37476), .Z(n37478) );
  XOR U40007 ( .A(n37479), .B(mreg[275]), .Z(n37476) );
  NAND U40008 ( .A(n37480), .B(mul_pow), .Z(n37479) );
  XOR U40009 ( .A(mreg[275]), .B(creg[275]), .Z(n37480) );
  XOR U40010 ( .A(n37481), .B(n37482), .Z(n37472) );
  ANDN U40011 ( .A(n37483), .B(n29099), .Z(n37482) );
  XOR U40012 ( .A(n37484), .B(\modmult_1/zin[0][273] ), .Z(n29099) );
  IV U40013 ( .A(n37481), .Z(n37484) );
  XNOR U40014 ( .A(n37481), .B(n29098), .Z(n37483) );
  XOR U40015 ( .A(n37485), .B(n37486), .Z(n29098) );
  AND U40016 ( .A(\modmult_1/xin[1023] ), .B(n37487), .Z(n37486) );
  IV U40017 ( .A(n37485), .Z(n37487) );
  XOR U40018 ( .A(n37488), .B(mreg[274]), .Z(n37485) );
  NAND U40019 ( .A(n37489), .B(mul_pow), .Z(n37488) );
  XOR U40020 ( .A(mreg[274]), .B(creg[274]), .Z(n37489) );
  XOR U40021 ( .A(n37490), .B(n37491), .Z(n37481) );
  ANDN U40022 ( .A(n37492), .B(n29105), .Z(n37491) );
  XOR U40023 ( .A(n37493), .B(\modmult_1/zin[0][272] ), .Z(n29105) );
  IV U40024 ( .A(n37490), .Z(n37493) );
  XNOR U40025 ( .A(n37490), .B(n29104), .Z(n37492) );
  XOR U40026 ( .A(n37494), .B(n37495), .Z(n29104) );
  AND U40027 ( .A(\modmult_1/xin[1023] ), .B(n37496), .Z(n37495) );
  IV U40028 ( .A(n37494), .Z(n37496) );
  XOR U40029 ( .A(n37497), .B(mreg[273]), .Z(n37494) );
  NAND U40030 ( .A(n37498), .B(mul_pow), .Z(n37497) );
  XOR U40031 ( .A(mreg[273]), .B(creg[273]), .Z(n37498) );
  XOR U40032 ( .A(n37499), .B(n37500), .Z(n37490) );
  ANDN U40033 ( .A(n37501), .B(n29111), .Z(n37500) );
  XOR U40034 ( .A(n37502), .B(\modmult_1/zin[0][271] ), .Z(n29111) );
  IV U40035 ( .A(n37499), .Z(n37502) );
  XNOR U40036 ( .A(n37499), .B(n29110), .Z(n37501) );
  XOR U40037 ( .A(n37503), .B(n37504), .Z(n29110) );
  AND U40038 ( .A(\modmult_1/xin[1023] ), .B(n37505), .Z(n37504) );
  IV U40039 ( .A(n37503), .Z(n37505) );
  XOR U40040 ( .A(n37506), .B(mreg[272]), .Z(n37503) );
  NAND U40041 ( .A(n37507), .B(mul_pow), .Z(n37506) );
  XOR U40042 ( .A(mreg[272]), .B(creg[272]), .Z(n37507) );
  XOR U40043 ( .A(n37508), .B(n37509), .Z(n37499) );
  ANDN U40044 ( .A(n37510), .B(n29117), .Z(n37509) );
  XOR U40045 ( .A(n37511), .B(\modmult_1/zin[0][270] ), .Z(n29117) );
  IV U40046 ( .A(n37508), .Z(n37511) );
  XNOR U40047 ( .A(n37508), .B(n29116), .Z(n37510) );
  XOR U40048 ( .A(n37512), .B(n37513), .Z(n29116) );
  AND U40049 ( .A(\modmult_1/xin[1023] ), .B(n37514), .Z(n37513) );
  IV U40050 ( .A(n37512), .Z(n37514) );
  XOR U40051 ( .A(n37515), .B(mreg[271]), .Z(n37512) );
  NAND U40052 ( .A(n37516), .B(mul_pow), .Z(n37515) );
  XOR U40053 ( .A(mreg[271]), .B(creg[271]), .Z(n37516) );
  XOR U40054 ( .A(n37517), .B(n37518), .Z(n37508) );
  ANDN U40055 ( .A(n37519), .B(n29123), .Z(n37518) );
  XOR U40056 ( .A(n37520), .B(\modmult_1/zin[0][269] ), .Z(n29123) );
  IV U40057 ( .A(n37517), .Z(n37520) );
  XNOR U40058 ( .A(n37517), .B(n29122), .Z(n37519) );
  XOR U40059 ( .A(n37521), .B(n37522), .Z(n29122) );
  AND U40060 ( .A(\modmult_1/xin[1023] ), .B(n37523), .Z(n37522) );
  IV U40061 ( .A(n37521), .Z(n37523) );
  XOR U40062 ( .A(n37524), .B(mreg[270]), .Z(n37521) );
  NAND U40063 ( .A(n37525), .B(mul_pow), .Z(n37524) );
  XOR U40064 ( .A(mreg[270]), .B(creg[270]), .Z(n37525) );
  XOR U40065 ( .A(n37526), .B(n37527), .Z(n37517) );
  ANDN U40066 ( .A(n37528), .B(n29129), .Z(n37527) );
  XOR U40067 ( .A(n37529), .B(\modmult_1/zin[0][268] ), .Z(n29129) );
  IV U40068 ( .A(n37526), .Z(n37529) );
  XNOR U40069 ( .A(n37526), .B(n29128), .Z(n37528) );
  XOR U40070 ( .A(n37530), .B(n37531), .Z(n29128) );
  AND U40071 ( .A(\modmult_1/xin[1023] ), .B(n37532), .Z(n37531) );
  IV U40072 ( .A(n37530), .Z(n37532) );
  XOR U40073 ( .A(n37533), .B(mreg[269]), .Z(n37530) );
  NAND U40074 ( .A(n37534), .B(mul_pow), .Z(n37533) );
  XOR U40075 ( .A(mreg[269]), .B(creg[269]), .Z(n37534) );
  XOR U40076 ( .A(n37535), .B(n37536), .Z(n37526) );
  ANDN U40077 ( .A(n37537), .B(n29135), .Z(n37536) );
  XOR U40078 ( .A(n37538), .B(\modmult_1/zin[0][267] ), .Z(n29135) );
  IV U40079 ( .A(n37535), .Z(n37538) );
  XNOR U40080 ( .A(n37535), .B(n29134), .Z(n37537) );
  XOR U40081 ( .A(n37539), .B(n37540), .Z(n29134) );
  AND U40082 ( .A(\modmult_1/xin[1023] ), .B(n37541), .Z(n37540) );
  IV U40083 ( .A(n37539), .Z(n37541) );
  XOR U40084 ( .A(n37542), .B(mreg[268]), .Z(n37539) );
  NAND U40085 ( .A(n37543), .B(mul_pow), .Z(n37542) );
  XOR U40086 ( .A(mreg[268]), .B(creg[268]), .Z(n37543) );
  XOR U40087 ( .A(n37544), .B(n37545), .Z(n37535) );
  ANDN U40088 ( .A(n37546), .B(n29141), .Z(n37545) );
  XOR U40089 ( .A(n37547), .B(\modmult_1/zin[0][266] ), .Z(n29141) );
  IV U40090 ( .A(n37544), .Z(n37547) );
  XNOR U40091 ( .A(n37544), .B(n29140), .Z(n37546) );
  XOR U40092 ( .A(n37548), .B(n37549), .Z(n29140) );
  AND U40093 ( .A(\modmult_1/xin[1023] ), .B(n37550), .Z(n37549) );
  IV U40094 ( .A(n37548), .Z(n37550) );
  XOR U40095 ( .A(n37551), .B(mreg[267]), .Z(n37548) );
  NAND U40096 ( .A(n37552), .B(mul_pow), .Z(n37551) );
  XOR U40097 ( .A(mreg[267]), .B(creg[267]), .Z(n37552) );
  XOR U40098 ( .A(n37553), .B(n37554), .Z(n37544) );
  ANDN U40099 ( .A(n37555), .B(n29147), .Z(n37554) );
  XOR U40100 ( .A(n37556), .B(\modmult_1/zin[0][265] ), .Z(n29147) );
  IV U40101 ( .A(n37553), .Z(n37556) );
  XNOR U40102 ( .A(n37553), .B(n29146), .Z(n37555) );
  XOR U40103 ( .A(n37557), .B(n37558), .Z(n29146) );
  AND U40104 ( .A(\modmult_1/xin[1023] ), .B(n37559), .Z(n37558) );
  IV U40105 ( .A(n37557), .Z(n37559) );
  XOR U40106 ( .A(n37560), .B(mreg[266]), .Z(n37557) );
  NAND U40107 ( .A(n37561), .B(mul_pow), .Z(n37560) );
  XOR U40108 ( .A(mreg[266]), .B(creg[266]), .Z(n37561) );
  XOR U40109 ( .A(n37562), .B(n37563), .Z(n37553) );
  ANDN U40110 ( .A(n37564), .B(n29153), .Z(n37563) );
  XOR U40111 ( .A(n37565), .B(\modmult_1/zin[0][264] ), .Z(n29153) );
  IV U40112 ( .A(n37562), .Z(n37565) );
  XNOR U40113 ( .A(n37562), .B(n29152), .Z(n37564) );
  XOR U40114 ( .A(n37566), .B(n37567), .Z(n29152) );
  AND U40115 ( .A(\modmult_1/xin[1023] ), .B(n37568), .Z(n37567) );
  IV U40116 ( .A(n37566), .Z(n37568) );
  XOR U40117 ( .A(n37569), .B(mreg[265]), .Z(n37566) );
  NAND U40118 ( .A(n37570), .B(mul_pow), .Z(n37569) );
  XOR U40119 ( .A(mreg[265]), .B(creg[265]), .Z(n37570) );
  XOR U40120 ( .A(n37571), .B(n37572), .Z(n37562) );
  ANDN U40121 ( .A(n37573), .B(n29159), .Z(n37572) );
  XOR U40122 ( .A(n37574), .B(\modmult_1/zin[0][263] ), .Z(n29159) );
  IV U40123 ( .A(n37571), .Z(n37574) );
  XNOR U40124 ( .A(n37571), .B(n29158), .Z(n37573) );
  XOR U40125 ( .A(n37575), .B(n37576), .Z(n29158) );
  AND U40126 ( .A(\modmult_1/xin[1023] ), .B(n37577), .Z(n37576) );
  IV U40127 ( .A(n37575), .Z(n37577) );
  XOR U40128 ( .A(n37578), .B(mreg[264]), .Z(n37575) );
  NAND U40129 ( .A(n37579), .B(mul_pow), .Z(n37578) );
  XOR U40130 ( .A(mreg[264]), .B(creg[264]), .Z(n37579) );
  XOR U40131 ( .A(n37580), .B(n37581), .Z(n37571) );
  ANDN U40132 ( .A(n37582), .B(n29165), .Z(n37581) );
  XOR U40133 ( .A(n37583), .B(\modmult_1/zin[0][262] ), .Z(n29165) );
  IV U40134 ( .A(n37580), .Z(n37583) );
  XNOR U40135 ( .A(n37580), .B(n29164), .Z(n37582) );
  XOR U40136 ( .A(n37584), .B(n37585), .Z(n29164) );
  AND U40137 ( .A(\modmult_1/xin[1023] ), .B(n37586), .Z(n37585) );
  IV U40138 ( .A(n37584), .Z(n37586) );
  XOR U40139 ( .A(n37587), .B(mreg[263]), .Z(n37584) );
  NAND U40140 ( .A(n37588), .B(mul_pow), .Z(n37587) );
  XOR U40141 ( .A(mreg[263]), .B(creg[263]), .Z(n37588) );
  XOR U40142 ( .A(n37589), .B(n37590), .Z(n37580) );
  ANDN U40143 ( .A(n37591), .B(n29171), .Z(n37590) );
  XOR U40144 ( .A(n37592), .B(\modmult_1/zin[0][261] ), .Z(n29171) );
  IV U40145 ( .A(n37589), .Z(n37592) );
  XNOR U40146 ( .A(n37589), .B(n29170), .Z(n37591) );
  XOR U40147 ( .A(n37593), .B(n37594), .Z(n29170) );
  AND U40148 ( .A(\modmult_1/xin[1023] ), .B(n37595), .Z(n37594) );
  IV U40149 ( .A(n37593), .Z(n37595) );
  XOR U40150 ( .A(n37596), .B(mreg[262]), .Z(n37593) );
  NAND U40151 ( .A(n37597), .B(mul_pow), .Z(n37596) );
  XOR U40152 ( .A(mreg[262]), .B(creg[262]), .Z(n37597) );
  XOR U40153 ( .A(n37598), .B(n37599), .Z(n37589) );
  ANDN U40154 ( .A(n37600), .B(n29177), .Z(n37599) );
  XOR U40155 ( .A(n37601), .B(\modmult_1/zin[0][260] ), .Z(n29177) );
  IV U40156 ( .A(n37598), .Z(n37601) );
  XNOR U40157 ( .A(n37598), .B(n29176), .Z(n37600) );
  XOR U40158 ( .A(n37602), .B(n37603), .Z(n29176) );
  AND U40159 ( .A(\modmult_1/xin[1023] ), .B(n37604), .Z(n37603) );
  IV U40160 ( .A(n37602), .Z(n37604) );
  XOR U40161 ( .A(n37605), .B(mreg[261]), .Z(n37602) );
  NAND U40162 ( .A(n37606), .B(mul_pow), .Z(n37605) );
  XOR U40163 ( .A(mreg[261]), .B(creg[261]), .Z(n37606) );
  XOR U40164 ( .A(n37607), .B(n37608), .Z(n37598) );
  ANDN U40165 ( .A(n37609), .B(n29183), .Z(n37608) );
  XOR U40166 ( .A(n37610), .B(\modmult_1/zin[0][259] ), .Z(n29183) );
  IV U40167 ( .A(n37607), .Z(n37610) );
  XNOR U40168 ( .A(n37607), .B(n29182), .Z(n37609) );
  XOR U40169 ( .A(n37611), .B(n37612), .Z(n29182) );
  AND U40170 ( .A(\modmult_1/xin[1023] ), .B(n37613), .Z(n37612) );
  IV U40171 ( .A(n37611), .Z(n37613) );
  XOR U40172 ( .A(n37614), .B(mreg[260]), .Z(n37611) );
  NAND U40173 ( .A(n37615), .B(mul_pow), .Z(n37614) );
  XOR U40174 ( .A(mreg[260]), .B(creg[260]), .Z(n37615) );
  XOR U40175 ( .A(n37616), .B(n37617), .Z(n37607) );
  ANDN U40176 ( .A(n37618), .B(n29189), .Z(n37617) );
  XOR U40177 ( .A(n37619), .B(\modmult_1/zin[0][258] ), .Z(n29189) );
  IV U40178 ( .A(n37616), .Z(n37619) );
  XNOR U40179 ( .A(n37616), .B(n29188), .Z(n37618) );
  XOR U40180 ( .A(n37620), .B(n37621), .Z(n29188) );
  AND U40181 ( .A(\modmult_1/xin[1023] ), .B(n37622), .Z(n37621) );
  IV U40182 ( .A(n37620), .Z(n37622) );
  XOR U40183 ( .A(n37623), .B(mreg[259]), .Z(n37620) );
  NAND U40184 ( .A(n37624), .B(mul_pow), .Z(n37623) );
  XOR U40185 ( .A(mreg[259]), .B(creg[259]), .Z(n37624) );
  XOR U40186 ( .A(n37625), .B(n37626), .Z(n37616) );
  ANDN U40187 ( .A(n37627), .B(n29195), .Z(n37626) );
  XOR U40188 ( .A(n37628), .B(\modmult_1/zin[0][257] ), .Z(n29195) );
  IV U40189 ( .A(n37625), .Z(n37628) );
  XNOR U40190 ( .A(n37625), .B(n29194), .Z(n37627) );
  XOR U40191 ( .A(n37629), .B(n37630), .Z(n29194) );
  AND U40192 ( .A(\modmult_1/xin[1023] ), .B(n37631), .Z(n37630) );
  IV U40193 ( .A(n37629), .Z(n37631) );
  XOR U40194 ( .A(n37632), .B(mreg[258]), .Z(n37629) );
  NAND U40195 ( .A(n37633), .B(mul_pow), .Z(n37632) );
  XOR U40196 ( .A(mreg[258]), .B(creg[258]), .Z(n37633) );
  XOR U40197 ( .A(n37634), .B(n37635), .Z(n37625) );
  ANDN U40198 ( .A(n37636), .B(n29201), .Z(n37635) );
  XOR U40199 ( .A(n37637), .B(\modmult_1/zin[0][256] ), .Z(n29201) );
  IV U40200 ( .A(n37634), .Z(n37637) );
  XNOR U40201 ( .A(n37634), .B(n29200), .Z(n37636) );
  XOR U40202 ( .A(n37638), .B(n37639), .Z(n29200) );
  AND U40203 ( .A(\modmult_1/xin[1023] ), .B(n37640), .Z(n37639) );
  IV U40204 ( .A(n37638), .Z(n37640) );
  XOR U40205 ( .A(n37641), .B(mreg[257]), .Z(n37638) );
  NAND U40206 ( .A(n37642), .B(mul_pow), .Z(n37641) );
  XOR U40207 ( .A(mreg[257]), .B(creg[257]), .Z(n37642) );
  XOR U40208 ( .A(n37643), .B(n37644), .Z(n37634) );
  ANDN U40209 ( .A(n37645), .B(n29207), .Z(n37644) );
  XOR U40210 ( .A(n37646), .B(\modmult_1/zin[0][255] ), .Z(n29207) );
  IV U40211 ( .A(n37643), .Z(n37646) );
  XNOR U40212 ( .A(n37643), .B(n29206), .Z(n37645) );
  XOR U40213 ( .A(n37647), .B(n37648), .Z(n29206) );
  AND U40214 ( .A(\modmult_1/xin[1023] ), .B(n37649), .Z(n37648) );
  IV U40215 ( .A(n37647), .Z(n37649) );
  XOR U40216 ( .A(n37650), .B(mreg[256]), .Z(n37647) );
  NAND U40217 ( .A(n37651), .B(mul_pow), .Z(n37650) );
  XOR U40218 ( .A(mreg[256]), .B(creg[256]), .Z(n37651) );
  XOR U40219 ( .A(n37652), .B(n37653), .Z(n37643) );
  ANDN U40220 ( .A(n37654), .B(n29213), .Z(n37653) );
  XOR U40221 ( .A(n37655), .B(\modmult_1/zin[0][254] ), .Z(n29213) );
  IV U40222 ( .A(n37652), .Z(n37655) );
  XNOR U40223 ( .A(n37652), .B(n29212), .Z(n37654) );
  XOR U40224 ( .A(n37656), .B(n37657), .Z(n29212) );
  AND U40225 ( .A(\modmult_1/xin[1023] ), .B(n37658), .Z(n37657) );
  IV U40226 ( .A(n37656), .Z(n37658) );
  XOR U40227 ( .A(n37659), .B(mreg[255]), .Z(n37656) );
  NAND U40228 ( .A(n37660), .B(mul_pow), .Z(n37659) );
  XOR U40229 ( .A(mreg[255]), .B(creg[255]), .Z(n37660) );
  XOR U40230 ( .A(n37661), .B(n37662), .Z(n37652) );
  ANDN U40231 ( .A(n37663), .B(n29219), .Z(n37662) );
  XOR U40232 ( .A(n37664), .B(\modmult_1/zin[0][253] ), .Z(n29219) );
  IV U40233 ( .A(n37661), .Z(n37664) );
  XNOR U40234 ( .A(n37661), .B(n29218), .Z(n37663) );
  XOR U40235 ( .A(n37665), .B(n37666), .Z(n29218) );
  AND U40236 ( .A(\modmult_1/xin[1023] ), .B(n37667), .Z(n37666) );
  IV U40237 ( .A(n37665), .Z(n37667) );
  XOR U40238 ( .A(n37668), .B(mreg[254]), .Z(n37665) );
  NAND U40239 ( .A(n37669), .B(mul_pow), .Z(n37668) );
  XOR U40240 ( .A(mreg[254]), .B(creg[254]), .Z(n37669) );
  XOR U40241 ( .A(n37670), .B(n37671), .Z(n37661) );
  ANDN U40242 ( .A(n37672), .B(n29225), .Z(n37671) );
  XOR U40243 ( .A(n37673), .B(\modmult_1/zin[0][252] ), .Z(n29225) );
  IV U40244 ( .A(n37670), .Z(n37673) );
  XNOR U40245 ( .A(n37670), .B(n29224), .Z(n37672) );
  XOR U40246 ( .A(n37674), .B(n37675), .Z(n29224) );
  AND U40247 ( .A(\modmult_1/xin[1023] ), .B(n37676), .Z(n37675) );
  IV U40248 ( .A(n37674), .Z(n37676) );
  XOR U40249 ( .A(n37677), .B(mreg[253]), .Z(n37674) );
  NAND U40250 ( .A(n37678), .B(mul_pow), .Z(n37677) );
  XOR U40251 ( .A(mreg[253]), .B(creg[253]), .Z(n37678) );
  XOR U40252 ( .A(n37679), .B(n37680), .Z(n37670) );
  ANDN U40253 ( .A(n37681), .B(n29231), .Z(n37680) );
  XOR U40254 ( .A(n37682), .B(\modmult_1/zin[0][251] ), .Z(n29231) );
  IV U40255 ( .A(n37679), .Z(n37682) );
  XNOR U40256 ( .A(n37679), .B(n29230), .Z(n37681) );
  XOR U40257 ( .A(n37683), .B(n37684), .Z(n29230) );
  AND U40258 ( .A(\modmult_1/xin[1023] ), .B(n37685), .Z(n37684) );
  IV U40259 ( .A(n37683), .Z(n37685) );
  XOR U40260 ( .A(n37686), .B(mreg[252]), .Z(n37683) );
  NAND U40261 ( .A(n37687), .B(mul_pow), .Z(n37686) );
  XOR U40262 ( .A(mreg[252]), .B(creg[252]), .Z(n37687) );
  XOR U40263 ( .A(n37688), .B(n37689), .Z(n37679) );
  ANDN U40264 ( .A(n37690), .B(n29237), .Z(n37689) );
  XOR U40265 ( .A(n37691), .B(\modmult_1/zin[0][250] ), .Z(n29237) );
  IV U40266 ( .A(n37688), .Z(n37691) );
  XNOR U40267 ( .A(n37688), .B(n29236), .Z(n37690) );
  XOR U40268 ( .A(n37692), .B(n37693), .Z(n29236) );
  AND U40269 ( .A(\modmult_1/xin[1023] ), .B(n37694), .Z(n37693) );
  IV U40270 ( .A(n37692), .Z(n37694) );
  XOR U40271 ( .A(n37695), .B(mreg[251]), .Z(n37692) );
  NAND U40272 ( .A(n37696), .B(mul_pow), .Z(n37695) );
  XOR U40273 ( .A(mreg[251]), .B(creg[251]), .Z(n37696) );
  XOR U40274 ( .A(n37697), .B(n37698), .Z(n37688) );
  ANDN U40275 ( .A(n37699), .B(n29243), .Z(n37698) );
  XOR U40276 ( .A(n37700), .B(\modmult_1/zin[0][249] ), .Z(n29243) );
  IV U40277 ( .A(n37697), .Z(n37700) );
  XNOR U40278 ( .A(n37697), .B(n29242), .Z(n37699) );
  XOR U40279 ( .A(n37701), .B(n37702), .Z(n29242) );
  AND U40280 ( .A(\modmult_1/xin[1023] ), .B(n37703), .Z(n37702) );
  IV U40281 ( .A(n37701), .Z(n37703) );
  XOR U40282 ( .A(n37704), .B(mreg[250]), .Z(n37701) );
  NAND U40283 ( .A(n37705), .B(mul_pow), .Z(n37704) );
  XOR U40284 ( .A(mreg[250]), .B(creg[250]), .Z(n37705) );
  XOR U40285 ( .A(n37706), .B(n37707), .Z(n37697) );
  ANDN U40286 ( .A(n37708), .B(n29249), .Z(n37707) );
  XOR U40287 ( .A(n37709), .B(\modmult_1/zin[0][248] ), .Z(n29249) );
  IV U40288 ( .A(n37706), .Z(n37709) );
  XNOR U40289 ( .A(n37706), .B(n29248), .Z(n37708) );
  XOR U40290 ( .A(n37710), .B(n37711), .Z(n29248) );
  AND U40291 ( .A(\modmult_1/xin[1023] ), .B(n37712), .Z(n37711) );
  IV U40292 ( .A(n37710), .Z(n37712) );
  XOR U40293 ( .A(n37713), .B(mreg[249]), .Z(n37710) );
  NAND U40294 ( .A(n37714), .B(mul_pow), .Z(n37713) );
  XOR U40295 ( .A(mreg[249]), .B(creg[249]), .Z(n37714) );
  XOR U40296 ( .A(n37715), .B(n37716), .Z(n37706) );
  ANDN U40297 ( .A(n37717), .B(n29255), .Z(n37716) );
  XOR U40298 ( .A(n37718), .B(\modmult_1/zin[0][247] ), .Z(n29255) );
  IV U40299 ( .A(n37715), .Z(n37718) );
  XNOR U40300 ( .A(n37715), .B(n29254), .Z(n37717) );
  XOR U40301 ( .A(n37719), .B(n37720), .Z(n29254) );
  AND U40302 ( .A(\modmult_1/xin[1023] ), .B(n37721), .Z(n37720) );
  IV U40303 ( .A(n37719), .Z(n37721) );
  XOR U40304 ( .A(n37722), .B(mreg[248]), .Z(n37719) );
  NAND U40305 ( .A(n37723), .B(mul_pow), .Z(n37722) );
  XOR U40306 ( .A(mreg[248]), .B(creg[248]), .Z(n37723) );
  XOR U40307 ( .A(n37724), .B(n37725), .Z(n37715) );
  ANDN U40308 ( .A(n37726), .B(n29261), .Z(n37725) );
  XOR U40309 ( .A(n37727), .B(\modmult_1/zin[0][246] ), .Z(n29261) );
  IV U40310 ( .A(n37724), .Z(n37727) );
  XNOR U40311 ( .A(n37724), .B(n29260), .Z(n37726) );
  XOR U40312 ( .A(n37728), .B(n37729), .Z(n29260) );
  AND U40313 ( .A(\modmult_1/xin[1023] ), .B(n37730), .Z(n37729) );
  IV U40314 ( .A(n37728), .Z(n37730) );
  XOR U40315 ( .A(n37731), .B(mreg[247]), .Z(n37728) );
  NAND U40316 ( .A(n37732), .B(mul_pow), .Z(n37731) );
  XOR U40317 ( .A(mreg[247]), .B(creg[247]), .Z(n37732) );
  XOR U40318 ( .A(n37733), .B(n37734), .Z(n37724) );
  ANDN U40319 ( .A(n37735), .B(n29267), .Z(n37734) );
  XOR U40320 ( .A(n37736), .B(\modmult_1/zin[0][245] ), .Z(n29267) );
  IV U40321 ( .A(n37733), .Z(n37736) );
  XNOR U40322 ( .A(n37733), .B(n29266), .Z(n37735) );
  XOR U40323 ( .A(n37737), .B(n37738), .Z(n29266) );
  AND U40324 ( .A(\modmult_1/xin[1023] ), .B(n37739), .Z(n37738) );
  IV U40325 ( .A(n37737), .Z(n37739) );
  XOR U40326 ( .A(n37740), .B(mreg[246]), .Z(n37737) );
  NAND U40327 ( .A(n37741), .B(mul_pow), .Z(n37740) );
  XOR U40328 ( .A(mreg[246]), .B(creg[246]), .Z(n37741) );
  XOR U40329 ( .A(n37742), .B(n37743), .Z(n37733) );
  ANDN U40330 ( .A(n37744), .B(n29273), .Z(n37743) );
  XOR U40331 ( .A(n37745), .B(\modmult_1/zin[0][244] ), .Z(n29273) );
  IV U40332 ( .A(n37742), .Z(n37745) );
  XNOR U40333 ( .A(n37742), .B(n29272), .Z(n37744) );
  XOR U40334 ( .A(n37746), .B(n37747), .Z(n29272) );
  AND U40335 ( .A(\modmult_1/xin[1023] ), .B(n37748), .Z(n37747) );
  IV U40336 ( .A(n37746), .Z(n37748) );
  XOR U40337 ( .A(n37749), .B(mreg[245]), .Z(n37746) );
  NAND U40338 ( .A(n37750), .B(mul_pow), .Z(n37749) );
  XOR U40339 ( .A(mreg[245]), .B(creg[245]), .Z(n37750) );
  XOR U40340 ( .A(n37751), .B(n37752), .Z(n37742) );
  ANDN U40341 ( .A(n37753), .B(n29279), .Z(n37752) );
  XOR U40342 ( .A(n37754), .B(\modmult_1/zin[0][243] ), .Z(n29279) );
  IV U40343 ( .A(n37751), .Z(n37754) );
  XNOR U40344 ( .A(n37751), .B(n29278), .Z(n37753) );
  XOR U40345 ( .A(n37755), .B(n37756), .Z(n29278) );
  AND U40346 ( .A(\modmult_1/xin[1023] ), .B(n37757), .Z(n37756) );
  IV U40347 ( .A(n37755), .Z(n37757) );
  XOR U40348 ( .A(n37758), .B(mreg[244]), .Z(n37755) );
  NAND U40349 ( .A(n37759), .B(mul_pow), .Z(n37758) );
  XOR U40350 ( .A(mreg[244]), .B(creg[244]), .Z(n37759) );
  XOR U40351 ( .A(n37760), .B(n37761), .Z(n37751) );
  ANDN U40352 ( .A(n37762), .B(n29285), .Z(n37761) );
  XOR U40353 ( .A(n37763), .B(\modmult_1/zin[0][242] ), .Z(n29285) );
  IV U40354 ( .A(n37760), .Z(n37763) );
  XNOR U40355 ( .A(n37760), .B(n29284), .Z(n37762) );
  XOR U40356 ( .A(n37764), .B(n37765), .Z(n29284) );
  AND U40357 ( .A(\modmult_1/xin[1023] ), .B(n37766), .Z(n37765) );
  IV U40358 ( .A(n37764), .Z(n37766) );
  XOR U40359 ( .A(n37767), .B(mreg[243]), .Z(n37764) );
  NAND U40360 ( .A(n37768), .B(mul_pow), .Z(n37767) );
  XOR U40361 ( .A(mreg[243]), .B(creg[243]), .Z(n37768) );
  XOR U40362 ( .A(n37769), .B(n37770), .Z(n37760) );
  ANDN U40363 ( .A(n37771), .B(n29291), .Z(n37770) );
  XOR U40364 ( .A(n37772), .B(\modmult_1/zin[0][241] ), .Z(n29291) );
  IV U40365 ( .A(n37769), .Z(n37772) );
  XNOR U40366 ( .A(n37769), .B(n29290), .Z(n37771) );
  XOR U40367 ( .A(n37773), .B(n37774), .Z(n29290) );
  AND U40368 ( .A(\modmult_1/xin[1023] ), .B(n37775), .Z(n37774) );
  IV U40369 ( .A(n37773), .Z(n37775) );
  XOR U40370 ( .A(n37776), .B(mreg[242]), .Z(n37773) );
  NAND U40371 ( .A(n37777), .B(mul_pow), .Z(n37776) );
  XOR U40372 ( .A(mreg[242]), .B(creg[242]), .Z(n37777) );
  XOR U40373 ( .A(n37778), .B(n37779), .Z(n37769) );
  ANDN U40374 ( .A(n37780), .B(n29297), .Z(n37779) );
  XOR U40375 ( .A(n37781), .B(\modmult_1/zin[0][240] ), .Z(n29297) );
  IV U40376 ( .A(n37778), .Z(n37781) );
  XNOR U40377 ( .A(n37778), .B(n29296), .Z(n37780) );
  XOR U40378 ( .A(n37782), .B(n37783), .Z(n29296) );
  AND U40379 ( .A(\modmult_1/xin[1023] ), .B(n37784), .Z(n37783) );
  IV U40380 ( .A(n37782), .Z(n37784) );
  XOR U40381 ( .A(n37785), .B(mreg[241]), .Z(n37782) );
  NAND U40382 ( .A(n37786), .B(mul_pow), .Z(n37785) );
  XOR U40383 ( .A(mreg[241]), .B(creg[241]), .Z(n37786) );
  XOR U40384 ( .A(n37787), .B(n37788), .Z(n37778) );
  ANDN U40385 ( .A(n37789), .B(n29303), .Z(n37788) );
  XOR U40386 ( .A(n37790), .B(\modmult_1/zin[0][239] ), .Z(n29303) );
  IV U40387 ( .A(n37787), .Z(n37790) );
  XNOR U40388 ( .A(n37787), .B(n29302), .Z(n37789) );
  XOR U40389 ( .A(n37791), .B(n37792), .Z(n29302) );
  AND U40390 ( .A(\modmult_1/xin[1023] ), .B(n37793), .Z(n37792) );
  IV U40391 ( .A(n37791), .Z(n37793) );
  XOR U40392 ( .A(n37794), .B(mreg[240]), .Z(n37791) );
  NAND U40393 ( .A(n37795), .B(mul_pow), .Z(n37794) );
  XOR U40394 ( .A(mreg[240]), .B(creg[240]), .Z(n37795) );
  XOR U40395 ( .A(n37796), .B(n37797), .Z(n37787) );
  ANDN U40396 ( .A(n37798), .B(n29309), .Z(n37797) );
  XOR U40397 ( .A(n37799), .B(\modmult_1/zin[0][238] ), .Z(n29309) );
  IV U40398 ( .A(n37796), .Z(n37799) );
  XNOR U40399 ( .A(n37796), .B(n29308), .Z(n37798) );
  XOR U40400 ( .A(n37800), .B(n37801), .Z(n29308) );
  AND U40401 ( .A(\modmult_1/xin[1023] ), .B(n37802), .Z(n37801) );
  IV U40402 ( .A(n37800), .Z(n37802) );
  XOR U40403 ( .A(n37803), .B(mreg[239]), .Z(n37800) );
  NAND U40404 ( .A(n37804), .B(mul_pow), .Z(n37803) );
  XOR U40405 ( .A(mreg[239]), .B(creg[239]), .Z(n37804) );
  XOR U40406 ( .A(n37805), .B(n37806), .Z(n37796) );
  ANDN U40407 ( .A(n37807), .B(n29315), .Z(n37806) );
  XOR U40408 ( .A(n37808), .B(\modmult_1/zin[0][237] ), .Z(n29315) );
  IV U40409 ( .A(n37805), .Z(n37808) );
  XNOR U40410 ( .A(n37805), .B(n29314), .Z(n37807) );
  XOR U40411 ( .A(n37809), .B(n37810), .Z(n29314) );
  AND U40412 ( .A(\modmult_1/xin[1023] ), .B(n37811), .Z(n37810) );
  IV U40413 ( .A(n37809), .Z(n37811) );
  XOR U40414 ( .A(n37812), .B(mreg[238]), .Z(n37809) );
  NAND U40415 ( .A(n37813), .B(mul_pow), .Z(n37812) );
  XOR U40416 ( .A(mreg[238]), .B(creg[238]), .Z(n37813) );
  XOR U40417 ( .A(n37814), .B(n37815), .Z(n37805) );
  ANDN U40418 ( .A(n37816), .B(n29321), .Z(n37815) );
  XOR U40419 ( .A(n37817), .B(\modmult_1/zin[0][236] ), .Z(n29321) );
  IV U40420 ( .A(n37814), .Z(n37817) );
  XNOR U40421 ( .A(n37814), .B(n29320), .Z(n37816) );
  XOR U40422 ( .A(n37818), .B(n37819), .Z(n29320) );
  AND U40423 ( .A(\modmult_1/xin[1023] ), .B(n37820), .Z(n37819) );
  IV U40424 ( .A(n37818), .Z(n37820) );
  XOR U40425 ( .A(n37821), .B(mreg[237]), .Z(n37818) );
  NAND U40426 ( .A(n37822), .B(mul_pow), .Z(n37821) );
  XOR U40427 ( .A(mreg[237]), .B(creg[237]), .Z(n37822) );
  XOR U40428 ( .A(n37823), .B(n37824), .Z(n37814) );
  ANDN U40429 ( .A(n37825), .B(n29327), .Z(n37824) );
  XOR U40430 ( .A(n37826), .B(\modmult_1/zin[0][235] ), .Z(n29327) );
  IV U40431 ( .A(n37823), .Z(n37826) );
  XNOR U40432 ( .A(n37823), .B(n29326), .Z(n37825) );
  XOR U40433 ( .A(n37827), .B(n37828), .Z(n29326) );
  AND U40434 ( .A(\modmult_1/xin[1023] ), .B(n37829), .Z(n37828) );
  IV U40435 ( .A(n37827), .Z(n37829) );
  XOR U40436 ( .A(n37830), .B(mreg[236]), .Z(n37827) );
  NAND U40437 ( .A(n37831), .B(mul_pow), .Z(n37830) );
  XOR U40438 ( .A(mreg[236]), .B(creg[236]), .Z(n37831) );
  XOR U40439 ( .A(n37832), .B(n37833), .Z(n37823) );
  ANDN U40440 ( .A(n37834), .B(n29333), .Z(n37833) );
  XOR U40441 ( .A(n37835), .B(\modmult_1/zin[0][234] ), .Z(n29333) );
  IV U40442 ( .A(n37832), .Z(n37835) );
  XNOR U40443 ( .A(n37832), .B(n29332), .Z(n37834) );
  XOR U40444 ( .A(n37836), .B(n37837), .Z(n29332) );
  AND U40445 ( .A(\modmult_1/xin[1023] ), .B(n37838), .Z(n37837) );
  IV U40446 ( .A(n37836), .Z(n37838) );
  XOR U40447 ( .A(n37839), .B(mreg[235]), .Z(n37836) );
  NAND U40448 ( .A(n37840), .B(mul_pow), .Z(n37839) );
  XOR U40449 ( .A(mreg[235]), .B(creg[235]), .Z(n37840) );
  XOR U40450 ( .A(n37841), .B(n37842), .Z(n37832) );
  ANDN U40451 ( .A(n37843), .B(n29339), .Z(n37842) );
  XOR U40452 ( .A(n37844), .B(\modmult_1/zin[0][233] ), .Z(n29339) );
  IV U40453 ( .A(n37841), .Z(n37844) );
  XNOR U40454 ( .A(n37841), .B(n29338), .Z(n37843) );
  XOR U40455 ( .A(n37845), .B(n37846), .Z(n29338) );
  AND U40456 ( .A(\modmult_1/xin[1023] ), .B(n37847), .Z(n37846) );
  IV U40457 ( .A(n37845), .Z(n37847) );
  XOR U40458 ( .A(n37848), .B(mreg[234]), .Z(n37845) );
  NAND U40459 ( .A(n37849), .B(mul_pow), .Z(n37848) );
  XOR U40460 ( .A(mreg[234]), .B(creg[234]), .Z(n37849) );
  XOR U40461 ( .A(n37850), .B(n37851), .Z(n37841) );
  ANDN U40462 ( .A(n37852), .B(n29345), .Z(n37851) );
  XOR U40463 ( .A(n37853), .B(\modmult_1/zin[0][232] ), .Z(n29345) );
  IV U40464 ( .A(n37850), .Z(n37853) );
  XNOR U40465 ( .A(n37850), .B(n29344), .Z(n37852) );
  XOR U40466 ( .A(n37854), .B(n37855), .Z(n29344) );
  AND U40467 ( .A(\modmult_1/xin[1023] ), .B(n37856), .Z(n37855) );
  IV U40468 ( .A(n37854), .Z(n37856) );
  XOR U40469 ( .A(n37857), .B(mreg[233]), .Z(n37854) );
  NAND U40470 ( .A(n37858), .B(mul_pow), .Z(n37857) );
  XOR U40471 ( .A(mreg[233]), .B(creg[233]), .Z(n37858) );
  XOR U40472 ( .A(n37859), .B(n37860), .Z(n37850) );
  ANDN U40473 ( .A(n37861), .B(n29351), .Z(n37860) );
  XOR U40474 ( .A(n37862), .B(\modmult_1/zin[0][231] ), .Z(n29351) );
  IV U40475 ( .A(n37859), .Z(n37862) );
  XNOR U40476 ( .A(n37859), .B(n29350), .Z(n37861) );
  XOR U40477 ( .A(n37863), .B(n37864), .Z(n29350) );
  AND U40478 ( .A(\modmult_1/xin[1023] ), .B(n37865), .Z(n37864) );
  IV U40479 ( .A(n37863), .Z(n37865) );
  XOR U40480 ( .A(n37866), .B(mreg[232]), .Z(n37863) );
  NAND U40481 ( .A(n37867), .B(mul_pow), .Z(n37866) );
  XOR U40482 ( .A(mreg[232]), .B(creg[232]), .Z(n37867) );
  XOR U40483 ( .A(n37868), .B(n37869), .Z(n37859) );
  ANDN U40484 ( .A(n37870), .B(n29357), .Z(n37869) );
  XOR U40485 ( .A(n37871), .B(\modmult_1/zin[0][230] ), .Z(n29357) );
  IV U40486 ( .A(n37868), .Z(n37871) );
  XNOR U40487 ( .A(n37868), .B(n29356), .Z(n37870) );
  XOR U40488 ( .A(n37872), .B(n37873), .Z(n29356) );
  AND U40489 ( .A(\modmult_1/xin[1023] ), .B(n37874), .Z(n37873) );
  IV U40490 ( .A(n37872), .Z(n37874) );
  XOR U40491 ( .A(n37875), .B(mreg[231]), .Z(n37872) );
  NAND U40492 ( .A(n37876), .B(mul_pow), .Z(n37875) );
  XOR U40493 ( .A(mreg[231]), .B(creg[231]), .Z(n37876) );
  XOR U40494 ( .A(n37877), .B(n37878), .Z(n37868) );
  ANDN U40495 ( .A(n37879), .B(n29363), .Z(n37878) );
  XOR U40496 ( .A(n37880), .B(\modmult_1/zin[0][229] ), .Z(n29363) );
  IV U40497 ( .A(n37877), .Z(n37880) );
  XNOR U40498 ( .A(n37877), .B(n29362), .Z(n37879) );
  XOR U40499 ( .A(n37881), .B(n37882), .Z(n29362) );
  AND U40500 ( .A(\modmult_1/xin[1023] ), .B(n37883), .Z(n37882) );
  IV U40501 ( .A(n37881), .Z(n37883) );
  XOR U40502 ( .A(n37884), .B(mreg[230]), .Z(n37881) );
  NAND U40503 ( .A(n37885), .B(mul_pow), .Z(n37884) );
  XOR U40504 ( .A(mreg[230]), .B(creg[230]), .Z(n37885) );
  XOR U40505 ( .A(n37886), .B(n37887), .Z(n37877) );
  ANDN U40506 ( .A(n37888), .B(n29369), .Z(n37887) );
  XOR U40507 ( .A(n37889), .B(\modmult_1/zin[0][228] ), .Z(n29369) );
  IV U40508 ( .A(n37886), .Z(n37889) );
  XNOR U40509 ( .A(n37886), .B(n29368), .Z(n37888) );
  XOR U40510 ( .A(n37890), .B(n37891), .Z(n29368) );
  AND U40511 ( .A(\modmult_1/xin[1023] ), .B(n37892), .Z(n37891) );
  IV U40512 ( .A(n37890), .Z(n37892) );
  XOR U40513 ( .A(n37893), .B(mreg[229]), .Z(n37890) );
  NAND U40514 ( .A(n37894), .B(mul_pow), .Z(n37893) );
  XOR U40515 ( .A(mreg[229]), .B(creg[229]), .Z(n37894) );
  XOR U40516 ( .A(n37895), .B(n37896), .Z(n37886) );
  ANDN U40517 ( .A(n37897), .B(n29375), .Z(n37896) );
  XOR U40518 ( .A(n37898), .B(\modmult_1/zin[0][227] ), .Z(n29375) );
  IV U40519 ( .A(n37895), .Z(n37898) );
  XNOR U40520 ( .A(n37895), .B(n29374), .Z(n37897) );
  XOR U40521 ( .A(n37899), .B(n37900), .Z(n29374) );
  AND U40522 ( .A(\modmult_1/xin[1023] ), .B(n37901), .Z(n37900) );
  IV U40523 ( .A(n37899), .Z(n37901) );
  XOR U40524 ( .A(n37902), .B(mreg[228]), .Z(n37899) );
  NAND U40525 ( .A(n37903), .B(mul_pow), .Z(n37902) );
  XOR U40526 ( .A(mreg[228]), .B(creg[228]), .Z(n37903) );
  XOR U40527 ( .A(n37904), .B(n37905), .Z(n37895) );
  ANDN U40528 ( .A(n37906), .B(n29381), .Z(n37905) );
  XOR U40529 ( .A(n37907), .B(\modmult_1/zin[0][226] ), .Z(n29381) );
  IV U40530 ( .A(n37904), .Z(n37907) );
  XNOR U40531 ( .A(n37904), .B(n29380), .Z(n37906) );
  XOR U40532 ( .A(n37908), .B(n37909), .Z(n29380) );
  AND U40533 ( .A(\modmult_1/xin[1023] ), .B(n37910), .Z(n37909) );
  IV U40534 ( .A(n37908), .Z(n37910) );
  XOR U40535 ( .A(n37911), .B(mreg[227]), .Z(n37908) );
  NAND U40536 ( .A(n37912), .B(mul_pow), .Z(n37911) );
  XOR U40537 ( .A(mreg[227]), .B(creg[227]), .Z(n37912) );
  XOR U40538 ( .A(n37913), .B(n37914), .Z(n37904) );
  ANDN U40539 ( .A(n37915), .B(n29387), .Z(n37914) );
  XOR U40540 ( .A(n37916), .B(\modmult_1/zin[0][225] ), .Z(n29387) );
  IV U40541 ( .A(n37913), .Z(n37916) );
  XNOR U40542 ( .A(n37913), .B(n29386), .Z(n37915) );
  XOR U40543 ( .A(n37917), .B(n37918), .Z(n29386) );
  AND U40544 ( .A(\modmult_1/xin[1023] ), .B(n37919), .Z(n37918) );
  IV U40545 ( .A(n37917), .Z(n37919) );
  XOR U40546 ( .A(n37920), .B(mreg[226]), .Z(n37917) );
  NAND U40547 ( .A(n37921), .B(mul_pow), .Z(n37920) );
  XOR U40548 ( .A(mreg[226]), .B(creg[226]), .Z(n37921) );
  XOR U40549 ( .A(n37922), .B(n37923), .Z(n37913) );
  ANDN U40550 ( .A(n37924), .B(n29393), .Z(n37923) );
  XOR U40551 ( .A(n37925), .B(\modmult_1/zin[0][224] ), .Z(n29393) );
  IV U40552 ( .A(n37922), .Z(n37925) );
  XNOR U40553 ( .A(n37922), .B(n29392), .Z(n37924) );
  XOR U40554 ( .A(n37926), .B(n37927), .Z(n29392) );
  AND U40555 ( .A(\modmult_1/xin[1023] ), .B(n37928), .Z(n37927) );
  IV U40556 ( .A(n37926), .Z(n37928) );
  XOR U40557 ( .A(n37929), .B(mreg[225]), .Z(n37926) );
  NAND U40558 ( .A(n37930), .B(mul_pow), .Z(n37929) );
  XOR U40559 ( .A(mreg[225]), .B(creg[225]), .Z(n37930) );
  XOR U40560 ( .A(n37931), .B(n37932), .Z(n37922) );
  ANDN U40561 ( .A(n37933), .B(n29399), .Z(n37932) );
  XOR U40562 ( .A(n37934), .B(\modmult_1/zin[0][223] ), .Z(n29399) );
  IV U40563 ( .A(n37931), .Z(n37934) );
  XNOR U40564 ( .A(n37931), .B(n29398), .Z(n37933) );
  XOR U40565 ( .A(n37935), .B(n37936), .Z(n29398) );
  AND U40566 ( .A(\modmult_1/xin[1023] ), .B(n37937), .Z(n37936) );
  IV U40567 ( .A(n37935), .Z(n37937) );
  XOR U40568 ( .A(n37938), .B(mreg[224]), .Z(n37935) );
  NAND U40569 ( .A(n37939), .B(mul_pow), .Z(n37938) );
  XOR U40570 ( .A(mreg[224]), .B(creg[224]), .Z(n37939) );
  XOR U40571 ( .A(n37940), .B(n37941), .Z(n37931) );
  ANDN U40572 ( .A(n37942), .B(n29405), .Z(n37941) );
  XOR U40573 ( .A(n37943), .B(\modmult_1/zin[0][222] ), .Z(n29405) );
  IV U40574 ( .A(n37940), .Z(n37943) );
  XNOR U40575 ( .A(n37940), .B(n29404), .Z(n37942) );
  XOR U40576 ( .A(n37944), .B(n37945), .Z(n29404) );
  AND U40577 ( .A(\modmult_1/xin[1023] ), .B(n37946), .Z(n37945) );
  IV U40578 ( .A(n37944), .Z(n37946) );
  XOR U40579 ( .A(n37947), .B(mreg[223]), .Z(n37944) );
  NAND U40580 ( .A(n37948), .B(mul_pow), .Z(n37947) );
  XOR U40581 ( .A(mreg[223]), .B(creg[223]), .Z(n37948) );
  XOR U40582 ( .A(n37949), .B(n37950), .Z(n37940) );
  ANDN U40583 ( .A(n37951), .B(n29411), .Z(n37950) );
  XOR U40584 ( .A(n37952), .B(\modmult_1/zin[0][221] ), .Z(n29411) );
  IV U40585 ( .A(n37949), .Z(n37952) );
  XNOR U40586 ( .A(n37949), .B(n29410), .Z(n37951) );
  XOR U40587 ( .A(n37953), .B(n37954), .Z(n29410) );
  AND U40588 ( .A(\modmult_1/xin[1023] ), .B(n37955), .Z(n37954) );
  IV U40589 ( .A(n37953), .Z(n37955) );
  XOR U40590 ( .A(n37956), .B(mreg[222]), .Z(n37953) );
  NAND U40591 ( .A(n37957), .B(mul_pow), .Z(n37956) );
  XOR U40592 ( .A(mreg[222]), .B(creg[222]), .Z(n37957) );
  XOR U40593 ( .A(n37958), .B(n37959), .Z(n37949) );
  ANDN U40594 ( .A(n37960), .B(n29417), .Z(n37959) );
  XOR U40595 ( .A(n37961), .B(\modmult_1/zin[0][220] ), .Z(n29417) );
  IV U40596 ( .A(n37958), .Z(n37961) );
  XNOR U40597 ( .A(n37958), .B(n29416), .Z(n37960) );
  XOR U40598 ( .A(n37962), .B(n37963), .Z(n29416) );
  AND U40599 ( .A(\modmult_1/xin[1023] ), .B(n37964), .Z(n37963) );
  IV U40600 ( .A(n37962), .Z(n37964) );
  XOR U40601 ( .A(n37965), .B(mreg[221]), .Z(n37962) );
  NAND U40602 ( .A(n37966), .B(mul_pow), .Z(n37965) );
  XOR U40603 ( .A(mreg[221]), .B(creg[221]), .Z(n37966) );
  XOR U40604 ( .A(n37967), .B(n37968), .Z(n37958) );
  ANDN U40605 ( .A(n37969), .B(n29423), .Z(n37968) );
  XOR U40606 ( .A(n37970), .B(\modmult_1/zin[0][219] ), .Z(n29423) );
  IV U40607 ( .A(n37967), .Z(n37970) );
  XNOR U40608 ( .A(n37967), .B(n29422), .Z(n37969) );
  XOR U40609 ( .A(n37971), .B(n37972), .Z(n29422) );
  AND U40610 ( .A(\modmult_1/xin[1023] ), .B(n37973), .Z(n37972) );
  IV U40611 ( .A(n37971), .Z(n37973) );
  XOR U40612 ( .A(n37974), .B(mreg[220]), .Z(n37971) );
  NAND U40613 ( .A(n37975), .B(mul_pow), .Z(n37974) );
  XOR U40614 ( .A(mreg[220]), .B(creg[220]), .Z(n37975) );
  XOR U40615 ( .A(n37976), .B(n37977), .Z(n37967) );
  ANDN U40616 ( .A(n37978), .B(n29429), .Z(n37977) );
  XOR U40617 ( .A(n37979), .B(\modmult_1/zin[0][218] ), .Z(n29429) );
  IV U40618 ( .A(n37976), .Z(n37979) );
  XNOR U40619 ( .A(n37976), .B(n29428), .Z(n37978) );
  XOR U40620 ( .A(n37980), .B(n37981), .Z(n29428) );
  AND U40621 ( .A(\modmult_1/xin[1023] ), .B(n37982), .Z(n37981) );
  IV U40622 ( .A(n37980), .Z(n37982) );
  XOR U40623 ( .A(n37983), .B(mreg[219]), .Z(n37980) );
  NAND U40624 ( .A(n37984), .B(mul_pow), .Z(n37983) );
  XOR U40625 ( .A(mreg[219]), .B(creg[219]), .Z(n37984) );
  XOR U40626 ( .A(n37985), .B(n37986), .Z(n37976) );
  ANDN U40627 ( .A(n37987), .B(n29435), .Z(n37986) );
  XOR U40628 ( .A(n37988), .B(\modmult_1/zin[0][217] ), .Z(n29435) );
  IV U40629 ( .A(n37985), .Z(n37988) );
  XNOR U40630 ( .A(n37985), .B(n29434), .Z(n37987) );
  XOR U40631 ( .A(n37989), .B(n37990), .Z(n29434) );
  AND U40632 ( .A(\modmult_1/xin[1023] ), .B(n37991), .Z(n37990) );
  IV U40633 ( .A(n37989), .Z(n37991) );
  XOR U40634 ( .A(n37992), .B(mreg[218]), .Z(n37989) );
  NAND U40635 ( .A(n37993), .B(mul_pow), .Z(n37992) );
  XOR U40636 ( .A(mreg[218]), .B(creg[218]), .Z(n37993) );
  XOR U40637 ( .A(n37994), .B(n37995), .Z(n37985) );
  ANDN U40638 ( .A(n37996), .B(n29441), .Z(n37995) );
  XOR U40639 ( .A(n37997), .B(\modmult_1/zin[0][216] ), .Z(n29441) );
  IV U40640 ( .A(n37994), .Z(n37997) );
  XNOR U40641 ( .A(n37994), .B(n29440), .Z(n37996) );
  XOR U40642 ( .A(n37998), .B(n37999), .Z(n29440) );
  AND U40643 ( .A(\modmult_1/xin[1023] ), .B(n38000), .Z(n37999) );
  IV U40644 ( .A(n37998), .Z(n38000) );
  XOR U40645 ( .A(n38001), .B(mreg[217]), .Z(n37998) );
  NAND U40646 ( .A(n38002), .B(mul_pow), .Z(n38001) );
  XOR U40647 ( .A(mreg[217]), .B(creg[217]), .Z(n38002) );
  XOR U40648 ( .A(n38003), .B(n38004), .Z(n37994) );
  ANDN U40649 ( .A(n38005), .B(n29447), .Z(n38004) );
  XOR U40650 ( .A(n38006), .B(\modmult_1/zin[0][215] ), .Z(n29447) );
  IV U40651 ( .A(n38003), .Z(n38006) );
  XNOR U40652 ( .A(n38003), .B(n29446), .Z(n38005) );
  XOR U40653 ( .A(n38007), .B(n38008), .Z(n29446) );
  AND U40654 ( .A(\modmult_1/xin[1023] ), .B(n38009), .Z(n38008) );
  IV U40655 ( .A(n38007), .Z(n38009) );
  XOR U40656 ( .A(n38010), .B(mreg[216]), .Z(n38007) );
  NAND U40657 ( .A(n38011), .B(mul_pow), .Z(n38010) );
  XOR U40658 ( .A(mreg[216]), .B(creg[216]), .Z(n38011) );
  XOR U40659 ( .A(n38012), .B(n38013), .Z(n38003) );
  ANDN U40660 ( .A(n38014), .B(n29453), .Z(n38013) );
  XOR U40661 ( .A(n38015), .B(\modmult_1/zin[0][214] ), .Z(n29453) );
  IV U40662 ( .A(n38012), .Z(n38015) );
  XNOR U40663 ( .A(n38012), .B(n29452), .Z(n38014) );
  XOR U40664 ( .A(n38016), .B(n38017), .Z(n29452) );
  AND U40665 ( .A(\modmult_1/xin[1023] ), .B(n38018), .Z(n38017) );
  IV U40666 ( .A(n38016), .Z(n38018) );
  XOR U40667 ( .A(n38019), .B(mreg[215]), .Z(n38016) );
  NAND U40668 ( .A(n38020), .B(mul_pow), .Z(n38019) );
  XOR U40669 ( .A(mreg[215]), .B(creg[215]), .Z(n38020) );
  XOR U40670 ( .A(n38021), .B(n38022), .Z(n38012) );
  ANDN U40671 ( .A(n38023), .B(n29459), .Z(n38022) );
  XOR U40672 ( .A(n38024), .B(\modmult_1/zin[0][213] ), .Z(n29459) );
  IV U40673 ( .A(n38021), .Z(n38024) );
  XNOR U40674 ( .A(n38021), .B(n29458), .Z(n38023) );
  XOR U40675 ( .A(n38025), .B(n38026), .Z(n29458) );
  AND U40676 ( .A(\modmult_1/xin[1023] ), .B(n38027), .Z(n38026) );
  IV U40677 ( .A(n38025), .Z(n38027) );
  XOR U40678 ( .A(n38028), .B(mreg[214]), .Z(n38025) );
  NAND U40679 ( .A(n38029), .B(mul_pow), .Z(n38028) );
  XOR U40680 ( .A(mreg[214]), .B(creg[214]), .Z(n38029) );
  XOR U40681 ( .A(n38030), .B(n38031), .Z(n38021) );
  ANDN U40682 ( .A(n38032), .B(n29465), .Z(n38031) );
  XOR U40683 ( .A(n38033), .B(\modmult_1/zin[0][212] ), .Z(n29465) );
  IV U40684 ( .A(n38030), .Z(n38033) );
  XNOR U40685 ( .A(n38030), .B(n29464), .Z(n38032) );
  XOR U40686 ( .A(n38034), .B(n38035), .Z(n29464) );
  AND U40687 ( .A(\modmult_1/xin[1023] ), .B(n38036), .Z(n38035) );
  IV U40688 ( .A(n38034), .Z(n38036) );
  XOR U40689 ( .A(n38037), .B(mreg[213]), .Z(n38034) );
  NAND U40690 ( .A(n38038), .B(mul_pow), .Z(n38037) );
  XOR U40691 ( .A(mreg[213]), .B(creg[213]), .Z(n38038) );
  XOR U40692 ( .A(n38039), .B(n38040), .Z(n38030) );
  ANDN U40693 ( .A(n38041), .B(n29471), .Z(n38040) );
  XOR U40694 ( .A(n38042), .B(\modmult_1/zin[0][211] ), .Z(n29471) );
  IV U40695 ( .A(n38039), .Z(n38042) );
  XNOR U40696 ( .A(n38039), .B(n29470), .Z(n38041) );
  XOR U40697 ( .A(n38043), .B(n38044), .Z(n29470) );
  AND U40698 ( .A(\modmult_1/xin[1023] ), .B(n38045), .Z(n38044) );
  IV U40699 ( .A(n38043), .Z(n38045) );
  XOR U40700 ( .A(n38046), .B(mreg[212]), .Z(n38043) );
  NAND U40701 ( .A(n38047), .B(mul_pow), .Z(n38046) );
  XOR U40702 ( .A(mreg[212]), .B(creg[212]), .Z(n38047) );
  XOR U40703 ( .A(n38048), .B(n38049), .Z(n38039) );
  ANDN U40704 ( .A(n38050), .B(n29477), .Z(n38049) );
  XOR U40705 ( .A(n38051), .B(\modmult_1/zin[0][210] ), .Z(n29477) );
  IV U40706 ( .A(n38048), .Z(n38051) );
  XNOR U40707 ( .A(n38048), .B(n29476), .Z(n38050) );
  XOR U40708 ( .A(n38052), .B(n38053), .Z(n29476) );
  AND U40709 ( .A(\modmult_1/xin[1023] ), .B(n38054), .Z(n38053) );
  IV U40710 ( .A(n38052), .Z(n38054) );
  XOR U40711 ( .A(n38055), .B(mreg[211]), .Z(n38052) );
  NAND U40712 ( .A(n38056), .B(mul_pow), .Z(n38055) );
  XOR U40713 ( .A(mreg[211]), .B(creg[211]), .Z(n38056) );
  XOR U40714 ( .A(n38057), .B(n38058), .Z(n38048) );
  ANDN U40715 ( .A(n38059), .B(n29483), .Z(n38058) );
  XOR U40716 ( .A(n38060), .B(\modmult_1/zin[0][209] ), .Z(n29483) );
  IV U40717 ( .A(n38057), .Z(n38060) );
  XNOR U40718 ( .A(n38057), .B(n29482), .Z(n38059) );
  XOR U40719 ( .A(n38061), .B(n38062), .Z(n29482) );
  AND U40720 ( .A(\modmult_1/xin[1023] ), .B(n38063), .Z(n38062) );
  IV U40721 ( .A(n38061), .Z(n38063) );
  XOR U40722 ( .A(n38064), .B(mreg[210]), .Z(n38061) );
  NAND U40723 ( .A(n38065), .B(mul_pow), .Z(n38064) );
  XOR U40724 ( .A(mreg[210]), .B(creg[210]), .Z(n38065) );
  XOR U40725 ( .A(n38066), .B(n38067), .Z(n38057) );
  ANDN U40726 ( .A(n38068), .B(n29489), .Z(n38067) );
  XOR U40727 ( .A(n38069), .B(\modmult_1/zin[0][208] ), .Z(n29489) );
  IV U40728 ( .A(n38066), .Z(n38069) );
  XNOR U40729 ( .A(n38066), .B(n29488), .Z(n38068) );
  XOR U40730 ( .A(n38070), .B(n38071), .Z(n29488) );
  AND U40731 ( .A(\modmult_1/xin[1023] ), .B(n38072), .Z(n38071) );
  IV U40732 ( .A(n38070), .Z(n38072) );
  XOR U40733 ( .A(n38073), .B(mreg[209]), .Z(n38070) );
  NAND U40734 ( .A(n38074), .B(mul_pow), .Z(n38073) );
  XOR U40735 ( .A(mreg[209]), .B(creg[209]), .Z(n38074) );
  XOR U40736 ( .A(n38075), .B(n38076), .Z(n38066) );
  ANDN U40737 ( .A(n38077), .B(n29495), .Z(n38076) );
  XOR U40738 ( .A(n38078), .B(\modmult_1/zin[0][207] ), .Z(n29495) );
  IV U40739 ( .A(n38075), .Z(n38078) );
  XNOR U40740 ( .A(n38075), .B(n29494), .Z(n38077) );
  XOR U40741 ( .A(n38079), .B(n38080), .Z(n29494) );
  AND U40742 ( .A(\modmult_1/xin[1023] ), .B(n38081), .Z(n38080) );
  IV U40743 ( .A(n38079), .Z(n38081) );
  XOR U40744 ( .A(n38082), .B(mreg[208]), .Z(n38079) );
  NAND U40745 ( .A(n38083), .B(mul_pow), .Z(n38082) );
  XOR U40746 ( .A(mreg[208]), .B(creg[208]), .Z(n38083) );
  XOR U40747 ( .A(n38084), .B(n38085), .Z(n38075) );
  ANDN U40748 ( .A(n38086), .B(n29501), .Z(n38085) );
  XOR U40749 ( .A(n38087), .B(\modmult_1/zin[0][206] ), .Z(n29501) );
  IV U40750 ( .A(n38084), .Z(n38087) );
  XNOR U40751 ( .A(n38084), .B(n29500), .Z(n38086) );
  XOR U40752 ( .A(n38088), .B(n38089), .Z(n29500) );
  AND U40753 ( .A(\modmult_1/xin[1023] ), .B(n38090), .Z(n38089) );
  IV U40754 ( .A(n38088), .Z(n38090) );
  XOR U40755 ( .A(n38091), .B(mreg[207]), .Z(n38088) );
  NAND U40756 ( .A(n38092), .B(mul_pow), .Z(n38091) );
  XOR U40757 ( .A(mreg[207]), .B(creg[207]), .Z(n38092) );
  XOR U40758 ( .A(n38093), .B(n38094), .Z(n38084) );
  ANDN U40759 ( .A(n38095), .B(n29507), .Z(n38094) );
  XOR U40760 ( .A(n38096), .B(\modmult_1/zin[0][205] ), .Z(n29507) );
  IV U40761 ( .A(n38093), .Z(n38096) );
  XNOR U40762 ( .A(n38093), .B(n29506), .Z(n38095) );
  XOR U40763 ( .A(n38097), .B(n38098), .Z(n29506) );
  AND U40764 ( .A(\modmult_1/xin[1023] ), .B(n38099), .Z(n38098) );
  IV U40765 ( .A(n38097), .Z(n38099) );
  XOR U40766 ( .A(n38100), .B(mreg[206]), .Z(n38097) );
  NAND U40767 ( .A(n38101), .B(mul_pow), .Z(n38100) );
  XOR U40768 ( .A(mreg[206]), .B(creg[206]), .Z(n38101) );
  XOR U40769 ( .A(n38102), .B(n38103), .Z(n38093) );
  ANDN U40770 ( .A(n38104), .B(n29513), .Z(n38103) );
  XOR U40771 ( .A(n38105), .B(\modmult_1/zin[0][204] ), .Z(n29513) );
  IV U40772 ( .A(n38102), .Z(n38105) );
  XNOR U40773 ( .A(n38102), .B(n29512), .Z(n38104) );
  XOR U40774 ( .A(n38106), .B(n38107), .Z(n29512) );
  AND U40775 ( .A(\modmult_1/xin[1023] ), .B(n38108), .Z(n38107) );
  IV U40776 ( .A(n38106), .Z(n38108) );
  XOR U40777 ( .A(n38109), .B(mreg[205]), .Z(n38106) );
  NAND U40778 ( .A(n38110), .B(mul_pow), .Z(n38109) );
  XOR U40779 ( .A(mreg[205]), .B(creg[205]), .Z(n38110) );
  XOR U40780 ( .A(n38111), .B(n38112), .Z(n38102) );
  ANDN U40781 ( .A(n38113), .B(n29519), .Z(n38112) );
  XOR U40782 ( .A(n38114), .B(\modmult_1/zin[0][203] ), .Z(n29519) );
  IV U40783 ( .A(n38111), .Z(n38114) );
  XNOR U40784 ( .A(n38111), .B(n29518), .Z(n38113) );
  XOR U40785 ( .A(n38115), .B(n38116), .Z(n29518) );
  AND U40786 ( .A(\modmult_1/xin[1023] ), .B(n38117), .Z(n38116) );
  IV U40787 ( .A(n38115), .Z(n38117) );
  XOR U40788 ( .A(n38118), .B(mreg[204]), .Z(n38115) );
  NAND U40789 ( .A(n38119), .B(mul_pow), .Z(n38118) );
  XOR U40790 ( .A(mreg[204]), .B(creg[204]), .Z(n38119) );
  XOR U40791 ( .A(n38120), .B(n38121), .Z(n38111) );
  ANDN U40792 ( .A(n38122), .B(n29525), .Z(n38121) );
  XOR U40793 ( .A(n38123), .B(\modmult_1/zin[0][202] ), .Z(n29525) );
  IV U40794 ( .A(n38120), .Z(n38123) );
  XNOR U40795 ( .A(n38120), .B(n29524), .Z(n38122) );
  XOR U40796 ( .A(n38124), .B(n38125), .Z(n29524) );
  AND U40797 ( .A(\modmult_1/xin[1023] ), .B(n38126), .Z(n38125) );
  IV U40798 ( .A(n38124), .Z(n38126) );
  XOR U40799 ( .A(n38127), .B(mreg[203]), .Z(n38124) );
  NAND U40800 ( .A(n38128), .B(mul_pow), .Z(n38127) );
  XOR U40801 ( .A(mreg[203]), .B(creg[203]), .Z(n38128) );
  XOR U40802 ( .A(n38129), .B(n38130), .Z(n38120) );
  ANDN U40803 ( .A(n38131), .B(n29531), .Z(n38130) );
  XOR U40804 ( .A(n38132), .B(\modmult_1/zin[0][201] ), .Z(n29531) );
  IV U40805 ( .A(n38129), .Z(n38132) );
  XNOR U40806 ( .A(n38129), .B(n29530), .Z(n38131) );
  XOR U40807 ( .A(n38133), .B(n38134), .Z(n29530) );
  AND U40808 ( .A(\modmult_1/xin[1023] ), .B(n38135), .Z(n38134) );
  IV U40809 ( .A(n38133), .Z(n38135) );
  XOR U40810 ( .A(n38136), .B(mreg[202]), .Z(n38133) );
  NAND U40811 ( .A(n38137), .B(mul_pow), .Z(n38136) );
  XOR U40812 ( .A(mreg[202]), .B(creg[202]), .Z(n38137) );
  XOR U40813 ( .A(n38138), .B(n38139), .Z(n38129) );
  ANDN U40814 ( .A(n38140), .B(n29537), .Z(n38139) );
  XOR U40815 ( .A(n38141), .B(\modmult_1/zin[0][200] ), .Z(n29537) );
  IV U40816 ( .A(n38138), .Z(n38141) );
  XNOR U40817 ( .A(n38138), .B(n29536), .Z(n38140) );
  XOR U40818 ( .A(n38142), .B(n38143), .Z(n29536) );
  AND U40819 ( .A(\modmult_1/xin[1023] ), .B(n38144), .Z(n38143) );
  IV U40820 ( .A(n38142), .Z(n38144) );
  XOR U40821 ( .A(n38145), .B(mreg[201]), .Z(n38142) );
  NAND U40822 ( .A(n38146), .B(mul_pow), .Z(n38145) );
  XOR U40823 ( .A(mreg[201]), .B(creg[201]), .Z(n38146) );
  XOR U40824 ( .A(n38147), .B(n38148), .Z(n38138) );
  ANDN U40825 ( .A(n38149), .B(n29543), .Z(n38148) );
  XOR U40826 ( .A(n38150), .B(\modmult_1/zin[0][199] ), .Z(n29543) );
  IV U40827 ( .A(n38147), .Z(n38150) );
  XNOR U40828 ( .A(n38147), .B(n29542), .Z(n38149) );
  XOR U40829 ( .A(n38151), .B(n38152), .Z(n29542) );
  AND U40830 ( .A(\modmult_1/xin[1023] ), .B(n38153), .Z(n38152) );
  IV U40831 ( .A(n38151), .Z(n38153) );
  XOR U40832 ( .A(n38154), .B(mreg[200]), .Z(n38151) );
  NAND U40833 ( .A(n38155), .B(mul_pow), .Z(n38154) );
  XOR U40834 ( .A(mreg[200]), .B(creg[200]), .Z(n38155) );
  XOR U40835 ( .A(n38156), .B(n38157), .Z(n38147) );
  ANDN U40836 ( .A(n38158), .B(n29549), .Z(n38157) );
  XOR U40837 ( .A(n38159), .B(\modmult_1/zin[0][198] ), .Z(n29549) );
  IV U40838 ( .A(n38156), .Z(n38159) );
  XNOR U40839 ( .A(n38156), .B(n29548), .Z(n38158) );
  XOR U40840 ( .A(n38160), .B(n38161), .Z(n29548) );
  AND U40841 ( .A(\modmult_1/xin[1023] ), .B(n38162), .Z(n38161) );
  IV U40842 ( .A(n38160), .Z(n38162) );
  XOR U40843 ( .A(n38163), .B(mreg[199]), .Z(n38160) );
  NAND U40844 ( .A(n38164), .B(mul_pow), .Z(n38163) );
  XOR U40845 ( .A(mreg[199]), .B(creg[199]), .Z(n38164) );
  XOR U40846 ( .A(n38165), .B(n38166), .Z(n38156) );
  ANDN U40847 ( .A(n38167), .B(n29555), .Z(n38166) );
  XOR U40848 ( .A(n38168), .B(\modmult_1/zin[0][197] ), .Z(n29555) );
  IV U40849 ( .A(n38165), .Z(n38168) );
  XNOR U40850 ( .A(n38165), .B(n29554), .Z(n38167) );
  XOR U40851 ( .A(n38169), .B(n38170), .Z(n29554) );
  AND U40852 ( .A(\modmult_1/xin[1023] ), .B(n38171), .Z(n38170) );
  IV U40853 ( .A(n38169), .Z(n38171) );
  XOR U40854 ( .A(n38172), .B(mreg[198]), .Z(n38169) );
  NAND U40855 ( .A(n38173), .B(mul_pow), .Z(n38172) );
  XOR U40856 ( .A(mreg[198]), .B(creg[198]), .Z(n38173) );
  XOR U40857 ( .A(n38174), .B(n38175), .Z(n38165) );
  ANDN U40858 ( .A(n38176), .B(n29561), .Z(n38175) );
  XOR U40859 ( .A(n38177), .B(\modmult_1/zin[0][196] ), .Z(n29561) );
  IV U40860 ( .A(n38174), .Z(n38177) );
  XNOR U40861 ( .A(n38174), .B(n29560), .Z(n38176) );
  XOR U40862 ( .A(n38178), .B(n38179), .Z(n29560) );
  AND U40863 ( .A(\modmult_1/xin[1023] ), .B(n38180), .Z(n38179) );
  IV U40864 ( .A(n38178), .Z(n38180) );
  XOR U40865 ( .A(n38181), .B(mreg[197]), .Z(n38178) );
  NAND U40866 ( .A(n38182), .B(mul_pow), .Z(n38181) );
  XOR U40867 ( .A(mreg[197]), .B(creg[197]), .Z(n38182) );
  XOR U40868 ( .A(n38183), .B(n38184), .Z(n38174) );
  ANDN U40869 ( .A(n38185), .B(n29567), .Z(n38184) );
  XOR U40870 ( .A(n38186), .B(\modmult_1/zin[0][195] ), .Z(n29567) );
  IV U40871 ( .A(n38183), .Z(n38186) );
  XNOR U40872 ( .A(n38183), .B(n29566), .Z(n38185) );
  XOR U40873 ( .A(n38187), .B(n38188), .Z(n29566) );
  AND U40874 ( .A(\modmult_1/xin[1023] ), .B(n38189), .Z(n38188) );
  IV U40875 ( .A(n38187), .Z(n38189) );
  XOR U40876 ( .A(n38190), .B(mreg[196]), .Z(n38187) );
  NAND U40877 ( .A(n38191), .B(mul_pow), .Z(n38190) );
  XOR U40878 ( .A(mreg[196]), .B(creg[196]), .Z(n38191) );
  XOR U40879 ( .A(n38192), .B(n38193), .Z(n38183) );
  ANDN U40880 ( .A(n38194), .B(n29573), .Z(n38193) );
  XOR U40881 ( .A(n38195), .B(\modmult_1/zin[0][194] ), .Z(n29573) );
  IV U40882 ( .A(n38192), .Z(n38195) );
  XNOR U40883 ( .A(n38192), .B(n29572), .Z(n38194) );
  XOR U40884 ( .A(n38196), .B(n38197), .Z(n29572) );
  AND U40885 ( .A(\modmult_1/xin[1023] ), .B(n38198), .Z(n38197) );
  IV U40886 ( .A(n38196), .Z(n38198) );
  XOR U40887 ( .A(n38199), .B(mreg[195]), .Z(n38196) );
  NAND U40888 ( .A(n38200), .B(mul_pow), .Z(n38199) );
  XOR U40889 ( .A(mreg[195]), .B(creg[195]), .Z(n38200) );
  XOR U40890 ( .A(n38201), .B(n38202), .Z(n38192) );
  ANDN U40891 ( .A(n38203), .B(n29579), .Z(n38202) );
  XOR U40892 ( .A(n38204), .B(\modmult_1/zin[0][193] ), .Z(n29579) );
  IV U40893 ( .A(n38201), .Z(n38204) );
  XNOR U40894 ( .A(n38201), .B(n29578), .Z(n38203) );
  XOR U40895 ( .A(n38205), .B(n38206), .Z(n29578) );
  AND U40896 ( .A(\modmult_1/xin[1023] ), .B(n38207), .Z(n38206) );
  IV U40897 ( .A(n38205), .Z(n38207) );
  XOR U40898 ( .A(n38208), .B(mreg[194]), .Z(n38205) );
  NAND U40899 ( .A(n38209), .B(mul_pow), .Z(n38208) );
  XOR U40900 ( .A(mreg[194]), .B(creg[194]), .Z(n38209) );
  XOR U40901 ( .A(n38210), .B(n38211), .Z(n38201) );
  ANDN U40902 ( .A(n38212), .B(n29585), .Z(n38211) );
  XOR U40903 ( .A(n38213), .B(\modmult_1/zin[0][192] ), .Z(n29585) );
  IV U40904 ( .A(n38210), .Z(n38213) );
  XNOR U40905 ( .A(n38210), .B(n29584), .Z(n38212) );
  XOR U40906 ( .A(n38214), .B(n38215), .Z(n29584) );
  AND U40907 ( .A(\modmult_1/xin[1023] ), .B(n38216), .Z(n38215) );
  IV U40908 ( .A(n38214), .Z(n38216) );
  XOR U40909 ( .A(n38217), .B(mreg[193]), .Z(n38214) );
  NAND U40910 ( .A(n38218), .B(mul_pow), .Z(n38217) );
  XOR U40911 ( .A(mreg[193]), .B(creg[193]), .Z(n38218) );
  XOR U40912 ( .A(n38219), .B(n38220), .Z(n38210) );
  ANDN U40913 ( .A(n38221), .B(n29591), .Z(n38220) );
  XOR U40914 ( .A(n38222), .B(\modmult_1/zin[0][191] ), .Z(n29591) );
  IV U40915 ( .A(n38219), .Z(n38222) );
  XNOR U40916 ( .A(n38219), .B(n29590), .Z(n38221) );
  XOR U40917 ( .A(n38223), .B(n38224), .Z(n29590) );
  AND U40918 ( .A(\modmult_1/xin[1023] ), .B(n38225), .Z(n38224) );
  IV U40919 ( .A(n38223), .Z(n38225) );
  XOR U40920 ( .A(n38226), .B(mreg[192]), .Z(n38223) );
  NAND U40921 ( .A(n38227), .B(mul_pow), .Z(n38226) );
  XOR U40922 ( .A(mreg[192]), .B(creg[192]), .Z(n38227) );
  XOR U40923 ( .A(n38228), .B(n38229), .Z(n38219) );
  ANDN U40924 ( .A(n38230), .B(n29597), .Z(n38229) );
  XOR U40925 ( .A(n38231), .B(\modmult_1/zin[0][190] ), .Z(n29597) );
  IV U40926 ( .A(n38228), .Z(n38231) );
  XNOR U40927 ( .A(n38228), .B(n29596), .Z(n38230) );
  XOR U40928 ( .A(n38232), .B(n38233), .Z(n29596) );
  AND U40929 ( .A(\modmult_1/xin[1023] ), .B(n38234), .Z(n38233) );
  IV U40930 ( .A(n38232), .Z(n38234) );
  XOR U40931 ( .A(n38235), .B(mreg[191]), .Z(n38232) );
  NAND U40932 ( .A(n38236), .B(mul_pow), .Z(n38235) );
  XOR U40933 ( .A(mreg[191]), .B(creg[191]), .Z(n38236) );
  XOR U40934 ( .A(n38237), .B(n38238), .Z(n38228) );
  ANDN U40935 ( .A(n38239), .B(n29603), .Z(n38238) );
  XOR U40936 ( .A(n38240), .B(\modmult_1/zin[0][189] ), .Z(n29603) );
  IV U40937 ( .A(n38237), .Z(n38240) );
  XNOR U40938 ( .A(n38237), .B(n29602), .Z(n38239) );
  XOR U40939 ( .A(n38241), .B(n38242), .Z(n29602) );
  AND U40940 ( .A(\modmult_1/xin[1023] ), .B(n38243), .Z(n38242) );
  IV U40941 ( .A(n38241), .Z(n38243) );
  XOR U40942 ( .A(n38244), .B(mreg[190]), .Z(n38241) );
  NAND U40943 ( .A(n38245), .B(mul_pow), .Z(n38244) );
  XOR U40944 ( .A(mreg[190]), .B(creg[190]), .Z(n38245) );
  XOR U40945 ( .A(n38246), .B(n38247), .Z(n38237) );
  ANDN U40946 ( .A(n38248), .B(n29609), .Z(n38247) );
  XOR U40947 ( .A(n38249), .B(\modmult_1/zin[0][188] ), .Z(n29609) );
  IV U40948 ( .A(n38246), .Z(n38249) );
  XNOR U40949 ( .A(n38246), .B(n29608), .Z(n38248) );
  XOR U40950 ( .A(n38250), .B(n38251), .Z(n29608) );
  AND U40951 ( .A(\modmult_1/xin[1023] ), .B(n38252), .Z(n38251) );
  IV U40952 ( .A(n38250), .Z(n38252) );
  XOR U40953 ( .A(n38253), .B(mreg[189]), .Z(n38250) );
  NAND U40954 ( .A(n38254), .B(mul_pow), .Z(n38253) );
  XOR U40955 ( .A(mreg[189]), .B(creg[189]), .Z(n38254) );
  XOR U40956 ( .A(n38255), .B(n38256), .Z(n38246) );
  ANDN U40957 ( .A(n38257), .B(n29615), .Z(n38256) );
  XOR U40958 ( .A(n38258), .B(\modmult_1/zin[0][187] ), .Z(n29615) );
  IV U40959 ( .A(n38255), .Z(n38258) );
  XNOR U40960 ( .A(n38255), .B(n29614), .Z(n38257) );
  XOR U40961 ( .A(n38259), .B(n38260), .Z(n29614) );
  AND U40962 ( .A(\modmult_1/xin[1023] ), .B(n38261), .Z(n38260) );
  IV U40963 ( .A(n38259), .Z(n38261) );
  XOR U40964 ( .A(n38262), .B(mreg[188]), .Z(n38259) );
  NAND U40965 ( .A(n38263), .B(mul_pow), .Z(n38262) );
  XOR U40966 ( .A(mreg[188]), .B(creg[188]), .Z(n38263) );
  XOR U40967 ( .A(n38264), .B(n38265), .Z(n38255) );
  ANDN U40968 ( .A(n38266), .B(n29621), .Z(n38265) );
  XOR U40969 ( .A(n38267), .B(\modmult_1/zin[0][186] ), .Z(n29621) );
  IV U40970 ( .A(n38264), .Z(n38267) );
  XNOR U40971 ( .A(n38264), .B(n29620), .Z(n38266) );
  XOR U40972 ( .A(n38268), .B(n38269), .Z(n29620) );
  AND U40973 ( .A(\modmult_1/xin[1023] ), .B(n38270), .Z(n38269) );
  IV U40974 ( .A(n38268), .Z(n38270) );
  XOR U40975 ( .A(n38271), .B(mreg[187]), .Z(n38268) );
  NAND U40976 ( .A(n38272), .B(mul_pow), .Z(n38271) );
  XOR U40977 ( .A(mreg[187]), .B(creg[187]), .Z(n38272) );
  XOR U40978 ( .A(n38273), .B(n38274), .Z(n38264) );
  ANDN U40979 ( .A(n38275), .B(n29627), .Z(n38274) );
  XOR U40980 ( .A(n38276), .B(\modmult_1/zin[0][185] ), .Z(n29627) );
  IV U40981 ( .A(n38273), .Z(n38276) );
  XNOR U40982 ( .A(n38273), .B(n29626), .Z(n38275) );
  XOR U40983 ( .A(n38277), .B(n38278), .Z(n29626) );
  AND U40984 ( .A(\modmult_1/xin[1023] ), .B(n38279), .Z(n38278) );
  IV U40985 ( .A(n38277), .Z(n38279) );
  XOR U40986 ( .A(n38280), .B(mreg[186]), .Z(n38277) );
  NAND U40987 ( .A(n38281), .B(mul_pow), .Z(n38280) );
  XOR U40988 ( .A(mreg[186]), .B(creg[186]), .Z(n38281) );
  XOR U40989 ( .A(n38282), .B(n38283), .Z(n38273) );
  ANDN U40990 ( .A(n38284), .B(n29633), .Z(n38283) );
  XOR U40991 ( .A(n38285), .B(\modmult_1/zin[0][184] ), .Z(n29633) );
  IV U40992 ( .A(n38282), .Z(n38285) );
  XNOR U40993 ( .A(n38282), .B(n29632), .Z(n38284) );
  XOR U40994 ( .A(n38286), .B(n38287), .Z(n29632) );
  AND U40995 ( .A(\modmult_1/xin[1023] ), .B(n38288), .Z(n38287) );
  IV U40996 ( .A(n38286), .Z(n38288) );
  XOR U40997 ( .A(n38289), .B(mreg[185]), .Z(n38286) );
  NAND U40998 ( .A(n38290), .B(mul_pow), .Z(n38289) );
  XOR U40999 ( .A(mreg[185]), .B(creg[185]), .Z(n38290) );
  XOR U41000 ( .A(n38291), .B(n38292), .Z(n38282) );
  ANDN U41001 ( .A(n38293), .B(n29639), .Z(n38292) );
  XOR U41002 ( .A(n38294), .B(\modmult_1/zin[0][183] ), .Z(n29639) );
  IV U41003 ( .A(n38291), .Z(n38294) );
  XNOR U41004 ( .A(n38291), .B(n29638), .Z(n38293) );
  XOR U41005 ( .A(n38295), .B(n38296), .Z(n29638) );
  AND U41006 ( .A(\modmult_1/xin[1023] ), .B(n38297), .Z(n38296) );
  IV U41007 ( .A(n38295), .Z(n38297) );
  XOR U41008 ( .A(n38298), .B(mreg[184]), .Z(n38295) );
  NAND U41009 ( .A(n38299), .B(mul_pow), .Z(n38298) );
  XOR U41010 ( .A(mreg[184]), .B(creg[184]), .Z(n38299) );
  XOR U41011 ( .A(n38300), .B(n38301), .Z(n38291) );
  ANDN U41012 ( .A(n38302), .B(n29645), .Z(n38301) );
  XOR U41013 ( .A(n38303), .B(\modmult_1/zin[0][182] ), .Z(n29645) );
  IV U41014 ( .A(n38300), .Z(n38303) );
  XNOR U41015 ( .A(n38300), .B(n29644), .Z(n38302) );
  XOR U41016 ( .A(n38304), .B(n38305), .Z(n29644) );
  AND U41017 ( .A(\modmult_1/xin[1023] ), .B(n38306), .Z(n38305) );
  IV U41018 ( .A(n38304), .Z(n38306) );
  XOR U41019 ( .A(n38307), .B(mreg[183]), .Z(n38304) );
  NAND U41020 ( .A(n38308), .B(mul_pow), .Z(n38307) );
  XOR U41021 ( .A(mreg[183]), .B(creg[183]), .Z(n38308) );
  XOR U41022 ( .A(n38309), .B(n38310), .Z(n38300) );
  ANDN U41023 ( .A(n38311), .B(n29651), .Z(n38310) );
  XOR U41024 ( .A(n38312), .B(\modmult_1/zin[0][181] ), .Z(n29651) );
  IV U41025 ( .A(n38309), .Z(n38312) );
  XNOR U41026 ( .A(n38309), .B(n29650), .Z(n38311) );
  XOR U41027 ( .A(n38313), .B(n38314), .Z(n29650) );
  AND U41028 ( .A(\modmult_1/xin[1023] ), .B(n38315), .Z(n38314) );
  IV U41029 ( .A(n38313), .Z(n38315) );
  XOR U41030 ( .A(n38316), .B(mreg[182]), .Z(n38313) );
  NAND U41031 ( .A(n38317), .B(mul_pow), .Z(n38316) );
  XOR U41032 ( .A(mreg[182]), .B(creg[182]), .Z(n38317) );
  XOR U41033 ( .A(n38318), .B(n38319), .Z(n38309) );
  ANDN U41034 ( .A(n38320), .B(n29657), .Z(n38319) );
  XOR U41035 ( .A(n38321), .B(\modmult_1/zin[0][180] ), .Z(n29657) );
  IV U41036 ( .A(n38318), .Z(n38321) );
  XNOR U41037 ( .A(n38318), .B(n29656), .Z(n38320) );
  XOR U41038 ( .A(n38322), .B(n38323), .Z(n29656) );
  AND U41039 ( .A(\modmult_1/xin[1023] ), .B(n38324), .Z(n38323) );
  IV U41040 ( .A(n38322), .Z(n38324) );
  XOR U41041 ( .A(n38325), .B(mreg[181]), .Z(n38322) );
  NAND U41042 ( .A(n38326), .B(mul_pow), .Z(n38325) );
  XOR U41043 ( .A(mreg[181]), .B(creg[181]), .Z(n38326) );
  XOR U41044 ( .A(n38327), .B(n38328), .Z(n38318) );
  ANDN U41045 ( .A(n38329), .B(n29663), .Z(n38328) );
  XOR U41046 ( .A(n38330), .B(\modmult_1/zin[0][179] ), .Z(n29663) );
  IV U41047 ( .A(n38327), .Z(n38330) );
  XNOR U41048 ( .A(n38327), .B(n29662), .Z(n38329) );
  XOR U41049 ( .A(n38331), .B(n38332), .Z(n29662) );
  AND U41050 ( .A(\modmult_1/xin[1023] ), .B(n38333), .Z(n38332) );
  IV U41051 ( .A(n38331), .Z(n38333) );
  XOR U41052 ( .A(n38334), .B(mreg[180]), .Z(n38331) );
  NAND U41053 ( .A(n38335), .B(mul_pow), .Z(n38334) );
  XOR U41054 ( .A(mreg[180]), .B(creg[180]), .Z(n38335) );
  XOR U41055 ( .A(n38336), .B(n38337), .Z(n38327) );
  ANDN U41056 ( .A(n38338), .B(n29669), .Z(n38337) );
  XOR U41057 ( .A(n38339), .B(\modmult_1/zin[0][178] ), .Z(n29669) );
  IV U41058 ( .A(n38336), .Z(n38339) );
  XNOR U41059 ( .A(n38336), .B(n29668), .Z(n38338) );
  XOR U41060 ( .A(n38340), .B(n38341), .Z(n29668) );
  AND U41061 ( .A(\modmult_1/xin[1023] ), .B(n38342), .Z(n38341) );
  IV U41062 ( .A(n38340), .Z(n38342) );
  XOR U41063 ( .A(n38343), .B(mreg[179]), .Z(n38340) );
  NAND U41064 ( .A(n38344), .B(mul_pow), .Z(n38343) );
  XOR U41065 ( .A(mreg[179]), .B(creg[179]), .Z(n38344) );
  XOR U41066 ( .A(n38345), .B(n38346), .Z(n38336) );
  ANDN U41067 ( .A(n38347), .B(n29675), .Z(n38346) );
  XOR U41068 ( .A(n38348), .B(\modmult_1/zin[0][177] ), .Z(n29675) );
  IV U41069 ( .A(n38345), .Z(n38348) );
  XNOR U41070 ( .A(n38345), .B(n29674), .Z(n38347) );
  XOR U41071 ( .A(n38349), .B(n38350), .Z(n29674) );
  AND U41072 ( .A(\modmult_1/xin[1023] ), .B(n38351), .Z(n38350) );
  IV U41073 ( .A(n38349), .Z(n38351) );
  XOR U41074 ( .A(n38352), .B(mreg[178]), .Z(n38349) );
  NAND U41075 ( .A(n38353), .B(mul_pow), .Z(n38352) );
  XOR U41076 ( .A(mreg[178]), .B(creg[178]), .Z(n38353) );
  XOR U41077 ( .A(n38354), .B(n38355), .Z(n38345) );
  ANDN U41078 ( .A(n38356), .B(n29681), .Z(n38355) );
  XOR U41079 ( .A(n38357), .B(\modmult_1/zin[0][176] ), .Z(n29681) );
  IV U41080 ( .A(n38354), .Z(n38357) );
  XNOR U41081 ( .A(n38354), .B(n29680), .Z(n38356) );
  XOR U41082 ( .A(n38358), .B(n38359), .Z(n29680) );
  AND U41083 ( .A(\modmult_1/xin[1023] ), .B(n38360), .Z(n38359) );
  IV U41084 ( .A(n38358), .Z(n38360) );
  XOR U41085 ( .A(n38361), .B(mreg[177]), .Z(n38358) );
  NAND U41086 ( .A(n38362), .B(mul_pow), .Z(n38361) );
  XOR U41087 ( .A(mreg[177]), .B(creg[177]), .Z(n38362) );
  XOR U41088 ( .A(n38363), .B(n38364), .Z(n38354) );
  ANDN U41089 ( .A(n38365), .B(n29687), .Z(n38364) );
  XOR U41090 ( .A(n38366), .B(\modmult_1/zin[0][175] ), .Z(n29687) );
  IV U41091 ( .A(n38363), .Z(n38366) );
  XNOR U41092 ( .A(n38363), .B(n29686), .Z(n38365) );
  XOR U41093 ( .A(n38367), .B(n38368), .Z(n29686) );
  AND U41094 ( .A(\modmult_1/xin[1023] ), .B(n38369), .Z(n38368) );
  IV U41095 ( .A(n38367), .Z(n38369) );
  XOR U41096 ( .A(n38370), .B(mreg[176]), .Z(n38367) );
  NAND U41097 ( .A(n38371), .B(mul_pow), .Z(n38370) );
  XOR U41098 ( .A(mreg[176]), .B(creg[176]), .Z(n38371) );
  XOR U41099 ( .A(n38372), .B(n38373), .Z(n38363) );
  ANDN U41100 ( .A(n38374), .B(n29693), .Z(n38373) );
  XOR U41101 ( .A(n38375), .B(\modmult_1/zin[0][174] ), .Z(n29693) );
  IV U41102 ( .A(n38372), .Z(n38375) );
  XNOR U41103 ( .A(n38372), .B(n29692), .Z(n38374) );
  XOR U41104 ( .A(n38376), .B(n38377), .Z(n29692) );
  AND U41105 ( .A(\modmult_1/xin[1023] ), .B(n38378), .Z(n38377) );
  IV U41106 ( .A(n38376), .Z(n38378) );
  XOR U41107 ( .A(n38379), .B(mreg[175]), .Z(n38376) );
  NAND U41108 ( .A(n38380), .B(mul_pow), .Z(n38379) );
  XOR U41109 ( .A(mreg[175]), .B(creg[175]), .Z(n38380) );
  XOR U41110 ( .A(n38381), .B(n38382), .Z(n38372) );
  ANDN U41111 ( .A(n38383), .B(n29699), .Z(n38382) );
  XOR U41112 ( .A(n38384), .B(\modmult_1/zin[0][173] ), .Z(n29699) );
  IV U41113 ( .A(n38381), .Z(n38384) );
  XNOR U41114 ( .A(n38381), .B(n29698), .Z(n38383) );
  XOR U41115 ( .A(n38385), .B(n38386), .Z(n29698) );
  AND U41116 ( .A(\modmult_1/xin[1023] ), .B(n38387), .Z(n38386) );
  IV U41117 ( .A(n38385), .Z(n38387) );
  XOR U41118 ( .A(n38388), .B(mreg[174]), .Z(n38385) );
  NAND U41119 ( .A(n38389), .B(mul_pow), .Z(n38388) );
  XOR U41120 ( .A(mreg[174]), .B(creg[174]), .Z(n38389) );
  XOR U41121 ( .A(n38390), .B(n38391), .Z(n38381) );
  ANDN U41122 ( .A(n38392), .B(n29705), .Z(n38391) );
  XOR U41123 ( .A(n38393), .B(\modmult_1/zin[0][172] ), .Z(n29705) );
  IV U41124 ( .A(n38390), .Z(n38393) );
  XNOR U41125 ( .A(n38390), .B(n29704), .Z(n38392) );
  XOR U41126 ( .A(n38394), .B(n38395), .Z(n29704) );
  AND U41127 ( .A(\modmult_1/xin[1023] ), .B(n38396), .Z(n38395) );
  IV U41128 ( .A(n38394), .Z(n38396) );
  XOR U41129 ( .A(n38397), .B(mreg[173]), .Z(n38394) );
  NAND U41130 ( .A(n38398), .B(mul_pow), .Z(n38397) );
  XOR U41131 ( .A(mreg[173]), .B(creg[173]), .Z(n38398) );
  XOR U41132 ( .A(n38399), .B(n38400), .Z(n38390) );
  ANDN U41133 ( .A(n38401), .B(n29711), .Z(n38400) );
  XOR U41134 ( .A(n38402), .B(\modmult_1/zin[0][171] ), .Z(n29711) );
  IV U41135 ( .A(n38399), .Z(n38402) );
  XNOR U41136 ( .A(n38399), .B(n29710), .Z(n38401) );
  XOR U41137 ( .A(n38403), .B(n38404), .Z(n29710) );
  AND U41138 ( .A(\modmult_1/xin[1023] ), .B(n38405), .Z(n38404) );
  IV U41139 ( .A(n38403), .Z(n38405) );
  XOR U41140 ( .A(n38406), .B(mreg[172]), .Z(n38403) );
  NAND U41141 ( .A(n38407), .B(mul_pow), .Z(n38406) );
  XOR U41142 ( .A(mreg[172]), .B(creg[172]), .Z(n38407) );
  XOR U41143 ( .A(n38408), .B(n38409), .Z(n38399) );
  ANDN U41144 ( .A(n38410), .B(n29717), .Z(n38409) );
  XOR U41145 ( .A(n38411), .B(\modmult_1/zin[0][170] ), .Z(n29717) );
  IV U41146 ( .A(n38408), .Z(n38411) );
  XNOR U41147 ( .A(n38408), .B(n29716), .Z(n38410) );
  XOR U41148 ( .A(n38412), .B(n38413), .Z(n29716) );
  AND U41149 ( .A(\modmult_1/xin[1023] ), .B(n38414), .Z(n38413) );
  IV U41150 ( .A(n38412), .Z(n38414) );
  XOR U41151 ( .A(n38415), .B(mreg[171]), .Z(n38412) );
  NAND U41152 ( .A(n38416), .B(mul_pow), .Z(n38415) );
  XOR U41153 ( .A(mreg[171]), .B(creg[171]), .Z(n38416) );
  XOR U41154 ( .A(n38417), .B(n38418), .Z(n38408) );
  ANDN U41155 ( .A(n38419), .B(n29723), .Z(n38418) );
  XOR U41156 ( .A(n38420), .B(\modmult_1/zin[0][169] ), .Z(n29723) );
  IV U41157 ( .A(n38417), .Z(n38420) );
  XNOR U41158 ( .A(n38417), .B(n29722), .Z(n38419) );
  XOR U41159 ( .A(n38421), .B(n38422), .Z(n29722) );
  AND U41160 ( .A(\modmult_1/xin[1023] ), .B(n38423), .Z(n38422) );
  IV U41161 ( .A(n38421), .Z(n38423) );
  XOR U41162 ( .A(n38424), .B(mreg[170]), .Z(n38421) );
  NAND U41163 ( .A(n38425), .B(mul_pow), .Z(n38424) );
  XOR U41164 ( .A(mreg[170]), .B(creg[170]), .Z(n38425) );
  XOR U41165 ( .A(n38426), .B(n38427), .Z(n38417) );
  ANDN U41166 ( .A(n38428), .B(n29729), .Z(n38427) );
  XOR U41167 ( .A(n38429), .B(\modmult_1/zin[0][168] ), .Z(n29729) );
  IV U41168 ( .A(n38426), .Z(n38429) );
  XNOR U41169 ( .A(n38426), .B(n29728), .Z(n38428) );
  XOR U41170 ( .A(n38430), .B(n38431), .Z(n29728) );
  AND U41171 ( .A(\modmult_1/xin[1023] ), .B(n38432), .Z(n38431) );
  IV U41172 ( .A(n38430), .Z(n38432) );
  XOR U41173 ( .A(n38433), .B(mreg[169]), .Z(n38430) );
  NAND U41174 ( .A(n38434), .B(mul_pow), .Z(n38433) );
  XOR U41175 ( .A(mreg[169]), .B(creg[169]), .Z(n38434) );
  XOR U41176 ( .A(n38435), .B(n38436), .Z(n38426) );
  ANDN U41177 ( .A(n38437), .B(n29735), .Z(n38436) );
  XOR U41178 ( .A(n38438), .B(\modmult_1/zin[0][167] ), .Z(n29735) );
  IV U41179 ( .A(n38435), .Z(n38438) );
  XNOR U41180 ( .A(n38435), .B(n29734), .Z(n38437) );
  XOR U41181 ( .A(n38439), .B(n38440), .Z(n29734) );
  AND U41182 ( .A(\modmult_1/xin[1023] ), .B(n38441), .Z(n38440) );
  IV U41183 ( .A(n38439), .Z(n38441) );
  XOR U41184 ( .A(n38442), .B(mreg[168]), .Z(n38439) );
  NAND U41185 ( .A(n38443), .B(mul_pow), .Z(n38442) );
  XOR U41186 ( .A(mreg[168]), .B(creg[168]), .Z(n38443) );
  XOR U41187 ( .A(n38444), .B(n38445), .Z(n38435) );
  ANDN U41188 ( .A(n38446), .B(n29741), .Z(n38445) );
  XOR U41189 ( .A(n38447), .B(\modmult_1/zin[0][166] ), .Z(n29741) );
  IV U41190 ( .A(n38444), .Z(n38447) );
  XNOR U41191 ( .A(n38444), .B(n29740), .Z(n38446) );
  XOR U41192 ( .A(n38448), .B(n38449), .Z(n29740) );
  AND U41193 ( .A(\modmult_1/xin[1023] ), .B(n38450), .Z(n38449) );
  IV U41194 ( .A(n38448), .Z(n38450) );
  XOR U41195 ( .A(n38451), .B(mreg[167]), .Z(n38448) );
  NAND U41196 ( .A(n38452), .B(mul_pow), .Z(n38451) );
  XOR U41197 ( .A(mreg[167]), .B(creg[167]), .Z(n38452) );
  XOR U41198 ( .A(n38453), .B(n38454), .Z(n38444) );
  ANDN U41199 ( .A(n38455), .B(n29747), .Z(n38454) );
  XOR U41200 ( .A(n38456), .B(\modmult_1/zin[0][165] ), .Z(n29747) );
  IV U41201 ( .A(n38453), .Z(n38456) );
  XNOR U41202 ( .A(n38453), .B(n29746), .Z(n38455) );
  XOR U41203 ( .A(n38457), .B(n38458), .Z(n29746) );
  AND U41204 ( .A(\modmult_1/xin[1023] ), .B(n38459), .Z(n38458) );
  IV U41205 ( .A(n38457), .Z(n38459) );
  XOR U41206 ( .A(n38460), .B(mreg[166]), .Z(n38457) );
  NAND U41207 ( .A(n38461), .B(mul_pow), .Z(n38460) );
  XOR U41208 ( .A(mreg[166]), .B(creg[166]), .Z(n38461) );
  XOR U41209 ( .A(n38462), .B(n38463), .Z(n38453) );
  ANDN U41210 ( .A(n38464), .B(n29753), .Z(n38463) );
  XOR U41211 ( .A(n38465), .B(\modmult_1/zin[0][164] ), .Z(n29753) );
  IV U41212 ( .A(n38462), .Z(n38465) );
  XNOR U41213 ( .A(n38462), .B(n29752), .Z(n38464) );
  XOR U41214 ( .A(n38466), .B(n38467), .Z(n29752) );
  AND U41215 ( .A(\modmult_1/xin[1023] ), .B(n38468), .Z(n38467) );
  IV U41216 ( .A(n38466), .Z(n38468) );
  XOR U41217 ( .A(n38469), .B(mreg[165]), .Z(n38466) );
  NAND U41218 ( .A(n38470), .B(mul_pow), .Z(n38469) );
  XOR U41219 ( .A(mreg[165]), .B(creg[165]), .Z(n38470) );
  XOR U41220 ( .A(n38471), .B(n38472), .Z(n38462) );
  ANDN U41221 ( .A(n38473), .B(n29759), .Z(n38472) );
  XOR U41222 ( .A(n38474), .B(\modmult_1/zin[0][163] ), .Z(n29759) );
  IV U41223 ( .A(n38471), .Z(n38474) );
  XNOR U41224 ( .A(n38471), .B(n29758), .Z(n38473) );
  XOR U41225 ( .A(n38475), .B(n38476), .Z(n29758) );
  AND U41226 ( .A(\modmult_1/xin[1023] ), .B(n38477), .Z(n38476) );
  IV U41227 ( .A(n38475), .Z(n38477) );
  XOR U41228 ( .A(n38478), .B(mreg[164]), .Z(n38475) );
  NAND U41229 ( .A(n38479), .B(mul_pow), .Z(n38478) );
  XOR U41230 ( .A(mreg[164]), .B(creg[164]), .Z(n38479) );
  XOR U41231 ( .A(n38480), .B(n38481), .Z(n38471) );
  ANDN U41232 ( .A(n38482), .B(n29765), .Z(n38481) );
  XOR U41233 ( .A(n38483), .B(\modmult_1/zin[0][162] ), .Z(n29765) );
  IV U41234 ( .A(n38480), .Z(n38483) );
  XNOR U41235 ( .A(n38480), .B(n29764), .Z(n38482) );
  XOR U41236 ( .A(n38484), .B(n38485), .Z(n29764) );
  AND U41237 ( .A(\modmult_1/xin[1023] ), .B(n38486), .Z(n38485) );
  IV U41238 ( .A(n38484), .Z(n38486) );
  XOR U41239 ( .A(n38487), .B(mreg[163]), .Z(n38484) );
  NAND U41240 ( .A(n38488), .B(mul_pow), .Z(n38487) );
  XOR U41241 ( .A(mreg[163]), .B(creg[163]), .Z(n38488) );
  XOR U41242 ( .A(n38489), .B(n38490), .Z(n38480) );
  ANDN U41243 ( .A(n38491), .B(n29771), .Z(n38490) );
  XOR U41244 ( .A(n38492), .B(\modmult_1/zin[0][161] ), .Z(n29771) );
  IV U41245 ( .A(n38489), .Z(n38492) );
  XNOR U41246 ( .A(n38489), .B(n29770), .Z(n38491) );
  XOR U41247 ( .A(n38493), .B(n38494), .Z(n29770) );
  AND U41248 ( .A(\modmult_1/xin[1023] ), .B(n38495), .Z(n38494) );
  IV U41249 ( .A(n38493), .Z(n38495) );
  XOR U41250 ( .A(n38496), .B(mreg[162]), .Z(n38493) );
  NAND U41251 ( .A(n38497), .B(mul_pow), .Z(n38496) );
  XOR U41252 ( .A(mreg[162]), .B(creg[162]), .Z(n38497) );
  XOR U41253 ( .A(n38498), .B(n38499), .Z(n38489) );
  ANDN U41254 ( .A(n38500), .B(n29777), .Z(n38499) );
  XOR U41255 ( .A(n38501), .B(\modmult_1/zin[0][160] ), .Z(n29777) );
  IV U41256 ( .A(n38498), .Z(n38501) );
  XNOR U41257 ( .A(n38498), .B(n29776), .Z(n38500) );
  XOR U41258 ( .A(n38502), .B(n38503), .Z(n29776) );
  AND U41259 ( .A(\modmult_1/xin[1023] ), .B(n38504), .Z(n38503) );
  IV U41260 ( .A(n38502), .Z(n38504) );
  XOR U41261 ( .A(n38505), .B(mreg[161]), .Z(n38502) );
  NAND U41262 ( .A(n38506), .B(mul_pow), .Z(n38505) );
  XOR U41263 ( .A(mreg[161]), .B(creg[161]), .Z(n38506) );
  XOR U41264 ( .A(n38507), .B(n38508), .Z(n38498) );
  ANDN U41265 ( .A(n38509), .B(n29783), .Z(n38508) );
  XOR U41266 ( .A(n38510), .B(\modmult_1/zin[0][159] ), .Z(n29783) );
  IV U41267 ( .A(n38507), .Z(n38510) );
  XNOR U41268 ( .A(n38507), .B(n29782), .Z(n38509) );
  XOR U41269 ( .A(n38511), .B(n38512), .Z(n29782) );
  AND U41270 ( .A(\modmult_1/xin[1023] ), .B(n38513), .Z(n38512) );
  IV U41271 ( .A(n38511), .Z(n38513) );
  XOR U41272 ( .A(n38514), .B(mreg[160]), .Z(n38511) );
  NAND U41273 ( .A(n38515), .B(mul_pow), .Z(n38514) );
  XOR U41274 ( .A(mreg[160]), .B(creg[160]), .Z(n38515) );
  XOR U41275 ( .A(n38516), .B(n38517), .Z(n38507) );
  ANDN U41276 ( .A(n38518), .B(n29789), .Z(n38517) );
  XOR U41277 ( .A(n38519), .B(\modmult_1/zin[0][158] ), .Z(n29789) );
  IV U41278 ( .A(n38516), .Z(n38519) );
  XNOR U41279 ( .A(n38516), .B(n29788), .Z(n38518) );
  XOR U41280 ( .A(n38520), .B(n38521), .Z(n29788) );
  AND U41281 ( .A(\modmult_1/xin[1023] ), .B(n38522), .Z(n38521) );
  IV U41282 ( .A(n38520), .Z(n38522) );
  XOR U41283 ( .A(n38523), .B(mreg[159]), .Z(n38520) );
  NAND U41284 ( .A(n38524), .B(mul_pow), .Z(n38523) );
  XOR U41285 ( .A(mreg[159]), .B(creg[159]), .Z(n38524) );
  XOR U41286 ( .A(n38525), .B(n38526), .Z(n38516) );
  ANDN U41287 ( .A(n38527), .B(n29795), .Z(n38526) );
  XOR U41288 ( .A(n38528), .B(\modmult_1/zin[0][157] ), .Z(n29795) );
  IV U41289 ( .A(n38525), .Z(n38528) );
  XNOR U41290 ( .A(n38525), .B(n29794), .Z(n38527) );
  XOR U41291 ( .A(n38529), .B(n38530), .Z(n29794) );
  AND U41292 ( .A(\modmult_1/xin[1023] ), .B(n38531), .Z(n38530) );
  IV U41293 ( .A(n38529), .Z(n38531) );
  XOR U41294 ( .A(n38532), .B(mreg[158]), .Z(n38529) );
  NAND U41295 ( .A(n38533), .B(mul_pow), .Z(n38532) );
  XOR U41296 ( .A(mreg[158]), .B(creg[158]), .Z(n38533) );
  XOR U41297 ( .A(n38534), .B(n38535), .Z(n38525) );
  ANDN U41298 ( .A(n38536), .B(n29801), .Z(n38535) );
  XOR U41299 ( .A(n38537), .B(\modmult_1/zin[0][156] ), .Z(n29801) );
  IV U41300 ( .A(n38534), .Z(n38537) );
  XNOR U41301 ( .A(n38534), .B(n29800), .Z(n38536) );
  XOR U41302 ( .A(n38538), .B(n38539), .Z(n29800) );
  AND U41303 ( .A(\modmult_1/xin[1023] ), .B(n38540), .Z(n38539) );
  IV U41304 ( .A(n38538), .Z(n38540) );
  XOR U41305 ( .A(n38541), .B(mreg[157]), .Z(n38538) );
  NAND U41306 ( .A(n38542), .B(mul_pow), .Z(n38541) );
  XOR U41307 ( .A(mreg[157]), .B(creg[157]), .Z(n38542) );
  XOR U41308 ( .A(n38543), .B(n38544), .Z(n38534) );
  ANDN U41309 ( .A(n38545), .B(n29807), .Z(n38544) );
  XOR U41310 ( .A(n38546), .B(\modmult_1/zin[0][155] ), .Z(n29807) );
  IV U41311 ( .A(n38543), .Z(n38546) );
  XNOR U41312 ( .A(n38543), .B(n29806), .Z(n38545) );
  XOR U41313 ( .A(n38547), .B(n38548), .Z(n29806) );
  AND U41314 ( .A(\modmult_1/xin[1023] ), .B(n38549), .Z(n38548) );
  IV U41315 ( .A(n38547), .Z(n38549) );
  XOR U41316 ( .A(n38550), .B(mreg[156]), .Z(n38547) );
  NAND U41317 ( .A(n38551), .B(mul_pow), .Z(n38550) );
  XOR U41318 ( .A(mreg[156]), .B(creg[156]), .Z(n38551) );
  XOR U41319 ( .A(n38552), .B(n38553), .Z(n38543) );
  ANDN U41320 ( .A(n38554), .B(n29813), .Z(n38553) );
  XOR U41321 ( .A(n38555), .B(\modmult_1/zin[0][154] ), .Z(n29813) );
  IV U41322 ( .A(n38552), .Z(n38555) );
  XNOR U41323 ( .A(n38552), .B(n29812), .Z(n38554) );
  XOR U41324 ( .A(n38556), .B(n38557), .Z(n29812) );
  AND U41325 ( .A(\modmult_1/xin[1023] ), .B(n38558), .Z(n38557) );
  IV U41326 ( .A(n38556), .Z(n38558) );
  XOR U41327 ( .A(n38559), .B(mreg[155]), .Z(n38556) );
  NAND U41328 ( .A(n38560), .B(mul_pow), .Z(n38559) );
  XOR U41329 ( .A(mreg[155]), .B(creg[155]), .Z(n38560) );
  XOR U41330 ( .A(n38561), .B(n38562), .Z(n38552) );
  ANDN U41331 ( .A(n38563), .B(n29819), .Z(n38562) );
  XOR U41332 ( .A(n38564), .B(\modmult_1/zin[0][153] ), .Z(n29819) );
  IV U41333 ( .A(n38561), .Z(n38564) );
  XNOR U41334 ( .A(n38561), .B(n29818), .Z(n38563) );
  XOR U41335 ( .A(n38565), .B(n38566), .Z(n29818) );
  AND U41336 ( .A(\modmult_1/xin[1023] ), .B(n38567), .Z(n38566) );
  IV U41337 ( .A(n38565), .Z(n38567) );
  XOR U41338 ( .A(n38568), .B(mreg[154]), .Z(n38565) );
  NAND U41339 ( .A(n38569), .B(mul_pow), .Z(n38568) );
  XOR U41340 ( .A(mreg[154]), .B(creg[154]), .Z(n38569) );
  XOR U41341 ( .A(n38570), .B(n38571), .Z(n38561) );
  ANDN U41342 ( .A(n38572), .B(n29825), .Z(n38571) );
  XOR U41343 ( .A(n38573), .B(\modmult_1/zin[0][152] ), .Z(n29825) );
  IV U41344 ( .A(n38570), .Z(n38573) );
  XNOR U41345 ( .A(n38570), .B(n29824), .Z(n38572) );
  XOR U41346 ( .A(n38574), .B(n38575), .Z(n29824) );
  AND U41347 ( .A(\modmult_1/xin[1023] ), .B(n38576), .Z(n38575) );
  IV U41348 ( .A(n38574), .Z(n38576) );
  XOR U41349 ( .A(n38577), .B(mreg[153]), .Z(n38574) );
  NAND U41350 ( .A(n38578), .B(mul_pow), .Z(n38577) );
  XOR U41351 ( .A(mreg[153]), .B(creg[153]), .Z(n38578) );
  XOR U41352 ( .A(n38579), .B(n38580), .Z(n38570) );
  ANDN U41353 ( .A(n38581), .B(n29831), .Z(n38580) );
  XOR U41354 ( .A(n38582), .B(\modmult_1/zin[0][151] ), .Z(n29831) );
  IV U41355 ( .A(n38579), .Z(n38582) );
  XNOR U41356 ( .A(n38579), .B(n29830), .Z(n38581) );
  XOR U41357 ( .A(n38583), .B(n38584), .Z(n29830) );
  AND U41358 ( .A(\modmult_1/xin[1023] ), .B(n38585), .Z(n38584) );
  IV U41359 ( .A(n38583), .Z(n38585) );
  XOR U41360 ( .A(n38586), .B(mreg[152]), .Z(n38583) );
  NAND U41361 ( .A(n38587), .B(mul_pow), .Z(n38586) );
  XOR U41362 ( .A(mreg[152]), .B(creg[152]), .Z(n38587) );
  XOR U41363 ( .A(n38588), .B(n38589), .Z(n38579) );
  ANDN U41364 ( .A(n38590), .B(n29837), .Z(n38589) );
  XOR U41365 ( .A(n38591), .B(\modmult_1/zin[0][150] ), .Z(n29837) );
  IV U41366 ( .A(n38588), .Z(n38591) );
  XNOR U41367 ( .A(n38588), .B(n29836), .Z(n38590) );
  XOR U41368 ( .A(n38592), .B(n38593), .Z(n29836) );
  AND U41369 ( .A(\modmult_1/xin[1023] ), .B(n38594), .Z(n38593) );
  IV U41370 ( .A(n38592), .Z(n38594) );
  XOR U41371 ( .A(n38595), .B(mreg[151]), .Z(n38592) );
  NAND U41372 ( .A(n38596), .B(mul_pow), .Z(n38595) );
  XOR U41373 ( .A(mreg[151]), .B(creg[151]), .Z(n38596) );
  XOR U41374 ( .A(n38597), .B(n38598), .Z(n38588) );
  ANDN U41375 ( .A(n38599), .B(n29843), .Z(n38598) );
  XOR U41376 ( .A(n38600), .B(\modmult_1/zin[0][149] ), .Z(n29843) );
  IV U41377 ( .A(n38597), .Z(n38600) );
  XNOR U41378 ( .A(n38597), .B(n29842), .Z(n38599) );
  XOR U41379 ( .A(n38601), .B(n38602), .Z(n29842) );
  AND U41380 ( .A(\modmult_1/xin[1023] ), .B(n38603), .Z(n38602) );
  IV U41381 ( .A(n38601), .Z(n38603) );
  XOR U41382 ( .A(n38604), .B(mreg[150]), .Z(n38601) );
  NAND U41383 ( .A(n38605), .B(mul_pow), .Z(n38604) );
  XOR U41384 ( .A(mreg[150]), .B(creg[150]), .Z(n38605) );
  XOR U41385 ( .A(n38606), .B(n38607), .Z(n38597) );
  ANDN U41386 ( .A(n38608), .B(n29849), .Z(n38607) );
  XOR U41387 ( .A(n38609), .B(\modmult_1/zin[0][148] ), .Z(n29849) );
  IV U41388 ( .A(n38606), .Z(n38609) );
  XNOR U41389 ( .A(n38606), .B(n29848), .Z(n38608) );
  XOR U41390 ( .A(n38610), .B(n38611), .Z(n29848) );
  AND U41391 ( .A(\modmult_1/xin[1023] ), .B(n38612), .Z(n38611) );
  IV U41392 ( .A(n38610), .Z(n38612) );
  XOR U41393 ( .A(n38613), .B(mreg[149]), .Z(n38610) );
  NAND U41394 ( .A(n38614), .B(mul_pow), .Z(n38613) );
  XOR U41395 ( .A(mreg[149]), .B(creg[149]), .Z(n38614) );
  XOR U41396 ( .A(n38615), .B(n38616), .Z(n38606) );
  ANDN U41397 ( .A(n38617), .B(n29855), .Z(n38616) );
  XOR U41398 ( .A(n38618), .B(\modmult_1/zin[0][147] ), .Z(n29855) );
  IV U41399 ( .A(n38615), .Z(n38618) );
  XNOR U41400 ( .A(n38615), .B(n29854), .Z(n38617) );
  XOR U41401 ( .A(n38619), .B(n38620), .Z(n29854) );
  AND U41402 ( .A(\modmult_1/xin[1023] ), .B(n38621), .Z(n38620) );
  IV U41403 ( .A(n38619), .Z(n38621) );
  XOR U41404 ( .A(n38622), .B(mreg[148]), .Z(n38619) );
  NAND U41405 ( .A(n38623), .B(mul_pow), .Z(n38622) );
  XOR U41406 ( .A(mreg[148]), .B(creg[148]), .Z(n38623) );
  XOR U41407 ( .A(n38624), .B(n38625), .Z(n38615) );
  ANDN U41408 ( .A(n38626), .B(n29861), .Z(n38625) );
  XOR U41409 ( .A(n38627), .B(\modmult_1/zin[0][146] ), .Z(n29861) );
  IV U41410 ( .A(n38624), .Z(n38627) );
  XNOR U41411 ( .A(n38624), .B(n29860), .Z(n38626) );
  XOR U41412 ( .A(n38628), .B(n38629), .Z(n29860) );
  AND U41413 ( .A(\modmult_1/xin[1023] ), .B(n38630), .Z(n38629) );
  IV U41414 ( .A(n38628), .Z(n38630) );
  XOR U41415 ( .A(n38631), .B(mreg[147]), .Z(n38628) );
  NAND U41416 ( .A(n38632), .B(mul_pow), .Z(n38631) );
  XOR U41417 ( .A(mreg[147]), .B(creg[147]), .Z(n38632) );
  XOR U41418 ( .A(n38633), .B(n38634), .Z(n38624) );
  ANDN U41419 ( .A(n38635), .B(n29867), .Z(n38634) );
  XOR U41420 ( .A(n38636), .B(\modmult_1/zin[0][145] ), .Z(n29867) );
  IV U41421 ( .A(n38633), .Z(n38636) );
  XNOR U41422 ( .A(n38633), .B(n29866), .Z(n38635) );
  XOR U41423 ( .A(n38637), .B(n38638), .Z(n29866) );
  AND U41424 ( .A(\modmult_1/xin[1023] ), .B(n38639), .Z(n38638) );
  IV U41425 ( .A(n38637), .Z(n38639) );
  XOR U41426 ( .A(n38640), .B(mreg[146]), .Z(n38637) );
  NAND U41427 ( .A(n38641), .B(mul_pow), .Z(n38640) );
  XOR U41428 ( .A(mreg[146]), .B(creg[146]), .Z(n38641) );
  XOR U41429 ( .A(n38642), .B(n38643), .Z(n38633) );
  ANDN U41430 ( .A(n38644), .B(n29873), .Z(n38643) );
  XOR U41431 ( .A(n38645), .B(\modmult_1/zin[0][144] ), .Z(n29873) );
  IV U41432 ( .A(n38642), .Z(n38645) );
  XNOR U41433 ( .A(n38642), .B(n29872), .Z(n38644) );
  XOR U41434 ( .A(n38646), .B(n38647), .Z(n29872) );
  AND U41435 ( .A(\modmult_1/xin[1023] ), .B(n38648), .Z(n38647) );
  IV U41436 ( .A(n38646), .Z(n38648) );
  XOR U41437 ( .A(n38649), .B(mreg[145]), .Z(n38646) );
  NAND U41438 ( .A(n38650), .B(mul_pow), .Z(n38649) );
  XOR U41439 ( .A(mreg[145]), .B(creg[145]), .Z(n38650) );
  XOR U41440 ( .A(n38651), .B(n38652), .Z(n38642) );
  ANDN U41441 ( .A(n38653), .B(n29879), .Z(n38652) );
  XOR U41442 ( .A(n38654), .B(\modmult_1/zin[0][143] ), .Z(n29879) );
  IV U41443 ( .A(n38651), .Z(n38654) );
  XNOR U41444 ( .A(n38651), .B(n29878), .Z(n38653) );
  XOR U41445 ( .A(n38655), .B(n38656), .Z(n29878) );
  AND U41446 ( .A(\modmult_1/xin[1023] ), .B(n38657), .Z(n38656) );
  IV U41447 ( .A(n38655), .Z(n38657) );
  XOR U41448 ( .A(n38658), .B(mreg[144]), .Z(n38655) );
  NAND U41449 ( .A(n38659), .B(mul_pow), .Z(n38658) );
  XOR U41450 ( .A(mreg[144]), .B(creg[144]), .Z(n38659) );
  XOR U41451 ( .A(n38660), .B(n38661), .Z(n38651) );
  ANDN U41452 ( .A(n38662), .B(n29885), .Z(n38661) );
  XOR U41453 ( .A(n38663), .B(\modmult_1/zin[0][142] ), .Z(n29885) );
  IV U41454 ( .A(n38660), .Z(n38663) );
  XNOR U41455 ( .A(n38660), .B(n29884), .Z(n38662) );
  XOR U41456 ( .A(n38664), .B(n38665), .Z(n29884) );
  AND U41457 ( .A(\modmult_1/xin[1023] ), .B(n38666), .Z(n38665) );
  IV U41458 ( .A(n38664), .Z(n38666) );
  XOR U41459 ( .A(n38667), .B(mreg[143]), .Z(n38664) );
  NAND U41460 ( .A(n38668), .B(mul_pow), .Z(n38667) );
  XOR U41461 ( .A(mreg[143]), .B(creg[143]), .Z(n38668) );
  XOR U41462 ( .A(n38669), .B(n38670), .Z(n38660) );
  ANDN U41463 ( .A(n38671), .B(n29891), .Z(n38670) );
  XOR U41464 ( .A(n38672), .B(\modmult_1/zin[0][141] ), .Z(n29891) );
  IV U41465 ( .A(n38669), .Z(n38672) );
  XNOR U41466 ( .A(n38669), .B(n29890), .Z(n38671) );
  XOR U41467 ( .A(n38673), .B(n38674), .Z(n29890) );
  AND U41468 ( .A(\modmult_1/xin[1023] ), .B(n38675), .Z(n38674) );
  IV U41469 ( .A(n38673), .Z(n38675) );
  XOR U41470 ( .A(n38676), .B(mreg[142]), .Z(n38673) );
  NAND U41471 ( .A(n38677), .B(mul_pow), .Z(n38676) );
  XOR U41472 ( .A(mreg[142]), .B(creg[142]), .Z(n38677) );
  XOR U41473 ( .A(n38678), .B(n38679), .Z(n38669) );
  ANDN U41474 ( .A(n38680), .B(n29897), .Z(n38679) );
  XOR U41475 ( .A(n38681), .B(\modmult_1/zin[0][140] ), .Z(n29897) );
  IV U41476 ( .A(n38678), .Z(n38681) );
  XNOR U41477 ( .A(n38678), .B(n29896), .Z(n38680) );
  XOR U41478 ( .A(n38682), .B(n38683), .Z(n29896) );
  AND U41479 ( .A(\modmult_1/xin[1023] ), .B(n38684), .Z(n38683) );
  IV U41480 ( .A(n38682), .Z(n38684) );
  XOR U41481 ( .A(n38685), .B(mreg[141]), .Z(n38682) );
  NAND U41482 ( .A(n38686), .B(mul_pow), .Z(n38685) );
  XOR U41483 ( .A(mreg[141]), .B(creg[141]), .Z(n38686) );
  XOR U41484 ( .A(n38687), .B(n38688), .Z(n38678) );
  ANDN U41485 ( .A(n38689), .B(n29903), .Z(n38688) );
  XOR U41486 ( .A(n38690), .B(\modmult_1/zin[0][139] ), .Z(n29903) );
  IV U41487 ( .A(n38687), .Z(n38690) );
  XNOR U41488 ( .A(n38687), .B(n29902), .Z(n38689) );
  XOR U41489 ( .A(n38691), .B(n38692), .Z(n29902) );
  AND U41490 ( .A(\modmult_1/xin[1023] ), .B(n38693), .Z(n38692) );
  IV U41491 ( .A(n38691), .Z(n38693) );
  XOR U41492 ( .A(n38694), .B(mreg[140]), .Z(n38691) );
  NAND U41493 ( .A(n38695), .B(mul_pow), .Z(n38694) );
  XOR U41494 ( .A(mreg[140]), .B(creg[140]), .Z(n38695) );
  XOR U41495 ( .A(n38696), .B(n38697), .Z(n38687) );
  ANDN U41496 ( .A(n38698), .B(n29909), .Z(n38697) );
  XOR U41497 ( .A(n38699), .B(\modmult_1/zin[0][138] ), .Z(n29909) );
  IV U41498 ( .A(n38696), .Z(n38699) );
  XNOR U41499 ( .A(n38696), .B(n29908), .Z(n38698) );
  XOR U41500 ( .A(n38700), .B(n38701), .Z(n29908) );
  AND U41501 ( .A(\modmult_1/xin[1023] ), .B(n38702), .Z(n38701) );
  IV U41502 ( .A(n38700), .Z(n38702) );
  XOR U41503 ( .A(n38703), .B(mreg[139]), .Z(n38700) );
  NAND U41504 ( .A(n38704), .B(mul_pow), .Z(n38703) );
  XOR U41505 ( .A(mreg[139]), .B(creg[139]), .Z(n38704) );
  XOR U41506 ( .A(n38705), .B(n38706), .Z(n38696) );
  ANDN U41507 ( .A(n38707), .B(n29915), .Z(n38706) );
  XOR U41508 ( .A(n38708), .B(\modmult_1/zin[0][137] ), .Z(n29915) );
  IV U41509 ( .A(n38705), .Z(n38708) );
  XNOR U41510 ( .A(n38705), .B(n29914), .Z(n38707) );
  XOR U41511 ( .A(n38709), .B(n38710), .Z(n29914) );
  AND U41512 ( .A(\modmult_1/xin[1023] ), .B(n38711), .Z(n38710) );
  IV U41513 ( .A(n38709), .Z(n38711) );
  XOR U41514 ( .A(n38712), .B(mreg[138]), .Z(n38709) );
  NAND U41515 ( .A(n38713), .B(mul_pow), .Z(n38712) );
  XOR U41516 ( .A(mreg[138]), .B(creg[138]), .Z(n38713) );
  XOR U41517 ( .A(n38714), .B(n38715), .Z(n38705) );
  ANDN U41518 ( .A(n38716), .B(n29921), .Z(n38715) );
  XOR U41519 ( .A(n38717), .B(\modmult_1/zin[0][136] ), .Z(n29921) );
  IV U41520 ( .A(n38714), .Z(n38717) );
  XNOR U41521 ( .A(n38714), .B(n29920), .Z(n38716) );
  XOR U41522 ( .A(n38718), .B(n38719), .Z(n29920) );
  AND U41523 ( .A(\modmult_1/xin[1023] ), .B(n38720), .Z(n38719) );
  IV U41524 ( .A(n38718), .Z(n38720) );
  XOR U41525 ( .A(n38721), .B(mreg[137]), .Z(n38718) );
  NAND U41526 ( .A(n38722), .B(mul_pow), .Z(n38721) );
  XOR U41527 ( .A(mreg[137]), .B(creg[137]), .Z(n38722) );
  XOR U41528 ( .A(n38723), .B(n38724), .Z(n38714) );
  ANDN U41529 ( .A(n38725), .B(n29927), .Z(n38724) );
  XOR U41530 ( .A(n38726), .B(\modmult_1/zin[0][135] ), .Z(n29927) );
  IV U41531 ( .A(n38723), .Z(n38726) );
  XNOR U41532 ( .A(n38723), .B(n29926), .Z(n38725) );
  XOR U41533 ( .A(n38727), .B(n38728), .Z(n29926) );
  AND U41534 ( .A(\modmult_1/xin[1023] ), .B(n38729), .Z(n38728) );
  IV U41535 ( .A(n38727), .Z(n38729) );
  XOR U41536 ( .A(n38730), .B(mreg[136]), .Z(n38727) );
  NAND U41537 ( .A(n38731), .B(mul_pow), .Z(n38730) );
  XOR U41538 ( .A(mreg[136]), .B(creg[136]), .Z(n38731) );
  XOR U41539 ( .A(n38732), .B(n38733), .Z(n38723) );
  ANDN U41540 ( .A(n38734), .B(n29933), .Z(n38733) );
  XOR U41541 ( .A(n38735), .B(\modmult_1/zin[0][134] ), .Z(n29933) );
  IV U41542 ( .A(n38732), .Z(n38735) );
  XNOR U41543 ( .A(n38732), .B(n29932), .Z(n38734) );
  XOR U41544 ( .A(n38736), .B(n38737), .Z(n29932) );
  AND U41545 ( .A(\modmult_1/xin[1023] ), .B(n38738), .Z(n38737) );
  IV U41546 ( .A(n38736), .Z(n38738) );
  XOR U41547 ( .A(n38739), .B(mreg[135]), .Z(n38736) );
  NAND U41548 ( .A(n38740), .B(mul_pow), .Z(n38739) );
  XOR U41549 ( .A(mreg[135]), .B(creg[135]), .Z(n38740) );
  XOR U41550 ( .A(n38741), .B(n38742), .Z(n38732) );
  ANDN U41551 ( .A(n38743), .B(n29939), .Z(n38742) );
  XOR U41552 ( .A(n38744), .B(\modmult_1/zin[0][133] ), .Z(n29939) );
  IV U41553 ( .A(n38741), .Z(n38744) );
  XNOR U41554 ( .A(n38741), .B(n29938), .Z(n38743) );
  XOR U41555 ( .A(n38745), .B(n38746), .Z(n29938) );
  AND U41556 ( .A(\modmult_1/xin[1023] ), .B(n38747), .Z(n38746) );
  IV U41557 ( .A(n38745), .Z(n38747) );
  XOR U41558 ( .A(n38748), .B(mreg[134]), .Z(n38745) );
  NAND U41559 ( .A(n38749), .B(mul_pow), .Z(n38748) );
  XOR U41560 ( .A(mreg[134]), .B(creg[134]), .Z(n38749) );
  XOR U41561 ( .A(n38750), .B(n38751), .Z(n38741) );
  ANDN U41562 ( .A(n38752), .B(n29945), .Z(n38751) );
  XOR U41563 ( .A(n38753), .B(\modmult_1/zin[0][132] ), .Z(n29945) );
  IV U41564 ( .A(n38750), .Z(n38753) );
  XNOR U41565 ( .A(n38750), .B(n29944), .Z(n38752) );
  XOR U41566 ( .A(n38754), .B(n38755), .Z(n29944) );
  AND U41567 ( .A(\modmult_1/xin[1023] ), .B(n38756), .Z(n38755) );
  IV U41568 ( .A(n38754), .Z(n38756) );
  XOR U41569 ( .A(n38757), .B(mreg[133]), .Z(n38754) );
  NAND U41570 ( .A(n38758), .B(mul_pow), .Z(n38757) );
  XOR U41571 ( .A(mreg[133]), .B(creg[133]), .Z(n38758) );
  XOR U41572 ( .A(n38759), .B(n38760), .Z(n38750) );
  ANDN U41573 ( .A(n38761), .B(n29951), .Z(n38760) );
  XOR U41574 ( .A(n38762), .B(\modmult_1/zin[0][131] ), .Z(n29951) );
  IV U41575 ( .A(n38759), .Z(n38762) );
  XNOR U41576 ( .A(n38759), .B(n29950), .Z(n38761) );
  XOR U41577 ( .A(n38763), .B(n38764), .Z(n29950) );
  AND U41578 ( .A(\modmult_1/xin[1023] ), .B(n38765), .Z(n38764) );
  IV U41579 ( .A(n38763), .Z(n38765) );
  XOR U41580 ( .A(n38766), .B(mreg[132]), .Z(n38763) );
  NAND U41581 ( .A(n38767), .B(mul_pow), .Z(n38766) );
  XOR U41582 ( .A(mreg[132]), .B(creg[132]), .Z(n38767) );
  XOR U41583 ( .A(n38768), .B(n38769), .Z(n38759) );
  ANDN U41584 ( .A(n38770), .B(n29957), .Z(n38769) );
  XOR U41585 ( .A(n38771), .B(\modmult_1/zin[0][130] ), .Z(n29957) );
  IV U41586 ( .A(n38768), .Z(n38771) );
  XNOR U41587 ( .A(n38768), .B(n29956), .Z(n38770) );
  XOR U41588 ( .A(n38772), .B(n38773), .Z(n29956) );
  AND U41589 ( .A(\modmult_1/xin[1023] ), .B(n38774), .Z(n38773) );
  IV U41590 ( .A(n38772), .Z(n38774) );
  XOR U41591 ( .A(n38775), .B(mreg[131]), .Z(n38772) );
  NAND U41592 ( .A(n38776), .B(mul_pow), .Z(n38775) );
  XOR U41593 ( .A(mreg[131]), .B(creg[131]), .Z(n38776) );
  XOR U41594 ( .A(n38777), .B(n38778), .Z(n38768) );
  ANDN U41595 ( .A(n38779), .B(n29963), .Z(n38778) );
  XOR U41596 ( .A(n38780), .B(\modmult_1/zin[0][129] ), .Z(n29963) );
  IV U41597 ( .A(n38777), .Z(n38780) );
  XNOR U41598 ( .A(n38777), .B(n29962), .Z(n38779) );
  XOR U41599 ( .A(n38781), .B(n38782), .Z(n29962) );
  AND U41600 ( .A(\modmult_1/xin[1023] ), .B(n38783), .Z(n38782) );
  IV U41601 ( .A(n38781), .Z(n38783) );
  XOR U41602 ( .A(n38784), .B(mreg[130]), .Z(n38781) );
  NAND U41603 ( .A(n38785), .B(mul_pow), .Z(n38784) );
  XOR U41604 ( .A(mreg[130]), .B(creg[130]), .Z(n38785) );
  XOR U41605 ( .A(n38786), .B(n38787), .Z(n38777) );
  ANDN U41606 ( .A(n38788), .B(n29969), .Z(n38787) );
  XOR U41607 ( .A(n38789), .B(\modmult_1/zin[0][128] ), .Z(n29969) );
  IV U41608 ( .A(n38786), .Z(n38789) );
  XNOR U41609 ( .A(n38786), .B(n29968), .Z(n38788) );
  XOR U41610 ( .A(n38790), .B(n38791), .Z(n29968) );
  AND U41611 ( .A(\modmult_1/xin[1023] ), .B(n38792), .Z(n38791) );
  IV U41612 ( .A(n38790), .Z(n38792) );
  XOR U41613 ( .A(n38793), .B(mreg[129]), .Z(n38790) );
  NAND U41614 ( .A(n38794), .B(mul_pow), .Z(n38793) );
  XOR U41615 ( .A(mreg[129]), .B(creg[129]), .Z(n38794) );
  XOR U41616 ( .A(n38795), .B(n38796), .Z(n38786) );
  ANDN U41617 ( .A(n38797), .B(n29975), .Z(n38796) );
  XOR U41618 ( .A(n38798), .B(\modmult_1/zin[0][127] ), .Z(n29975) );
  IV U41619 ( .A(n38795), .Z(n38798) );
  XNOR U41620 ( .A(n38795), .B(n29974), .Z(n38797) );
  XOR U41621 ( .A(n38799), .B(n38800), .Z(n29974) );
  AND U41622 ( .A(\modmult_1/xin[1023] ), .B(n38801), .Z(n38800) );
  IV U41623 ( .A(n38799), .Z(n38801) );
  XOR U41624 ( .A(n38802), .B(mreg[128]), .Z(n38799) );
  NAND U41625 ( .A(n38803), .B(mul_pow), .Z(n38802) );
  XOR U41626 ( .A(mreg[128]), .B(creg[128]), .Z(n38803) );
  XOR U41627 ( .A(n38804), .B(n38805), .Z(n38795) );
  ANDN U41628 ( .A(n38806), .B(n29981), .Z(n38805) );
  XOR U41629 ( .A(n38807), .B(\modmult_1/zin[0][126] ), .Z(n29981) );
  IV U41630 ( .A(n38804), .Z(n38807) );
  XNOR U41631 ( .A(n38804), .B(n29980), .Z(n38806) );
  XOR U41632 ( .A(n38808), .B(n38809), .Z(n29980) );
  AND U41633 ( .A(\modmult_1/xin[1023] ), .B(n38810), .Z(n38809) );
  IV U41634 ( .A(n38808), .Z(n38810) );
  XOR U41635 ( .A(n38811), .B(mreg[127]), .Z(n38808) );
  NAND U41636 ( .A(n38812), .B(mul_pow), .Z(n38811) );
  XOR U41637 ( .A(mreg[127]), .B(creg[127]), .Z(n38812) );
  XOR U41638 ( .A(n38813), .B(n38814), .Z(n38804) );
  ANDN U41639 ( .A(n38815), .B(n29987), .Z(n38814) );
  XOR U41640 ( .A(n38816), .B(\modmult_1/zin[0][125] ), .Z(n29987) );
  IV U41641 ( .A(n38813), .Z(n38816) );
  XNOR U41642 ( .A(n38813), .B(n29986), .Z(n38815) );
  XOR U41643 ( .A(n38817), .B(n38818), .Z(n29986) );
  AND U41644 ( .A(\modmult_1/xin[1023] ), .B(n38819), .Z(n38818) );
  IV U41645 ( .A(n38817), .Z(n38819) );
  XOR U41646 ( .A(n38820), .B(mreg[126]), .Z(n38817) );
  NAND U41647 ( .A(n38821), .B(mul_pow), .Z(n38820) );
  XOR U41648 ( .A(mreg[126]), .B(creg[126]), .Z(n38821) );
  XOR U41649 ( .A(n38822), .B(n38823), .Z(n38813) );
  ANDN U41650 ( .A(n38824), .B(n29993), .Z(n38823) );
  XOR U41651 ( .A(n38825), .B(\modmult_1/zin[0][124] ), .Z(n29993) );
  IV U41652 ( .A(n38822), .Z(n38825) );
  XNOR U41653 ( .A(n38822), .B(n29992), .Z(n38824) );
  XOR U41654 ( .A(n38826), .B(n38827), .Z(n29992) );
  AND U41655 ( .A(\modmult_1/xin[1023] ), .B(n38828), .Z(n38827) );
  IV U41656 ( .A(n38826), .Z(n38828) );
  XOR U41657 ( .A(n38829), .B(mreg[125]), .Z(n38826) );
  NAND U41658 ( .A(n38830), .B(mul_pow), .Z(n38829) );
  XOR U41659 ( .A(mreg[125]), .B(creg[125]), .Z(n38830) );
  XOR U41660 ( .A(n38831), .B(n38832), .Z(n38822) );
  ANDN U41661 ( .A(n38833), .B(n29999), .Z(n38832) );
  XOR U41662 ( .A(n38834), .B(\modmult_1/zin[0][123] ), .Z(n29999) );
  IV U41663 ( .A(n38831), .Z(n38834) );
  XNOR U41664 ( .A(n38831), .B(n29998), .Z(n38833) );
  XOR U41665 ( .A(n38835), .B(n38836), .Z(n29998) );
  AND U41666 ( .A(\modmult_1/xin[1023] ), .B(n38837), .Z(n38836) );
  IV U41667 ( .A(n38835), .Z(n38837) );
  XOR U41668 ( .A(n38838), .B(mreg[124]), .Z(n38835) );
  NAND U41669 ( .A(n38839), .B(mul_pow), .Z(n38838) );
  XOR U41670 ( .A(mreg[124]), .B(creg[124]), .Z(n38839) );
  XOR U41671 ( .A(n38840), .B(n38841), .Z(n38831) );
  ANDN U41672 ( .A(n38842), .B(n30005), .Z(n38841) );
  XOR U41673 ( .A(n38843), .B(\modmult_1/zin[0][122] ), .Z(n30005) );
  IV U41674 ( .A(n38840), .Z(n38843) );
  XNOR U41675 ( .A(n38840), .B(n30004), .Z(n38842) );
  XOR U41676 ( .A(n38844), .B(n38845), .Z(n30004) );
  AND U41677 ( .A(\modmult_1/xin[1023] ), .B(n38846), .Z(n38845) );
  IV U41678 ( .A(n38844), .Z(n38846) );
  XOR U41679 ( .A(n38847), .B(mreg[123]), .Z(n38844) );
  NAND U41680 ( .A(n38848), .B(mul_pow), .Z(n38847) );
  XOR U41681 ( .A(mreg[123]), .B(creg[123]), .Z(n38848) );
  XOR U41682 ( .A(n38849), .B(n38850), .Z(n38840) );
  ANDN U41683 ( .A(n38851), .B(n30011), .Z(n38850) );
  XOR U41684 ( .A(n38852), .B(\modmult_1/zin[0][121] ), .Z(n30011) );
  IV U41685 ( .A(n38849), .Z(n38852) );
  XNOR U41686 ( .A(n38849), .B(n30010), .Z(n38851) );
  XOR U41687 ( .A(n38853), .B(n38854), .Z(n30010) );
  AND U41688 ( .A(\modmult_1/xin[1023] ), .B(n38855), .Z(n38854) );
  IV U41689 ( .A(n38853), .Z(n38855) );
  XOR U41690 ( .A(n38856), .B(mreg[122]), .Z(n38853) );
  NAND U41691 ( .A(n38857), .B(mul_pow), .Z(n38856) );
  XOR U41692 ( .A(mreg[122]), .B(creg[122]), .Z(n38857) );
  XOR U41693 ( .A(n38858), .B(n38859), .Z(n38849) );
  ANDN U41694 ( .A(n38860), .B(n30017), .Z(n38859) );
  XOR U41695 ( .A(n38861), .B(\modmult_1/zin[0][120] ), .Z(n30017) );
  IV U41696 ( .A(n38858), .Z(n38861) );
  XNOR U41697 ( .A(n38858), .B(n30016), .Z(n38860) );
  XOR U41698 ( .A(n38862), .B(n38863), .Z(n30016) );
  AND U41699 ( .A(\modmult_1/xin[1023] ), .B(n38864), .Z(n38863) );
  IV U41700 ( .A(n38862), .Z(n38864) );
  XOR U41701 ( .A(n38865), .B(mreg[121]), .Z(n38862) );
  NAND U41702 ( .A(n38866), .B(mul_pow), .Z(n38865) );
  XOR U41703 ( .A(mreg[121]), .B(creg[121]), .Z(n38866) );
  XOR U41704 ( .A(n38867), .B(n38868), .Z(n38858) );
  ANDN U41705 ( .A(n38869), .B(n30023), .Z(n38868) );
  XOR U41706 ( .A(n38870), .B(\modmult_1/zin[0][119] ), .Z(n30023) );
  IV U41707 ( .A(n38867), .Z(n38870) );
  XNOR U41708 ( .A(n38867), .B(n30022), .Z(n38869) );
  XOR U41709 ( .A(n38871), .B(n38872), .Z(n30022) );
  AND U41710 ( .A(\modmult_1/xin[1023] ), .B(n38873), .Z(n38872) );
  IV U41711 ( .A(n38871), .Z(n38873) );
  XOR U41712 ( .A(n38874), .B(mreg[120]), .Z(n38871) );
  NAND U41713 ( .A(n38875), .B(mul_pow), .Z(n38874) );
  XOR U41714 ( .A(mreg[120]), .B(creg[120]), .Z(n38875) );
  XOR U41715 ( .A(n38876), .B(n38877), .Z(n38867) );
  ANDN U41716 ( .A(n38878), .B(n30029), .Z(n38877) );
  XOR U41717 ( .A(n38879), .B(\modmult_1/zin[0][118] ), .Z(n30029) );
  IV U41718 ( .A(n38876), .Z(n38879) );
  XNOR U41719 ( .A(n38876), .B(n30028), .Z(n38878) );
  XOR U41720 ( .A(n38880), .B(n38881), .Z(n30028) );
  AND U41721 ( .A(\modmult_1/xin[1023] ), .B(n38882), .Z(n38881) );
  IV U41722 ( .A(n38880), .Z(n38882) );
  XOR U41723 ( .A(n38883), .B(mreg[119]), .Z(n38880) );
  NAND U41724 ( .A(n38884), .B(mul_pow), .Z(n38883) );
  XOR U41725 ( .A(mreg[119]), .B(creg[119]), .Z(n38884) );
  XOR U41726 ( .A(n38885), .B(n38886), .Z(n38876) );
  ANDN U41727 ( .A(n38887), .B(n30035), .Z(n38886) );
  XOR U41728 ( .A(n38888), .B(\modmult_1/zin[0][117] ), .Z(n30035) );
  IV U41729 ( .A(n38885), .Z(n38888) );
  XNOR U41730 ( .A(n38885), .B(n30034), .Z(n38887) );
  XOR U41731 ( .A(n38889), .B(n38890), .Z(n30034) );
  AND U41732 ( .A(\modmult_1/xin[1023] ), .B(n38891), .Z(n38890) );
  IV U41733 ( .A(n38889), .Z(n38891) );
  XOR U41734 ( .A(n38892), .B(mreg[118]), .Z(n38889) );
  NAND U41735 ( .A(n38893), .B(mul_pow), .Z(n38892) );
  XOR U41736 ( .A(mreg[118]), .B(creg[118]), .Z(n38893) );
  XOR U41737 ( .A(n38894), .B(n38895), .Z(n38885) );
  ANDN U41738 ( .A(n38896), .B(n30041), .Z(n38895) );
  XOR U41739 ( .A(n38897), .B(\modmult_1/zin[0][116] ), .Z(n30041) );
  IV U41740 ( .A(n38894), .Z(n38897) );
  XNOR U41741 ( .A(n38894), .B(n30040), .Z(n38896) );
  XOR U41742 ( .A(n38898), .B(n38899), .Z(n30040) );
  AND U41743 ( .A(\modmult_1/xin[1023] ), .B(n38900), .Z(n38899) );
  IV U41744 ( .A(n38898), .Z(n38900) );
  XOR U41745 ( .A(n38901), .B(mreg[117]), .Z(n38898) );
  NAND U41746 ( .A(n38902), .B(mul_pow), .Z(n38901) );
  XOR U41747 ( .A(mreg[117]), .B(creg[117]), .Z(n38902) );
  XOR U41748 ( .A(n38903), .B(n38904), .Z(n38894) );
  ANDN U41749 ( .A(n38905), .B(n30047), .Z(n38904) );
  XOR U41750 ( .A(n38906), .B(\modmult_1/zin[0][115] ), .Z(n30047) );
  IV U41751 ( .A(n38903), .Z(n38906) );
  XNOR U41752 ( .A(n38903), .B(n30046), .Z(n38905) );
  XOR U41753 ( .A(n38907), .B(n38908), .Z(n30046) );
  AND U41754 ( .A(\modmult_1/xin[1023] ), .B(n38909), .Z(n38908) );
  IV U41755 ( .A(n38907), .Z(n38909) );
  XOR U41756 ( .A(n38910), .B(mreg[116]), .Z(n38907) );
  NAND U41757 ( .A(n38911), .B(mul_pow), .Z(n38910) );
  XOR U41758 ( .A(mreg[116]), .B(creg[116]), .Z(n38911) );
  XOR U41759 ( .A(n38912), .B(n38913), .Z(n38903) );
  ANDN U41760 ( .A(n38914), .B(n30053), .Z(n38913) );
  XOR U41761 ( .A(n38915), .B(\modmult_1/zin[0][114] ), .Z(n30053) );
  IV U41762 ( .A(n38912), .Z(n38915) );
  XNOR U41763 ( .A(n38912), .B(n30052), .Z(n38914) );
  XOR U41764 ( .A(n38916), .B(n38917), .Z(n30052) );
  AND U41765 ( .A(\modmult_1/xin[1023] ), .B(n38918), .Z(n38917) );
  IV U41766 ( .A(n38916), .Z(n38918) );
  XOR U41767 ( .A(n38919), .B(mreg[115]), .Z(n38916) );
  NAND U41768 ( .A(n38920), .B(mul_pow), .Z(n38919) );
  XOR U41769 ( .A(mreg[115]), .B(creg[115]), .Z(n38920) );
  XOR U41770 ( .A(n38921), .B(n38922), .Z(n38912) );
  ANDN U41771 ( .A(n38923), .B(n30059), .Z(n38922) );
  XOR U41772 ( .A(n38924), .B(\modmult_1/zin[0][113] ), .Z(n30059) );
  IV U41773 ( .A(n38921), .Z(n38924) );
  XNOR U41774 ( .A(n38921), .B(n30058), .Z(n38923) );
  XOR U41775 ( .A(n38925), .B(n38926), .Z(n30058) );
  AND U41776 ( .A(\modmult_1/xin[1023] ), .B(n38927), .Z(n38926) );
  IV U41777 ( .A(n38925), .Z(n38927) );
  XOR U41778 ( .A(n38928), .B(mreg[114]), .Z(n38925) );
  NAND U41779 ( .A(n38929), .B(mul_pow), .Z(n38928) );
  XOR U41780 ( .A(mreg[114]), .B(creg[114]), .Z(n38929) );
  XOR U41781 ( .A(n38930), .B(n38931), .Z(n38921) );
  ANDN U41782 ( .A(n38932), .B(n30065), .Z(n38931) );
  XOR U41783 ( .A(n38933), .B(\modmult_1/zin[0][112] ), .Z(n30065) );
  IV U41784 ( .A(n38930), .Z(n38933) );
  XNOR U41785 ( .A(n38930), .B(n30064), .Z(n38932) );
  XOR U41786 ( .A(n38934), .B(n38935), .Z(n30064) );
  AND U41787 ( .A(\modmult_1/xin[1023] ), .B(n38936), .Z(n38935) );
  IV U41788 ( .A(n38934), .Z(n38936) );
  XOR U41789 ( .A(n38937), .B(mreg[113]), .Z(n38934) );
  NAND U41790 ( .A(n38938), .B(mul_pow), .Z(n38937) );
  XOR U41791 ( .A(mreg[113]), .B(creg[113]), .Z(n38938) );
  XOR U41792 ( .A(n38939), .B(n38940), .Z(n38930) );
  ANDN U41793 ( .A(n38941), .B(n30071), .Z(n38940) );
  XOR U41794 ( .A(n38942), .B(\modmult_1/zin[0][111] ), .Z(n30071) );
  IV U41795 ( .A(n38939), .Z(n38942) );
  XNOR U41796 ( .A(n38939), .B(n30070), .Z(n38941) );
  XOR U41797 ( .A(n38943), .B(n38944), .Z(n30070) );
  AND U41798 ( .A(\modmult_1/xin[1023] ), .B(n38945), .Z(n38944) );
  IV U41799 ( .A(n38943), .Z(n38945) );
  XOR U41800 ( .A(n38946), .B(mreg[112]), .Z(n38943) );
  NAND U41801 ( .A(n38947), .B(mul_pow), .Z(n38946) );
  XOR U41802 ( .A(mreg[112]), .B(creg[112]), .Z(n38947) );
  XOR U41803 ( .A(n38948), .B(n38949), .Z(n38939) );
  ANDN U41804 ( .A(n38950), .B(n30077), .Z(n38949) );
  XOR U41805 ( .A(n38951), .B(\modmult_1/zin[0][110] ), .Z(n30077) );
  IV U41806 ( .A(n38948), .Z(n38951) );
  XNOR U41807 ( .A(n38948), .B(n30076), .Z(n38950) );
  XOR U41808 ( .A(n38952), .B(n38953), .Z(n30076) );
  AND U41809 ( .A(\modmult_1/xin[1023] ), .B(n38954), .Z(n38953) );
  IV U41810 ( .A(n38952), .Z(n38954) );
  XOR U41811 ( .A(n38955), .B(mreg[111]), .Z(n38952) );
  NAND U41812 ( .A(n38956), .B(mul_pow), .Z(n38955) );
  XOR U41813 ( .A(mreg[111]), .B(creg[111]), .Z(n38956) );
  XOR U41814 ( .A(n38957), .B(n38958), .Z(n38948) );
  ANDN U41815 ( .A(n38959), .B(n30083), .Z(n38958) );
  XOR U41816 ( .A(n38960), .B(\modmult_1/zin[0][109] ), .Z(n30083) );
  IV U41817 ( .A(n38957), .Z(n38960) );
  XNOR U41818 ( .A(n38957), .B(n30082), .Z(n38959) );
  XOR U41819 ( .A(n38961), .B(n38962), .Z(n30082) );
  AND U41820 ( .A(\modmult_1/xin[1023] ), .B(n38963), .Z(n38962) );
  IV U41821 ( .A(n38961), .Z(n38963) );
  XOR U41822 ( .A(n38964), .B(mreg[110]), .Z(n38961) );
  NAND U41823 ( .A(n38965), .B(mul_pow), .Z(n38964) );
  XOR U41824 ( .A(mreg[110]), .B(creg[110]), .Z(n38965) );
  XOR U41825 ( .A(n38966), .B(n38967), .Z(n38957) );
  ANDN U41826 ( .A(n38968), .B(n30089), .Z(n38967) );
  XOR U41827 ( .A(n38969), .B(\modmult_1/zin[0][108] ), .Z(n30089) );
  IV U41828 ( .A(n38966), .Z(n38969) );
  XNOR U41829 ( .A(n38966), .B(n30088), .Z(n38968) );
  XOR U41830 ( .A(n38970), .B(n38971), .Z(n30088) );
  AND U41831 ( .A(\modmult_1/xin[1023] ), .B(n38972), .Z(n38971) );
  IV U41832 ( .A(n38970), .Z(n38972) );
  XOR U41833 ( .A(n38973), .B(mreg[109]), .Z(n38970) );
  NAND U41834 ( .A(n38974), .B(mul_pow), .Z(n38973) );
  XOR U41835 ( .A(mreg[109]), .B(creg[109]), .Z(n38974) );
  XOR U41836 ( .A(n38975), .B(n38976), .Z(n38966) );
  ANDN U41837 ( .A(n38977), .B(n30095), .Z(n38976) );
  XOR U41838 ( .A(n38978), .B(\modmult_1/zin[0][107] ), .Z(n30095) );
  IV U41839 ( .A(n38975), .Z(n38978) );
  XNOR U41840 ( .A(n38975), .B(n30094), .Z(n38977) );
  XOR U41841 ( .A(n38979), .B(n38980), .Z(n30094) );
  AND U41842 ( .A(\modmult_1/xin[1023] ), .B(n38981), .Z(n38980) );
  IV U41843 ( .A(n38979), .Z(n38981) );
  XOR U41844 ( .A(n38982), .B(mreg[108]), .Z(n38979) );
  NAND U41845 ( .A(n38983), .B(mul_pow), .Z(n38982) );
  XOR U41846 ( .A(mreg[108]), .B(creg[108]), .Z(n38983) );
  XOR U41847 ( .A(n38984), .B(n38985), .Z(n38975) );
  ANDN U41848 ( .A(n38986), .B(n30101), .Z(n38985) );
  XOR U41849 ( .A(n38987), .B(\modmult_1/zin[0][106] ), .Z(n30101) );
  IV U41850 ( .A(n38984), .Z(n38987) );
  XNOR U41851 ( .A(n38984), .B(n30100), .Z(n38986) );
  XOR U41852 ( .A(n38988), .B(n38989), .Z(n30100) );
  AND U41853 ( .A(\modmult_1/xin[1023] ), .B(n38990), .Z(n38989) );
  IV U41854 ( .A(n38988), .Z(n38990) );
  XOR U41855 ( .A(n38991), .B(mreg[107]), .Z(n38988) );
  NAND U41856 ( .A(n38992), .B(mul_pow), .Z(n38991) );
  XOR U41857 ( .A(mreg[107]), .B(creg[107]), .Z(n38992) );
  XOR U41858 ( .A(n38993), .B(n38994), .Z(n38984) );
  ANDN U41859 ( .A(n38995), .B(n30107), .Z(n38994) );
  XOR U41860 ( .A(n38996), .B(\modmult_1/zin[0][105] ), .Z(n30107) );
  IV U41861 ( .A(n38993), .Z(n38996) );
  XNOR U41862 ( .A(n38993), .B(n30106), .Z(n38995) );
  XOR U41863 ( .A(n38997), .B(n38998), .Z(n30106) );
  AND U41864 ( .A(\modmult_1/xin[1023] ), .B(n38999), .Z(n38998) );
  IV U41865 ( .A(n38997), .Z(n38999) );
  XOR U41866 ( .A(n39000), .B(mreg[106]), .Z(n38997) );
  NAND U41867 ( .A(n39001), .B(mul_pow), .Z(n39000) );
  XOR U41868 ( .A(mreg[106]), .B(creg[106]), .Z(n39001) );
  XOR U41869 ( .A(n39002), .B(n39003), .Z(n38993) );
  ANDN U41870 ( .A(n39004), .B(n30113), .Z(n39003) );
  XOR U41871 ( .A(n39005), .B(\modmult_1/zin[0][104] ), .Z(n30113) );
  IV U41872 ( .A(n39002), .Z(n39005) );
  XNOR U41873 ( .A(n39002), .B(n30112), .Z(n39004) );
  XOR U41874 ( .A(n39006), .B(n39007), .Z(n30112) );
  AND U41875 ( .A(\modmult_1/xin[1023] ), .B(n39008), .Z(n39007) );
  IV U41876 ( .A(n39006), .Z(n39008) );
  XOR U41877 ( .A(n39009), .B(mreg[105]), .Z(n39006) );
  NAND U41878 ( .A(n39010), .B(mul_pow), .Z(n39009) );
  XOR U41879 ( .A(mreg[105]), .B(creg[105]), .Z(n39010) );
  XOR U41880 ( .A(n39011), .B(n39012), .Z(n39002) );
  ANDN U41881 ( .A(n39013), .B(n30119), .Z(n39012) );
  XOR U41882 ( .A(n39014), .B(\modmult_1/zin[0][103] ), .Z(n30119) );
  IV U41883 ( .A(n39011), .Z(n39014) );
  XNOR U41884 ( .A(n39011), .B(n30118), .Z(n39013) );
  XOR U41885 ( .A(n39015), .B(n39016), .Z(n30118) );
  AND U41886 ( .A(\modmult_1/xin[1023] ), .B(n39017), .Z(n39016) );
  IV U41887 ( .A(n39015), .Z(n39017) );
  XOR U41888 ( .A(n39018), .B(mreg[104]), .Z(n39015) );
  NAND U41889 ( .A(n39019), .B(mul_pow), .Z(n39018) );
  XOR U41890 ( .A(mreg[104]), .B(creg[104]), .Z(n39019) );
  XOR U41891 ( .A(n39020), .B(n39021), .Z(n39011) );
  ANDN U41892 ( .A(n39022), .B(n30125), .Z(n39021) );
  XOR U41893 ( .A(n39023), .B(\modmult_1/zin[0][102] ), .Z(n30125) );
  IV U41894 ( .A(n39020), .Z(n39023) );
  XNOR U41895 ( .A(n39020), .B(n30124), .Z(n39022) );
  XOR U41896 ( .A(n39024), .B(n39025), .Z(n30124) );
  AND U41897 ( .A(\modmult_1/xin[1023] ), .B(n39026), .Z(n39025) );
  IV U41898 ( .A(n39024), .Z(n39026) );
  XOR U41899 ( .A(n39027), .B(mreg[103]), .Z(n39024) );
  NAND U41900 ( .A(n39028), .B(mul_pow), .Z(n39027) );
  XOR U41901 ( .A(mreg[103]), .B(creg[103]), .Z(n39028) );
  XOR U41902 ( .A(n39029), .B(n39030), .Z(n39020) );
  ANDN U41903 ( .A(n39031), .B(n30131), .Z(n39030) );
  XOR U41904 ( .A(n39032), .B(\modmult_1/zin[0][101] ), .Z(n30131) );
  IV U41905 ( .A(n39029), .Z(n39032) );
  XNOR U41906 ( .A(n39029), .B(n30130), .Z(n39031) );
  XOR U41907 ( .A(n39033), .B(n39034), .Z(n30130) );
  AND U41908 ( .A(\modmult_1/xin[1023] ), .B(n39035), .Z(n39034) );
  IV U41909 ( .A(n39033), .Z(n39035) );
  XOR U41910 ( .A(n39036), .B(mreg[102]), .Z(n39033) );
  NAND U41911 ( .A(n39037), .B(mul_pow), .Z(n39036) );
  XOR U41912 ( .A(mreg[102]), .B(creg[102]), .Z(n39037) );
  XOR U41913 ( .A(n39038), .B(n39039), .Z(n39029) );
  ANDN U41914 ( .A(n39040), .B(n30137), .Z(n39039) );
  XOR U41915 ( .A(n39041), .B(\modmult_1/zin[0][100] ), .Z(n30137) );
  IV U41916 ( .A(n39038), .Z(n39041) );
  XNOR U41917 ( .A(n39038), .B(n30136), .Z(n39040) );
  XOR U41918 ( .A(n39042), .B(n39043), .Z(n30136) );
  AND U41919 ( .A(\modmult_1/xin[1023] ), .B(n39044), .Z(n39043) );
  IV U41920 ( .A(n39042), .Z(n39044) );
  XOR U41921 ( .A(n39045), .B(mreg[101]), .Z(n39042) );
  NAND U41922 ( .A(n39046), .B(mul_pow), .Z(n39045) );
  XOR U41923 ( .A(mreg[101]), .B(creg[101]), .Z(n39046) );
  XOR U41924 ( .A(n39047), .B(n39048), .Z(n39038) );
  ANDN U41925 ( .A(n39049), .B(n30143), .Z(n39048) );
  XOR U41926 ( .A(n39050), .B(\modmult_1/zin[0][99] ), .Z(n30143) );
  IV U41927 ( .A(n39047), .Z(n39050) );
  XNOR U41928 ( .A(n39047), .B(n30142), .Z(n39049) );
  XOR U41929 ( .A(n39051), .B(n39052), .Z(n30142) );
  AND U41930 ( .A(\modmult_1/xin[1023] ), .B(n39053), .Z(n39052) );
  IV U41931 ( .A(n39051), .Z(n39053) );
  XOR U41932 ( .A(n39054), .B(mreg[100]), .Z(n39051) );
  NAND U41933 ( .A(n39055), .B(mul_pow), .Z(n39054) );
  XOR U41934 ( .A(mreg[100]), .B(creg[100]), .Z(n39055) );
  XOR U41935 ( .A(n39056), .B(n39057), .Z(n39047) );
  ANDN U41936 ( .A(n39058), .B(n30149), .Z(n39057) );
  XOR U41937 ( .A(n39059), .B(\modmult_1/zin[0][98] ), .Z(n30149) );
  IV U41938 ( .A(n39056), .Z(n39059) );
  XNOR U41939 ( .A(n39056), .B(n30148), .Z(n39058) );
  XOR U41940 ( .A(n39060), .B(n39061), .Z(n30148) );
  AND U41941 ( .A(\modmult_1/xin[1023] ), .B(n39062), .Z(n39061) );
  IV U41942 ( .A(n39060), .Z(n39062) );
  XOR U41943 ( .A(n39063), .B(mreg[99]), .Z(n39060) );
  NAND U41944 ( .A(n39064), .B(mul_pow), .Z(n39063) );
  XOR U41945 ( .A(mreg[99]), .B(creg[99]), .Z(n39064) );
  XOR U41946 ( .A(n39065), .B(n39066), .Z(n39056) );
  ANDN U41947 ( .A(n39067), .B(n30155), .Z(n39066) );
  XOR U41948 ( .A(n39068), .B(\modmult_1/zin[0][97] ), .Z(n30155) );
  IV U41949 ( .A(n39065), .Z(n39068) );
  XNOR U41950 ( .A(n39065), .B(n30154), .Z(n39067) );
  XOR U41951 ( .A(n39069), .B(n39070), .Z(n30154) );
  AND U41952 ( .A(\modmult_1/xin[1023] ), .B(n39071), .Z(n39070) );
  IV U41953 ( .A(n39069), .Z(n39071) );
  XOR U41954 ( .A(n39072), .B(mreg[98]), .Z(n39069) );
  NAND U41955 ( .A(n39073), .B(mul_pow), .Z(n39072) );
  XOR U41956 ( .A(mreg[98]), .B(creg[98]), .Z(n39073) );
  XOR U41957 ( .A(n39074), .B(n39075), .Z(n39065) );
  ANDN U41958 ( .A(n39076), .B(n30161), .Z(n39075) );
  XOR U41959 ( .A(n39077), .B(\modmult_1/zin[0][96] ), .Z(n30161) );
  IV U41960 ( .A(n39074), .Z(n39077) );
  XNOR U41961 ( .A(n39074), .B(n30160), .Z(n39076) );
  XOR U41962 ( .A(n39078), .B(n39079), .Z(n30160) );
  AND U41963 ( .A(\modmult_1/xin[1023] ), .B(n39080), .Z(n39079) );
  IV U41964 ( .A(n39078), .Z(n39080) );
  XOR U41965 ( .A(n39081), .B(mreg[97]), .Z(n39078) );
  NAND U41966 ( .A(n39082), .B(mul_pow), .Z(n39081) );
  XOR U41967 ( .A(mreg[97]), .B(creg[97]), .Z(n39082) );
  XOR U41968 ( .A(n39083), .B(n39084), .Z(n39074) );
  ANDN U41969 ( .A(n39085), .B(n30167), .Z(n39084) );
  XOR U41970 ( .A(n39086), .B(\modmult_1/zin[0][95] ), .Z(n30167) );
  IV U41971 ( .A(n39083), .Z(n39086) );
  XNOR U41972 ( .A(n39083), .B(n30166), .Z(n39085) );
  XOR U41973 ( .A(n39087), .B(n39088), .Z(n30166) );
  AND U41974 ( .A(\modmult_1/xin[1023] ), .B(n39089), .Z(n39088) );
  IV U41975 ( .A(n39087), .Z(n39089) );
  XOR U41976 ( .A(n39090), .B(mreg[96]), .Z(n39087) );
  NAND U41977 ( .A(n39091), .B(mul_pow), .Z(n39090) );
  XOR U41978 ( .A(mreg[96]), .B(creg[96]), .Z(n39091) );
  XOR U41979 ( .A(n39092), .B(n39093), .Z(n39083) );
  ANDN U41980 ( .A(n39094), .B(n30173), .Z(n39093) );
  XOR U41981 ( .A(n39095), .B(\modmult_1/zin[0][94] ), .Z(n30173) );
  IV U41982 ( .A(n39092), .Z(n39095) );
  XNOR U41983 ( .A(n39092), .B(n30172), .Z(n39094) );
  XOR U41984 ( .A(n39096), .B(n39097), .Z(n30172) );
  AND U41985 ( .A(\modmult_1/xin[1023] ), .B(n39098), .Z(n39097) );
  IV U41986 ( .A(n39096), .Z(n39098) );
  XOR U41987 ( .A(n39099), .B(mreg[95]), .Z(n39096) );
  NAND U41988 ( .A(n39100), .B(mul_pow), .Z(n39099) );
  XOR U41989 ( .A(mreg[95]), .B(creg[95]), .Z(n39100) );
  XOR U41990 ( .A(n39101), .B(n39102), .Z(n39092) );
  ANDN U41991 ( .A(n39103), .B(n30179), .Z(n39102) );
  XOR U41992 ( .A(n39104), .B(\modmult_1/zin[0][93] ), .Z(n30179) );
  IV U41993 ( .A(n39101), .Z(n39104) );
  XNOR U41994 ( .A(n39101), .B(n30178), .Z(n39103) );
  XOR U41995 ( .A(n39105), .B(n39106), .Z(n30178) );
  AND U41996 ( .A(\modmult_1/xin[1023] ), .B(n39107), .Z(n39106) );
  IV U41997 ( .A(n39105), .Z(n39107) );
  XOR U41998 ( .A(n39108), .B(mreg[94]), .Z(n39105) );
  NAND U41999 ( .A(n39109), .B(mul_pow), .Z(n39108) );
  XOR U42000 ( .A(mreg[94]), .B(creg[94]), .Z(n39109) );
  XOR U42001 ( .A(n39110), .B(n39111), .Z(n39101) );
  ANDN U42002 ( .A(n39112), .B(n30185), .Z(n39111) );
  XOR U42003 ( .A(n39113), .B(\modmult_1/zin[0][92] ), .Z(n30185) );
  IV U42004 ( .A(n39110), .Z(n39113) );
  XNOR U42005 ( .A(n39110), .B(n30184), .Z(n39112) );
  XOR U42006 ( .A(n39114), .B(n39115), .Z(n30184) );
  AND U42007 ( .A(\modmult_1/xin[1023] ), .B(n39116), .Z(n39115) );
  IV U42008 ( .A(n39114), .Z(n39116) );
  XOR U42009 ( .A(n39117), .B(mreg[93]), .Z(n39114) );
  NAND U42010 ( .A(n39118), .B(mul_pow), .Z(n39117) );
  XOR U42011 ( .A(mreg[93]), .B(creg[93]), .Z(n39118) );
  XOR U42012 ( .A(n39119), .B(n39120), .Z(n39110) );
  ANDN U42013 ( .A(n39121), .B(n30191), .Z(n39120) );
  XOR U42014 ( .A(n39122), .B(\modmult_1/zin[0][91] ), .Z(n30191) );
  IV U42015 ( .A(n39119), .Z(n39122) );
  XNOR U42016 ( .A(n39119), .B(n30190), .Z(n39121) );
  XOR U42017 ( .A(n39123), .B(n39124), .Z(n30190) );
  AND U42018 ( .A(\modmult_1/xin[1023] ), .B(n39125), .Z(n39124) );
  IV U42019 ( .A(n39123), .Z(n39125) );
  XOR U42020 ( .A(n39126), .B(mreg[92]), .Z(n39123) );
  NAND U42021 ( .A(n39127), .B(mul_pow), .Z(n39126) );
  XOR U42022 ( .A(mreg[92]), .B(creg[92]), .Z(n39127) );
  XOR U42023 ( .A(n39128), .B(n39129), .Z(n39119) );
  ANDN U42024 ( .A(n39130), .B(n30197), .Z(n39129) );
  XOR U42025 ( .A(n39131), .B(\modmult_1/zin[0][90] ), .Z(n30197) );
  IV U42026 ( .A(n39128), .Z(n39131) );
  XNOR U42027 ( .A(n39128), .B(n30196), .Z(n39130) );
  XOR U42028 ( .A(n39132), .B(n39133), .Z(n30196) );
  AND U42029 ( .A(\modmult_1/xin[1023] ), .B(n39134), .Z(n39133) );
  IV U42030 ( .A(n39132), .Z(n39134) );
  XOR U42031 ( .A(n39135), .B(mreg[91]), .Z(n39132) );
  NAND U42032 ( .A(n39136), .B(mul_pow), .Z(n39135) );
  XOR U42033 ( .A(mreg[91]), .B(creg[91]), .Z(n39136) );
  XOR U42034 ( .A(n39137), .B(n39138), .Z(n39128) );
  ANDN U42035 ( .A(n39139), .B(n30203), .Z(n39138) );
  XOR U42036 ( .A(n39140), .B(\modmult_1/zin[0][89] ), .Z(n30203) );
  IV U42037 ( .A(n39137), .Z(n39140) );
  XNOR U42038 ( .A(n39137), .B(n30202), .Z(n39139) );
  XOR U42039 ( .A(n39141), .B(n39142), .Z(n30202) );
  AND U42040 ( .A(\modmult_1/xin[1023] ), .B(n39143), .Z(n39142) );
  IV U42041 ( .A(n39141), .Z(n39143) );
  XOR U42042 ( .A(n39144), .B(mreg[90]), .Z(n39141) );
  NAND U42043 ( .A(n39145), .B(mul_pow), .Z(n39144) );
  XOR U42044 ( .A(mreg[90]), .B(creg[90]), .Z(n39145) );
  XOR U42045 ( .A(n39146), .B(n39147), .Z(n39137) );
  ANDN U42046 ( .A(n39148), .B(n30209), .Z(n39147) );
  XOR U42047 ( .A(n39149), .B(\modmult_1/zin[0][88] ), .Z(n30209) );
  IV U42048 ( .A(n39146), .Z(n39149) );
  XNOR U42049 ( .A(n39146), .B(n30208), .Z(n39148) );
  XOR U42050 ( .A(n39150), .B(n39151), .Z(n30208) );
  AND U42051 ( .A(\modmult_1/xin[1023] ), .B(n39152), .Z(n39151) );
  IV U42052 ( .A(n39150), .Z(n39152) );
  XOR U42053 ( .A(n39153), .B(mreg[89]), .Z(n39150) );
  NAND U42054 ( .A(n39154), .B(mul_pow), .Z(n39153) );
  XOR U42055 ( .A(mreg[89]), .B(creg[89]), .Z(n39154) );
  XOR U42056 ( .A(n39155), .B(n39156), .Z(n39146) );
  ANDN U42057 ( .A(n39157), .B(n30215), .Z(n39156) );
  XOR U42058 ( .A(n39158), .B(\modmult_1/zin[0][87] ), .Z(n30215) );
  IV U42059 ( .A(n39155), .Z(n39158) );
  XNOR U42060 ( .A(n39155), .B(n30214), .Z(n39157) );
  XOR U42061 ( .A(n39159), .B(n39160), .Z(n30214) );
  AND U42062 ( .A(\modmult_1/xin[1023] ), .B(n39161), .Z(n39160) );
  IV U42063 ( .A(n39159), .Z(n39161) );
  XOR U42064 ( .A(n39162), .B(mreg[88]), .Z(n39159) );
  NAND U42065 ( .A(n39163), .B(mul_pow), .Z(n39162) );
  XOR U42066 ( .A(mreg[88]), .B(creg[88]), .Z(n39163) );
  XOR U42067 ( .A(n39164), .B(n39165), .Z(n39155) );
  ANDN U42068 ( .A(n39166), .B(n30221), .Z(n39165) );
  XOR U42069 ( .A(n39167), .B(\modmult_1/zin[0][86] ), .Z(n30221) );
  IV U42070 ( .A(n39164), .Z(n39167) );
  XNOR U42071 ( .A(n39164), .B(n30220), .Z(n39166) );
  XOR U42072 ( .A(n39168), .B(n39169), .Z(n30220) );
  AND U42073 ( .A(\modmult_1/xin[1023] ), .B(n39170), .Z(n39169) );
  IV U42074 ( .A(n39168), .Z(n39170) );
  XOR U42075 ( .A(n39171), .B(mreg[87]), .Z(n39168) );
  NAND U42076 ( .A(n39172), .B(mul_pow), .Z(n39171) );
  XOR U42077 ( .A(mreg[87]), .B(creg[87]), .Z(n39172) );
  XOR U42078 ( .A(n39173), .B(n39174), .Z(n39164) );
  ANDN U42079 ( .A(n39175), .B(n30227), .Z(n39174) );
  XOR U42080 ( .A(n39176), .B(\modmult_1/zin[0][85] ), .Z(n30227) );
  IV U42081 ( .A(n39173), .Z(n39176) );
  XNOR U42082 ( .A(n39173), .B(n30226), .Z(n39175) );
  XOR U42083 ( .A(n39177), .B(n39178), .Z(n30226) );
  AND U42084 ( .A(\modmult_1/xin[1023] ), .B(n39179), .Z(n39178) );
  IV U42085 ( .A(n39177), .Z(n39179) );
  XOR U42086 ( .A(n39180), .B(mreg[86]), .Z(n39177) );
  NAND U42087 ( .A(n39181), .B(mul_pow), .Z(n39180) );
  XOR U42088 ( .A(mreg[86]), .B(creg[86]), .Z(n39181) );
  XOR U42089 ( .A(n39182), .B(n39183), .Z(n39173) );
  ANDN U42090 ( .A(n39184), .B(n30233), .Z(n39183) );
  XOR U42091 ( .A(n39185), .B(\modmult_1/zin[0][84] ), .Z(n30233) );
  IV U42092 ( .A(n39182), .Z(n39185) );
  XNOR U42093 ( .A(n39182), .B(n30232), .Z(n39184) );
  XOR U42094 ( .A(n39186), .B(n39187), .Z(n30232) );
  AND U42095 ( .A(\modmult_1/xin[1023] ), .B(n39188), .Z(n39187) );
  IV U42096 ( .A(n39186), .Z(n39188) );
  XOR U42097 ( .A(n39189), .B(mreg[85]), .Z(n39186) );
  NAND U42098 ( .A(n39190), .B(mul_pow), .Z(n39189) );
  XOR U42099 ( .A(mreg[85]), .B(creg[85]), .Z(n39190) );
  XOR U42100 ( .A(n39191), .B(n39192), .Z(n39182) );
  ANDN U42101 ( .A(n39193), .B(n30239), .Z(n39192) );
  XOR U42102 ( .A(n39194), .B(\modmult_1/zin[0][83] ), .Z(n30239) );
  IV U42103 ( .A(n39191), .Z(n39194) );
  XNOR U42104 ( .A(n39191), .B(n30238), .Z(n39193) );
  XOR U42105 ( .A(n39195), .B(n39196), .Z(n30238) );
  AND U42106 ( .A(\modmult_1/xin[1023] ), .B(n39197), .Z(n39196) );
  IV U42107 ( .A(n39195), .Z(n39197) );
  XOR U42108 ( .A(n39198), .B(mreg[84]), .Z(n39195) );
  NAND U42109 ( .A(n39199), .B(mul_pow), .Z(n39198) );
  XOR U42110 ( .A(mreg[84]), .B(creg[84]), .Z(n39199) );
  XOR U42111 ( .A(n39200), .B(n39201), .Z(n39191) );
  ANDN U42112 ( .A(n39202), .B(n30245), .Z(n39201) );
  XOR U42113 ( .A(n39203), .B(\modmult_1/zin[0][82] ), .Z(n30245) );
  IV U42114 ( .A(n39200), .Z(n39203) );
  XNOR U42115 ( .A(n39200), .B(n30244), .Z(n39202) );
  XOR U42116 ( .A(n39204), .B(n39205), .Z(n30244) );
  AND U42117 ( .A(\modmult_1/xin[1023] ), .B(n39206), .Z(n39205) );
  IV U42118 ( .A(n39204), .Z(n39206) );
  XOR U42119 ( .A(n39207), .B(mreg[83]), .Z(n39204) );
  NAND U42120 ( .A(n39208), .B(mul_pow), .Z(n39207) );
  XOR U42121 ( .A(mreg[83]), .B(creg[83]), .Z(n39208) );
  XOR U42122 ( .A(n39209), .B(n39210), .Z(n39200) );
  ANDN U42123 ( .A(n39211), .B(n30251), .Z(n39210) );
  XOR U42124 ( .A(n39212), .B(\modmult_1/zin[0][81] ), .Z(n30251) );
  IV U42125 ( .A(n39209), .Z(n39212) );
  XNOR U42126 ( .A(n39209), .B(n30250), .Z(n39211) );
  XOR U42127 ( .A(n39213), .B(n39214), .Z(n30250) );
  AND U42128 ( .A(\modmult_1/xin[1023] ), .B(n39215), .Z(n39214) );
  IV U42129 ( .A(n39213), .Z(n39215) );
  XOR U42130 ( .A(n39216), .B(mreg[82]), .Z(n39213) );
  NAND U42131 ( .A(n39217), .B(mul_pow), .Z(n39216) );
  XOR U42132 ( .A(mreg[82]), .B(creg[82]), .Z(n39217) );
  XOR U42133 ( .A(n39218), .B(n39219), .Z(n39209) );
  ANDN U42134 ( .A(n39220), .B(n30257), .Z(n39219) );
  XOR U42135 ( .A(n39221), .B(\modmult_1/zin[0][80] ), .Z(n30257) );
  IV U42136 ( .A(n39218), .Z(n39221) );
  XNOR U42137 ( .A(n39218), .B(n30256), .Z(n39220) );
  XOR U42138 ( .A(n39222), .B(n39223), .Z(n30256) );
  AND U42139 ( .A(\modmult_1/xin[1023] ), .B(n39224), .Z(n39223) );
  IV U42140 ( .A(n39222), .Z(n39224) );
  XOR U42141 ( .A(n39225), .B(mreg[81]), .Z(n39222) );
  NAND U42142 ( .A(n39226), .B(mul_pow), .Z(n39225) );
  XOR U42143 ( .A(mreg[81]), .B(creg[81]), .Z(n39226) );
  XOR U42144 ( .A(n39227), .B(n39228), .Z(n39218) );
  ANDN U42145 ( .A(n39229), .B(n30263), .Z(n39228) );
  XOR U42146 ( .A(n39230), .B(\modmult_1/zin[0][79] ), .Z(n30263) );
  IV U42147 ( .A(n39227), .Z(n39230) );
  XNOR U42148 ( .A(n39227), .B(n30262), .Z(n39229) );
  XOR U42149 ( .A(n39231), .B(n39232), .Z(n30262) );
  AND U42150 ( .A(\modmult_1/xin[1023] ), .B(n39233), .Z(n39232) );
  IV U42151 ( .A(n39231), .Z(n39233) );
  XOR U42152 ( .A(n39234), .B(mreg[80]), .Z(n39231) );
  NAND U42153 ( .A(n39235), .B(mul_pow), .Z(n39234) );
  XOR U42154 ( .A(mreg[80]), .B(creg[80]), .Z(n39235) );
  XOR U42155 ( .A(n39236), .B(n39237), .Z(n39227) );
  ANDN U42156 ( .A(n39238), .B(n30269), .Z(n39237) );
  XOR U42157 ( .A(n39239), .B(\modmult_1/zin[0][78] ), .Z(n30269) );
  IV U42158 ( .A(n39236), .Z(n39239) );
  XNOR U42159 ( .A(n39236), .B(n30268), .Z(n39238) );
  XOR U42160 ( .A(n39240), .B(n39241), .Z(n30268) );
  AND U42161 ( .A(\modmult_1/xin[1023] ), .B(n39242), .Z(n39241) );
  IV U42162 ( .A(n39240), .Z(n39242) );
  XOR U42163 ( .A(n39243), .B(mreg[79]), .Z(n39240) );
  NAND U42164 ( .A(n39244), .B(mul_pow), .Z(n39243) );
  XOR U42165 ( .A(mreg[79]), .B(creg[79]), .Z(n39244) );
  XOR U42166 ( .A(n39245), .B(n39246), .Z(n39236) );
  ANDN U42167 ( .A(n39247), .B(n30275), .Z(n39246) );
  XOR U42168 ( .A(n39248), .B(\modmult_1/zin[0][77] ), .Z(n30275) );
  IV U42169 ( .A(n39245), .Z(n39248) );
  XNOR U42170 ( .A(n39245), .B(n30274), .Z(n39247) );
  XOR U42171 ( .A(n39249), .B(n39250), .Z(n30274) );
  AND U42172 ( .A(\modmult_1/xin[1023] ), .B(n39251), .Z(n39250) );
  IV U42173 ( .A(n39249), .Z(n39251) );
  XOR U42174 ( .A(n39252), .B(mreg[78]), .Z(n39249) );
  NAND U42175 ( .A(n39253), .B(mul_pow), .Z(n39252) );
  XOR U42176 ( .A(mreg[78]), .B(creg[78]), .Z(n39253) );
  XOR U42177 ( .A(n39254), .B(n39255), .Z(n39245) );
  ANDN U42178 ( .A(n39256), .B(n30281), .Z(n39255) );
  XOR U42179 ( .A(n39257), .B(\modmult_1/zin[0][76] ), .Z(n30281) );
  IV U42180 ( .A(n39254), .Z(n39257) );
  XNOR U42181 ( .A(n39254), .B(n30280), .Z(n39256) );
  XOR U42182 ( .A(n39258), .B(n39259), .Z(n30280) );
  AND U42183 ( .A(\modmult_1/xin[1023] ), .B(n39260), .Z(n39259) );
  IV U42184 ( .A(n39258), .Z(n39260) );
  XOR U42185 ( .A(n39261), .B(mreg[77]), .Z(n39258) );
  NAND U42186 ( .A(n39262), .B(mul_pow), .Z(n39261) );
  XOR U42187 ( .A(mreg[77]), .B(creg[77]), .Z(n39262) );
  XOR U42188 ( .A(n39263), .B(n39264), .Z(n39254) );
  ANDN U42189 ( .A(n39265), .B(n30287), .Z(n39264) );
  XOR U42190 ( .A(n39266), .B(\modmult_1/zin[0][75] ), .Z(n30287) );
  IV U42191 ( .A(n39263), .Z(n39266) );
  XNOR U42192 ( .A(n39263), .B(n30286), .Z(n39265) );
  XOR U42193 ( .A(n39267), .B(n39268), .Z(n30286) );
  AND U42194 ( .A(\modmult_1/xin[1023] ), .B(n39269), .Z(n39268) );
  IV U42195 ( .A(n39267), .Z(n39269) );
  XOR U42196 ( .A(n39270), .B(mreg[76]), .Z(n39267) );
  NAND U42197 ( .A(n39271), .B(mul_pow), .Z(n39270) );
  XOR U42198 ( .A(mreg[76]), .B(creg[76]), .Z(n39271) );
  XOR U42199 ( .A(n39272), .B(n39273), .Z(n39263) );
  ANDN U42200 ( .A(n39274), .B(n30293), .Z(n39273) );
  XOR U42201 ( .A(n39275), .B(\modmult_1/zin[0][74] ), .Z(n30293) );
  IV U42202 ( .A(n39272), .Z(n39275) );
  XNOR U42203 ( .A(n39272), .B(n30292), .Z(n39274) );
  XOR U42204 ( .A(n39276), .B(n39277), .Z(n30292) );
  AND U42205 ( .A(\modmult_1/xin[1023] ), .B(n39278), .Z(n39277) );
  IV U42206 ( .A(n39276), .Z(n39278) );
  XOR U42207 ( .A(n39279), .B(mreg[75]), .Z(n39276) );
  NAND U42208 ( .A(n39280), .B(mul_pow), .Z(n39279) );
  XOR U42209 ( .A(mreg[75]), .B(creg[75]), .Z(n39280) );
  XOR U42210 ( .A(n39281), .B(n39282), .Z(n39272) );
  ANDN U42211 ( .A(n39283), .B(n30299), .Z(n39282) );
  XOR U42212 ( .A(n39284), .B(\modmult_1/zin[0][73] ), .Z(n30299) );
  IV U42213 ( .A(n39281), .Z(n39284) );
  XNOR U42214 ( .A(n39281), .B(n30298), .Z(n39283) );
  XOR U42215 ( .A(n39285), .B(n39286), .Z(n30298) );
  AND U42216 ( .A(\modmult_1/xin[1023] ), .B(n39287), .Z(n39286) );
  IV U42217 ( .A(n39285), .Z(n39287) );
  XOR U42218 ( .A(n39288), .B(mreg[74]), .Z(n39285) );
  NAND U42219 ( .A(n39289), .B(mul_pow), .Z(n39288) );
  XOR U42220 ( .A(mreg[74]), .B(creg[74]), .Z(n39289) );
  XOR U42221 ( .A(n39290), .B(n39291), .Z(n39281) );
  ANDN U42222 ( .A(n39292), .B(n30305), .Z(n39291) );
  XOR U42223 ( .A(n39293), .B(\modmult_1/zin[0][72] ), .Z(n30305) );
  IV U42224 ( .A(n39290), .Z(n39293) );
  XNOR U42225 ( .A(n39290), .B(n30304), .Z(n39292) );
  XOR U42226 ( .A(n39294), .B(n39295), .Z(n30304) );
  AND U42227 ( .A(\modmult_1/xin[1023] ), .B(n39296), .Z(n39295) );
  IV U42228 ( .A(n39294), .Z(n39296) );
  XOR U42229 ( .A(n39297), .B(mreg[73]), .Z(n39294) );
  NAND U42230 ( .A(n39298), .B(mul_pow), .Z(n39297) );
  XOR U42231 ( .A(mreg[73]), .B(creg[73]), .Z(n39298) );
  XOR U42232 ( .A(n39299), .B(n39300), .Z(n39290) );
  ANDN U42233 ( .A(n39301), .B(n30311), .Z(n39300) );
  XOR U42234 ( .A(n39302), .B(\modmult_1/zin[0][71] ), .Z(n30311) );
  IV U42235 ( .A(n39299), .Z(n39302) );
  XNOR U42236 ( .A(n39299), .B(n30310), .Z(n39301) );
  XOR U42237 ( .A(n39303), .B(n39304), .Z(n30310) );
  AND U42238 ( .A(\modmult_1/xin[1023] ), .B(n39305), .Z(n39304) );
  IV U42239 ( .A(n39303), .Z(n39305) );
  XOR U42240 ( .A(n39306), .B(mreg[72]), .Z(n39303) );
  NAND U42241 ( .A(n39307), .B(mul_pow), .Z(n39306) );
  XOR U42242 ( .A(mreg[72]), .B(creg[72]), .Z(n39307) );
  XOR U42243 ( .A(n39308), .B(n39309), .Z(n39299) );
  ANDN U42244 ( .A(n39310), .B(n30317), .Z(n39309) );
  XOR U42245 ( .A(n39311), .B(\modmult_1/zin[0][70] ), .Z(n30317) );
  IV U42246 ( .A(n39308), .Z(n39311) );
  XNOR U42247 ( .A(n39308), .B(n30316), .Z(n39310) );
  XOR U42248 ( .A(n39312), .B(n39313), .Z(n30316) );
  AND U42249 ( .A(\modmult_1/xin[1023] ), .B(n39314), .Z(n39313) );
  IV U42250 ( .A(n39312), .Z(n39314) );
  XOR U42251 ( .A(n39315), .B(mreg[71]), .Z(n39312) );
  NAND U42252 ( .A(n39316), .B(mul_pow), .Z(n39315) );
  XOR U42253 ( .A(mreg[71]), .B(creg[71]), .Z(n39316) );
  XOR U42254 ( .A(n39317), .B(n39318), .Z(n39308) );
  ANDN U42255 ( .A(n39319), .B(n30323), .Z(n39318) );
  XOR U42256 ( .A(n39320), .B(\modmult_1/zin[0][69] ), .Z(n30323) );
  IV U42257 ( .A(n39317), .Z(n39320) );
  XNOR U42258 ( .A(n39317), .B(n30322), .Z(n39319) );
  XOR U42259 ( .A(n39321), .B(n39322), .Z(n30322) );
  AND U42260 ( .A(\modmult_1/xin[1023] ), .B(n39323), .Z(n39322) );
  IV U42261 ( .A(n39321), .Z(n39323) );
  XOR U42262 ( .A(n39324), .B(mreg[70]), .Z(n39321) );
  NAND U42263 ( .A(n39325), .B(mul_pow), .Z(n39324) );
  XOR U42264 ( .A(mreg[70]), .B(creg[70]), .Z(n39325) );
  XOR U42265 ( .A(n39326), .B(n39327), .Z(n39317) );
  ANDN U42266 ( .A(n39328), .B(n30329), .Z(n39327) );
  XOR U42267 ( .A(n39329), .B(\modmult_1/zin[0][68] ), .Z(n30329) );
  IV U42268 ( .A(n39326), .Z(n39329) );
  XNOR U42269 ( .A(n39326), .B(n30328), .Z(n39328) );
  XOR U42270 ( .A(n39330), .B(n39331), .Z(n30328) );
  AND U42271 ( .A(\modmult_1/xin[1023] ), .B(n39332), .Z(n39331) );
  IV U42272 ( .A(n39330), .Z(n39332) );
  XOR U42273 ( .A(n39333), .B(mreg[69]), .Z(n39330) );
  NAND U42274 ( .A(n39334), .B(mul_pow), .Z(n39333) );
  XOR U42275 ( .A(mreg[69]), .B(creg[69]), .Z(n39334) );
  XOR U42276 ( .A(n39335), .B(n39336), .Z(n39326) );
  ANDN U42277 ( .A(n39337), .B(n30335), .Z(n39336) );
  XOR U42278 ( .A(n39338), .B(\modmult_1/zin[0][67] ), .Z(n30335) );
  IV U42279 ( .A(n39335), .Z(n39338) );
  XNOR U42280 ( .A(n39335), .B(n30334), .Z(n39337) );
  XOR U42281 ( .A(n39339), .B(n39340), .Z(n30334) );
  AND U42282 ( .A(\modmult_1/xin[1023] ), .B(n39341), .Z(n39340) );
  IV U42283 ( .A(n39339), .Z(n39341) );
  XOR U42284 ( .A(n39342), .B(mreg[68]), .Z(n39339) );
  NAND U42285 ( .A(n39343), .B(mul_pow), .Z(n39342) );
  XOR U42286 ( .A(mreg[68]), .B(creg[68]), .Z(n39343) );
  XOR U42287 ( .A(n39344), .B(n39345), .Z(n39335) );
  ANDN U42288 ( .A(n39346), .B(n30341), .Z(n39345) );
  XOR U42289 ( .A(n39347), .B(\modmult_1/zin[0][66] ), .Z(n30341) );
  IV U42290 ( .A(n39344), .Z(n39347) );
  XNOR U42291 ( .A(n39344), .B(n30340), .Z(n39346) );
  XOR U42292 ( .A(n39348), .B(n39349), .Z(n30340) );
  AND U42293 ( .A(\modmult_1/xin[1023] ), .B(n39350), .Z(n39349) );
  IV U42294 ( .A(n39348), .Z(n39350) );
  XOR U42295 ( .A(n39351), .B(mreg[67]), .Z(n39348) );
  NAND U42296 ( .A(n39352), .B(mul_pow), .Z(n39351) );
  XOR U42297 ( .A(mreg[67]), .B(creg[67]), .Z(n39352) );
  XOR U42298 ( .A(n39353), .B(n39354), .Z(n39344) );
  ANDN U42299 ( .A(n39355), .B(n30347), .Z(n39354) );
  XOR U42300 ( .A(n39356), .B(\modmult_1/zin[0][65] ), .Z(n30347) );
  IV U42301 ( .A(n39353), .Z(n39356) );
  XNOR U42302 ( .A(n39353), .B(n30346), .Z(n39355) );
  XOR U42303 ( .A(n39357), .B(n39358), .Z(n30346) );
  AND U42304 ( .A(\modmult_1/xin[1023] ), .B(n39359), .Z(n39358) );
  IV U42305 ( .A(n39357), .Z(n39359) );
  XOR U42306 ( .A(n39360), .B(mreg[66]), .Z(n39357) );
  NAND U42307 ( .A(n39361), .B(mul_pow), .Z(n39360) );
  XOR U42308 ( .A(mreg[66]), .B(creg[66]), .Z(n39361) );
  XOR U42309 ( .A(n39362), .B(n39363), .Z(n39353) );
  ANDN U42310 ( .A(n39364), .B(n30353), .Z(n39363) );
  XOR U42311 ( .A(n39365), .B(\modmult_1/zin[0][64] ), .Z(n30353) );
  IV U42312 ( .A(n39362), .Z(n39365) );
  XNOR U42313 ( .A(n39362), .B(n30352), .Z(n39364) );
  XOR U42314 ( .A(n39366), .B(n39367), .Z(n30352) );
  AND U42315 ( .A(\modmult_1/xin[1023] ), .B(n39368), .Z(n39367) );
  IV U42316 ( .A(n39366), .Z(n39368) );
  XOR U42317 ( .A(n39369), .B(mreg[65]), .Z(n39366) );
  NAND U42318 ( .A(n39370), .B(mul_pow), .Z(n39369) );
  XOR U42319 ( .A(mreg[65]), .B(creg[65]), .Z(n39370) );
  XOR U42320 ( .A(n39371), .B(n39372), .Z(n39362) );
  ANDN U42321 ( .A(n39373), .B(n30359), .Z(n39372) );
  XOR U42322 ( .A(n39374), .B(\modmult_1/zin[0][63] ), .Z(n30359) );
  IV U42323 ( .A(n39371), .Z(n39374) );
  XNOR U42324 ( .A(n39371), .B(n30358), .Z(n39373) );
  XOR U42325 ( .A(n39375), .B(n39376), .Z(n30358) );
  AND U42326 ( .A(\modmult_1/xin[1023] ), .B(n39377), .Z(n39376) );
  IV U42327 ( .A(n39375), .Z(n39377) );
  XOR U42328 ( .A(n39378), .B(mreg[64]), .Z(n39375) );
  NAND U42329 ( .A(n39379), .B(mul_pow), .Z(n39378) );
  XOR U42330 ( .A(mreg[64]), .B(creg[64]), .Z(n39379) );
  XOR U42331 ( .A(n39380), .B(n39381), .Z(n39371) );
  ANDN U42332 ( .A(n39382), .B(n30365), .Z(n39381) );
  XOR U42333 ( .A(n39383), .B(\modmult_1/zin[0][62] ), .Z(n30365) );
  IV U42334 ( .A(n39380), .Z(n39383) );
  XNOR U42335 ( .A(n39380), .B(n30364), .Z(n39382) );
  XOR U42336 ( .A(n39384), .B(n39385), .Z(n30364) );
  AND U42337 ( .A(\modmult_1/xin[1023] ), .B(n39386), .Z(n39385) );
  IV U42338 ( .A(n39384), .Z(n39386) );
  XOR U42339 ( .A(n39387), .B(mreg[63]), .Z(n39384) );
  NAND U42340 ( .A(n39388), .B(mul_pow), .Z(n39387) );
  XOR U42341 ( .A(mreg[63]), .B(creg[63]), .Z(n39388) );
  XOR U42342 ( .A(n39389), .B(n39390), .Z(n39380) );
  ANDN U42343 ( .A(n39391), .B(n30371), .Z(n39390) );
  XOR U42344 ( .A(n39392), .B(\modmult_1/zin[0][61] ), .Z(n30371) );
  IV U42345 ( .A(n39389), .Z(n39392) );
  XNOR U42346 ( .A(n39389), .B(n30370), .Z(n39391) );
  XOR U42347 ( .A(n39393), .B(n39394), .Z(n30370) );
  AND U42348 ( .A(\modmult_1/xin[1023] ), .B(n39395), .Z(n39394) );
  IV U42349 ( .A(n39393), .Z(n39395) );
  XOR U42350 ( .A(n39396), .B(mreg[62]), .Z(n39393) );
  NAND U42351 ( .A(n39397), .B(mul_pow), .Z(n39396) );
  XOR U42352 ( .A(mreg[62]), .B(creg[62]), .Z(n39397) );
  XOR U42353 ( .A(n39398), .B(n39399), .Z(n39389) );
  ANDN U42354 ( .A(n39400), .B(n30377), .Z(n39399) );
  XOR U42355 ( .A(n39401), .B(\modmult_1/zin[0][60] ), .Z(n30377) );
  IV U42356 ( .A(n39398), .Z(n39401) );
  XNOR U42357 ( .A(n39398), .B(n30376), .Z(n39400) );
  XOR U42358 ( .A(n39402), .B(n39403), .Z(n30376) );
  AND U42359 ( .A(\modmult_1/xin[1023] ), .B(n39404), .Z(n39403) );
  IV U42360 ( .A(n39402), .Z(n39404) );
  XOR U42361 ( .A(n39405), .B(mreg[61]), .Z(n39402) );
  NAND U42362 ( .A(n39406), .B(mul_pow), .Z(n39405) );
  XOR U42363 ( .A(mreg[61]), .B(creg[61]), .Z(n39406) );
  XOR U42364 ( .A(n39407), .B(n39408), .Z(n39398) );
  ANDN U42365 ( .A(n39409), .B(n30383), .Z(n39408) );
  XOR U42366 ( .A(n39410), .B(\modmult_1/zin[0][59] ), .Z(n30383) );
  IV U42367 ( .A(n39407), .Z(n39410) );
  XNOR U42368 ( .A(n39407), .B(n30382), .Z(n39409) );
  XOR U42369 ( .A(n39411), .B(n39412), .Z(n30382) );
  AND U42370 ( .A(\modmult_1/xin[1023] ), .B(n39413), .Z(n39412) );
  IV U42371 ( .A(n39411), .Z(n39413) );
  XOR U42372 ( .A(n39414), .B(mreg[60]), .Z(n39411) );
  NAND U42373 ( .A(n39415), .B(mul_pow), .Z(n39414) );
  XOR U42374 ( .A(mreg[60]), .B(creg[60]), .Z(n39415) );
  XOR U42375 ( .A(n39416), .B(n39417), .Z(n39407) );
  ANDN U42376 ( .A(n39418), .B(n30389), .Z(n39417) );
  XOR U42377 ( .A(n39419), .B(\modmult_1/zin[0][58] ), .Z(n30389) );
  IV U42378 ( .A(n39416), .Z(n39419) );
  XNOR U42379 ( .A(n39416), .B(n30388), .Z(n39418) );
  XOR U42380 ( .A(n39420), .B(n39421), .Z(n30388) );
  AND U42381 ( .A(\modmult_1/xin[1023] ), .B(n39422), .Z(n39421) );
  IV U42382 ( .A(n39420), .Z(n39422) );
  XOR U42383 ( .A(n39423), .B(mreg[59]), .Z(n39420) );
  NAND U42384 ( .A(n39424), .B(mul_pow), .Z(n39423) );
  XOR U42385 ( .A(mreg[59]), .B(creg[59]), .Z(n39424) );
  XOR U42386 ( .A(n39425), .B(n39426), .Z(n39416) );
  ANDN U42387 ( .A(n39427), .B(n30395), .Z(n39426) );
  XOR U42388 ( .A(n39428), .B(\modmult_1/zin[0][57] ), .Z(n30395) );
  IV U42389 ( .A(n39425), .Z(n39428) );
  XNOR U42390 ( .A(n39425), .B(n30394), .Z(n39427) );
  XOR U42391 ( .A(n39429), .B(n39430), .Z(n30394) );
  AND U42392 ( .A(\modmult_1/xin[1023] ), .B(n39431), .Z(n39430) );
  IV U42393 ( .A(n39429), .Z(n39431) );
  XOR U42394 ( .A(n39432), .B(mreg[58]), .Z(n39429) );
  NAND U42395 ( .A(n39433), .B(mul_pow), .Z(n39432) );
  XOR U42396 ( .A(mreg[58]), .B(creg[58]), .Z(n39433) );
  XOR U42397 ( .A(n39434), .B(n39435), .Z(n39425) );
  ANDN U42398 ( .A(n39436), .B(n30401), .Z(n39435) );
  XOR U42399 ( .A(n39437), .B(\modmult_1/zin[0][56] ), .Z(n30401) );
  IV U42400 ( .A(n39434), .Z(n39437) );
  XNOR U42401 ( .A(n39434), .B(n30400), .Z(n39436) );
  XOR U42402 ( .A(n39438), .B(n39439), .Z(n30400) );
  AND U42403 ( .A(\modmult_1/xin[1023] ), .B(n39440), .Z(n39439) );
  IV U42404 ( .A(n39438), .Z(n39440) );
  XOR U42405 ( .A(n39441), .B(mreg[57]), .Z(n39438) );
  NAND U42406 ( .A(n39442), .B(mul_pow), .Z(n39441) );
  XOR U42407 ( .A(mreg[57]), .B(creg[57]), .Z(n39442) );
  XOR U42408 ( .A(n39443), .B(n39444), .Z(n39434) );
  ANDN U42409 ( .A(n39445), .B(n30407), .Z(n39444) );
  XOR U42410 ( .A(n39446), .B(\modmult_1/zin[0][55] ), .Z(n30407) );
  IV U42411 ( .A(n39443), .Z(n39446) );
  XNOR U42412 ( .A(n39443), .B(n30406), .Z(n39445) );
  XOR U42413 ( .A(n39447), .B(n39448), .Z(n30406) );
  AND U42414 ( .A(\modmult_1/xin[1023] ), .B(n39449), .Z(n39448) );
  IV U42415 ( .A(n39447), .Z(n39449) );
  XOR U42416 ( .A(n39450), .B(mreg[56]), .Z(n39447) );
  NAND U42417 ( .A(n39451), .B(mul_pow), .Z(n39450) );
  XOR U42418 ( .A(mreg[56]), .B(creg[56]), .Z(n39451) );
  XOR U42419 ( .A(n39452), .B(n39453), .Z(n39443) );
  ANDN U42420 ( .A(n39454), .B(n30413), .Z(n39453) );
  XOR U42421 ( .A(n39455), .B(\modmult_1/zin[0][54] ), .Z(n30413) );
  IV U42422 ( .A(n39452), .Z(n39455) );
  XNOR U42423 ( .A(n39452), .B(n30412), .Z(n39454) );
  XOR U42424 ( .A(n39456), .B(n39457), .Z(n30412) );
  AND U42425 ( .A(\modmult_1/xin[1023] ), .B(n39458), .Z(n39457) );
  IV U42426 ( .A(n39456), .Z(n39458) );
  XOR U42427 ( .A(n39459), .B(mreg[55]), .Z(n39456) );
  NAND U42428 ( .A(n39460), .B(mul_pow), .Z(n39459) );
  XOR U42429 ( .A(mreg[55]), .B(creg[55]), .Z(n39460) );
  XOR U42430 ( .A(n39461), .B(n39462), .Z(n39452) );
  ANDN U42431 ( .A(n39463), .B(n30419), .Z(n39462) );
  XOR U42432 ( .A(n39464), .B(\modmult_1/zin[0][53] ), .Z(n30419) );
  IV U42433 ( .A(n39461), .Z(n39464) );
  XNOR U42434 ( .A(n39461), .B(n30418), .Z(n39463) );
  XOR U42435 ( .A(n39465), .B(n39466), .Z(n30418) );
  AND U42436 ( .A(\modmult_1/xin[1023] ), .B(n39467), .Z(n39466) );
  IV U42437 ( .A(n39465), .Z(n39467) );
  XOR U42438 ( .A(n39468), .B(mreg[54]), .Z(n39465) );
  NAND U42439 ( .A(n39469), .B(mul_pow), .Z(n39468) );
  XOR U42440 ( .A(mreg[54]), .B(creg[54]), .Z(n39469) );
  XOR U42441 ( .A(n39470), .B(n39471), .Z(n39461) );
  ANDN U42442 ( .A(n39472), .B(n30425), .Z(n39471) );
  XOR U42443 ( .A(n39473), .B(\modmult_1/zin[0][52] ), .Z(n30425) );
  IV U42444 ( .A(n39470), .Z(n39473) );
  XNOR U42445 ( .A(n39470), .B(n30424), .Z(n39472) );
  XOR U42446 ( .A(n39474), .B(n39475), .Z(n30424) );
  AND U42447 ( .A(\modmult_1/xin[1023] ), .B(n39476), .Z(n39475) );
  IV U42448 ( .A(n39474), .Z(n39476) );
  XOR U42449 ( .A(n39477), .B(mreg[53]), .Z(n39474) );
  NAND U42450 ( .A(n39478), .B(mul_pow), .Z(n39477) );
  XOR U42451 ( .A(mreg[53]), .B(creg[53]), .Z(n39478) );
  XOR U42452 ( .A(n39479), .B(n39480), .Z(n39470) );
  ANDN U42453 ( .A(n39481), .B(n30431), .Z(n39480) );
  XOR U42454 ( .A(n39482), .B(\modmult_1/zin[0][51] ), .Z(n30431) );
  IV U42455 ( .A(n39479), .Z(n39482) );
  XNOR U42456 ( .A(n39479), .B(n30430), .Z(n39481) );
  XOR U42457 ( .A(n39483), .B(n39484), .Z(n30430) );
  AND U42458 ( .A(\modmult_1/xin[1023] ), .B(n39485), .Z(n39484) );
  IV U42459 ( .A(n39483), .Z(n39485) );
  XOR U42460 ( .A(n39486), .B(mreg[52]), .Z(n39483) );
  NAND U42461 ( .A(n39487), .B(mul_pow), .Z(n39486) );
  XOR U42462 ( .A(mreg[52]), .B(creg[52]), .Z(n39487) );
  XOR U42463 ( .A(n39488), .B(n39489), .Z(n39479) );
  ANDN U42464 ( .A(n39490), .B(n30437), .Z(n39489) );
  XOR U42465 ( .A(n39491), .B(\modmult_1/zin[0][50] ), .Z(n30437) );
  IV U42466 ( .A(n39488), .Z(n39491) );
  XNOR U42467 ( .A(n39488), .B(n30436), .Z(n39490) );
  XOR U42468 ( .A(n39492), .B(n39493), .Z(n30436) );
  AND U42469 ( .A(\modmult_1/xin[1023] ), .B(n39494), .Z(n39493) );
  IV U42470 ( .A(n39492), .Z(n39494) );
  XOR U42471 ( .A(n39495), .B(mreg[51]), .Z(n39492) );
  NAND U42472 ( .A(n39496), .B(mul_pow), .Z(n39495) );
  XOR U42473 ( .A(mreg[51]), .B(creg[51]), .Z(n39496) );
  XOR U42474 ( .A(n39497), .B(n39498), .Z(n39488) );
  ANDN U42475 ( .A(n39499), .B(n30443), .Z(n39498) );
  XOR U42476 ( .A(n39500), .B(\modmult_1/zin[0][49] ), .Z(n30443) );
  IV U42477 ( .A(n39497), .Z(n39500) );
  XNOR U42478 ( .A(n39497), .B(n30442), .Z(n39499) );
  XOR U42479 ( .A(n39501), .B(n39502), .Z(n30442) );
  AND U42480 ( .A(\modmult_1/xin[1023] ), .B(n39503), .Z(n39502) );
  IV U42481 ( .A(n39501), .Z(n39503) );
  XOR U42482 ( .A(n39504), .B(mreg[50]), .Z(n39501) );
  NAND U42483 ( .A(n39505), .B(mul_pow), .Z(n39504) );
  XOR U42484 ( .A(mreg[50]), .B(creg[50]), .Z(n39505) );
  XOR U42485 ( .A(n39506), .B(n39507), .Z(n39497) );
  ANDN U42486 ( .A(n39508), .B(n30449), .Z(n39507) );
  XOR U42487 ( .A(n39509), .B(\modmult_1/zin[0][48] ), .Z(n30449) );
  IV U42488 ( .A(n39506), .Z(n39509) );
  XNOR U42489 ( .A(n39506), .B(n30448), .Z(n39508) );
  XOR U42490 ( .A(n39510), .B(n39511), .Z(n30448) );
  AND U42491 ( .A(\modmult_1/xin[1023] ), .B(n39512), .Z(n39511) );
  IV U42492 ( .A(n39510), .Z(n39512) );
  XOR U42493 ( .A(n39513), .B(mreg[49]), .Z(n39510) );
  NAND U42494 ( .A(n39514), .B(mul_pow), .Z(n39513) );
  XOR U42495 ( .A(mreg[49]), .B(creg[49]), .Z(n39514) );
  XOR U42496 ( .A(n39515), .B(n39516), .Z(n39506) );
  ANDN U42497 ( .A(n39517), .B(n30455), .Z(n39516) );
  XOR U42498 ( .A(n39518), .B(\modmult_1/zin[0][47] ), .Z(n30455) );
  IV U42499 ( .A(n39515), .Z(n39518) );
  XNOR U42500 ( .A(n39515), .B(n30454), .Z(n39517) );
  XOR U42501 ( .A(n39519), .B(n39520), .Z(n30454) );
  AND U42502 ( .A(\modmult_1/xin[1023] ), .B(n39521), .Z(n39520) );
  IV U42503 ( .A(n39519), .Z(n39521) );
  XOR U42504 ( .A(n39522), .B(mreg[48]), .Z(n39519) );
  NAND U42505 ( .A(n39523), .B(mul_pow), .Z(n39522) );
  XOR U42506 ( .A(mreg[48]), .B(creg[48]), .Z(n39523) );
  XOR U42507 ( .A(n39524), .B(n39525), .Z(n39515) );
  ANDN U42508 ( .A(n39526), .B(n30461), .Z(n39525) );
  XOR U42509 ( .A(n39527), .B(\modmult_1/zin[0][46] ), .Z(n30461) );
  IV U42510 ( .A(n39524), .Z(n39527) );
  XNOR U42511 ( .A(n39524), .B(n30460), .Z(n39526) );
  XOR U42512 ( .A(n39528), .B(n39529), .Z(n30460) );
  AND U42513 ( .A(\modmult_1/xin[1023] ), .B(n39530), .Z(n39529) );
  IV U42514 ( .A(n39528), .Z(n39530) );
  XOR U42515 ( .A(n39531), .B(mreg[47]), .Z(n39528) );
  NAND U42516 ( .A(n39532), .B(mul_pow), .Z(n39531) );
  XOR U42517 ( .A(mreg[47]), .B(creg[47]), .Z(n39532) );
  XOR U42518 ( .A(n39533), .B(n39534), .Z(n39524) );
  ANDN U42519 ( .A(n39535), .B(n30467), .Z(n39534) );
  XOR U42520 ( .A(n39536), .B(\modmult_1/zin[0][45] ), .Z(n30467) );
  IV U42521 ( .A(n39533), .Z(n39536) );
  XNOR U42522 ( .A(n39533), .B(n30466), .Z(n39535) );
  XOR U42523 ( .A(n39537), .B(n39538), .Z(n30466) );
  AND U42524 ( .A(\modmult_1/xin[1023] ), .B(n39539), .Z(n39538) );
  IV U42525 ( .A(n39537), .Z(n39539) );
  XOR U42526 ( .A(n39540), .B(mreg[46]), .Z(n39537) );
  NAND U42527 ( .A(n39541), .B(mul_pow), .Z(n39540) );
  XOR U42528 ( .A(mreg[46]), .B(creg[46]), .Z(n39541) );
  XOR U42529 ( .A(n39542), .B(n39543), .Z(n39533) );
  ANDN U42530 ( .A(n39544), .B(n30473), .Z(n39543) );
  XOR U42531 ( .A(n39545), .B(\modmult_1/zin[0][44] ), .Z(n30473) );
  IV U42532 ( .A(n39542), .Z(n39545) );
  XNOR U42533 ( .A(n39542), .B(n30472), .Z(n39544) );
  XOR U42534 ( .A(n39546), .B(n39547), .Z(n30472) );
  AND U42535 ( .A(\modmult_1/xin[1023] ), .B(n39548), .Z(n39547) );
  IV U42536 ( .A(n39546), .Z(n39548) );
  XOR U42537 ( .A(n39549), .B(mreg[45]), .Z(n39546) );
  NAND U42538 ( .A(n39550), .B(mul_pow), .Z(n39549) );
  XOR U42539 ( .A(mreg[45]), .B(creg[45]), .Z(n39550) );
  XOR U42540 ( .A(n39551), .B(n39552), .Z(n39542) );
  ANDN U42541 ( .A(n39553), .B(n30479), .Z(n39552) );
  XOR U42542 ( .A(n39554), .B(\modmult_1/zin[0][43] ), .Z(n30479) );
  IV U42543 ( .A(n39551), .Z(n39554) );
  XNOR U42544 ( .A(n39551), .B(n30478), .Z(n39553) );
  XOR U42545 ( .A(n39555), .B(n39556), .Z(n30478) );
  AND U42546 ( .A(\modmult_1/xin[1023] ), .B(n39557), .Z(n39556) );
  IV U42547 ( .A(n39555), .Z(n39557) );
  XOR U42548 ( .A(n39558), .B(mreg[44]), .Z(n39555) );
  NAND U42549 ( .A(n39559), .B(mul_pow), .Z(n39558) );
  XOR U42550 ( .A(mreg[44]), .B(creg[44]), .Z(n39559) );
  XOR U42551 ( .A(n39560), .B(n39561), .Z(n39551) );
  ANDN U42552 ( .A(n39562), .B(n30485), .Z(n39561) );
  XOR U42553 ( .A(n39563), .B(\modmult_1/zin[0][42] ), .Z(n30485) );
  IV U42554 ( .A(n39560), .Z(n39563) );
  XNOR U42555 ( .A(n39560), .B(n30484), .Z(n39562) );
  XOR U42556 ( .A(n39564), .B(n39565), .Z(n30484) );
  AND U42557 ( .A(\modmult_1/xin[1023] ), .B(n39566), .Z(n39565) );
  IV U42558 ( .A(n39564), .Z(n39566) );
  XOR U42559 ( .A(n39567), .B(mreg[43]), .Z(n39564) );
  NAND U42560 ( .A(n39568), .B(mul_pow), .Z(n39567) );
  XOR U42561 ( .A(mreg[43]), .B(creg[43]), .Z(n39568) );
  XOR U42562 ( .A(n39569), .B(n39570), .Z(n39560) );
  ANDN U42563 ( .A(n39571), .B(n30491), .Z(n39570) );
  XOR U42564 ( .A(n39572), .B(\modmult_1/zin[0][41] ), .Z(n30491) );
  IV U42565 ( .A(n39569), .Z(n39572) );
  XNOR U42566 ( .A(n39569), .B(n30490), .Z(n39571) );
  XOR U42567 ( .A(n39573), .B(n39574), .Z(n30490) );
  AND U42568 ( .A(\modmult_1/xin[1023] ), .B(n39575), .Z(n39574) );
  IV U42569 ( .A(n39573), .Z(n39575) );
  XOR U42570 ( .A(n39576), .B(mreg[42]), .Z(n39573) );
  NAND U42571 ( .A(n39577), .B(mul_pow), .Z(n39576) );
  XOR U42572 ( .A(mreg[42]), .B(creg[42]), .Z(n39577) );
  XOR U42573 ( .A(n39578), .B(n39579), .Z(n39569) );
  ANDN U42574 ( .A(n39580), .B(n30497), .Z(n39579) );
  XOR U42575 ( .A(n39581), .B(\modmult_1/zin[0][40] ), .Z(n30497) );
  IV U42576 ( .A(n39578), .Z(n39581) );
  XNOR U42577 ( .A(n39578), .B(n30496), .Z(n39580) );
  XOR U42578 ( .A(n39582), .B(n39583), .Z(n30496) );
  AND U42579 ( .A(\modmult_1/xin[1023] ), .B(n39584), .Z(n39583) );
  IV U42580 ( .A(n39582), .Z(n39584) );
  XOR U42581 ( .A(n39585), .B(mreg[41]), .Z(n39582) );
  NAND U42582 ( .A(n39586), .B(mul_pow), .Z(n39585) );
  XOR U42583 ( .A(mreg[41]), .B(creg[41]), .Z(n39586) );
  XOR U42584 ( .A(n39587), .B(n39588), .Z(n39578) );
  ANDN U42585 ( .A(n39589), .B(n30503), .Z(n39588) );
  XOR U42586 ( .A(n39590), .B(\modmult_1/zin[0][39] ), .Z(n30503) );
  IV U42587 ( .A(n39587), .Z(n39590) );
  XNOR U42588 ( .A(n39587), .B(n30502), .Z(n39589) );
  XOR U42589 ( .A(n39591), .B(n39592), .Z(n30502) );
  AND U42590 ( .A(\modmult_1/xin[1023] ), .B(n39593), .Z(n39592) );
  IV U42591 ( .A(n39591), .Z(n39593) );
  XOR U42592 ( .A(n39594), .B(mreg[40]), .Z(n39591) );
  NAND U42593 ( .A(n39595), .B(mul_pow), .Z(n39594) );
  XOR U42594 ( .A(mreg[40]), .B(creg[40]), .Z(n39595) );
  XOR U42595 ( .A(n39596), .B(n39597), .Z(n39587) );
  ANDN U42596 ( .A(n39598), .B(n30509), .Z(n39597) );
  XOR U42597 ( .A(n39599), .B(\modmult_1/zin[0][38] ), .Z(n30509) );
  IV U42598 ( .A(n39596), .Z(n39599) );
  XNOR U42599 ( .A(n39596), .B(n30508), .Z(n39598) );
  XOR U42600 ( .A(n39600), .B(n39601), .Z(n30508) );
  AND U42601 ( .A(\modmult_1/xin[1023] ), .B(n39602), .Z(n39601) );
  IV U42602 ( .A(n39600), .Z(n39602) );
  XOR U42603 ( .A(n39603), .B(mreg[39]), .Z(n39600) );
  NAND U42604 ( .A(n39604), .B(mul_pow), .Z(n39603) );
  XOR U42605 ( .A(mreg[39]), .B(creg[39]), .Z(n39604) );
  XOR U42606 ( .A(n39605), .B(n39606), .Z(n39596) );
  ANDN U42607 ( .A(n39607), .B(n30515), .Z(n39606) );
  XOR U42608 ( .A(n39608), .B(\modmult_1/zin[0][37] ), .Z(n30515) );
  IV U42609 ( .A(n39605), .Z(n39608) );
  XNOR U42610 ( .A(n39605), .B(n30514), .Z(n39607) );
  XOR U42611 ( .A(n39609), .B(n39610), .Z(n30514) );
  AND U42612 ( .A(\modmult_1/xin[1023] ), .B(n39611), .Z(n39610) );
  IV U42613 ( .A(n39609), .Z(n39611) );
  XOR U42614 ( .A(n39612), .B(mreg[38]), .Z(n39609) );
  NAND U42615 ( .A(n39613), .B(mul_pow), .Z(n39612) );
  XOR U42616 ( .A(mreg[38]), .B(creg[38]), .Z(n39613) );
  XOR U42617 ( .A(n39614), .B(n39615), .Z(n39605) );
  ANDN U42618 ( .A(n39616), .B(n30521), .Z(n39615) );
  XOR U42619 ( .A(n39617), .B(\modmult_1/zin[0][36] ), .Z(n30521) );
  IV U42620 ( .A(n39614), .Z(n39617) );
  XNOR U42621 ( .A(n39614), .B(n30520), .Z(n39616) );
  XOR U42622 ( .A(n39618), .B(n39619), .Z(n30520) );
  AND U42623 ( .A(\modmult_1/xin[1023] ), .B(n39620), .Z(n39619) );
  IV U42624 ( .A(n39618), .Z(n39620) );
  XOR U42625 ( .A(n39621), .B(mreg[37]), .Z(n39618) );
  NAND U42626 ( .A(n39622), .B(mul_pow), .Z(n39621) );
  XOR U42627 ( .A(mreg[37]), .B(creg[37]), .Z(n39622) );
  XOR U42628 ( .A(n39623), .B(n39624), .Z(n39614) );
  ANDN U42629 ( .A(n39625), .B(n30527), .Z(n39624) );
  XOR U42630 ( .A(n39626), .B(\modmult_1/zin[0][35] ), .Z(n30527) );
  IV U42631 ( .A(n39623), .Z(n39626) );
  XNOR U42632 ( .A(n39623), .B(n30526), .Z(n39625) );
  XOR U42633 ( .A(n39627), .B(n39628), .Z(n30526) );
  AND U42634 ( .A(\modmult_1/xin[1023] ), .B(n39629), .Z(n39628) );
  IV U42635 ( .A(n39627), .Z(n39629) );
  XOR U42636 ( .A(n39630), .B(mreg[36]), .Z(n39627) );
  NAND U42637 ( .A(n39631), .B(mul_pow), .Z(n39630) );
  XOR U42638 ( .A(mreg[36]), .B(creg[36]), .Z(n39631) );
  XOR U42639 ( .A(n39632), .B(n39633), .Z(n39623) );
  ANDN U42640 ( .A(n39634), .B(n30533), .Z(n39633) );
  XOR U42641 ( .A(n39635), .B(\modmult_1/zin[0][34] ), .Z(n30533) );
  IV U42642 ( .A(n39632), .Z(n39635) );
  XNOR U42643 ( .A(n39632), .B(n30532), .Z(n39634) );
  XOR U42644 ( .A(n39636), .B(n39637), .Z(n30532) );
  AND U42645 ( .A(\modmult_1/xin[1023] ), .B(n39638), .Z(n39637) );
  IV U42646 ( .A(n39636), .Z(n39638) );
  XOR U42647 ( .A(n39639), .B(mreg[35]), .Z(n39636) );
  NAND U42648 ( .A(n39640), .B(mul_pow), .Z(n39639) );
  XOR U42649 ( .A(mreg[35]), .B(creg[35]), .Z(n39640) );
  XOR U42650 ( .A(n39641), .B(n39642), .Z(n39632) );
  ANDN U42651 ( .A(n39643), .B(n30539), .Z(n39642) );
  XOR U42652 ( .A(n39644), .B(\modmult_1/zin[0][33] ), .Z(n30539) );
  IV U42653 ( .A(n39641), .Z(n39644) );
  XNOR U42654 ( .A(n39641), .B(n30538), .Z(n39643) );
  XOR U42655 ( .A(n39645), .B(n39646), .Z(n30538) );
  AND U42656 ( .A(\modmult_1/xin[1023] ), .B(n39647), .Z(n39646) );
  IV U42657 ( .A(n39645), .Z(n39647) );
  XOR U42658 ( .A(n39648), .B(mreg[34]), .Z(n39645) );
  NAND U42659 ( .A(n39649), .B(mul_pow), .Z(n39648) );
  XOR U42660 ( .A(mreg[34]), .B(creg[34]), .Z(n39649) );
  XOR U42661 ( .A(n39650), .B(n39651), .Z(n39641) );
  ANDN U42662 ( .A(n39652), .B(n30545), .Z(n39651) );
  XOR U42663 ( .A(n39653), .B(\modmult_1/zin[0][32] ), .Z(n30545) );
  IV U42664 ( .A(n39650), .Z(n39653) );
  XNOR U42665 ( .A(n39650), .B(n30544), .Z(n39652) );
  XOR U42666 ( .A(n39654), .B(n39655), .Z(n30544) );
  AND U42667 ( .A(\modmult_1/xin[1023] ), .B(n39656), .Z(n39655) );
  IV U42668 ( .A(n39654), .Z(n39656) );
  XOR U42669 ( .A(n39657), .B(mreg[33]), .Z(n39654) );
  NAND U42670 ( .A(n39658), .B(mul_pow), .Z(n39657) );
  XOR U42671 ( .A(mreg[33]), .B(creg[33]), .Z(n39658) );
  XOR U42672 ( .A(n39659), .B(n39660), .Z(n39650) );
  ANDN U42673 ( .A(n39661), .B(n30551), .Z(n39660) );
  XOR U42674 ( .A(n39662), .B(\modmult_1/zin[0][31] ), .Z(n30551) );
  IV U42675 ( .A(n39659), .Z(n39662) );
  XNOR U42676 ( .A(n39659), .B(n30550), .Z(n39661) );
  XOR U42677 ( .A(n39663), .B(n39664), .Z(n30550) );
  AND U42678 ( .A(\modmult_1/xin[1023] ), .B(n39665), .Z(n39664) );
  IV U42679 ( .A(n39663), .Z(n39665) );
  XOR U42680 ( .A(n39666), .B(mreg[32]), .Z(n39663) );
  NAND U42681 ( .A(n39667), .B(mul_pow), .Z(n39666) );
  XOR U42682 ( .A(mreg[32]), .B(creg[32]), .Z(n39667) );
  XOR U42683 ( .A(n39668), .B(n39669), .Z(n39659) );
  ANDN U42684 ( .A(n39670), .B(n30557), .Z(n39669) );
  XOR U42685 ( .A(n39671), .B(\modmult_1/zin[0][30] ), .Z(n30557) );
  IV U42686 ( .A(n39668), .Z(n39671) );
  XNOR U42687 ( .A(n39668), .B(n30556), .Z(n39670) );
  XOR U42688 ( .A(n39672), .B(n39673), .Z(n30556) );
  AND U42689 ( .A(\modmult_1/xin[1023] ), .B(n39674), .Z(n39673) );
  IV U42690 ( .A(n39672), .Z(n39674) );
  XOR U42691 ( .A(n39675), .B(mreg[31]), .Z(n39672) );
  NAND U42692 ( .A(n39676), .B(mul_pow), .Z(n39675) );
  XOR U42693 ( .A(mreg[31]), .B(creg[31]), .Z(n39676) );
  XOR U42694 ( .A(n39677), .B(n39678), .Z(n39668) );
  ANDN U42695 ( .A(n39679), .B(n30563), .Z(n39678) );
  XOR U42696 ( .A(n39680), .B(\modmult_1/zin[0][29] ), .Z(n30563) );
  IV U42697 ( .A(n39677), .Z(n39680) );
  XNOR U42698 ( .A(n39677), .B(n30562), .Z(n39679) );
  XOR U42699 ( .A(n39681), .B(n39682), .Z(n30562) );
  AND U42700 ( .A(\modmult_1/xin[1023] ), .B(n39683), .Z(n39682) );
  IV U42701 ( .A(n39681), .Z(n39683) );
  XOR U42702 ( .A(n39684), .B(mreg[30]), .Z(n39681) );
  NAND U42703 ( .A(n39685), .B(mul_pow), .Z(n39684) );
  XOR U42704 ( .A(mreg[30]), .B(creg[30]), .Z(n39685) );
  XOR U42705 ( .A(n39686), .B(n39687), .Z(n39677) );
  ANDN U42706 ( .A(n39688), .B(n30569), .Z(n39687) );
  XOR U42707 ( .A(n39689), .B(\modmult_1/zin[0][28] ), .Z(n30569) );
  IV U42708 ( .A(n39686), .Z(n39689) );
  XNOR U42709 ( .A(n39686), .B(n30568), .Z(n39688) );
  XOR U42710 ( .A(n39690), .B(n39691), .Z(n30568) );
  AND U42711 ( .A(\modmult_1/xin[1023] ), .B(n39692), .Z(n39691) );
  IV U42712 ( .A(n39690), .Z(n39692) );
  XOR U42713 ( .A(n39693), .B(mreg[29]), .Z(n39690) );
  NAND U42714 ( .A(n39694), .B(mul_pow), .Z(n39693) );
  XOR U42715 ( .A(mreg[29]), .B(creg[29]), .Z(n39694) );
  XOR U42716 ( .A(n39695), .B(n39696), .Z(n39686) );
  ANDN U42717 ( .A(n39697), .B(n30575), .Z(n39696) );
  XOR U42718 ( .A(n39698), .B(\modmult_1/zin[0][27] ), .Z(n30575) );
  IV U42719 ( .A(n39695), .Z(n39698) );
  XNOR U42720 ( .A(n39695), .B(n30574), .Z(n39697) );
  XOR U42721 ( .A(n39699), .B(n39700), .Z(n30574) );
  AND U42722 ( .A(\modmult_1/xin[1023] ), .B(n39701), .Z(n39700) );
  IV U42723 ( .A(n39699), .Z(n39701) );
  XOR U42724 ( .A(n39702), .B(mreg[28]), .Z(n39699) );
  NAND U42725 ( .A(n39703), .B(mul_pow), .Z(n39702) );
  XOR U42726 ( .A(mreg[28]), .B(creg[28]), .Z(n39703) );
  XOR U42727 ( .A(n39704), .B(n39705), .Z(n39695) );
  ANDN U42728 ( .A(n39706), .B(n30581), .Z(n39705) );
  XOR U42729 ( .A(n39707), .B(\modmult_1/zin[0][26] ), .Z(n30581) );
  IV U42730 ( .A(n39704), .Z(n39707) );
  XNOR U42731 ( .A(n39704), .B(n30580), .Z(n39706) );
  XOR U42732 ( .A(n39708), .B(n39709), .Z(n30580) );
  AND U42733 ( .A(\modmult_1/xin[1023] ), .B(n39710), .Z(n39709) );
  IV U42734 ( .A(n39708), .Z(n39710) );
  XOR U42735 ( .A(n39711), .B(mreg[27]), .Z(n39708) );
  NAND U42736 ( .A(n39712), .B(mul_pow), .Z(n39711) );
  XOR U42737 ( .A(mreg[27]), .B(creg[27]), .Z(n39712) );
  XOR U42738 ( .A(n39713), .B(n39714), .Z(n39704) );
  ANDN U42739 ( .A(n39715), .B(n30587), .Z(n39714) );
  XOR U42740 ( .A(n39716), .B(\modmult_1/zin[0][25] ), .Z(n30587) );
  IV U42741 ( .A(n39713), .Z(n39716) );
  XNOR U42742 ( .A(n39713), .B(n30586), .Z(n39715) );
  XOR U42743 ( .A(n39717), .B(n39718), .Z(n30586) );
  AND U42744 ( .A(\modmult_1/xin[1023] ), .B(n39719), .Z(n39718) );
  IV U42745 ( .A(n39717), .Z(n39719) );
  XOR U42746 ( .A(n39720), .B(mreg[26]), .Z(n39717) );
  NAND U42747 ( .A(n39721), .B(mul_pow), .Z(n39720) );
  XOR U42748 ( .A(mreg[26]), .B(creg[26]), .Z(n39721) );
  XOR U42749 ( .A(n39722), .B(n39723), .Z(n39713) );
  ANDN U42750 ( .A(n39724), .B(n30593), .Z(n39723) );
  XOR U42751 ( .A(n39725), .B(\modmult_1/zin[0][24] ), .Z(n30593) );
  IV U42752 ( .A(n39722), .Z(n39725) );
  XNOR U42753 ( .A(n39722), .B(n30592), .Z(n39724) );
  XOR U42754 ( .A(n39726), .B(n39727), .Z(n30592) );
  AND U42755 ( .A(\modmult_1/xin[1023] ), .B(n39728), .Z(n39727) );
  IV U42756 ( .A(n39726), .Z(n39728) );
  XOR U42757 ( .A(n39729), .B(mreg[25]), .Z(n39726) );
  NAND U42758 ( .A(n39730), .B(mul_pow), .Z(n39729) );
  XOR U42759 ( .A(mreg[25]), .B(creg[25]), .Z(n39730) );
  XOR U42760 ( .A(n39731), .B(n39732), .Z(n39722) );
  ANDN U42761 ( .A(n39733), .B(n30599), .Z(n39732) );
  XOR U42762 ( .A(n39734), .B(\modmult_1/zin[0][23] ), .Z(n30599) );
  IV U42763 ( .A(n39731), .Z(n39734) );
  XNOR U42764 ( .A(n39731), .B(n30598), .Z(n39733) );
  XOR U42765 ( .A(n39735), .B(n39736), .Z(n30598) );
  AND U42766 ( .A(\modmult_1/xin[1023] ), .B(n39737), .Z(n39736) );
  IV U42767 ( .A(n39735), .Z(n39737) );
  XOR U42768 ( .A(n39738), .B(mreg[24]), .Z(n39735) );
  NAND U42769 ( .A(n39739), .B(mul_pow), .Z(n39738) );
  XOR U42770 ( .A(mreg[24]), .B(creg[24]), .Z(n39739) );
  XOR U42771 ( .A(n39740), .B(n39741), .Z(n39731) );
  ANDN U42772 ( .A(n39742), .B(n30605), .Z(n39741) );
  XOR U42773 ( .A(n39743), .B(\modmult_1/zin[0][22] ), .Z(n30605) );
  IV U42774 ( .A(n39740), .Z(n39743) );
  XNOR U42775 ( .A(n39740), .B(n30604), .Z(n39742) );
  XOR U42776 ( .A(n39744), .B(n39745), .Z(n30604) );
  AND U42777 ( .A(\modmult_1/xin[1023] ), .B(n39746), .Z(n39745) );
  IV U42778 ( .A(n39744), .Z(n39746) );
  XOR U42779 ( .A(n39747), .B(mreg[23]), .Z(n39744) );
  NAND U42780 ( .A(n39748), .B(mul_pow), .Z(n39747) );
  XOR U42781 ( .A(mreg[23]), .B(creg[23]), .Z(n39748) );
  XOR U42782 ( .A(n39749), .B(n39750), .Z(n39740) );
  ANDN U42783 ( .A(n39751), .B(n30611), .Z(n39750) );
  XOR U42784 ( .A(n39752), .B(\modmult_1/zin[0][21] ), .Z(n30611) );
  IV U42785 ( .A(n39749), .Z(n39752) );
  XNOR U42786 ( .A(n39749), .B(n30610), .Z(n39751) );
  XOR U42787 ( .A(n39753), .B(n39754), .Z(n30610) );
  AND U42788 ( .A(\modmult_1/xin[1023] ), .B(n39755), .Z(n39754) );
  IV U42789 ( .A(n39753), .Z(n39755) );
  XOR U42790 ( .A(n39756), .B(mreg[22]), .Z(n39753) );
  NAND U42791 ( .A(n39757), .B(mul_pow), .Z(n39756) );
  XOR U42792 ( .A(mreg[22]), .B(creg[22]), .Z(n39757) );
  XOR U42793 ( .A(n39758), .B(n39759), .Z(n39749) );
  ANDN U42794 ( .A(n39760), .B(n30617), .Z(n39759) );
  XOR U42795 ( .A(n39761), .B(\modmult_1/zin[0][20] ), .Z(n30617) );
  IV U42796 ( .A(n39758), .Z(n39761) );
  XNOR U42797 ( .A(n39758), .B(n30616), .Z(n39760) );
  XOR U42798 ( .A(n39762), .B(n39763), .Z(n30616) );
  AND U42799 ( .A(\modmult_1/xin[1023] ), .B(n39764), .Z(n39763) );
  IV U42800 ( .A(n39762), .Z(n39764) );
  XOR U42801 ( .A(n39765), .B(mreg[21]), .Z(n39762) );
  NAND U42802 ( .A(n39766), .B(mul_pow), .Z(n39765) );
  XOR U42803 ( .A(mreg[21]), .B(creg[21]), .Z(n39766) );
  XOR U42804 ( .A(n39767), .B(n39768), .Z(n39758) );
  ANDN U42805 ( .A(n39769), .B(n30623), .Z(n39768) );
  XOR U42806 ( .A(n39770), .B(\modmult_1/zin[0][19] ), .Z(n30623) );
  IV U42807 ( .A(n39767), .Z(n39770) );
  XNOR U42808 ( .A(n39767), .B(n30622), .Z(n39769) );
  XOR U42809 ( .A(n39771), .B(n39772), .Z(n30622) );
  AND U42810 ( .A(\modmult_1/xin[1023] ), .B(n39773), .Z(n39772) );
  IV U42811 ( .A(n39771), .Z(n39773) );
  XOR U42812 ( .A(n39774), .B(mreg[20]), .Z(n39771) );
  NAND U42813 ( .A(n39775), .B(mul_pow), .Z(n39774) );
  XOR U42814 ( .A(mreg[20]), .B(creg[20]), .Z(n39775) );
  XOR U42815 ( .A(n39776), .B(n39777), .Z(n39767) );
  ANDN U42816 ( .A(n39778), .B(n30629), .Z(n39777) );
  XOR U42817 ( .A(n39779), .B(\modmult_1/zin[0][18] ), .Z(n30629) );
  IV U42818 ( .A(n39776), .Z(n39779) );
  XNOR U42819 ( .A(n39776), .B(n30628), .Z(n39778) );
  XOR U42820 ( .A(n39780), .B(n39781), .Z(n30628) );
  AND U42821 ( .A(\modmult_1/xin[1023] ), .B(n39782), .Z(n39781) );
  IV U42822 ( .A(n39780), .Z(n39782) );
  XOR U42823 ( .A(n39783), .B(mreg[19]), .Z(n39780) );
  NAND U42824 ( .A(n39784), .B(mul_pow), .Z(n39783) );
  XOR U42825 ( .A(mreg[19]), .B(creg[19]), .Z(n39784) );
  XOR U42826 ( .A(n39785), .B(n39786), .Z(n39776) );
  ANDN U42827 ( .A(n39787), .B(n30635), .Z(n39786) );
  XOR U42828 ( .A(n39788), .B(\modmult_1/zin[0][17] ), .Z(n30635) );
  IV U42829 ( .A(n39785), .Z(n39788) );
  XNOR U42830 ( .A(n39785), .B(n30634), .Z(n39787) );
  XOR U42831 ( .A(n39789), .B(n39790), .Z(n30634) );
  AND U42832 ( .A(\modmult_1/xin[1023] ), .B(n39791), .Z(n39790) );
  IV U42833 ( .A(n39789), .Z(n39791) );
  XOR U42834 ( .A(n39792), .B(mreg[18]), .Z(n39789) );
  NAND U42835 ( .A(n39793), .B(mul_pow), .Z(n39792) );
  XOR U42836 ( .A(mreg[18]), .B(creg[18]), .Z(n39793) );
  XOR U42837 ( .A(n39794), .B(n39795), .Z(n39785) );
  ANDN U42838 ( .A(n39796), .B(n30641), .Z(n39795) );
  XOR U42839 ( .A(n39797), .B(\modmult_1/zin[0][16] ), .Z(n30641) );
  IV U42840 ( .A(n39794), .Z(n39797) );
  XNOR U42841 ( .A(n39794), .B(n30640), .Z(n39796) );
  XOR U42842 ( .A(n39798), .B(n39799), .Z(n30640) );
  AND U42843 ( .A(\modmult_1/xin[1023] ), .B(n39800), .Z(n39799) );
  IV U42844 ( .A(n39798), .Z(n39800) );
  XOR U42845 ( .A(n39801), .B(mreg[17]), .Z(n39798) );
  NAND U42846 ( .A(n39802), .B(mul_pow), .Z(n39801) );
  XOR U42847 ( .A(mreg[17]), .B(creg[17]), .Z(n39802) );
  XOR U42848 ( .A(n39803), .B(n39804), .Z(n39794) );
  ANDN U42849 ( .A(n39805), .B(n30647), .Z(n39804) );
  XOR U42850 ( .A(n39806), .B(\modmult_1/zin[0][15] ), .Z(n30647) );
  IV U42851 ( .A(n39803), .Z(n39806) );
  XNOR U42852 ( .A(n39803), .B(n30646), .Z(n39805) );
  XOR U42853 ( .A(n39807), .B(n39808), .Z(n30646) );
  AND U42854 ( .A(\modmult_1/xin[1023] ), .B(n39809), .Z(n39808) );
  IV U42855 ( .A(n39807), .Z(n39809) );
  XOR U42856 ( .A(n39810), .B(mreg[16]), .Z(n39807) );
  NAND U42857 ( .A(n39811), .B(mul_pow), .Z(n39810) );
  XOR U42858 ( .A(mreg[16]), .B(creg[16]), .Z(n39811) );
  XOR U42859 ( .A(n39812), .B(n39813), .Z(n39803) );
  ANDN U42860 ( .A(n39814), .B(n30653), .Z(n39813) );
  XOR U42861 ( .A(n39815), .B(\modmult_1/zin[0][14] ), .Z(n30653) );
  IV U42862 ( .A(n39812), .Z(n39815) );
  XNOR U42863 ( .A(n39812), .B(n30652), .Z(n39814) );
  XOR U42864 ( .A(n39816), .B(n39817), .Z(n30652) );
  AND U42865 ( .A(\modmult_1/xin[1023] ), .B(n39818), .Z(n39817) );
  IV U42866 ( .A(n39816), .Z(n39818) );
  XOR U42867 ( .A(n39819), .B(mreg[15]), .Z(n39816) );
  NAND U42868 ( .A(n39820), .B(mul_pow), .Z(n39819) );
  XOR U42869 ( .A(mreg[15]), .B(creg[15]), .Z(n39820) );
  XOR U42870 ( .A(n39821), .B(n39822), .Z(n39812) );
  ANDN U42871 ( .A(n39823), .B(n30659), .Z(n39822) );
  XOR U42872 ( .A(n39824), .B(\modmult_1/zin[0][13] ), .Z(n30659) );
  IV U42873 ( .A(n39821), .Z(n39824) );
  XNOR U42874 ( .A(n39821), .B(n30658), .Z(n39823) );
  XOR U42875 ( .A(n39825), .B(n39826), .Z(n30658) );
  AND U42876 ( .A(\modmult_1/xin[1023] ), .B(n39827), .Z(n39826) );
  IV U42877 ( .A(n39825), .Z(n39827) );
  XOR U42878 ( .A(n39828), .B(mreg[14]), .Z(n39825) );
  NAND U42879 ( .A(n39829), .B(mul_pow), .Z(n39828) );
  XOR U42880 ( .A(mreg[14]), .B(creg[14]), .Z(n39829) );
  XOR U42881 ( .A(n39830), .B(n39831), .Z(n39821) );
  ANDN U42882 ( .A(n39832), .B(n30665), .Z(n39831) );
  XOR U42883 ( .A(n39833), .B(\modmult_1/zin[0][12] ), .Z(n30665) );
  IV U42884 ( .A(n39830), .Z(n39833) );
  XNOR U42885 ( .A(n39830), .B(n30664), .Z(n39832) );
  XOR U42886 ( .A(n39834), .B(n39835), .Z(n30664) );
  AND U42887 ( .A(\modmult_1/xin[1023] ), .B(n39836), .Z(n39835) );
  IV U42888 ( .A(n39834), .Z(n39836) );
  XOR U42889 ( .A(n39837), .B(mreg[13]), .Z(n39834) );
  NAND U42890 ( .A(n39838), .B(mul_pow), .Z(n39837) );
  XOR U42891 ( .A(mreg[13]), .B(creg[13]), .Z(n39838) );
  XOR U42892 ( .A(n39839), .B(n39840), .Z(n39830) );
  ANDN U42893 ( .A(n39841), .B(n30671), .Z(n39840) );
  XOR U42894 ( .A(n39842), .B(\modmult_1/zin[0][11] ), .Z(n30671) );
  IV U42895 ( .A(n39839), .Z(n39842) );
  XNOR U42896 ( .A(n39839), .B(n30670), .Z(n39841) );
  XOR U42897 ( .A(n39843), .B(n39844), .Z(n30670) );
  AND U42898 ( .A(\modmult_1/xin[1023] ), .B(n39845), .Z(n39844) );
  IV U42899 ( .A(n39843), .Z(n39845) );
  XOR U42900 ( .A(n39846), .B(mreg[12]), .Z(n39843) );
  NAND U42901 ( .A(n39847), .B(mul_pow), .Z(n39846) );
  XOR U42902 ( .A(mreg[12]), .B(creg[12]), .Z(n39847) );
  XOR U42903 ( .A(n39848), .B(n39849), .Z(n39839) );
  ANDN U42904 ( .A(n39850), .B(n30677), .Z(n39849) );
  XOR U42905 ( .A(n39851), .B(\modmult_1/zin[0][10] ), .Z(n30677) );
  IV U42906 ( .A(n39848), .Z(n39851) );
  XNOR U42907 ( .A(n39848), .B(n30676), .Z(n39850) );
  XOR U42908 ( .A(n39852), .B(n39853), .Z(n30676) );
  AND U42909 ( .A(\modmult_1/xin[1023] ), .B(n39854), .Z(n39853) );
  IV U42910 ( .A(n39852), .Z(n39854) );
  XOR U42911 ( .A(n39855), .B(mreg[11]), .Z(n39852) );
  NAND U42912 ( .A(n39856), .B(mul_pow), .Z(n39855) );
  XOR U42913 ( .A(mreg[11]), .B(creg[11]), .Z(n39856) );
  XOR U42914 ( .A(n39857), .B(n39858), .Z(n39848) );
  ANDN U42915 ( .A(n39859), .B(n30683), .Z(n39858) );
  XOR U42916 ( .A(n39860), .B(\modmult_1/zin[0][9] ), .Z(n30683) );
  IV U42917 ( .A(n39857), .Z(n39860) );
  XNOR U42918 ( .A(n39857), .B(n30682), .Z(n39859) );
  XOR U42919 ( .A(n39861), .B(n39862), .Z(n30682) );
  AND U42920 ( .A(\modmult_1/xin[1023] ), .B(n39863), .Z(n39862) );
  IV U42921 ( .A(n39861), .Z(n39863) );
  XOR U42922 ( .A(n39864), .B(mreg[10]), .Z(n39861) );
  NAND U42923 ( .A(n39865), .B(mul_pow), .Z(n39864) );
  XOR U42924 ( .A(mreg[10]), .B(creg[10]), .Z(n39865) );
  XOR U42925 ( .A(n39866), .B(n39867), .Z(n39857) );
  ANDN U42926 ( .A(n39868), .B(n30689), .Z(n39867) );
  XOR U42927 ( .A(n39869), .B(\modmult_1/zin[0][8] ), .Z(n30689) );
  IV U42928 ( .A(n39866), .Z(n39869) );
  XNOR U42929 ( .A(n39866), .B(n30688), .Z(n39868) );
  XOR U42930 ( .A(n39870), .B(n39871), .Z(n30688) );
  AND U42931 ( .A(\modmult_1/xin[1023] ), .B(n39872), .Z(n39871) );
  IV U42932 ( .A(n39870), .Z(n39872) );
  XOR U42933 ( .A(n39873), .B(mreg[9]), .Z(n39870) );
  NAND U42934 ( .A(n39874), .B(mul_pow), .Z(n39873) );
  XOR U42935 ( .A(mreg[9]), .B(creg[9]), .Z(n39874) );
  XOR U42936 ( .A(n39875), .B(n39876), .Z(n39866) );
  ANDN U42937 ( .A(n39877), .B(n30695), .Z(n39876) );
  XOR U42938 ( .A(n39878), .B(\modmult_1/zin[0][7] ), .Z(n30695) );
  IV U42939 ( .A(n39875), .Z(n39878) );
  XNOR U42940 ( .A(n39875), .B(n30694), .Z(n39877) );
  XOR U42941 ( .A(n39879), .B(n39880), .Z(n30694) );
  AND U42942 ( .A(\modmult_1/xin[1023] ), .B(n39881), .Z(n39880) );
  IV U42943 ( .A(n39879), .Z(n39881) );
  XOR U42944 ( .A(n39882), .B(mreg[8]), .Z(n39879) );
  NAND U42945 ( .A(n39883), .B(mul_pow), .Z(n39882) );
  XOR U42946 ( .A(mreg[8]), .B(creg[8]), .Z(n39883) );
  XOR U42947 ( .A(n39884), .B(n39885), .Z(n39875) );
  ANDN U42948 ( .A(n39886), .B(n30701), .Z(n39885) );
  XOR U42949 ( .A(n39887), .B(\modmult_1/zin[0][6] ), .Z(n30701) );
  IV U42950 ( .A(n39884), .Z(n39887) );
  XNOR U42951 ( .A(n39884), .B(n30700), .Z(n39886) );
  XOR U42952 ( .A(n39888), .B(n39889), .Z(n30700) );
  AND U42953 ( .A(\modmult_1/xin[1023] ), .B(n39890), .Z(n39889) );
  IV U42954 ( .A(n39888), .Z(n39890) );
  XOR U42955 ( .A(n39891), .B(mreg[7]), .Z(n39888) );
  NAND U42956 ( .A(n39892), .B(mul_pow), .Z(n39891) );
  XOR U42957 ( .A(mreg[7]), .B(creg[7]), .Z(n39892) );
  XOR U42958 ( .A(n39893), .B(n39894), .Z(n39884) );
  ANDN U42959 ( .A(n39895), .B(n30707), .Z(n39894) );
  XOR U42960 ( .A(n39896), .B(\modmult_1/zin[0][5] ), .Z(n30707) );
  IV U42961 ( .A(n39893), .Z(n39896) );
  XNOR U42962 ( .A(n39893), .B(n30706), .Z(n39895) );
  XOR U42963 ( .A(n39897), .B(n39898), .Z(n30706) );
  AND U42964 ( .A(\modmult_1/xin[1023] ), .B(n39899), .Z(n39898) );
  IV U42965 ( .A(n39897), .Z(n39899) );
  XOR U42966 ( .A(n39900), .B(mreg[6]), .Z(n39897) );
  NAND U42967 ( .A(n39901), .B(mul_pow), .Z(n39900) );
  XOR U42968 ( .A(mreg[6]), .B(creg[6]), .Z(n39901) );
  XOR U42969 ( .A(n39902), .B(n39903), .Z(n39893) );
  ANDN U42970 ( .A(n39904), .B(n30713), .Z(n39903) );
  XOR U42971 ( .A(n39905), .B(\modmult_1/zin[0][4] ), .Z(n30713) );
  IV U42972 ( .A(n39902), .Z(n39905) );
  XNOR U42973 ( .A(n39902), .B(n30712), .Z(n39904) );
  XOR U42974 ( .A(n39906), .B(n39907), .Z(n30712) );
  AND U42975 ( .A(\modmult_1/xin[1023] ), .B(n39908), .Z(n39907) );
  IV U42976 ( .A(n39906), .Z(n39908) );
  XOR U42977 ( .A(n39909), .B(mreg[5]), .Z(n39906) );
  NAND U42978 ( .A(n39910), .B(mul_pow), .Z(n39909) );
  XOR U42979 ( .A(mreg[5]), .B(creg[5]), .Z(n39910) );
  XOR U42980 ( .A(n39911), .B(n39912), .Z(n39902) );
  ANDN U42981 ( .A(n39913), .B(n30719), .Z(n39912) );
  XOR U42982 ( .A(n39914), .B(\modmult_1/zin[0][3] ), .Z(n30719) );
  IV U42983 ( .A(n39911), .Z(n39914) );
  XNOR U42984 ( .A(n39911), .B(n30718), .Z(n39913) );
  XOR U42985 ( .A(n39915), .B(n39916), .Z(n30718) );
  AND U42986 ( .A(\modmult_1/xin[1023] ), .B(n39917), .Z(n39916) );
  IV U42987 ( .A(n39915), .Z(n39917) );
  XOR U42988 ( .A(n39918), .B(mreg[4]), .Z(n39915) );
  NAND U42989 ( .A(n39919), .B(mul_pow), .Z(n39918) );
  XOR U42990 ( .A(mreg[4]), .B(creg[4]), .Z(n39919) );
  XNOR U42991 ( .A(n39920), .B(n39921), .Z(n39911) );
  ANDN U42992 ( .A(n39922), .B(n30725), .Z(n39921) );
  XOR U42993 ( .A(n39920), .B(\modmult_1/zin[0][2] ), .Z(n30725) );
  XOR U42994 ( .A(n39920), .B(n30724), .Z(n39922) );
  XOR U42995 ( .A(n39923), .B(n39924), .Z(n30724) );
  AND U42996 ( .A(\modmult_1/xin[1023] ), .B(n39925), .Z(n39924) );
  IV U42997 ( .A(n39923), .Z(n39925) );
  XOR U42998 ( .A(n39926), .B(mreg[3]), .Z(n39923) );
  NAND U42999 ( .A(n39927), .B(mul_pow), .Z(n39926) );
  XOR U43000 ( .A(mreg[3]), .B(creg[3]), .Z(n39927) );
  XOR U43001 ( .A(n39928), .B(n39929), .Z(n39920) );
  NAND U43002 ( .A(n39930), .B(n30731), .Z(n39928) );
  XNOR U43003 ( .A(n39931), .B(\modmult_1/zin[0][1] ), .Z(n30731) );
  IV U43004 ( .A(n39929), .Z(n39931) );
  XNOR U43005 ( .A(n39929), .B(n30730), .Z(n39930) );
  XOR U43006 ( .A(n39932), .B(n39933), .Z(n30730) );
  AND U43007 ( .A(\modmult_1/xin[1023] ), .B(n39934), .Z(n39933) );
  IV U43008 ( .A(n39932), .Z(n39934) );
  XOR U43009 ( .A(n39935), .B(mreg[2]), .Z(n39932) );
  NAND U43010 ( .A(n39936), .B(mul_pow), .Z(n39935) );
  XOR U43011 ( .A(mreg[2]), .B(creg[2]), .Z(n39936) );
  ANDN U43012 ( .A(\modmult_1/zin[0][0] ), .B(n39937), .Z(n39929) );
  XOR U43013 ( .A(n39938), .B(n39939), .Z(n24589) );
  AND U43014 ( .A(n39938), .B(\modmult_1/xin[1023] ), .Z(n39939) );
  XNOR U43015 ( .A(n39940), .B(mreg[0]), .Z(n39938) );
  NAND U43016 ( .A(n39941), .B(mul_pow), .Z(n39940) );
  XOR U43017 ( .A(mreg[0]), .B(creg[0]), .Z(n39941) );
  XNOR U43018 ( .A(n39937), .B(\modmult_1/zin[0][0] ), .Z(n24592) );
  XOR U43019 ( .A(n39942), .B(n39943), .Z(n39937) );
  AND U43020 ( .A(\modmult_1/xin[1023] ), .B(n39944), .Z(n39943) );
  IV U43021 ( .A(n39942), .Z(n39944) );
  XOR U43022 ( .A(n39945), .B(mreg[1]), .Z(n39942) );
  NAND U43023 ( .A(n39946), .B(mul_pow), .Z(n39945) );
  XOR U43024 ( .A(mreg[1]), .B(creg[1]), .Z(n39946) );
  IV U43025 ( .A(start_in[0]), .Z(n4110) );
  XOR U43026 ( .A(ein[8]), .B(n39947), .Z(ereg_next[9]) );
  AND U43027 ( .A(mul_pow), .B(n39948), .Z(n39947) );
  XOR U43028 ( .A(ein[9]), .B(ein[8]), .Z(n39948) );
  XOR U43029 ( .A(ein[98]), .B(n39949), .Z(ereg_next[99]) );
  AND U43030 ( .A(mul_pow), .B(n39950), .Z(n39949) );
  XOR U43031 ( .A(ein[99]), .B(ein[98]), .Z(n39950) );
  XOR U43032 ( .A(ein[998]), .B(n39951), .Z(ereg_next[999]) );
  AND U43033 ( .A(mul_pow), .B(n39952), .Z(n39951) );
  XOR U43034 ( .A(ein[999]), .B(ein[998]), .Z(n39952) );
  XOR U43035 ( .A(ein[997]), .B(n39953), .Z(ereg_next[998]) );
  AND U43036 ( .A(mul_pow), .B(n39954), .Z(n39953) );
  XOR U43037 ( .A(ein[998]), .B(ein[997]), .Z(n39954) );
  XOR U43038 ( .A(ein[996]), .B(n39955), .Z(ereg_next[997]) );
  AND U43039 ( .A(mul_pow), .B(n39956), .Z(n39955) );
  XOR U43040 ( .A(ein[997]), .B(ein[996]), .Z(n39956) );
  XOR U43041 ( .A(ein[995]), .B(n39957), .Z(ereg_next[996]) );
  AND U43042 ( .A(mul_pow), .B(n39958), .Z(n39957) );
  XOR U43043 ( .A(ein[996]), .B(ein[995]), .Z(n39958) );
  XOR U43044 ( .A(ein[994]), .B(n39959), .Z(ereg_next[995]) );
  AND U43045 ( .A(mul_pow), .B(n39960), .Z(n39959) );
  XOR U43046 ( .A(ein[995]), .B(ein[994]), .Z(n39960) );
  XOR U43047 ( .A(ein[993]), .B(n39961), .Z(ereg_next[994]) );
  AND U43048 ( .A(mul_pow), .B(n39962), .Z(n39961) );
  XOR U43049 ( .A(ein[994]), .B(ein[993]), .Z(n39962) );
  XOR U43050 ( .A(ein[992]), .B(n39963), .Z(ereg_next[993]) );
  AND U43051 ( .A(mul_pow), .B(n39964), .Z(n39963) );
  XOR U43052 ( .A(ein[993]), .B(ein[992]), .Z(n39964) );
  XOR U43053 ( .A(ein[991]), .B(n39965), .Z(ereg_next[992]) );
  AND U43054 ( .A(mul_pow), .B(n39966), .Z(n39965) );
  XOR U43055 ( .A(ein[992]), .B(ein[991]), .Z(n39966) );
  XOR U43056 ( .A(ein[990]), .B(n39967), .Z(ereg_next[991]) );
  AND U43057 ( .A(mul_pow), .B(n39968), .Z(n39967) );
  XOR U43058 ( .A(ein[991]), .B(ein[990]), .Z(n39968) );
  XOR U43059 ( .A(ein[989]), .B(n39969), .Z(ereg_next[990]) );
  AND U43060 ( .A(mul_pow), .B(n39970), .Z(n39969) );
  XOR U43061 ( .A(ein[990]), .B(ein[989]), .Z(n39970) );
  XOR U43062 ( .A(ein[97]), .B(n39971), .Z(ereg_next[98]) );
  AND U43063 ( .A(mul_pow), .B(n39972), .Z(n39971) );
  XOR U43064 ( .A(ein[98]), .B(ein[97]), .Z(n39972) );
  XOR U43065 ( .A(ein[988]), .B(n39973), .Z(ereg_next[989]) );
  AND U43066 ( .A(mul_pow), .B(n39974), .Z(n39973) );
  XOR U43067 ( .A(ein[989]), .B(ein[988]), .Z(n39974) );
  XOR U43068 ( .A(ein[987]), .B(n39975), .Z(ereg_next[988]) );
  AND U43069 ( .A(mul_pow), .B(n39976), .Z(n39975) );
  XOR U43070 ( .A(ein[988]), .B(ein[987]), .Z(n39976) );
  XOR U43071 ( .A(ein[986]), .B(n39977), .Z(ereg_next[987]) );
  AND U43072 ( .A(mul_pow), .B(n39978), .Z(n39977) );
  XOR U43073 ( .A(ein[987]), .B(ein[986]), .Z(n39978) );
  XOR U43074 ( .A(ein[985]), .B(n39979), .Z(ereg_next[986]) );
  AND U43075 ( .A(mul_pow), .B(n39980), .Z(n39979) );
  XOR U43076 ( .A(ein[986]), .B(ein[985]), .Z(n39980) );
  XOR U43077 ( .A(ein[984]), .B(n39981), .Z(ereg_next[985]) );
  AND U43078 ( .A(mul_pow), .B(n39982), .Z(n39981) );
  XOR U43079 ( .A(ein[985]), .B(ein[984]), .Z(n39982) );
  XOR U43080 ( .A(ein[983]), .B(n39983), .Z(ereg_next[984]) );
  AND U43081 ( .A(mul_pow), .B(n39984), .Z(n39983) );
  XOR U43082 ( .A(ein[984]), .B(ein[983]), .Z(n39984) );
  XOR U43083 ( .A(ein[982]), .B(n39985), .Z(ereg_next[983]) );
  AND U43084 ( .A(mul_pow), .B(n39986), .Z(n39985) );
  XOR U43085 ( .A(ein[983]), .B(ein[982]), .Z(n39986) );
  XOR U43086 ( .A(ein[981]), .B(n39987), .Z(ereg_next[982]) );
  AND U43087 ( .A(mul_pow), .B(n39988), .Z(n39987) );
  XOR U43088 ( .A(ein[982]), .B(ein[981]), .Z(n39988) );
  XOR U43089 ( .A(ein[980]), .B(n39989), .Z(ereg_next[981]) );
  AND U43090 ( .A(mul_pow), .B(n39990), .Z(n39989) );
  XOR U43091 ( .A(ein[981]), .B(ein[980]), .Z(n39990) );
  XOR U43092 ( .A(ein[979]), .B(n39991), .Z(ereg_next[980]) );
  AND U43093 ( .A(mul_pow), .B(n39992), .Z(n39991) );
  XOR U43094 ( .A(ein[980]), .B(ein[979]), .Z(n39992) );
  XOR U43095 ( .A(ein[96]), .B(n39993), .Z(ereg_next[97]) );
  AND U43096 ( .A(mul_pow), .B(n39994), .Z(n39993) );
  XOR U43097 ( .A(ein[97]), .B(ein[96]), .Z(n39994) );
  XOR U43098 ( .A(ein[978]), .B(n39995), .Z(ereg_next[979]) );
  AND U43099 ( .A(mul_pow), .B(n39996), .Z(n39995) );
  XOR U43100 ( .A(ein[979]), .B(ein[978]), .Z(n39996) );
  XOR U43101 ( .A(ein[977]), .B(n39997), .Z(ereg_next[978]) );
  AND U43102 ( .A(mul_pow), .B(n39998), .Z(n39997) );
  XOR U43103 ( .A(ein[978]), .B(ein[977]), .Z(n39998) );
  XOR U43104 ( .A(ein[976]), .B(n39999), .Z(ereg_next[977]) );
  AND U43105 ( .A(mul_pow), .B(n40000), .Z(n39999) );
  XOR U43106 ( .A(ein[977]), .B(ein[976]), .Z(n40000) );
  XOR U43107 ( .A(ein[975]), .B(n40001), .Z(ereg_next[976]) );
  AND U43108 ( .A(mul_pow), .B(n40002), .Z(n40001) );
  XOR U43109 ( .A(ein[976]), .B(ein[975]), .Z(n40002) );
  XOR U43110 ( .A(ein[974]), .B(n40003), .Z(ereg_next[975]) );
  AND U43111 ( .A(mul_pow), .B(n40004), .Z(n40003) );
  XOR U43112 ( .A(ein[975]), .B(ein[974]), .Z(n40004) );
  XOR U43113 ( .A(ein[973]), .B(n40005), .Z(ereg_next[974]) );
  AND U43114 ( .A(mul_pow), .B(n40006), .Z(n40005) );
  XOR U43115 ( .A(ein[974]), .B(ein[973]), .Z(n40006) );
  XOR U43116 ( .A(ein[972]), .B(n40007), .Z(ereg_next[973]) );
  AND U43117 ( .A(mul_pow), .B(n40008), .Z(n40007) );
  XOR U43118 ( .A(ein[973]), .B(ein[972]), .Z(n40008) );
  XOR U43119 ( .A(ein[971]), .B(n40009), .Z(ereg_next[972]) );
  AND U43120 ( .A(mul_pow), .B(n40010), .Z(n40009) );
  XOR U43121 ( .A(ein[972]), .B(ein[971]), .Z(n40010) );
  XOR U43122 ( .A(ein[970]), .B(n40011), .Z(ereg_next[971]) );
  AND U43123 ( .A(mul_pow), .B(n40012), .Z(n40011) );
  XOR U43124 ( .A(ein[971]), .B(ein[970]), .Z(n40012) );
  XOR U43125 ( .A(ein[969]), .B(n40013), .Z(ereg_next[970]) );
  AND U43126 ( .A(mul_pow), .B(n40014), .Z(n40013) );
  XOR U43127 ( .A(ein[970]), .B(ein[969]), .Z(n40014) );
  XOR U43128 ( .A(ein[95]), .B(n40015), .Z(ereg_next[96]) );
  AND U43129 ( .A(mul_pow), .B(n40016), .Z(n40015) );
  XOR U43130 ( .A(ein[96]), .B(ein[95]), .Z(n40016) );
  XOR U43131 ( .A(ein[968]), .B(n40017), .Z(ereg_next[969]) );
  AND U43132 ( .A(mul_pow), .B(n40018), .Z(n40017) );
  XOR U43133 ( .A(ein[969]), .B(ein[968]), .Z(n40018) );
  XOR U43134 ( .A(ein[967]), .B(n40019), .Z(ereg_next[968]) );
  AND U43135 ( .A(mul_pow), .B(n40020), .Z(n40019) );
  XOR U43136 ( .A(ein[968]), .B(ein[967]), .Z(n40020) );
  XOR U43137 ( .A(ein[966]), .B(n40021), .Z(ereg_next[967]) );
  AND U43138 ( .A(mul_pow), .B(n40022), .Z(n40021) );
  XOR U43139 ( .A(ein[967]), .B(ein[966]), .Z(n40022) );
  XOR U43140 ( .A(ein[965]), .B(n40023), .Z(ereg_next[966]) );
  AND U43141 ( .A(mul_pow), .B(n40024), .Z(n40023) );
  XOR U43142 ( .A(ein[966]), .B(ein[965]), .Z(n40024) );
  XOR U43143 ( .A(ein[964]), .B(n40025), .Z(ereg_next[965]) );
  AND U43144 ( .A(mul_pow), .B(n40026), .Z(n40025) );
  XOR U43145 ( .A(ein[965]), .B(ein[964]), .Z(n40026) );
  XOR U43146 ( .A(ein[963]), .B(n40027), .Z(ereg_next[964]) );
  AND U43147 ( .A(mul_pow), .B(n40028), .Z(n40027) );
  XOR U43148 ( .A(ein[964]), .B(ein[963]), .Z(n40028) );
  XOR U43149 ( .A(ein[962]), .B(n40029), .Z(ereg_next[963]) );
  AND U43150 ( .A(mul_pow), .B(n40030), .Z(n40029) );
  XOR U43151 ( .A(ein[963]), .B(ein[962]), .Z(n40030) );
  XOR U43152 ( .A(ein[961]), .B(n40031), .Z(ereg_next[962]) );
  AND U43153 ( .A(mul_pow), .B(n40032), .Z(n40031) );
  XOR U43154 ( .A(ein[962]), .B(ein[961]), .Z(n40032) );
  XOR U43155 ( .A(ein[960]), .B(n40033), .Z(ereg_next[961]) );
  AND U43156 ( .A(mul_pow), .B(n40034), .Z(n40033) );
  XOR U43157 ( .A(ein[961]), .B(ein[960]), .Z(n40034) );
  XOR U43158 ( .A(ein[959]), .B(n40035), .Z(ereg_next[960]) );
  AND U43159 ( .A(mul_pow), .B(n40036), .Z(n40035) );
  XOR U43160 ( .A(ein[960]), .B(ein[959]), .Z(n40036) );
  XOR U43161 ( .A(ein[94]), .B(n40037), .Z(ereg_next[95]) );
  AND U43162 ( .A(mul_pow), .B(n40038), .Z(n40037) );
  XOR U43163 ( .A(ein[95]), .B(ein[94]), .Z(n40038) );
  XOR U43164 ( .A(ein[958]), .B(n40039), .Z(ereg_next[959]) );
  AND U43165 ( .A(mul_pow), .B(n40040), .Z(n40039) );
  XOR U43166 ( .A(ein[959]), .B(ein[958]), .Z(n40040) );
  XOR U43167 ( .A(ein[957]), .B(n40041), .Z(ereg_next[958]) );
  AND U43168 ( .A(mul_pow), .B(n40042), .Z(n40041) );
  XOR U43169 ( .A(ein[958]), .B(ein[957]), .Z(n40042) );
  XOR U43170 ( .A(ein[956]), .B(n40043), .Z(ereg_next[957]) );
  AND U43171 ( .A(mul_pow), .B(n40044), .Z(n40043) );
  XOR U43172 ( .A(ein[957]), .B(ein[956]), .Z(n40044) );
  XOR U43173 ( .A(ein[955]), .B(n40045), .Z(ereg_next[956]) );
  AND U43174 ( .A(mul_pow), .B(n40046), .Z(n40045) );
  XOR U43175 ( .A(ein[956]), .B(ein[955]), .Z(n40046) );
  XOR U43176 ( .A(ein[954]), .B(n40047), .Z(ereg_next[955]) );
  AND U43177 ( .A(mul_pow), .B(n40048), .Z(n40047) );
  XOR U43178 ( .A(ein[955]), .B(ein[954]), .Z(n40048) );
  XOR U43179 ( .A(ein[953]), .B(n40049), .Z(ereg_next[954]) );
  AND U43180 ( .A(mul_pow), .B(n40050), .Z(n40049) );
  XOR U43181 ( .A(ein[954]), .B(ein[953]), .Z(n40050) );
  XOR U43182 ( .A(ein[952]), .B(n40051), .Z(ereg_next[953]) );
  AND U43183 ( .A(mul_pow), .B(n40052), .Z(n40051) );
  XOR U43184 ( .A(ein[953]), .B(ein[952]), .Z(n40052) );
  XOR U43185 ( .A(ein[951]), .B(n40053), .Z(ereg_next[952]) );
  AND U43186 ( .A(mul_pow), .B(n40054), .Z(n40053) );
  XOR U43187 ( .A(ein[952]), .B(ein[951]), .Z(n40054) );
  XOR U43188 ( .A(ein[950]), .B(n40055), .Z(ereg_next[951]) );
  AND U43189 ( .A(mul_pow), .B(n40056), .Z(n40055) );
  XOR U43190 ( .A(ein[951]), .B(ein[950]), .Z(n40056) );
  XOR U43191 ( .A(ein[949]), .B(n40057), .Z(ereg_next[950]) );
  AND U43192 ( .A(mul_pow), .B(n40058), .Z(n40057) );
  XOR U43193 ( .A(ein[950]), .B(ein[949]), .Z(n40058) );
  XOR U43194 ( .A(ein[93]), .B(n40059), .Z(ereg_next[94]) );
  AND U43195 ( .A(mul_pow), .B(n40060), .Z(n40059) );
  XOR U43196 ( .A(ein[94]), .B(ein[93]), .Z(n40060) );
  XOR U43197 ( .A(ein[948]), .B(n40061), .Z(ereg_next[949]) );
  AND U43198 ( .A(mul_pow), .B(n40062), .Z(n40061) );
  XOR U43199 ( .A(ein[949]), .B(ein[948]), .Z(n40062) );
  XOR U43200 ( .A(ein[947]), .B(n40063), .Z(ereg_next[948]) );
  AND U43201 ( .A(mul_pow), .B(n40064), .Z(n40063) );
  XOR U43202 ( .A(ein[948]), .B(ein[947]), .Z(n40064) );
  XOR U43203 ( .A(ein[946]), .B(n40065), .Z(ereg_next[947]) );
  AND U43204 ( .A(mul_pow), .B(n40066), .Z(n40065) );
  XOR U43205 ( .A(ein[947]), .B(ein[946]), .Z(n40066) );
  XOR U43206 ( .A(ein[945]), .B(n40067), .Z(ereg_next[946]) );
  AND U43207 ( .A(mul_pow), .B(n40068), .Z(n40067) );
  XOR U43208 ( .A(ein[946]), .B(ein[945]), .Z(n40068) );
  XOR U43209 ( .A(ein[944]), .B(n40069), .Z(ereg_next[945]) );
  AND U43210 ( .A(mul_pow), .B(n40070), .Z(n40069) );
  XOR U43211 ( .A(ein[945]), .B(ein[944]), .Z(n40070) );
  XOR U43212 ( .A(ein[943]), .B(n40071), .Z(ereg_next[944]) );
  AND U43213 ( .A(mul_pow), .B(n40072), .Z(n40071) );
  XOR U43214 ( .A(ein[944]), .B(ein[943]), .Z(n40072) );
  XOR U43215 ( .A(ein[942]), .B(n40073), .Z(ereg_next[943]) );
  AND U43216 ( .A(mul_pow), .B(n40074), .Z(n40073) );
  XOR U43217 ( .A(ein[943]), .B(ein[942]), .Z(n40074) );
  XOR U43218 ( .A(ein[941]), .B(n40075), .Z(ereg_next[942]) );
  AND U43219 ( .A(mul_pow), .B(n40076), .Z(n40075) );
  XOR U43220 ( .A(ein[942]), .B(ein[941]), .Z(n40076) );
  XOR U43221 ( .A(ein[940]), .B(n40077), .Z(ereg_next[941]) );
  AND U43222 ( .A(mul_pow), .B(n40078), .Z(n40077) );
  XOR U43223 ( .A(ein[941]), .B(ein[940]), .Z(n40078) );
  XOR U43224 ( .A(ein[939]), .B(n40079), .Z(ereg_next[940]) );
  AND U43225 ( .A(mul_pow), .B(n40080), .Z(n40079) );
  XOR U43226 ( .A(ein[940]), .B(ein[939]), .Z(n40080) );
  XOR U43227 ( .A(ein[92]), .B(n40081), .Z(ereg_next[93]) );
  AND U43228 ( .A(mul_pow), .B(n40082), .Z(n40081) );
  XOR U43229 ( .A(ein[93]), .B(ein[92]), .Z(n40082) );
  XOR U43230 ( .A(ein[938]), .B(n40083), .Z(ereg_next[939]) );
  AND U43231 ( .A(mul_pow), .B(n40084), .Z(n40083) );
  XOR U43232 ( .A(ein[939]), .B(ein[938]), .Z(n40084) );
  XOR U43233 ( .A(ein[937]), .B(n40085), .Z(ereg_next[938]) );
  AND U43234 ( .A(mul_pow), .B(n40086), .Z(n40085) );
  XOR U43235 ( .A(ein[938]), .B(ein[937]), .Z(n40086) );
  XOR U43236 ( .A(ein[936]), .B(n40087), .Z(ereg_next[937]) );
  AND U43237 ( .A(mul_pow), .B(n40088), .Z(n40087) );
  XOR U43238 ( .A(ein[937]), .B(ein[936]), .Z(n40088) );
  XOR U43239 ( .A(ein[935]), .B(n40089), .Z(ereg_next[936]) );
  AND U43240 ( .A(mul_pow), .B(n40090), .Z(n40089) );
  XOR U43241 ( .A(ein[936]), .B(ein[935]), .Z(n40090) );
  XOR U43242 ( .A(ein[934]), .B(n40091), .Z(ereg_next[935]) );
  AND U43243 ( .A(mul_pow), .B(n40092), .Z(n40091) );
  XOR U43244 ( .A(ein[935]), .B(ein[934]), .Z(n40092) );
  XOR U43245 ( .A(ein[933]), .B(n40093), .Z(ereg_next[934]) );
  AND U43246 ( .A(mul_pow), .B(n40094), .Z(n40093) );
  XOR U43247 ( .A(ein[934]), .B(ein[933]), .Z(n40094) );
  XOR U43248 ( .A(ein[932]), .B(n40095), .Z(ereg_next[933]) );
  AND U43249 ( .A(mul_pow), .B(n40096), .Z(n40095) );
  XOR U43250 ( .A(ein[933]), .B(ein[932]), .Z(n40096) );
  XOR U43251 ( .A(ein[931]), .B(n40097), .Z(ereg_next[932]) );
  AND U43252 ( .A(mul_pow), .B(n40098), .Z(n40097) );
  XOR U43253 ( .A(ein[932]), .B(ein[931]), .Z(n40098) );
  XOR U43254 ( .A(ein[930]), .B(n40099), .Z(ereg_next[931]) );
  AND U43255 ( .A(mul_pow), .B(n40100), .Z(n40099) );
  XOR U43256 ( .A(ein[931]), .B(ein[930]), .Z(n40100) );
  XOR U43257 ( .A(ein[929]), .B(n40101), .Z(ereg_next[930]) );
  AND U43258 ( .A(mul_pow), .B(n40102), .Z(n40101) );
  XOR U43259 ( .A(ein[930]), .B(ein[929]), .Z(n40102) );
  XOR U43260 ( .A(ein[91]), .B(n40103), .Z(ereg_next[92]) );
  AND U43261 ( .A(mul_pow), .B(n40104), .Z(n40103) );
  XOR U43262 ( .A(ein[92]), .B(ein[91]), .Z(n40104) );
  XOR U43263 ( .A(ein[928]), .B(n40105), .Z(ereg_next[929]) );
  AND U43264 ( .A(mul_pow), .B(n40106), .Z(n40105) );
  XOR U43265 ( .A(ein[929]), .B(ein[928]), .Z(n40106) );
  XOR U43266 ( .A(ein[927]), .B(n40107), .Z(ereg_next[928]) );
  AND U43267 ( .A(mul_pow), .B(n40108), .Z(n40107) );
  XOR U43268 ( .A(ein[928]), .B(ein[927]), .Z(n40108) );
  XOR U43269 ( .A(ein[926]), .B(n40109), .Z(ereg_next[927]) );
  AND U43270 ( .A(mul_pow), .B(n40110), .Z(n40109) );
  XOR U43271 ( .A(ein[927]), .B(ein[926]), .Z(n40110) );
  XOR U43272 ( .A(ein[925]), .B(n40111), .Z(ereg_next[926]) );
  AND U43273 ( .A(mul_pow), .B(n40112), .Z(n40111) );
  XOR U43274 ( .A(ein[926]), .B(ein[925]), .Z(n40112) );
  XOR U43275 ( .A(ein[924]), .B(n40113), .Z(ereg_next[925]) );
  AND U43276 ( .A(mul_pow), .B(n40114), .Z(n40113) );
  XOR U43277 ( .A(ein[925]), .B(ein[924]), .Z(n40114) );
  XOR U43278 ( .A(ein[923]), .B(n40115), .Z(ereg_next[924]) );
  AND U43279 ( .A(mul_pow), .B(n40116), .Z(n40115) );
  XOR U43280 ( .A(ein[924]), .B(ein[923]), .Z(n40116) );
  XOR U43281 ( .A(ein[922]), .B(n40117), .Z(ereg_next[923]) );
  AND U43282 ( .A(mul_pow), .B(n40118), .Z(n40117) );
  XOR U43283 ( .A(ein[923]), .B(ein[922]), .Z(n40118) );
  XOR U43284 ( .A(ein[921]), .B(n40119), .Z(ereg_next[922]) );
  AND U43285 ( .A(mul_pow), .B(n40120), .Z(n40119) );
  XOR U43286 ( .A(ein[922]), .B(ein[921]), .Z(n40120) );
  XOR U43287 ( .A(ein[920]), .B(n40121), .Z(ereg_next[921]) );
  AND U43288 ( .A(mul_pow), .B(n40122), .Z(n40121) );
  XOR U43289 ( .A(ein[921]), .B(ein[920]), .Z(n40122) );
  XOR U43290 ( .A(ein[919]), .B(n40123), .Z(ereg_next[920]) );
  AND U43291 ( .A(mul_pow), .B(n40124), .Z(n40123) );
  XOR U43292 ( .A(ein[920]), .B(ein[919]), .Z(n40124) );
  XOR U43293 ( .A(ein[90]), .B(n40125), .Z(ereg_next[91]) );
  AND U43294 ( .A(mul_pow), .B(n40126), .Z(n40125) );
  XOR U43295 ( .A(ein[91]), .B(ein[90]), .Z(n40126) );
  XOR U43296 ( .A(ein[918]), .B(n40127), .Z(ereg_next[919]) );
  AND U43297 ( .A(mul_pow), .B(n40128), .Z(n40127) );
  XOR U43298 ( .A(ein[919]), .B(ein[918]), .Z(n40128) );
  XOR U43299 ( .A(ein[917]), .B(n40129), .Z(ereg_next[918]) );
  AND U43300 ( .A(mul_pow), .B(n40130), .Z(n40129) );
  XOR U43301 ( .A(ein[918]), .B(ein[917]), .Z(n40130) );
  XOR U43302 ( .A(ein[916]), .B(n40131), .Z(ereg_next[917]) );
  AND U43303 ( .A(mul_pow), .B(n40132), .Z(n40131) );
  XOR U43304 ( .A(ein[917]), .B(ein[916]), .Z(n40132) );
  XOR U43305 ( .A(ein[915]), .B(n40133), .Z(ereg_next[916]) );
  AND U43306 ( .A(mul_pow), .B(n40134), .Z(n40133) );
  XOR U43307 ( .A(ein[916]), .B(ein[915]), .Z(n40134) );
  XOR U43308 ( .A(ein[914]), .B(n40135), .Z(ereg_next[915]) );
  AND U43309 ( .A(mul_pow), .B(n40136), .Z(n40135) );
  XOR U43310 ( .A(ein[915]), .B(ein[914]), .Z(n40136) );
  XOR U43311 ( .A(ein[913]), .B(n40137), .Z(ereg_next[914]) );
  AND U43312 ( .A(mul_pow), .B(n40138), .Z(n40137) );
  XOR U43313 ( .A(ein[914]), .B(ein[913]), .Z(n40138) );
  XOR U43314 ( .A(ein[912]), .B(n40139), .Z(ereg_next[913]) );
  AND U43315 ( .A(mul_pow), .B(n40140), .Z(n40139) );
  XOR U43316 ( .A(ein[913]), .B(ein[912]), .Z(n40140) );
  XOR U43317 ( .A(ein[911]), .B(n40141), .Z(ereg_next[912]) );
  AND U43318 ( .A(mul_pow), .B(n40142), .Z(n40141) );
  XOR U43319 ( .A(ein[912]), .B(ein[911]), .Z(n40142) );
  XOR U43320 ( .A(ein[910]), .B(n40143), .Z(ereg_next[911]) );
  AND U43321 ( .A(mul_pow), .B(n40144), .Z(n40143) );
  XOR U43322 ( .A(ein[911]), .B(ein[910]), .Z(n40144) );
  XOR U43323 ( .A(ein[909]), .B(n40145), .Z(ereg_next[910]) );
  AND U43324 ( .A(mul_pow), .B(n40146), .Z(n40145) );
  XOR U43325 ( .A(ein[910]), .B(ein[909]), .Z(n40146) );
  XOR U43326 ( .A(ein[89]), .B(n40147), .Z(ereg_next[90]) );
  AND U43327 ( .A(mul_pow), .B(n40148), .Z(n40147) );
  XOR U43328 ( .A(ein[90]), .B(ein[89]), .Z(n40148) );
  XOR U43329 ( .A(ein[908]), .B(n40149), .Z(ereg_next[909]) );
  AND U43330 ( .A(mul_pow), .B(n40150), .Z(n40149) );
  XOR U43331 ( .A(ein[909]), .B(ein[908]), .Z(n40150) );
  XOR U43332 ( .A(ein[907]), .B(n40151), .Z(ereg_next[908]) );
  AND U43333 ( .A(mul_pow), .B(n40152), .Z(n40151) );
  XOR U43334 ( .A(ein[908]), .B(ein[907]), .Z(n40152) );
  XOR U43335 ( .A(ein[906]), .B(n40153), .Z(ereg_next[907]) );
  AND U43336 ( .A(mul_pow), .B(n40154), .Z(n40153) );
  XOR U43337 ( .A(ein[907]), .B(ein[906]), .Z(n40154) );
  XOR U43338 ( .A(ein[905]), .B(n40155), .Z(ereg_next[906]) );
  AND U43339 ( .A(mul_pow), .B(n40156), .Z(n40155) );
  XOR U43340 ( .A(ein[906]), .B(ein[905]), .Z(n40156) );
  XOR U43341 ( .A(ein[904]), .B(n40157), .Z(ereg_next[905]) );
  AND U43342 ( .A(mul_pow), .B(n40158), .Z(n40157) );
  XOR U43343 ( .A(ein[905]), .B(ein[904]), .Z(n40158) );
  XOR U43344 ( .A(ein[903]), .B(n40159), .Z(ereg_next[904]) );
  AND U43345 ( .A(mul_pow), .B(n40160), .Z(n40159) );
  XOR U43346 ( .A(ein[904]), .B(ein[903]), .Z(n40160) );
  XOR U43347 ( .A(ein[902]), .B(n40161), .Z(ereg_next[903]) );
  AND U43348 ( .A(mul_pow), .B(n40162), .Z(n40161) );
  XOR U43349 ( .A(ein[903]), .B(ein[902]), .Z(n40162) );
  XOR U43350 ( .A(ein[901]), .B(n40163), .Z(ereg_next[902]) );
  AND U43351 ( .A(mul_pow), .B(n40164), .Z(n40163) );
  XOR U43352 ( .A(ein[902]), .B(ein[901]), .Z(n40164) );
  XOR U43353 ( .A(ein[900]), .B(n40165), .Z(ereg_next[901]) );
  AND U43354 ( .A(mul_pow), .B(n40166), .Z(n40165) );
  XOR U43355 ( .A(ein[901]), .B(ein[900]), .Z(n40166) );
  XOR U43356 ( .A(ein[899]), .B(n40167), .Z(ereg_next[900]) );
  AND U43357 ( .A(mul_pow), .B(n40168), .Z(n40167) );
  XOR U43358 ( .A(ein[900]), .B(ein[899]), .Z(n40168) );
  XOR U43359 ( .A(ein[7]), .B(n40169), .Z(ereg_next[8]) );
  AND U43360 ( .A(mul_pow), .B(n40170), .Z(n40169) );
  XOR U43361 ( .A(ein[8]), .B(ein[7]), .Z(n40170) );
  XOR U43362 ( .A(ein[88]), .B(n40171), .Z(ereg_next[89]) );
  AND U43363 ( .A(mul_pow), .B(n40172), .Z(n40171) );
  XOR U43364 ( .A(ein[89]), .B(ein[88]), .Z(n40172) );
  XOR U43365 ( .A(ein[898]), .B(n40173), .Z(ereg_next[899]) );
  AND U43366 ( .A(mul_pow), .B(n40174), .Z(n40173) );
  XOR U43367 ( .A(ein[899]), .B(ein[898]), .Z(n40174) );
  XOR U43368 ( .A(ein[897]), .B(n40175), .Z(ereg_next[898]) );
  AND U43369 ( .A(mul_pow), .B(n40176), .Z(n40175) );
  XOR U43370 ( .A(ein[898]), .B(ein[897]), .Z(n40176) );
  XOR U43371 ( .A(ein[896]), .B(n40177), .Z(ereg_next[897]) );
  AND U43372 ( .A(mul_pow), .B(n40178), .Z(n40177) );
  XOR U43373 ( .A(ein[897]), .B(ein[896]), .Z(n40178) );
  XOR U43374 ( .A(ein[895]), .B(n40179), .Z(ereg_next[896]) );
  AND U43375 ( .A(mul_pow), .B(n40180), .Z(n40179) );
  XOR U43376 ( .A(ein[896]), .B(ein[895]), .Z(n40180) );
  XOR U43377 ( .A(ein[894]), .B(n40181), .Z(ereg_next[895]) );
  AND U43378 ( .A(mul_pow), .B(n40182), .Z(n40181) );
  XOR U43379 ( .A(ein[895]), .B(ein[894]), .Z(n40182) );
  XOR U43380 ( .A(ein[893]), .B(n40183), .Z(ereg_next[894]) );
  AND U43381 ( .A(mul_pow), .B(n40184), .Z(n40183) );
  XOR U43382 ( .A(ein[894]), .B(ein[893]), .Z(n40184) );
  XOR U43383 ( .A(ein[892]), .B(n40185), .Z(ereg_next[893]) );
  AND U43384 ( .A(mul_pow), .B(n40186), .Z(n40185) );
  XOR U43385 ( .A(ein[893]), .B(ein[892]), .Z(n40186) );
  XOR U43386 ( .A(ein[891]), .B(n40187), .Z(ereg_next[892]) );
  AND U43387 ( .A(mul_pow), .B(n40188), .Z(n40187) );
  XOR U43388 ( .A(ein[892]), .B(ein[891]), .Z(n40188) );
  XOR U43389 ( .A(ein[890]), .B(n40189), .Z(ereg_next[891]) );
  AND U43390 ( .A(mul_pow), .B(n40190), .Z(n40189) );
  XOR U43391 ( .A(ein[891]), .B(ein[890]), .Z(n40190) );
  XOR U43392 ( .A(ein[889]), .B(n40191), .Z(ereg_next[890]) );
  AND U43393 ( .A(mul_pow), .B(n40192), .Z(n40191) );
  XOR U43394 ( .A(ein[890]), .B(ein[889]), .Z(n40192) );
  XOR U43395 ( .A(ein[87]), .B(n40193), .Z(ereg_next[88]) );
  AND U43396 ( .A(mul_pow), .B(n40194), .Z(n40193) );
  XOR U43397 ( .A(ein[88]), .B(ein[87]), .Z(n40194) );
  XOR U43398 ( .A(ein[888]), .B(n40195), .Z(ereg_next[889]) );
  AND U43399 ( .A(mul_pow), .B(n40196), .Z(n40195) );
  XOR U43400 ( .A(ein[889]), .B(ein[888]), .Z(n40196) );
  XOR U43401 ( .A(ein[887]), .B(n40197), .Z(ereg_next[888]) );
  AND U43402 ( .A(mul_pow), .B(n40198), .Z(n40197) );
  XOR U43403 ( .A(ein[888]), .B(ein[887]), .Z(n40198) );
  XOR U43404 ( .A(ein[886]), .B(n40199), .Z(ereg_next[887]) );
  AND U43405 ( .A(mul_pow), .B(n40200), .Z(n40199) );
  XOR U43406 ( .A(ein[887]), .B(ein[886]), .Z(n40200) );
  XOR U43407 ( .A(ein[885]), .B(n40201), .Z(ereg_next[886]) );
  AND U43408 ( .A(mul_pow), .B(n40202), .Z(n40201) );
  XOR U43409 ( .A(ein[886]), .B(ein[885]), .Z(n40202) );
  XOR U43410 ( .A(ein[884]), .B(n40203), .Z(ereg_next[885]) );
  AND U43411 ( .A(mul_pow), .B(n40204), .Z(n40203) );
  XOR U43412 ( .A(ein[885]), .B(ein[884]), .Z(n40204) );
  XOR U43413 ( .A(ein[883]), .B(n40205), .Z(ereg_next[884]) );
  AND U43414 ( .A(mul_pow), .B(n40206), .Z(n40205) );
  XOR U43415 ( .A(ein[884]), .B(ein[883]), .Z(n40206) );
  XOR U43416 ( .A(ein[882]), .B(n40207), .Z(ereg_next[883]) );
  AND U43417 ( .A(mul_pow), .B(n40208), .Z(n40207) );
  XOR U43418 ( .A(ein[883]), .B(ein[882]), .Z(n40208) );
  XOR U43419 ( .A(ein[881]), .B(n40209), .Z(ereg_next[882]) );
  AND U43420 ( .A(mul_pow), .B(n40210), .Z(n40209) );
  XOR U43421 ( .A(ein[882]), .B(ein[881]), .Z(n40210) );
  XOR U43422 ( .A(ein[880]), .B(n40211), .Z(ereg_next[881]) );
  AND U43423 ( .A(mul_pow), .B(n40212), .Z(n40211) );
  XOR U43424 ( .A(ein[881]), .B(ein[880]), .Z(n40212) );
  XOR U43425 ( .A(ein[879]), .B(n40213), .Z(ereg_next[880]) );
  AND U43426 ( .A(mul_pow), .B(n40214), .Z(n40213) );
  XOR U43427 ( .A(ein[880]), .B(ein[879]), .Z(n40214) );
  XOR U43428 ( .A(ein[86]), .B(n40215), .Z(ereg_next[87]) );
  AND U43429 ( .A(mul_pow), .B(n40216), .Z(n40215) );
  XOR U43430 ( .A(ein[87]), .B(ein[86]), .Z(n40216) );
  XOR U43431 ( .A(ein[878]), .B(n40217), .Z(ereg_next[879]) );
  AND U43432 ( .A(mul_pow), .B(n40218), .Z(n40217) );
  XOR U43433 ( .A(ein[879]), .B(ein[878]), .Z(n40218) );
  XOR U43434 ( .A(ein[877]), .B(n40219), .Z(ereg_next[878]) );
  AND U43435 ( .A(mul_pow), .B(n40220), .Z(n40219) );
  XOR U43436 ( .A(ein[878]), .B(ein[877]), .Z(n40220) );
  XOR U43437 ( .A(ein[876]), .B(n40221), .Z(ereg_next[877]) );
  AND U43438 ( .A(mul_pow), .B(n40222), .Z(n40221) );
  XOR U43439 ( .A(ein[877]), .B(ein[876]), .Z(n40222) );
  XOR U43440 ( .A(ein[875]), .B(n40223), .Z(ereg_next[876]) );
  AND U43441 ( .A(mul_pow), .B(n40224), .Z(n40223) );
  XOR U43442 ( .A(ein[876]), .B(ein[875]), .Z(n40224) );
  XOR U43443 ( .A(ein[874]), .B(n40225), .Z(ereg_next[875]) );
  AND U43444 ( .A(mul_pow), .B(n40226), .Z(n40225) );
  XOR U43445 ( .A(ein[875]), .B(ein[874]), .Z(n40226) );
  XOR U43446 ( .A(ein[873]), .B(n40227), .Z(ereg_next[874]) );
  AND U43447 ( .A(mul_pow), .B(n40228), .Z(n40227) );
  XOR U43448 ( .A(ein[874]), .B(ein[873]), .Z(n40228) );
  XOR U43449 ( .A(ein[872]), .B(n40229), .Z(ereg_next[873]) );
  AND U43450 ( .A(mul_pow), .B(n40230), .Z(n40229) );
  XOR U43451 ( .A(ein[873]), .B(ein[872]), .Z(n40230) );
  XOR U43452 ( .A(ein[871]), .B(n40231), .Z(ereg_next[872]) );
  AND U43453 ( .A(mul_pow), .B(n40232), .Z(n40231) );
  XOR U43454 ( .A(ein[872]), .B(ein[871]), .Z(n40232) );
  XOR U43455 ( .A(ein[870]), .B(n40233), .Z(ereg_next[871]) );
  AND U43456 ( .A(mul_pow), .B(n40234), .Z(n40233) );
  XOR U43457 ( .A(ein[871]), .B(ein[870]), .Z(n40234) );
  XOR U43458 ( .A(ein[869]), .B(n40235), .Z(ereg_next[870]) );
  AND U43459 ( .A(mul_pow), .B(n40236), .Z(n40235) );
  XOR U43460 ( .A(ein[870]), .B(ein[869]), .Z(n40236) );
  XOR U43461 ( .A(ein[85]), .B(n40237), .Z(ereg_next[86]) );
  AND U43462 ( .A(mul_pow), .B(n40238), .Z(n40237) );
  XOR U43463 ( .A(ein[86]), .B(ein[85]), .Z(n40238) );
  XOR U43464 ( .A(ein[868]), .B(n40239), .Z(ereg_next[869]) );
  AND U43465 ( .A(mul_pow), .B(n40240), .Z(n40239) );
  XOR U43466 ( .A(ein[869]), .B(ein[868]), .Z(n40240) );
  XOR U43467 ( .A(ein[867]), .B(n40241), .Z(ereg_next[868]) );
  AND U43468 ( .A(mul_pow), .B(n40242), .Z(n40241) );
  XOR U43469 ( .A(ein[868]), .B(ein[867]), .Z(n40242) );
  XOR U43470 ( .A(ein[866]), .B(n40243), .Z(ereg_next[867]) );
  AND U43471 ( .A(mul_pow), .B(n40244), .Z(n40243) );
  XOR U43472 ( .A(ein[867]), .B(ein[866]), .Z(n40244) );
  XOR U43473 ( .A(ein[865]), .B(n40245), .Z(ereg_next[866]) );
  AND U43474 ( .A(mul_pow), .B(n40246), .Z(n40245) );
  XOR U43475 ( .A(ein[866]), .B(ein[865]), .Z(n40246) );
  XOR U43476 ( .A(ein[864]), .B(n40247), .Z(ereg_next[865]) );
  AND U43477 ( .A(mul_pow), .B(n40248), .Z(n40247) );
  XOR U43478 ( .A(ein[865]), .B(ein[864]), .Z(n40248) );
  XOR U43479 ( .A(ein[863]), .B(n40249), .Z(ereg_next[864]) );
  AND U43480 ( .A(mul_pow), .B(n40250), .Z(n40249) );
  XOR U43481 ( .A(ein[864]), .B(ein[863]), .Z(n40250) );
  XOR U43482 ( .A(ein[862]), .B(n40251), .Z(ereg_next[863]) );
  AND U43483 ( .A(mul_pow), .B(n40252), .Z(n40251) );
  XOR U43484 ( .A(ein[863]), .B(ein[862]), .Z(n40252) );
  XOR U43485 ( .A(ein[861]), .B(n40253), .Z(ereg_next[862]) );
  AND U43486 ( .A(mul_pow), .B(n40254), .Z(n40253) );
  XOR U43487 ( .A(ein[862]), .B(ein[861]), .Z(n40254) );
  XOR U43488 ( .A(ein[860]), .B(n40255), .Z(ereg_next[861]) );
  AND U43489 ( .A(mul_pow), .B(n40256), .Z(n40255) );
  XOR U43490 ( .A(ein[861]), .B(ein[860]), .Z(n40256) );
  XOR U43491 ( .A(ein[859]), .B(n40257), .Z(ereg_next[860]) );
  AND U43492 ( .A(mul_pow), .B(n40258), .Z(n40257) );
  XOR U43493 ( .A(ein[860]), .B(ein[859]), .Z(n40258) );
  XOR U43494 ( .A(ein[84]), .B(n40259), .Z(ereg_next[85]) );
  AND U43495 ( .A(mul_pow), .B(n40260), .Z(n40259) );
  XOR U43496 ( .A(ein[85]), .B(ein[84]), .Z(n40260) );
  XOR U43497 ( .A(ein[858]), .B(n40261), .Z(ereg_next[859]) );
  AND U43498 ( .A(mul_pow), .B(n40262), .Z(n40261) );
  XOR U43499 ( .A(ein[859]), .B(ein[858]), .Z(n40262) );
  XOR U43500 ( .A(ein[857]), .B(n40263), .Z(ereg_next[858]) );
  AND U43501 ( .A(mul_pow), .B(n40264), .Z(n40263) );
  XOR U43502 ( .A(ein[858]), .B(ein[857]), .Z(n40264) );
  XOR U43503 ( .A(ein[856]), .B(n40265), .Z(ereg_next[857]) );
  AND U43504 ( .A(mul_pow), .B(n40266), .Z(n40265) );
  XOR U43505 ( .A(ein[857]), .B(ein[856]), .Z(n40266) );
  XOR U43506 ( .A(ein[855]), .B(n40267), .Z(ereg_next[856]) );
  AND U43507 ( .A(mul_pow), .B(n40268), .Z(n40267) );
  XOR U43508 ( .A(ein[856]), .B(ein[855]), .Z(n40268) );
  XOR U43509 ( .A(ein[854]), .B(n40269), .Z(ereg_next[855]) );
  AND U43510 ( .A(mul_pow), .B(n40270), .Z(n40269) );
  XOR U43511 ( .A(ein[855]), .B(ein[854]), .Z(n40270) );
  XOR U43512 ( .A(ein[853]), .B(n40271), .Z(ereg_next[854]) );
  AND U43513 ( .A(mul_pow), .B(n40272), .Z(n40271) );
  XOR U43514 ( .A(ein[854]), .B(ein[853]), .Z(n40272) );
  XOR U43515 ( .A(ein[852]), .B(n40273), .Z(ereg_next[853]) );
  AND U43516 ( .A(mul_pow), .B(n40274), .Z(n40273) );
  XOR U43517 ( .A(ein[853]), .B(ein[852]), .Z(n40274) );
  XOR U43518 ( .A(ein[851]), .B(n40275), .Z(ereg_next[852]) );
  AND U43519 ( .A(mul_pow), .B(n40276), .Z(n40275) );
  XOR U43520 ( .A(ein[852]), .B(ein[851]), .Z(n40276) );
  XOR U43521 ( .A(ein[850]), .B(n40277), .Z(ereg_next[851]) );
  AND U43522 ( .A(mul_pow), .B(n40278), .Z(n40277) );
  XOR U43523 ( .A(ein[851]), .B(ein[850]), .Z(n40278) );
  XOR U43524 ( .A(ein[849]), .B(n40279), .Z(ereg_next[850]) );
  AND U43525 ( .A(mul_pow), .B(n40280), .Z(n40279) );
  XOR U43526 ( .A(ein[850]), .B(ein[849]), .Z(n40280) );
  XOR U43527 ( .A(ein[83]), .B(n40281), .Z(ereg_next[84]) );
  AND U43528 ( .A(mul_pow), .B(n40282), .Z(n40281) );
  XOR U43529 ( .A(ein[84]), .B(ein[83]), .Z(n40282) );
  XOR U43530 ( .A(ein[848]), .B(n40283), .Z(ereg_next[849]) );
  AND U43531 ( .A(mul_pow), .B(n40284), .Z(n40283) );
  XOR U43532 ( .A(ein[849]), .B(ein[848]), .Z(n40284) );
  XOR U43533 ( .A(ein[847]), .B(n40285), .Z(ereg_next[848]) );
  AND U43534 ( .A(mul_pow), .B(n40286), .Z(n40285) );
  XOR U43535 ( .A(ein[848]), .B(ein[847]), .Z(n40286) );
  XOR U43536 ( .A(ein[846]), .B(n40287), .Z(ereg_next[847]) );
  AND U43537 ( .A(mul_pow), .B(n40288), .Z(n40287) );
  XOR U43538 ( .A(ein[847]), .B(ein[846]), .Z(n40288) );
  XOR U43539 ( .A(ein[845]), .B(n40289), .Z(ereg_next[846]) );
  AND U43540 ( .A(mul_pow), .B(n40290), .Z(n40289) );
  XOR U43541 ( .A(ein[846]), .B(ein[845]), .Z(n40290) );
  XOR U43542 ( .A(ein[844]), .B(n40291), .Z(ereg_next[845]) );
  AND U43543 ( .A(mul_pow), .B(n40292), .Z(n40291) );
  XOR U43544 ( .A(ein[845]), .B(ein[844]), .Z(n40292) );
  XOR U43545 ( .A(ein[843]), .B(n40293), .Z(ereg_next[844]) );
  AND U43546 ( .A(mul_pow), .B(n40294), .Z(n40293) );
  XOR U43547 ( .A(ein[844]), .B(ein[843]), .Z(n40294) );
  XOR U43548 ( .A(ein[842]), .B(n40295), .Z(ereg_next[843]) );
  AND U43549 ( .A(mul_pow), .B(n40296), .Z(n40295) );
  XOR U43550 ( .A(ein[843]), .B(ein[842]), .Z(n40296) );
  XOR U43551 ( .A(ein[841]), .B(n40297), .Z(ereg_next[842]) );
  AND U43552 ( .A(mul_pow), .B(n40298), .Z(n40297) );
  XOR U43553 ( .A(ein[842]), .B(ein[841]), .Z(n40298) );
  XOR U43554 ( .A(ein[840]), .B(n40299), .Z(ereg_next[841]) );
  AND U43555 ( .A(mul_pow), .B(n40300), .Z(n40299) );
  XOR U43556 ( .A(ein[841]), .B(ein[840]), .Z(n40300) );
  XOR U43557 ( .A(ein[839]), .B(n40301), .Z(ereg_next[840]) );
  AND U43558 ( .A(mul_pow), .B(n40302), .Z(n40301) );
  XOR U43559 ( .A(ein[840]), .B(ein[839]), .Z(n40302) );
  XOR U43560 ( .A(ein[82]), .B(n40303), .Z(ereg_next[83]) );
  AND U43561 ( .A(mul_pow), .B(n40304), .Z(n40303) );
  XOR U43562 ( .A(ein[83]), .B(ein[82]), .Z(n40304) );
  XOR U43563 ( .A(ein[838]), .B(n40305), .Z(ereg_next[839]) );
  AND U43564 ( .A(mul_pow), .B(n40306), .Z(n40305) );
  XOR U43565 ( .A(ein[839]), .B(ein[838]), .Z(n40306) );
  XOR U43566 ( .A(ein[837]), .B(n40307), .Z(ereg_next[838]) );
  AND U43567 ( .A(mul_pow), .B(n40308), .Z(n40307) );
  XOR U43568 ( .A(ein[838]), .B(ein[837]), .Z(n40308) );
  XOR U43569 ( .A(ein[836]), .B(n40309), .Z(ereg_next[837]) );
  AND U43570 ( .A(mul_pow), .B(n40310), .Z(n40309) );
  XOR U43571 ( .A(ein[837]), .B(ein[836]), .Z(n40310) );
  XOR U43572 ( .A(ein[835]), .B(n40311), .Z(ereg_next[836]) );
  AND U43573 ( .A(mul_pow), .B(n40312), .Z(n40311) );
  XOR U43574 ( .A(ein[836]), .B(ein[835]), .Z(n40312) );
  XOR U43575 ( .A(ein[834]), .B(n40313), .Z(ereg_next[835]) );
  AND U43576 ( .A(mul_pow), .B(n40314), .Z(n40313) );
  XOR U43577 ( .A(ein[835]), .B(ein[834]), .Z(n40314) );
  XOR U43578 ( .A(ein[833]), .B(n40315), .Z(ereg_next[834]) );
  AND U43579 ( .A(mul_pow), .B(n40316), .Z(n40315) );
  XOR U43580 ( .A(ein[834]), .B(ein[833]), .Z(n40316) );
  XOR U43581 ( .A(ein[832]), .B(n40317), .Z(ereg_next[833]) );
  AND U43582 ( .A(mul_pow), .B(n40318), .Z(n40317) );
  XOR U43583 ( .A(ein[833]), .B(ein[832]), .Z(n40318) );
  XOR U43584 ( .A(ein[831]), .B(n40319), .Z(ereg_next[832]) );
  AND U43585 ( .A(mul_pow), .B(n40320), .Z(n40319) );
  XOR U43586 ( .A(ein[832]), .B(ein[831]), .Z(n40320) );
  XOR U43587 ( .A(ein[830]), .B(n40321), .Z(ereg_next[831]) );
  AND U43588 ( .A(mul_pow), .B(n40322), .Z(n40321) );
  XOR U43589 ( .A(ein[831]), .B(ein[830]), .Z(n40322) );
  XOR U43590 ( .A(ein[829]), .B(n40323), .Z(ereg_next[830]) );
  AND U43591 ( .A(mul_pow), .B(n40324), .Z(n40323) );
  XOR U43592 ( .A(ein[830]), .B(ein[829]), .Z(n40324) );
  XOR U43593 ( .A(ein[81]), .B(n40325), .Z(ereg_next[82]) );
  AND U43594 ( .A(mul_pow), .B(n40326), .Z(n40325) );
  XOR U43595 ( .A(ein[82]), .B(ein[81]), .Z(n40326) );
  XOR U43596 ( .A(ein[828]), .B(n40327), .Z(ereg_next[829]) );
  AND U43597 ( .A(mul_pow), .B(n40328), .Z(n40327) );
  XOR U43598 ( .A(ein[829]), .B(ein[828]), .Z(n40328) );
  XOR U43599 ( .A(ein[827]), .B(n40329), .Z(ereg_next[828]) );
  AND U43600 ( .A(mul_pow), .B(n40330), .Z(n40329) );
  XOR U43601 ( .A(ein[828]), .B(ein[827]), .Z(n40330) );
  XOR U43602 ( .A(ein[826]), .B(n40331), .Z(ereg_next[827]) );
  AND U43603 ( .A(mul_pow), .B(n40332), .Z(n40331) );
  XOR U43604 ( .A(ein[827]), .B(ein[826]), .Z(n40332) );
  XOR U43605 ( .A(ein[825]), .B(n40333), .Z(ereg_next[826]) );
  AND U43606 ( .A(mul_pow), .B(n40334), .Z(n40333) );
  XOR U43607 ( .A(ein[826]), .B(ein[825]), .Z(n40334) );
  XOR U43608 ( .A(ein[824]), .B(n40335), .Z(ereg_next[825]) );
  AND U43609 ( .A(mul_pow), .B(n40336), .Z(n40335) );
  XOR U43610 ( .A(ein[825]), .B(ein[824]), .Z(n40336) );
  XOR U43611 ( .A(ein[823]), .B(n40337), .Z(ereg_next[824]) );
  AND U43612 ( .A(mul_pow), .B(n40338), .Z(n40337) );
  XOR U43613 ( .A(ein[824]), .B(ein[823]), .Z(n40338) );
  XOR U43614 ( .A(ein[822]), .B(n40339), .Z(ereg_next[823]) );
  AND U43615 ( .A(mul_pow), .B(n40340), .Z(n40339) );
  XOR U43616 ( .A(ein[823]), .B(ein[822]), .Z(n40340) );
  XOR U43617 ( .A(ein[821]), .B(n40341), .Z(ereg_next[822]) );
  AND U43618 ( .A(mul_pow), .B(n40342), .Z(n40341) );
  XOR U43619 ( .A(ein[822]), .B(ein[821]), .Z(n40342) );
  XOR U43620 ( .A(ein[820]), .B(n40343), .Z(ereg_next[821]) );
  AND U43621 ( .A(mul_pow), .B(n40344), .Z(n40343) );
  XOR U43622 ( .A(ein[821]), .B(ein[820]), .Z(n40344) );
  XOR U43623 ( .A(ein[819]), .B(n40345), .Z(ereg_next[820]) );
  AND U43624 ( .A(mul_pow), .B(n40346), .Z(n40345) );
  XOR U43625 ( .A(ein[820]), .B(ein[819]), .Z(n40346) );
  XOR U43626 ( .A(ein[80]), .B(n40347), .Z(ereg_next[81]) );
  AND U43627 ( .A(mul_pow), .B(n40348), .Z(n40347) );
  XOR U43628 ( .A(ein[81]), .B(ein[80]), .Z(n40348) );
  XOR U43629 ( .A(ein[818]), .B(n40349), .Z(ereg_next[819]) );
  AND U43630 ( .A(mul_pow), .B(n40350), .Z(n40349) );
  XOR U43631 ( .A(ein[819]), .B(ein[818]), .Z(n40350) );
  XOR U43632 ( .A(ein[817]), .B(n40351), .Z(ereg_next[818]) );
  AND U43633 ( .A(mul_pow), .B(n40352), .Z(n40351) );
  XOR U43634 ( .A(ein[818]), .B(ein[817]), .Z(n40352) );
  XOR U43635 ( .A(ein[816]), .B(n40353), .Z(ereg_next[817]) );
  AND U43636 ( .A(mul_pow), .B(n40354), .Z(n40353) );
  XOR U43637 ( .A(ein[817]), .B(ein[816]), .Z(n40354) );
  XOR U43638 ( .A(ein[815]), .B(n40355), .Z(ereg_next[816]) );
  AND U43639 ( .A(mul_pow), .B(n40356), .Z(n40355) );
  XOR U43640 ( .A(ein[816]), .B(ein[815]), .Z(n40356) );
  XOR U43641 ( .A(ein[814]), .B(n40357), .Z(ereg_next[815]) );
  AND U43642 ( .A(mul_pow), .B(n40358), .Z(n40357) );
  XOR U43643 ( .A(ein[815]), .B(ein[814]), .Z(n40358) );
  XOR U43644 ( .A(ein[813]), .B(n40359), .Z(ereg_next[814]) );
  AND U43645 ( .A(mul_pow), .B(n40360), .Z(n40359) );
  XOR U43646 ( .A(ein[814]), .B(ein[813]), .Z(n40360) );
  XOR U43647 ( .A(ein[812]), .B(n40361), .Z(ereg_next[813]) );
  AND U43648 ( .A(mul_pow), .B(n40362), .Z(n40361) );
  XOR U43649 ( .A(ein[813]), .B(ein[812]), .Z(n40362) );
  XOR U43650 ( .A(ein[811]), .B(n40363), .Z(ereg_next[812]) );
  AND U43651 ( .A(mul_pow), .B(n40364), .Z(n40363) );
  XOR U43652 ( .A(ein[812]), .B(ein[811]), .Z(n40364) );
  XOR U43653 ( .A(ein[810]), .B(n40365), .Z(ereg_next[811]) );
  AND U43654 ( .A(mul_pow), .B(n40366), .Z(n40365) );
  XOR U43655 ( .A(ein[811]), .B(ein[810]), .Z(n40366) );
  XOR U43656 ( .A(ein[809]), .B(n40367), .Z(ereg_next[810]) );
  AND U43657 ( .A(mul_pow), .B(n40368), .Z(n40367) );
  XOR U43658 ( .A(ein[810]), .B(ein[809]), .Z(n40368) );
  XOR U43659 ( .A(ein[79]), .B(n40369), .Z(ereg_next[80]) );
  AND U43660 ( .A(mul_pow), .B(n40370), .Z(n40369) );
  XOR U43661 ( .A(ein[80]), .B(ein[79]), .Z(n40370) );
  XOR U43662 ( .A(ein[808]), .B(n40371), .Z(ereg_next[809]) );
  AND U43663 ( .A(mul_pow), .B(n40372), .Z(n40371) );
  XOR U43664 ( .A(ein[809]), .B(ein[808]), .Z(n40372) );
  XOR U43665 ( .A(ein[807]), .B(n40373), .Z(ereg_next[808]) );
  AND U43666 ( .A(mul_pow), .B(n40374), .Z(n40373) );
  XOR U43667 ( .A(ein[808]), .B(ein[807]), .Z(n40374) );
  XOR U43668 ( .A(ein[806]), .B(n40375), .Z(ereg_next[807]) );
  AND U43669 ( .A(mul_pow), .B(n40376), .Z(n40375) );
  XOR U43670 ( .A(ein[807]), .B(ein[806]), .Z(n40376) );
  XOR U43671 ( .A(ein[805]), .B(n40377), .Z(ereg_next[806]) );
  AND U43672 ( .A(mul_pow), .B(n40378), .Z(n40377) );
  XOR U43673 ( .A(ein[806]), .B(ein[805]), .Z(n40378) );
  XOR U43674 ( .A(ein[804]), .B(n40379), .Z(ereg_next[805]) );
  AND U43675 ( .A(mul_pow), .B(n40380), .Z(n40379) );
  XOR U43676 ( .A(ein[805]), .B(ein[804]), .Z(n40380) );
  XOR U43677 ( .A(ein[803]), .B(n40381), .Z(ereg_next[804]) );
  AND U43678 ( .A(mul_pow), .B(n40382), .Z(n40381) );
  XOR U43679 ( .A(ein[804]), .B(ein[803]), .Z(n40382) );
  XOR U43680 ( .A(ein[802]), .B(n40383), .Z(ereg_next[803]) );
  AND U43681 ( .A(mul_pow), .B(n40384), .Z(n40383) );
  XOR U43682 ( .A(ein[803]), .B(ein[802]), .Z(n40384) );
  XOR U43683 ( .A(ein[801]), .B(n40385), .Z(ereg_next[802]) );
  AND U43684 ( .A(mul_pow), .B(n40386), .Z(n40385) );
  XOR U43685 ( .A(ein[802]), .B(ein[801]), .Z(n40386) );
  XOR U43686 ( .A(ein[800]), .B(n40387), .Z(ereg_next[801]) );
  AND U43687 ( .A(mul_pow), .B(n40388), .Z(n40387) );
  XOR U43688 ( .A(ein[801]), .B(ein[800]), .Z(n40388) );
  XOR U43689 ( .A(ein[799]), .B(n40389), .Z(ereg_next[800]) );
  AND U43690 ( .A(mul_pow), .B(n40390), .Z(n40389) );
  XOR U43691 ( .A(ein[800]), .B(ein[799]), .Z(n40390) );
  XOR U43692 ( .A(ein[6]), .B(n40391), .Z(ereg_next[7]) );
  AND U43693 ( .A(mul_pow), .B(n40392), .Z(n40391) );
  XOR U43694 ( .A(ein[7]), .B(ein[6]), .Z(n40392) );
  XOR U43695 ( .A(ein[78]), .B(n40393), .Z(ereg_next[79]) );
  AND U43696 ( .A(mul_pow), .B(n40394), .Z(n40393) );
  XOR U43697 ( .A(ein[79]), .B(ein[78]), .Z(n40394) );
  XOR U43698 ( .A(ein[798]), .B(n40395), .Z(ereg_next[799]) );
  AND U43699 ( .A(mul_pow), .B(n40396), .Z(n40395) );
  XOR U43700 ( .A(ein[799]), .B(ein[798]), .Z(n40396) );
  XOR U43701 ( .A(ein[797]), .B(n40397), .Z(ereg_next[798]) );
  AND U43702 ( .A(mul_pow), .B(n40398), .Z(n40397) );
  XOR U43703 ( .A(ein[798]), .B(ein[797]), .Z(n40398) );
  XOR U43704 ( .A(ein[796]), .B(n40399), .Z(ereg_next[797]) );
  AND U43705 ( .A(mul_pow), .B(n40400), .Z(n40399) );
  XOR U43706 ( .A(ein[797]), .B(ein[796]), .Z(n40400) );
  XOR U43707 ( .A(ein[795]), .B(n40401), .Z(ereg_next[796]) );
  AND U43708 ( .A(mul_pow), .B(n40402), .Z(n40401) );
  XOR U43709 ( .A(ein[796]), .B(ein[795]), .Z(n40402) );
  XOR U43710 ( .A(ein[794]), .B(n40403), .Z(ereg_next[795]) );
  AND U43711 ( .A(mul_pow), .B(n40404), .Z(n40403) );
  XOR U43712 ( .A(ein[795]), .B(ein[794]), .Z(n40404) );
  XOR U43713 ( .A(ein[793]), .B(n40405), .Z(ereg_next[794]) );
  AND U43714 ( .A(mul_pow), .B(n40406), .Z(n40405) );
  XOR U43715 ( .A(ein[794]), .B(ein[793]), .Z(n40406) );
  XOR U43716 ( .A(ein[792]), .B(n40407), .Z(ereg_next[793]) );
  AND U43717 ( .A(mul_pow), .B(n40408), .Z(n40407) );
  XOR U43718 ( .A(ein[793]), .B(ein[792]), .Z(n40408) );
  XOR U43719 ( .A(ein[791]), .B(n40409), .Z(ereg_next[792]) );
  AND U43720 ( .A(mul_pow), .B(n40410), .Z(n40409) );
  XOR U43721 ( .A(ein[792]), .B(ein[791]), .Z(n40410) );
  XOR U43722 ( .A(ein[790]), .B(n40411), .Z(ereg_next[791]) );
  AND U43723 ( .A(mul_pow), .B(n40412), .Z(n40411) );
  XOR U43724 ( .A(ein[791]), .B(ein[790]), .Z(n40412) );
  XOR U43725 ( .A(ein[789]), .B(n40413), .Z(ereg_next[790]) );
  AND U43726 ( .A(mul_pow), .B(n40414), .Z(n40413) );
  XOR U43727 ( .A(ein[790]), .B(ein[789]), .Z(n40414) );
  XOR U43728 ( .A(ein[77]), .B(n40415), .Z(ereg_next[78]) );
  AND U43729 ( .A(mul_pow), .B(n40416), .Z(n40415) );
  XOR U43730 ( .A(ein[78]), .B(ein[77]), .Z(n40416) );
  XOR U43731 ( .A(ein[788]), .B(n40417), .Z(ereg_next[789]) );
  AND U43732 ( .A(mul_pow), .B(n40418), .Z(n40417) );
  XOR U43733 ( .A(ein[789]), .B(ein[788]), .Z(n40418) );
  XOR U43734 ( .A(ein[787]), .B(n40419), .Z(ereg_next[788]) );
  AND U43735 ( .A(mul_pow), .B(n40420), .Z(n40419) );
  XOR U43736 ( .A(ein[788]), .B(ein[787]), .Z(n40420) );
  XOR U43737 ( .A(ein[786]), .B(n40421), .Z(ereg_next[787]) );
  AND U43738 ( .A(mul_pow), .B(n40422), .Z(n40421) );
  XOR U43739 ( .A(ein[787]), .B(ein[786]), .Z(n40422) );
  XOR U43740 ( .A(ein[785]), .B(n40423), .Z(ereg_next[786]) );
  AND U43741 ( .A(mul_pow), .B(n40424), .Z(n40423) );
  XOR U43742 ( .A(ein[786]), .B(ein[785]), .Z(n40424) );
  XOR U43743 ( .A(ein[784]), .B(n40425), .Z(ereg_next[785]) );
  AND U43744 ( .A(mul_pow), .B(n40426), .Z(n40425) );
  XOR U43745 ( .A(ein[785]), .B(ein[784]), .Z(n40426) );
  XOR U43746 ( .A(ein[783]), .B(n40427), .Z(ereg_next[784]) );
  AND U43747 ( .A(mul_pow), .B(n40428), .Z(n40427) );
  XOR U43748 ( .A(ein[784]), .B(ein[783]), .Z(n40428) );
  XOR U43749 ( .A(ein[782]), .B(n40429), .Z(ereg_next[783]) );
  AND U43750 ( .A(mul_pow), .B(n40430), .Z(n40429) );
  XOR U43751 ( .A(ein[783]), .B(ein[782]), .Z(n40430) );
  XOR U43752 ( .A(ein[781]), .B(n40431), .Z(ereg_next[782]) );
  AND U43753 ( .A(mul_pow), .B(n40432), .Z(n40431) );
  XOR U43754 ( .A(ein[782]), .B(ein[781]), .Z(n40432) );
  XOR U43755 ( .A(ein[780]), .B(n40433), .Z(ereg_next[781]) );
  AND U43756 ( .A(mul_pow), .B(n40434), .Z(n40433) );
  XOR U43757 ( .A(ein[781]), .B(ein[780]), .Z(n40434) );
  XOR U43758 ( .A(ein[779]), .B(n40435), .Z(ereg_next[780]) );
  AND U43759 ( .A(mul_pow), .B(n40436), .Z(n40435) );
  XOR U43760 ( .A(ein[780]), .B(ein[779]), .Z(n40436) );
  XOR U43761 ( .A(ein[76]), .B(n40437), .Z(ereg_next[77]) );
  AND U43762 ( .A(mul_pow), .B(n40438), .Z(n40437) );
  XOR U43763 ( .A(ein[77]), .B(ein[76]), .Z(n40438) );
  XOR U43764 ( .A(ein[778]), .B(n40439), .Z(ereg_next[779]) );
  AND U43765 ( .A(mul_pow), .B(n40440), .Z(n40439) );
  XOR U43766 ( .A(ein[779]), .B(ein[778]), .Z(n40440) );
  XOR U43767 ( .A(ein[777]), .B(n40441), .Z(ereg_next[778]) );
  AND U43768 ( .A(mul_pow), .B(n40442), .Z(n40441) );
  XOR U43769 ( .A(ein[778]), .B(ein[777]), .Z(n40442) );
  XOR U43770 ( .A(ein[776]), .B(n40443), .Z(ereg_next[777]) );
  AND U43771 ( .A(mul_pow), .B(n40444), .Z(n40443) );
  XOR U43772 ( .A(ein[777]), .B(ein[776]), .Z(n40444) );
  XOR U43773 ( .A(ein[775]), .B(n40445), .Z(ereg_next[776]) );
  AND U43774 ( .A(mul_pow), .B(n40446), .Z(n40445) );
  XOR U43775 ( .A(ein[776]), .B(ein[775]), .Z(n40446) );
  XOR U43776 ( .A(ein[774]), .B(n40447), .Z(ereg_next[775]) );
  AND U43777 ( .A(mul_pow), .B(n40448), .Z(n40447) );
  XOR U43778 ( .A(ein[775]), .B(ein[774]), .Z(n40448) );
  XOR U43779 ( .A(ein[773]), .B(n40449), .Z(ereg_next[774]) );
  AND U43780 ( .A(mul_pow), .B(n40450), .Z(n40449) );
  XOR U43781 ( .A(ein[774]), .B(ein[773]), .Z(n40450) );
  XOR U43782 ( .A(ein[772]), .B(n40451), .Z(ereg_next[773]) );
  AND U43783 ( .A(mul_pow), .B(n40452), .Z(n40451) );
  XOR U43784 ( .A(ein[773]), .B(ein[772]), .Z(n40452) );
  XOR U43785 ( .A(ein[771]), .B(n40453), .Z(ereg_next[772]) );
  AND U43786 ( .A(mul_pow), .B(n40454), .Z(n40453) );
  XOR U43787 ( .A(ein[772]), .B(ein[771]), .Z(n40454) );
  XOR U43788 ( .A(ein[770]), .B(n40455), .Z(ereg_next[771]) );
  AND U43789 ( .A(mul_pow), .B(n40456), .Z(n40455) );
  XOR U43790 ( .A(ein[771]), .B(ein[770]), .Z(n40456) );
  XOR U43791 ( .A(ein[769]), .B(n40457), .Z(ereg_next[770]) );
  AND U43792 ( .A(mul_pow), .B(n40458), .Z(n40457) );
  XOR U43793 ( .A(ein[770]), .B(ein[769]), .Z(n40458) );
  XOR U43794 ( .A(ein[75]), .B(n40459), .Z(ereg_next[76]) );
  AND U43795 ( .A(mul_pow), .B(n40460), .Z(n40459) );
  XOR U43796 ( .A(ein[76]), .B(ein[75]), .Z(n40460) );
  XOR U43797 ( .A(ein[768]), .B(n40461), .Z(ereg_next[769]) );
  AND U43798 ( .A(mul_pow), .B(n40462), .Z(n40461) );
  XOR U43799 ( .A(ein[769]), .B(ein[768]), .Z(n40462) );
  XOR U43800 ( .A(ein[767]), .B(n40463), .Z(ereg_next[768]) );
  AND U43801 ( .A(mul_pow), .B(n40464), .Z(n40463) );
  XOR U43802 ( .A(ein[768]), .B(ein[767]), .Z(n40464) );
  XOR U43803 ( .A(ein[766]), .B(n40465), .Z(ereg_next[767]) );
  AND U43804 ( .A(mul_pow), .B(n40466), .Z(n40465) );
  XOR U43805 ( .A(ein[767]), .B(ein[766]), .Z(n40466) );
  XOR U43806 ( .A(ein[765]), .B(n40467), .Z(ereg_next[766]) );
  AND U43807 ( .A(mul_pow), .B(n40468), .Z(n40467) );
  XOR U43808 ( .A(ein[766]), .B(ein[765]), .Z(n40468) );
  XOR U43809 ( .A(ein[764]), .B(n40469), .Z(ereg_next[765]) );
  AND U43810 ( .A(mul_pow), .B(n40470), .Z(n40469) );
  XOR U43811 ( .A(ein[765]), .B(ein[764]), .Z(n40470) );
  XOR U43812 ( .A(ein[763]), .B(n40471), .Z(ereg_next[764]) );
  AND U43813 ( .A(mul_pow), .B(n40472), .Z(n40471) );
  XOR U43814 ( .A(ein[764]), .B(ein[763]), .Z(n40472) );
  XOR U43815 ( .A(ein[762]), .B(n40473), .Z(ereg_next[763]) );
  AND U43816 ( .A(mul_pow), .B(n40474), .Z(n40473) );
  XOR U43817 ( .A(ein[763]), .B(ein[762]), .Z(n40474) );
  XOR U43818 ( .A(ein[761]), .B(n40475), .Z(ereg_next[762]) );
  AND U43819 ( .A(mul_pow), .B(n40476), .Z(n40475) );
  XOR U43820 ( .A(ein[762]), .B(ein[761]), .Z(n40476) );
  XOR U43821 ( .A(ein[760]), .B(n40477), .Z(ereg_next[761]) );
  AND U43822 ( .A(mul_pow), .B(n40478), .Z(n40477) );
  XOR U43823 ( .A(ein[761]), .B(ein[760]), .Z(n40478) );
  XOR U43824 ( .A(ein[759]), .B(n40479), .Z(ereg_next[760]) );
  AND U43825 ( .A(mul_pow), .B(n40480), .Z(n40479) );
  XOR U43826 ( .A(ein[760]), .B(ein[759]), .Z(n40480) );
  XOR U43827 ( .A(ein[74]), .B(n40481), .Z(ereg_next[75]) );
  AND U43828 ( .A(mul_pow), .B(n40482), .Z(n40481) );
  XOR U43829 ( .A(ein[75]), .B(ein[74]), .Z(n40482) );
  XOR U43830 ( .A(ein[758]), .B(n40483), .Z(ereg_next[759]) );
  AND U43831 ( .A(mul_pow), .B(n40484), .Z(n40483) );
  XOR U43832 ( .A(ein[759]), .B(ein[758]), .Z(n40484) );
  XOR U43833 ( .A(ein[757]), .B(n40485), .Z(ereg_next[758]) );
  AND U43834 ( .A(mul_pow), .B(n40486), .Z(n40485) );
  XOR U43835 ( .A(ein[758]), .B(ein[757]), .Z(n40486) );
  XOR U43836 ( .A(ein[756]), .B(n40487), .Z(ereg_next[757]) );
  AND U43837 ( .A(mul_pow), .B(n40488), .Z(n40487) );
  XOR U43838 ( .A(ein[757]), .B(ein[756]), .Z(n40488) );
  XOR U43839 ( .A(ein[755]), .B(n40489), .Z(ereg_next[756]) );
  AND U43840 ( .A(mul_pow), .B(n40490), .Z(n40489) );
  XOR U43841 ( .A(ein[756]), .B(ein[755]), .Z(n40490) );
  XOR U43842 ( .A(ein[754]), .B(n40491), .Z(ereg_next[755]) );
  AND U43843 ( .A(mul_pow), .B(n40492), .Z(n40491) );
  XOR U43844 ( .A(ein[755]), .B(ein[754]), .Z(n40492) );
  XOR U43845 ( .A(ein[753]), .B(n40493), .Z(ereg_next[754]) );
  AND U43846 ( .A(mul_pow), .B(n40494), .Z(n40493) );
  XOR U43847 ( .A(ein[754]), .B(ein[753]), .Z(n40494) );
  XOR U43848 ( .A(ein[752]), .B(n40495), .Z(ereg_next[753]) );
  AND U43849 ( .A(mul_pow), .B(n40496), .Z(n40495) );
  XOR U43850 ( .A(ein[753]), .B(ein[752]), .Z(n40496) );
  XOR U43851 ( .A(ein[751]), .B(n40497), .Z(ereg_next[752]) );
  AND U43852 ( .A(mul_pow), .B(n40498), .Z(n40497) );
  XOR U43853 ( .A(ein[752]), .B(ein[751]), .Z(n40498) );
  XOR U43854 ( .A(ein[750]), .B(n40499), .Z(ereg_next[751]) );
  AND U43855 ( .A(mul_pow), .B(n40500), .Z(n40499) );
  XOR U43856 ( .A(ein[751]), .B(ein[750]), .Z(n40500) );
  XOR U43857 ( .A(ein[749]), .B(n40501), .Z(ereg_next[750]) );
  AND U43858 ( .A(mul_pow), .B(n40502), .Z(n40501) );
  XOR U43859 ( .A(ein[750]), .B(ein[749]), .Z(n40502) );
  XOR U43860 ( .A(ein[73]), .B(n40503), .Z(ereg_next[74]) );
  AND U43861 ( .A(mul_pow), .B(n40504), .Z(n40503) );
  XOR U43862 ( .A(ein[74]), .B(ein[73]), .Z(n40504) );
  XOR U43863 ( .A(ein[748]), .B(n40505), .Z(ereg_next[749]) );
  AND U43864 ( .A(mul_pow), .B(n40506), .Z(n40505) );
  XOR U43865 ( .A(ein[749]), .B(ein[748]), .Z(n40506) );
  XOR U43866 ( .A(ein[747]), .B(n40507), .Z(ereg_next[748]) );
  AND U43867 ( .A(mul_pow), .B(n40508), .Z(n40507) );
  XOR U43868 ( .A(ein[748]), .B(ein[747]), .Z(n40508) );
  XOR U43869 ( .A(ein[746]), .B(n40509), .Z(ereg_next[747]) );
  AND U43870 ( .A(mul_pow), .B(n40510), .Z(n40509) );
  XOR U43871 ( .A(ein[747]), .B(ein[746]), .Z(n40510) );
  XOR U43872 ( .A(ein[745]), .B(n40511), .Z(ereg_next[746]) );
  AND U43873 ( .A(mul_pow), .B(n40512), .Z(n40511) );
  XOR U43874 ( .A(ein[746]), .B(ein[745]), .Z(n40512) );
  XOR U43875 ( .A(ein[744]), .B(n40513), .Z(ereg_next[745]) );
  AND U43876 ( .A(mul_pow), .B(n40514), .Z(n40513) );
  XOR U43877 ( .A(ein[745]), .B(ein[744]), .Z(n40514) );
  XOR U43878 ( .A(ein[743]), .B(n40515), .Z(ereg_next[744]) );
  AND U43879 ( .A(mul_pow), .B(n40516), .Z(n40515) );
  XOR U43880 ( .A(ein[744]), .B(ein[743]), .Z(n40516) );
  XOR U43881 ( .A(ein[742]), .B(n40517), .Z(ereg_next[743]) );
  AND U43882 ( .A(mul_pow), .B(n40518), .Z(n40517) );
  XOR U43883 ( .A(ein[743]), .B(ein[742]), .Z(n40518) );
  XOR U43884 ( .A(ein[741]), .B(n40519), .Z(ereg_next[742]) );
  AND U43885 ( .A(mul_pow), .B(n40520), .Z(n40519) );
  XOR U43886 ( .A(ein[742]), .B(ein[741]), .Z(n40520) );
  XOR U43887 ( .A(ein[740]), .B(n40521), .Z(ereg_next[741]) );
  AND U43888 ( .A(mul_pow), .B(n40522), .Z(n40521) );
  XOR U43889 ( .A(ein[741]), .B(ein[740]), .Z(n40522) );
  XOR U43890 ( .A(ein[739]), .B(n40523), .Z(ereg_next[740]) );
  AND U43891 ( .A(mul_pow), .B(n40524), .Z(n40523) );
  XOR U43892 ( .A(ein[740]), .B(ein[739]), .Z(n40524) );
  XOR U43893 ( .A(ein[72]), .B(n40525), .Z(ereg_next[73]) );
  AND U43894 ( .A(mul_pow), .B(n40526), .Z(n40525) );
  XOR U43895 ( .A(ein[73]), .B(ein[72]), .Z(n40526) );
  XOR U43896 ( .A(ein[738]), .B(n40527), .Z(ereg_next[739]) );
  AND U43897 ( .A(mul_pow), .B(n40528), .Z(n40527) );
  XOR U43898 ( .A(ein[739]), .B(ein[738]), .Z(n40528) );
  XOR U43899 ( .A(ein[737]), .B(n40529), .Z(ereg_next[738]) );
  AND U43900 ( .A(mul_pow), .B(n40530), .Z(n40529) );
  XOR U43901 ( .A(ein[738]), .B(ein[737]), .Z(n40530) );
  XOR U43902 ( .A(ein[736]), .B(n40531), .Z(ereg_next[737]) );
  AND U43903 ( .A(mul_pow), .B(n40532), .Z(n40531) );
  XOR U43904 ( .A(ein[737]), .B(ein[736]), .Z(n40532) );
  XOR U43905 ( .A(ein[735]), .B(n40533), .Z(ereg_next[736]) );
  AND U43906 ( .A(mul_pow), .B(n40534), .Z(n40533) );
  XOR U43907 ( .A(ein[736]), .B(ein[735]), .Z(n40534) );
  XOR U43908 ( .A(ein[734]), .B(n40535), .Z(ereg_next[735]) );
  AND U43909 ( .A(mul_pow), .B(n40536), .Z(n40535) );
  XOR U43910 ( .A(ein[735]), .B(ein[734]), .Z(n40536) );
  XOR U43911 ( .A(ein[733]), .B(n40537), .Z(ereg_next[734]) );
  AND U43912 ( .A(mul_pow), .B(n40538), .Z(n40537) );
  XOR U43913 ( .A(ein[734]), .B(ein[733]), .Z(n40538) );
  XOR U43914 ( .A(ein[732]), .B(n40539), .Z(ereg_next[733]) );
  AND U43915 ( .A(mul_pow), .B(n40540), .Z(n40539) );
  XOR U43916 ( .A(ein[733]), .B(ein[732]), .Z(n40540) );
  XOR U43917 ( .A(ein[731]), .B(n40541), .Z(ereg_next[732]) );
  AND U43918 ( .A(mul_pow), .B(n40542), .Z(n40541) );
  XOR U43919 ( .A(ein[732]), .B(ein[731]), .Z(n40542) );
  XOR U43920 ( .A(ein[730]), .B(n40543), .Z(ereg_next[731]) );
  AND U43921 ( .A(mul_pow), .B(n40544), .Z(n40543) );
  XOR U43922 ( .A(ein[731]), .B(ein[730]), .Z(n40544) );
  XOR U43923 ( .A(ein[729]), .B(n40545), .Z(ereg_next[730]) );
  AND U43924 ( .A(mul_pow), .B(n40546), .Z(n40545) );
  XOR U43925 ( .A(ein[730]), .B(ein[729]), .Z(n40546) );
  XOR U43926 ( .A(ein[71]), .B(n40547), .Z(ereg_next[72]) );
  AND U43927 ( .A(mul_pow), .B(n40548), .Z(n40547) );
  XOR U43928 ( .A(ein[72]), .B(ein[71]), .Z(n40548) );
  XOR U43929 ( .A(ein[728]), .B(n40549), .Z(ereg_next[729]) );
  AND U43930 ( .A(mul_pow), .B(n40550), .Z(n40549) );
  XOR U43931 ( .A(ein[729]), .B(ein[728]), .Z(n40550) );
  XOR U43932 ( .A(ein[727]), .B(n40551), .Z(ereg_next[728]) );
  AND U43933 ( .A(mul_pow), .B(n40552), .Z(n40551) );
  XOR U43934 ( .A(ein[728]), .B(ein[727]), .Z(n40552) );
  XOR U43935 ( .A(ein[726]), .B(n40553), .Z(ereg_next[727]) );
  AND U43936 ( .A(mul_pow), .B(n40554), .Z(n40553) );
  XOR U43937 ( .A(ein[727]), .B(ein[726]), .Z(n40554) );
  XOR U43938 ( .A(ein[725]), .B(n40555), .Z(ereg_next[726]) );
  AND U43939 ( .A(mul_pow), .B(n40556), .Z(n40555) );
  XOR U43940 ( .A(ein[726]), .B(ein[725]), .Z(n40556) );
  XOR U43941 ( .A(ein[724]), .B(n40557), .Z(ereg_next[725]) );
  AND U43942 ( .A(mul_pow), .B(n40558), .Z(n40557) );
  XOR U43943 ( .A(ein[725]), .B(ein[724]), .Z(n40558) );
  XOR U43944 ( .A(ein[723]), .B(n40559), .Z(ereg_next[724]) );
  AND U43945 ( .A(mul_pow), .B(n40560), .Z(n40559) );
  XOR U43946 ( .A(ein[724]), .B(ein[723]), .Z(n40560) );
  XOR U43947 ( .A(ein[722]), .B(n40561), .Z(ereg_next[723]) );
  AND U43948 ( .A(mul_pow), .B(n40562), .Z(n40561) );
  XOR U43949 ( .A(ein[723]), .B(ein[722]), .Z(n40562) );
  XOR U43950 ( .A(ein[721]), .B(n40563), .Z(ereg_next[722]) );
  AND U43951 ( .A(mul_pow), .B(n40564), .Z(n40563) );
  XOR U43952 ( .A(ein[722]), .B(ein[721]), .Z(n40564) );
  XOR U43953 ( .A(ein[720]), .B(n40565), .Z(ereg_next[721]) );
  AND U43954 ( .A(mul_pow), .B(n40566), .Z(n40565) );
  XOR U43955 ( .A(ein[721]), .B(ein[720]), .Z(n40566) );
  XOR U43956 ( .A(ein[719]), .B(n40567), .Z(ereg_next[720]) );
  AND U43957 ( .A(mul_pow), .B(n40568), .Z(n40567) );
  XOR U43958 ( .A(ein[720]), .B(ein[719]), .Z(n40568) );
  XOR U43959 ( .A(ein[70]), .B(n40569), .Z(ereg_next[71]) );
  AND U43960 ( .A(mul_pow), .B(n40570), .Z(n40569) );
  XOR U43961 ( .A(ein[71]), .B(ein[70]), .Z(n40570) );
  XOR U43962 ( .A(ein[718]), .B(n40571), .Z(ereg_next[719]) );
  AND U43963 ( .A(mul_pow), .B(n40572), .Z(n40571) );
  XOR U43964 ( .A(ein[719]), .B(ein[718]), .Z(n40572) );
  XOR U43965 ( .A(ein[717]), .B(n40573), .Z(ereg_next[718]) );
  AND U43966 ( .A(mul_pow), .B(n40574), .Z(n40573) );
  XOR U43967 ( .A(ein[718]), .B(ein[717]), .Z(n40574) );
  XOR U43968 ( .A(ein[716]), .B(n40575), .Z(ereg_next[717]) );
  AND U43969 ( .A(mul_pow), .B(n40576), .Z(n40575) );
  XOR U43970 ( .A(ein[717]), .B(ein[716]), .Z(n40576) );
  XOR U43971 ( .A(ein[715]), .B(n40577), .Z(ereg_next[716]) );
  AND U43972 ( .A(mul_pow), .B(n40578), .Z(n40577) );
  XOR U43973 ( .A(ein[716]), .B(ein[715]), .Z(n40578) );
  XOR U43974 ( .A(ein[714]), .B(n40579), .Z(ereg_next[715]) );
  AND U43975 ( .A(mul_pow), .B(n40580), .Z(n40579) );
  XOR U43976 ( .A(ein[715]), .B(ein[714]), .Z(n40580) );
  XOR U43977 ( .A(ein[713]), .B(n40581), .Z(ereg_next[714]) );
  AND U43978 ( .A(mul_pow), .B(n40582), .Z(n40581) );
  XOR U43979 ( .A(ein[714]), .B(ein[713]), .Z(n40582) );
  XOR U43980 ( .A(ein[712]), .B(n40583), .Z(ereg_next[713]) );
  AND U43981 ( .A(mul_pow), .B(n40584), .Z(n40583) );
  XOR U43982 ( .A(ein[713]), .B(ein[712]), .Z(n40584) );
  XOR U43983 ( .A(ein[711]), .B(n40585), .Z(ereg_next[712]) );
  AND U43984 ( .A(mul_pow), .B(n40586), .Z(n40585) );
  XOR U43985 ( .A(ein[712]), .B(ein[711]), .Z(n40586) );
  XOR U43986 ( .A(ein[710]), .B(n40587), .Z(ereg_next[711]) );
  AND U43987 ( .A(mul_pow), .B(n40588), .Z(n40587) );
  XOR U43988 ( .A(ein[711]), .B(ein[710]), .Z(n40588) );
  XOR U43989 ( .A(ein[709]), .B(n40589), .Z(ereg_next[710]) );
  AND U43990 ( .A(mul_pow), .B(n40590), .Z(n40589) );
  XOR U43991 ( .A(ein[710]), .B(ein[709]), .Z(n40590) );
  XOR U43992 ( .A(ein[69]), .B(n40591), .Z(ereg_next[70]) );
  AND U43993 ( .A(mul_pow), .B(n40592), .Z(n40591) );
  XOR U43994 ( .A(ein[70]), .B(ein[69]), .Z(n40592) );
  XOR U43995 ( .A(ein[708]), .B(n40593), .Z(ereg_next[709]) );
  AND U43996 ( .A(mul_pow), .B(n40594), .Z(n40593) );
  XOR U43997 ( .A(ein[709]), .B(ein[708]), .Z(n40594) );
  XOR U43998 ( .A(ein[707]), .B(n40595), .Z(ereg_next[708]) );
  AND U43999 ( .A(mul_pow), .B(n40596), .Z(n40595) );
  XOR U44000 ( .A(ein[708]), .B(ein[707]), .Z(n40596) );
  XOR U44001 ( .A(ein[706]), .B(n40597), .Z(ereg_next[707]) );
  AND U44002 ( .A(mul_pow), .B(n40598), .Z(n40597) );
  XOR U44003 ( .A(ein[707]), .B(ein[706]), .Z(n40598) );
  XOR U44004 ( .A(ein[705]), .B(n40599), .Z(ereg_next[706]) );
  AND U44005 ( .A(mul_pow), .B(n40600), .Z(n40599) );
  XOR U44006 ( .A(ein[706]), .B(ein[705]), .Z(n40600) );
  XOR U44007 ( .A(ein[704]), .B(n40601), .Z(ereg_next[705]) );
  AND U44008 ( .A(mul_pow), .B(n40602), .Z(n40601) );
  XOR U44009 ( .A(ein[705]), .B(ein[704]), .Z(n40602) );
  XOR U44010 ( .A(ein[703]), .B(n40603), .Z(ereg_next[704]) );
  AND U44011 ( .A(mul_pow), .B(n40604), .Z(n40603) );
  XOR U44012 ( .A(ein[704]), .B(ein[703]), .Z(n40604) );
  XOR U44013 ( .A(ein[702]), .B(n40605), .Z(ereg_next[703]) );
  AND U44014 ( .A(mul_pow), .B(n40606), .Z(n40605) );
  XOR U44015 ( .A(ein[703]), .B(ein[702]), .Z(n40606) );
  XOR U44016 ( .A(ein[701]), .B(n40607), .Z(ereg_next[702]) );
  AND U44017 ( .A(mul_pow), .B(n40608), .Z(n40607) );
  XOR U44018 ( .A(ein[702]), .B(ein[701]), .Z(n40608) );
  XOR U44019 ( .A(ein[700]), .B(n40609), .Z(ereg_next[701]) );
  AND U44020 ( .A(mul_pow), .B(n40610), .Z(n40609) );
  XOR U44021 ( .A(ein[701]), .B(ein[700]), .Z(n40610) );
  XOR U44022 ( .A(ein[699]), .B(n40611), .Z(ereg_next[700]) );
  AND U44023 ( .A(mul_pow), .B(n40612), .Z(n40611) );
  XOR U44024 ( .A(ein[700]), .B(ein[699]), .Z(n40612) );
  XOR U44025 ( .A(ein[5]), .B(n40613), .Z(ereg_next[6]) );
  AND U44026 ( .A(mul_pow), .B(n40614), .Z(n40613) );
  XOR U44027 ( .A(ein[6]), .B(ein[5]), .Z(n40614) );
  XOR U44028 ( .A(ein[68]), .B(n40615), .Z(ereg_next[69]) );
  AND U44029 ( .A(mul_pow), .B(n40616), .Z(n40615) );
  XOR U44030 ( .A(ein[69]), .B(ein[68]), .Z(n40616) );
  XOR U44031 ( .A(ein[698]), .B(n40617), .Z(ereg_next[699]) );
  AND U44032 ( .A(mul_pow), .B(n40618), .Z(n40617) );
  XOR U44033 ( .A(ein[699]), .B(ein[698]), .Z(n40618) );
  XOR U44034 ( .A(ein[697]), .B(n40619), .Z(ereg_next[698]) );
  AND U44035 ( .A(mul_pow), .B(n40620), .Z(n40619) );
  XOR U44036 ( .A(ein[698]), .B(ein[697]), .Z(n40620) );
  XOR U44037 ( .A(ein[696]), .B(n40621), .Z(ereg_next[697]) );
  AND U44038 ( .A(mul_pow), .B(n40622), .Z(n40621) );
  XOR U44039 ( .A(ein[697]), .B(ein[696]), .Z(n40622) );
  XOR U44040 ( .A(ein[695]), .B(n40623), .Z(ereg_next[696]) );
  AND U44041 ( .A(mul_pow), .B(n40624), .Z(n40623) );
  XOR U44042 ( .A(ein[696]), .B(ein[695]), .Z(n40624) );
  XOR U44043 ( .A(ein[694]), .B(n40625), .Z(ereg_next[695]) );
  AND U44044 ( .A(mul_pow), .B(n40626), .Z(n40625) );
  XOR U44045 ( .A(ein[695]), .B(ein[694]), .Z(n40626) );
  XOR U44046 ( .A(ein[693]), .B(n40627), .Z(ereg_next[694]) );
  AND U44047 ( .A(mul_pow), .B(n40628), .Z(n40627) );
  XOR U44048 ( .A(ein[694]), .B(ein[693]), .Z(n40628) );
  XOR U44049 ( .A(ein[692]), .B(n40629), .Z(ereg_next[693]) );
  AND U44050 ( .A(mul_pow), .B(n40630), .Z(n40629) );
  XOR U44051 ( .A(ein[693]), .B(ein[692]), .Z(n40630) );
  XOR U44052 ( .A(ein[691]), .B(n40631), .Z(ereg_next[692]) );
  AND U44053 ( .A(mul_pow), .B(n40632), .Z(n40631) );
  XOR U44054 ( .A(ein[692]), .B(ein[691]), .Z(n40632) );
  XOR U44055 ( .A(ein[690]), .B(n40633), .Z(ereg_next[691]) );
  AND U44056 ( .A(mul_pow), .B(n40634), .Z(n40633) );
  XOR U44057 ( .A(ein[691]), .B(ein[690]), .Z(n40634) );
  XOR U44058 ( .A(ein[689]), .B(n40635), .Z(ereg_next[690]) );
  AND U44059 ( .A(mul_pow), .B(n40636), .Z(n40635) );
  XOR U44060 ( .A(ein[690]), .B(ein[689]), .Z(n40636) );
  XOR U44061 ( .A(ein[67]), .B(n40637), .Z(ereg_next[68]) );
  AND U44062 ( .A(mul_pow), .B(n40638), .Z(n40637) );
  XOR U44063 ( .A(ein[68]), .B(ein[67]), .Z(n40638) );
  XOR U44064 ( .A(ein[688]), .B(n40639), .Z(ereg_next[689]) );
  AND U44065 ( .A(mul_pow), .B(n40640), .Z(n40639) );
  XOR U44066 ( .A(ein[689]), .B(ein[688]), .Z(n40640) );
  XOR U44067 ( .A(ein[687]), .B(n40641), .Z(ereg_next[688]) );
  AND U44068 ( .A(mul_pow), .B(n40642), .Z(n40641) );
  XOR U44069 ( .A(ein[688]), .B(ein[687]), .Z(n40642) );
  XOR U44070 ( .A(ein[686]), .B(n40643), .Z(ereg_next[687]) );
  AND U44071 ( .A(mul_pow), .B(n40644), .Z(n40643) );
  XOR U44072 ( .A(ein[687]), .B(ein[686]), .Z(n40644) );
  XOR U44073 ( .A(ein[685]), .B(n40645), .Z(ereg_next[686]) );
  AND U44074 ( .A(mul_pow), .B(n40646), .Z(n40645) );
  XOR U44075 ( .A(ein[686]), .B(ein[685]), .Z(n40646) );
  XOR U44076 ( .A(ein[684]), .B(n40647), .Z(ereg_next[685]) );
  AND U44077 ( .A(mul_pow), .B(n40648), .Z(n40647) );
  XOR U44078 ( .A(ein[685]), .B(ein[684]), .Z(n40648) );
  XOR U44079 ( .A(ein[683]), .B(n40649), .Z(ereg_next[684]) );
  AND U44080 ( .A(mul_pow), .B(n40650), .Z(n40649) );
  XOR U44081 ( .A(ein[684]), .B(ein[683]), .Z(n40650) );
  XOR U44082 ( .A(ein[682]), .B(n40651), .Z(ereg_next[683]) );
  AND U44083 ( .A(mul_pow), .B(n40652), .Z(n40651) );
  XOR U44084 ( .A(ein[683]), .B(ein[682]), .Z(n40652) );
  XOR U44085 ( .A(ein[681]), .B(n40653), .Z(ereg_next[682]) );
  AND U44086 ( .A(mul_pow), .B(n40654), .Z(n40653) );
  XOR U44087 ( .A(ein[682]), .B(ein[681]), .Z(n40654) );
  XOR U44088 ( .A(ein[680]), .B(n40655), .Z(ereg_next[681]) );
  AND U44089 ( .A(mul_pow), .B(n40656), .Z(n40655) );
  XOR U44090 ( .A(ein[681]), .B(ein[680]), .Z(n40656) );
  XOR U44091 ( .A(ein[679]), .B(n40657), .Z(ereg_next[680]) );
  AND U44092 ( .A(mul_pow), .B(n40658), .Z(n40657) );
  XOR U44093 ( .A(ein[680]), .B(ein[679]), .Z(n40658) );
  XOR U44094 ( .A(ein[66]), .B(n40659), .Z(ereg_next[67]) );
  AND U44095 ( .A(mul_pow), .B(n40660), .Z(n40659) );
  XOR U44096 ( .A(ein[67]), .B(ein[66]), .Z(n40660) );
  XOR U44097 ( .A(ein[678]), .B(n40661), .Z(ereg_next[679]) );
  AND U44098 ( .A(mul_pow), .B(n40662), .Z(n40661) );
  XOR U44099 ( .A(ein[679]), .B(ein[678]), .Z(n40662) );
  XOR U44100 ( .A(ein[677]), .B(n40663), .Z(ereg_next[678]) );
  AND U44101 ( .A(mul_pow), .B(n40664), .Z(n40663) );
  XOR U44102 ( .A(ein[678]), .B(ein[677]), .Z(n40664) );
  XOR U44103 ( .A(ein[676]), .B(n40665), .Z(ereg_next[677]) );
  AND U44104 ( .A(mul_pow), .B(n40666), .Z(n40665) );
  XOR U44105 ( .A(ein[677]), .B(ein[676]), .Z(n40666) );
  XOR U44106 ( .A(ein[675]), .B(n40667), .Z(ereg_next[676]) );
  AND U44107 ( .A(mul_pow), .B(n40668), .Z(n40667) );
  XOR U44108 ( .A(ein[676]), .B(ein[675]), .Z(n40668) );
  XOR U44109 ( .A(ein[674]), .B(n40669), .Z(ereg_next[675]) );
  AND U44110 ( .A(mul_pow), .B(n40670), .Z(n40669) );
  XOR U44111 ( .A(ein[675]), .B(ein[674]), .Z(n40670) );
  XOR U44112 ( .A(ein[673]), .B(n40671), .Z(ereg_next[674]) );
  AND U44113 ( .A(mul_pow), .B(n40672), .Z(n40671) );
  XOR U44114 ( .A(ein[674]), .B(ein[673]), .Z(n40672) );
  XOR U44115 ( .A(ein[672]), .B(n40673), .Z(ereg_next[673]) );
  AND U44116 ( .A(mul_pow), .B(n40674), .Z(n40673) );
  XOR U44117 ( .A(ein[673]), .B(ein[672]), .Z(n40674) );
  XOR U44118 ( .A(ein[671]), .B(n40675), .Z(ereg_next[672]) );
  AND U44119 ( .A(mul_pow), .B(n40676), .Z(n40675) );
  XOR U44120 ( .A(ein[672]), .B(ein[671]), .Z(n40676) );
  XOR U44121 ( .A(ein[670]), .B(n40677), .Z(ereg_next[671]) );
  AND U44122 ( .A(mul_pow), .B(n40678), .Z(n40677) );
  XOR U44123 ( .A(ein[671]), .B(ein[670]), .Z(n40678) );
  XOR U44124 ( .A(ein[669]), .B(n40679), .Z(ereg_next[670]) );
  AND U44125 ( .A(mul_pow), .B(n40680), .Z(n40679) );
  XOR U44126 ( .A(ein[670]), .B(ein[669]), .Z(n40680) );
  XOR U44127 ( .A(ein[65]), .B(n40681), .Z(ereg_next[66]) );
  AND U44128 ( .A(mul_pow), .B(n40682), .Z(n40681) );
  XOR U44129 ( .A(ein[66]), .B(ein[65]), .Z(n40682) );
  XOR U44130 ( .A(ein[668]), .B(n40683), .Z(ereg_next[669]) );
  AND U44131 ( .A(mul_pow), .B(n40684), .Z(n40683) );
  XOR U44132 ( .A(ein[669]), .B(ein[668]), .Z(n40684) );
  XOR U44133 ( .A(ein[667]), .B(n40685), .Z(ereg_next[668]) );
  AND U44134 ( .A(mul_pow), .B(n40686), .Z(n40685) );
  XOR U44135 ( .A(ein[668]), .B(ein[667]), .Z(n40686) );
  XOR U44136 ( .A(ein[666]), .B(n40687), .Z(ereg_next[667]) );
  AND U44137 ( .A(mul_pow), .B(n40688), .Z(n40687) );
  XOR U44138 ( .A(ein[667]), .B(ein[666]), .Z(n40688) );
  XOR U44139 ( .A(ein[665]), .B(n40689), .Z(ereg_next[666]) );
  AND U44140 ( .A(mul_pow), .B(n40690), .Z(n40689) );
  XOR U44141 ( .A(ein[666]), .B(ein[665]), .Z(n40690) );
  XOR U44142 ( .A(ein[664]), .B(n40691), .Z(ereg_next[665]) );
  AND U44143 ( .A(mul_pow), .B(n40692), .Z(n40691) );
  XOR U44144 ( .A(ein[665]), .B(ein[664]), .Z(n40692) );
  XOR U44145 ( .A(ein[663]), .B(n40693), .Z(ereg_next[664]) );
  AND U44146 ( .A(mul_pow), .B(n40694), .Z(n40693) );
  XOR U44147 ( .A(ein[664]), .B(ein[663]), .Z(n40694) );
  XOR U44148 ( .A(ein[662]), .B(n40695), .Z(ereg_next[663]) );
  AND U44149 ( .A(mul_pow), .B(n40696), .Z(n40695) );
  XOR U44150 ( .A(ein[663]), .B(ein[662]), .Z(n40696) );
  XOR U44151 ( .A(ein[661]), .B(n40697), .Z(ereg_next[662]) );
  AND U44152 ( .A(mul_pow), .B(n40698), .Z(n40697) );
  XOR U44153 ( .A(ein[662]), .B(ein[661]), .Z(n40698) );
  XOR U44154 ( .A(ein[660]), .B(n40699), .Z(ereg_next[661]) );
  AND U44155 ( .A(mul_pow), .B(n40700), .Z(n40699) );
  XOR U44156 ( .A(ein[661]), .B(ein[660]), .Z(n40700) );
  XOR U44157 ( .A(ein[659]), .B(n40701), .Z(ereg_next[660]) );
  AND U44158 ( .A(mul_pow), .B(n40702), .Z(n40701) );
  XOR U44159 ( .A(ein[660]), .B(ein[659]), .Z(n40702) );
  XOR U44160 ( .A(ein[64]), .B(n40703), .Z(ereg_next[65]) );
  AND U44161 ( .A(mul_pow), .B(n40704), .Z(n40703) );
  XOR U44162 ( .A(ein[65]), .B(ein[64]), .Z(n40704) );
  XOR U44163 ( .A(ein[658]), .B(n40705), .Z(ereg_next[659]) );
  AND U44164 ( .A(mul_pow), .B(n40706), .Z(n40705) );
  XOR U44165 ( .A(ein[659]), .B(ein[658]), .Z(n40706) );
  XOR U44166 ( .A(ein[657]), .B(n40707), .Z(ereg_next[658]) );
  AND U44167 ( .A(mul_pow), .B(n40708), .Z(n40707) );
  XOR U44168 ( .A(ein[658]), .B(ein[657]), .Z(n40708) );
  XOR U44169 ( .A(ein[656]), .B(n40709), .Z(ereg_next[657]) );
  AND U44170 ( .A(mul_pow), .B(n40710), .Z(n40709) );
  XOR U44171 ( .A(ein[657]), .B(ein[656]), .Z(n40710) );
  XOR U44172 ( .A(ein[655]), .B(n40711), .Z(ereg_next[656]) );
  AND U44173 ( .A(mul_pow), .B(n40712), .Z(n40711) );
  XOR U44174 ( .A(ein[656]), .B(ein[655]), .Z(n40712) );
  XOR U44175 ( .A(ein[654]), .B(n40713), .Z(ereg_next[655]) );
  AND U44176 ( .A(mul_pow), .B(n40714), .Z(n40713) );
  XOR U44177 ( .A(ein[655]), .B(ein[654]), .Z(n40714) );
  XOR U44178 ( .A(ein[653]), .B(n40715), .Z(ereg_next[654]) );
  AND U44179 ( .A(mul_pow), .B(n40716), .Z(n40715) );
  XOR U44180 ( .A(ein[654]), .B(ein[653]), .Z(n40716) );
  XOR U44181 ( .A(ein[652]), .B(n40717), .Z(ereg_next[653]) );
  AND U44182 ( .A(mul_pow), .B(n40718), .Z(n40717) );
  XOR U44183 ( .A(ein[653]), .B(ein[652]), .Z(n40718) );
  XOR U44184 ( .A(ein[651]), .B(n40719), .Z(ereg_next[652]) );
  AND U44185 ( .A(mul_pow), .B(n40720), .Z(n40719) );
  XOR U44186 ( .A(ein[652]), .B(ein[651]), .Z(n40720) );
  XOR U44187 ( .A(ein[650]), .B(n40721), .Z(ereg_next[651]) );
  AND U44188 ( .A(mul_pow), .B(n40722), .Z(n40721) );
  XOR U44189 ( .A(ein[651]), .B(ein[650]), .Z(n40722) );
  XOR U44190 ( .A(ein[649]), .B(n40723), .Z(ereg_next[650]) );
  AND U44191 ( .A(mul_pow), .B(n40724), .Z(n40723) );
  XOR U44192 ( .A(ein[650]), .B(ein[649]), .Z(n40724) );
  XOR U44193 ( .A(ein[63]), .B(n40725), .Z(ereg_next[64]) );
  AND U44194 ( .A(mul_pow), .B(n40726), .Z(n40725) );
  XOR U44195 ( .A(ein[64]), .B(ein[63]), .Z(n40726) );
  XOR U44196 ( .A(ein[648]), .B(n40727), .Z(ereg_next[649]) );
  AND U44197 ( .A(mul_pow), .B(n40728), .Z(n40727) );
  XOR U44198 ( .A(ein[649]), .B(ein[648]), .Z(n40728) );
  XOR U44199 ( .A(ein[647]), .B(n40729), .Z(ereg_next[648]) );
  AND U44200 ( .A(mul_pow), .B(n40730), .Z(n40729) );
  XOR U44201 ( .A(ein[648]), .B(ein[647]), .Z(n40730) );
  XOR U44202 ( .A(ein[646]), .B(n40731), .Z(ereg_next[647]) );
  AND U44203 ( .A(mul_pow), .B(n40732), .Z(n40731) );
  XOR U44204 ( .A(ein[647]), .B(ein[646]), .Z(n40732) );
  XOR U44205 ( .A(ein[645]), .B(n40733), .Z(ereg_next[646]) );
  AND U44206 ( .A(mul_pow), .B(n40734), .Z(n40733) );
  XOR U44207 ( .A(ein[646]), .B(ein[645]), .Z(n40734) );
  XOR U44208 ( .A(ein[644]), .B(n40735), .Z(ereg_next[645]) );
  AND U44209 ( .A(mul_pow), .B(n40736), .Z(n40735) );
  XOR U44210 ( .A(ein[645]), .B(ein[644]), .Z(n40736) );
  XOR U44211 ( .A(ein[643]), .B(n40737), .Z(ereg_next[644]) );
  AND U44212 ( .A(mul_pow), .B(n40738), .Z(n40737) );
  XOR U44213 ( .A(ein[644]), .B(ein[643]), .Z(n40738) );
  XOR U44214 ( .A(ein[642]), .B(n40739), .Z(ereg_next[643]) );
  AND U44215 ( .A(mul_pow), .B(n40740), .Z(n40739) );
  XOR U44216 ( .A(ein[643]), .B(ein[642]), .Z(n40740) );
  XOR U44217 ( .A(ein[641]), .B(n40741), .Z(ereg_next[642]) );
  AND U44218 ( .A(mul_pow), .B(n40742), .Z(n40741) );
  XOR U44219 ( .A(ein[642]), .B(ein[641]), .Z(n40742) );
  XOR U44220 ( .A(ein[640]), .B(n40743), .Z(ereg_next[641]) );
  AND U44221 ( .A(mul_pow), .B(n40744), .Z(n40743) );
  XOR U44222 ( .A(ein[641]), .B(ein[640]), .Z(n40744) );
  XOR U44223 ( .A(ein[639]), .B(n40745), .Z(ereg_next[640]) );
  AND U44224 ( .A(mul_pow), .B(n40746), .Z(n40745) );
  XOR U44225 ( .A(ein[640]), .B(ein[639]), .Z(n40746) );
  XOR U44226 ( .A(ein[62]), .B(n40747), .Z(ereg_next[63]) );
  AND U44227 ( .A(mul_pow), .B(n40748), .Z(n40747) );
  XOR U44228 ( .A(ein[63]), .B(ein[62]), .Z(n40748) );
  XOR U44229 ( .A(ein[638]), .B(n40749), .Z(ereg_next[639]) );
  AND U44230 ( .A(mul_pow), .B(n40750), .Z(n40749) );
  XOR U44231 ( .A(ein[639]), .B(ein[638]), .Z(n40750) );
  XOR U44232 ( .A(ein[637]), .B(n40751), .Z(ereg_next[638]) );
  AND U44233 ( .A(mul_pow), .B(n40752), .Z(n40751) );
  XOR U44234 ( .A(ein[638]), .B(ein[637]), .Z(n40752) );
  XOR U44235 ( .A(ein[636]), .B(n40753), .Z(ereg_next[637]) );
  AND U44236 ( .A(mul_pow), .B(n40754), .Z(n40753) );
  XOR U44237 ( .A(ein[637]), .B(ein[636]), .Z(n40754) );
  XOR U44238 ( .A(ein[635]), .B(n40755), .Z(ereg_next[636]) );
  AND U44239 ( .A(mul_pow), .B(n40756), .Z(n40755) );
  XOR U44240 ( .A(ein[636]), .B(ein[635]), .Z(n40756) );
  XOR U44241 ( .A(ein[634]), .B(n40757), .Z(ereg_next[635]) );
  AND U44242 ( .A(mul_pow), .B(n40758), .Z(n40757) );
  XOR U44243 ( .A(ein[635]), .B(ein[634]), .Z(n40758) );
  XOR U44244 ( .A(ein[633]), .B(n40759), .Z(ereg_next[634]) );
  AND U44245 ( .A(mul_pow), .B(n40760), .Z(n40759) );
  XOR U44246 ( .A(ein[634]), .B(ein[633]), .Z(n40760) );
  XOR U44247 ( .A(ein[632]), .B(n40761), .Z(ereg_next[633]) );
  AND U44248 ( .A(mul_pow), .B(n40762), .Z(n40761) );
  XOR U44249 ( .A(ein[633]), .B(ein[632]), .Z(n40762) );
  XOR U44250 ( .A(ein[631]), .B(n40763), .Z(ereg_next[632]) );
  AND U44251 ( .A(mul_pow), .B(n40764), .Z(n40763) );
  XOR U44252 ( .A(ein[632]), .B(ein[631]), .Z(n40764) );
  XOR U44253 ( .A(ein[630]), .B(n40765), .Z(ereg_next[631]) );
  AND U44254 ( .A(mul_pow), .B(n40766), .Z(n40765) );
  XOR U44255 ( .A(ein[631]), .B(ein[630]), .Z(n40766) );
  XOR U44256 ( .A(ein[629]), .B(n40767), .Z(ereg_next[630]) );
  AND U44257 ( .A(mul_pow), .B(n40768), .Z(n40767) );
  XOR U44258 ( .A(ein[630]), .B(ein[629]), .Z(n40768) );
  XOR U44259 ( .A(ein[61]), .B(n40769), .Z(ereg_next[62]) );
  AND U44260 ( .A(mul_pow), .B(n40770), .Z(n40769) );
  XOR U44261 ( .A(ein[62]), .B(ein[61]), .Z(n40770) );
  XOR U44262 ( .A(ein[628]), .B(n40771), .Z(ereg_next[629]) );
  AND U44263 ( .A(mul_pow), .B(n40772), .Z(n40771) );
  XOR U44264 ( .A(ein[629]), .B(ein[628]), .Z(n40772) );
  XOR U44265 ( .A(ein[627]), .B(n40773), .Z(ereg_next[628]) );
  AND U44266 ( .A(mul_pow), .B(n40774), .Z(n40773) );
  XOR U44267 ( .A(ein[628]), .B(ein[627]), .Z(n40774) );
  XOR U44268 ( .A(ein[626]), .B(n40775), .Z(ereg_next[627]) );
  AND U44269 ( .A(mul_pow), .B(n40776), .Z(n40775) );
  XOR U44270 ( .A(ein[627]), .B(ein[626]), .Z(n40776) );
  XOR U44271 ( .A(ein[625]), .B(n40777), .Z(ereg_next[626]) );
  AND U44272 ( .A(mul_pow), .B(n40778), .Z(n40777) );
  XOR U44273 ( .A(ein[626]), .B(ein[625]), .Z(n40778) );
  XOR U44274 ( .A(ein[624]), .B(n40779), .Z(ereg_next[625]) );
  AND U44275 ( .A(mul_pow), .B(n40780), .Z(n40779) );
  XOR U44276 ( .A(ein[625]), .B(ein[624]), .Z(n40780) );
  XOR U44277 ( .A(ein[623]), .B(n40781), .Z(ereg_next[624]) );
  AND U44278 ( .A(mul_pow), .B(n40782), .Z(n40781) );
  XOR U44279 ( .A(ein[624]), .B(ein[623]), .Z(n40782) );
  XOR U44280 ( .A(ein[622]), .B(n40783), .Z(ereg_next[623]) );
  AND U44281 ( .A(mul_pow), .B(n40784), .Z(n40783) );
  XOR U44282 ( .A(ein[623]), .B(ein[622]), .Z(n40784) );
  XOR U44283 ( .A(ein[621]), .B(n40785), .Z(ereg_next[622]) );
  AND U44284 ( .A(mul_pow), .B(n40786), .Z(n40785) );
  XOR U44285 ( .A(ein[622]), .B(ein[621]), .Z(n40786) );
  XOR U44286 ( .A(ein[620]), .B(n40787), .Z(ereg_next[621]) );
  AND U44287 ( .A(mul_pow), .B(n40788), .Z(n40787) );
  XOR U44288 ( .A(ein[621]), .B(ein[620]), .Z(n40788) );
  XOR U44289 ( .A(ein[619]), .B(n40789), .Z(ereg_next[620]) );
  AND U44290 ( .A(mul_pow), .B(n40790), .Z(n40789) );
  XOR U44291 ( .A(ein[620]), .B(ein[619]), .Z(n40790) );
  XOR U44292 ( .A(ein[60]), .B(n40791), .Z(ereg_next[61]) );
  AND U44293 ( .A(mul_pow), .B(n40792), .Z(n40791) );
  XOR U44294 ( .A(ein[61]), .B(ein[60]), .Z(n40792) );
  XOR U44295 ( .A(ein[618]), .B(n40793), .Z(ereg_next[619]) );
  AND U44296 ( .A(mul_pow), .B(n40794), .Z(n40793) );
  XOR U44297 ( .A(ein[619]), .B(ein[618]), .Z(n40794) );
  XOR U44298 ( .A(ein[617]), .B(n40795), .Z(ereg_next[618]) );
  AND U44299 ( .A(mul_pow), .B(n40796), .Z(n40795) );
  XOR U44300 ( .A(ein[618]), .B(ein[617]), .Z(n40796) );
  XOR U44301 ( .A(ein[616]), .B(n40797), .Z(ereg_next[617]) );
  AND U44302 ( .A(mul_pow), .B(n40798), .Z(n40797) );
  XOR U44303 ( .A(ein[617]), .B(ein[616]), .Z(n40798) );
  XOR U44304 ( .A(ein[615]), .B(n40799), .Z(ereg_next[616]) );
  AND U44305 ( .A(mul_pow), .B(n40800), .Z(n40799) );
  XOR U44306 ( .A(ein[616]), .B(ein[615]), .Z(n40800) );
  XOR U44307 ( .A(ein[614]), .B(n40801), .Z(ereg_next[615]) );
  AND U44308 ( .A(mul_pow), .B(n40802), .Z(n40801) );
  XOR U44309 ( .A(ein[615]), .B(ein[614]), .Z(n40802) );
  XOR U44310 ( .A(ein[613]), .B(n40803), .Z(ereg_next[614]) );
  AND U44311 ( .A(mul_pow), .B(n40804), .Z(n40803) );
  XOR U44312 ( .A(ein[614]), .B(ein[613]), .Z(n40804) );
  XOR U44313 ( .A(ein[612]), .B(n40805), .Z(ereg_next[613]) );
  AND U44314 ( .A(mul_pow), .B(n40806), .Z(n40805) );
  XOR U44315 ( .A(ein[613]), .B(ein[612]), .Z(n40806) );
  XOR U44316 ( .A(ein[611]), .B(n40807), .Z(ereg_next[612]) );
  AND U44317 ( .A(mul_pow), .B(n40808), .Z(n40807) );
  XOR U44318 ( .A(ein[612]), .B(ein[611]), .Z(n40808) );
  XOR U44319 ( .A(ein[610]), .B(n40809), .Z(ereg_next[611]) );
  AND U44320 ( .A(mul_pow), .B(n40810), .Z(n40809) );
  XOR U44321 ( .A(ein[611]), .B(ein[610]), .Z(n40810) );
  XOR U44322 ( .A(ein[609]), .B(n40811), .Z(ereg_next[610]) );
  AND U44323 ( .A(mul_pow), .B(n40812), .Z(n40811) );
  XOR U44324 ( .A(ein[610]), .B(ein[609]), .Z(n40812) );
  XOR U44325 ( .A(ein[59]), .B(n40813), .Z(ereg_next[60]) );
  AND U44326 ( .A(mul_pow), .B(n40814), .Z(n40813) );
  XOR U44327 ( .A(ein[60]), .B(ein[59]), .Z(n40814) );
  XOR U44328 ( .A(ein[608]), .B(n40815), .Z(ereg_next[609]) );
  AND U44329 ( .A(mul_pow), .B(n40816), .Z(n40815) );
  XOR U44330 ( .A(ein[609]), .B(ein[608]), .Z(n40816) );
  XOR U44331 ( .A(ein[607]), .B(n40817), .Z(ereg_next[608]) );
  AND U44332 ( .A(mul_pow), .B(n40818), .Z(n40817) );
  XOR U44333 ( .A(ein[608]), .B(ein[607]), .Z(n40818) );
  XOR U44334 ( .A(ein[606]), .B(n40819), .Z(ereg_next[607]) );
  AND U44335 ( .A(mul_pow), .B(n40820), .Z(n40819) );
  XOR U44336 ( .A(ein[607]), .B(ein[606]), .Z(n40820) );
  XOR U44337 ( .A(ein[605]), .B(n40821), .Z(ereg_next[606]) );
  AND U44338 ( .A(mul_pow), .B(n40822), .Z(n40821) );
  XOR U44339 ( .A(ein[606]), .B(ein[605]), .Z(n40822) );
  XOR U44340 ( .A(ein[604]), .B(n40823), .Z(ereg_next[605]) );
  AND U44341 ( .A(mul_pow), .B(n40824), .Z(n40823) );
  XOR U44342 ( .A(ein[605]), .B(ein[604]), .Z(n40824) );
  XOR U44343 ( .A(ein[603]), .B(n40825), .Z(ereg_next[604]) );
  AND U44344 ( .A(mul_pow), .B(n40826), .Z(n40825) );
  XOR U44345 ( .A(ein[604]), .B(ein[603]), .Z(n40826) );
  XOR U44346 ( .A(ein[602]), .B(n40827), .Z(ereg_next[603]) );
  AND U44347 ( .A(mul_pow), .B(n40828), .Z(n40827) );
  XOR U44348 ( .A(ein[603]), .B(ein[602]), .Z(n40828) );
  XOR U44349 ( .A(ein[601]), .B(n40829), .Z(ereg_next[602]) );
  AND U44350 ( .A(mul_pow), .B(n40830), .Z(n40829) );
  XOR U44351 ( .A(ein[602]), .B(ein[601]), .Z(n40830) );
  XOR U44352 ( .A(ein[600]), .B(n40831), .Z(ereg_next[601]) );
  AND U44353 ( .A(mul_pow), .B(n40832), .Z(n40831) );
  XOR U44354 ( .A(ein[601]), .B(ein[600]), .Z(n40832) );
  XOR U44355 ( .A(ein[599]), .B(n40833), .Z(ereg_next[600]) );
  AND U44356 ( .A(mul_pow), .B(n40834), .Z(n40833) );
  XOR U44357 ( .A(ein[600]), .B(ein[599]), .Z(n40834) );
  XOR U44358 ( .A(ein[4]), .B(n40835), .Z(ereg_next[5]) );
  AND U44359 ( .A(mul_pow), .B(n40836), .Z(n40835) );
  XOR U44360 ( .A(ein[5]), .B(ein[4]), .Z(n40836) );
  XOR U44361 ( .A(ein[58]), .B(n40837), .Z(ereg_next[59]) );
  AND U44362 ( .A(mul_pow), .B(n40838), .Z(n40837) );
  XOR U44363 ( .A(ein[59]), .B(ein[58]), .Z(n40838) );
  XOR U44364 ( .A(ein[598]), .B(n40839), .Z(ereg_next[599]) );
  AND U44365 ( .A(mul_pow), .B(n40840), .Z(n40839) );
  XOR U44366 ( .A(ein[599]), .B(ein[598]), .Z(n40840) );
  XOR U44367 ( .A(ein[597]), .B(n40841), .Z(ereg_next[598]) );
  AND U44368 ( .A(mul_pow), .B(n40842), .Z(n40841) );
  XOR U44369 ( .A(ein[598]), .B(ein[597]), .Z(n40842) );
  XOR U44370 ( .A(ein[596]), .B(n40843), .Z(ereg_next[597]) );
  AND U44371 ( .A(mul_pow), .B(n40844), .Z(n40843) );
  XOR U44372 ( .A(ein[597]), .B(ein[596]), .Z(n40844) );
  XOR U44373 ( .A(ein[595]), .B(n40845), .Z(ereg_next[596]) );
  AND U44374 ( .A(mul_pow), .B(n40846), .Z(n40845) );
  XOR U44375 ( .A(ein[596]), .B(ein[595]), .Z(n40846) );
  XOR U44376 ( .A(ein[594]), .B(n40847), .Z(ereg_next[595]) );
  AND U44377 ( .A(mul_pow), .B(n40848), .Z(n40847) );
  XOR U44378 ( .A(ein[595]), .B(ein[594]), .Z(n40848) );
  XOR U44379 ( .A(ein[593]), .B(n40849), .Z(ereg_next[594]) );
  AND U44380 ( .A(mul_pow), .B(n40850), .Z(n40849) );
  XOR U44381 ( .A(ein[594]), .B(ein[593]), .Z(n40850) );
  XOR U44382 ( .A(ein[592]), .B(n40851), .Z(ereg_next[593]) );
  AND U44383 ( .A(mul_pow), .B(n40852), .Z(n40851) );
  XOR U44384 ( .A(ein[593]), .B(ein[592]), .Z(n40852) );
  XOR U44385 ( .A(ein[591]), .B(n40853), .Z(ereg_next[592]) );
  AND U44386 ( .A(mul_pow), .B(n40854), .Z(n40853) );
  XOR U44387 ( .A(ein[592]), .B(ein[591]), .Z(n40854) );
  XOR U44388 ( .A(ein[590]), .B(n40855), .Z(ereg_next[591]) );
  AND U44389 ( .A(mul_pow), .B(n40856), .Z(n40855) );
  XOR U44390 ( .A(ein[591]), .B(ein[590]), .Z(n40856) );
  XOR U44391 ( .A(ein[589]), .B(n40857), .Z(ereg_next[590]) );
  AND U44392 ( .A(mul_pow), .B(n40858), .Z(n40857) );
  XOR U44393 ( .A(ein[590]), .B(ein[589]), .Z(n40858) );
  XOR U44394 ( .A(ein[57]), .B(n40859), .Z(ereg_next[58]) );
  AND U44395 ( .A(mul_pow), .B(n40860), .Z(n40859) );
  XOR U44396 ( .A(ein[58]), .B(ein[57]), .Z(n40860) );
  XOR U44397 ( .A(ein[588]), .B(n40861), .Z(ereg_next[589]) );
  AND U44398 ( .A(mul_pow), .B(n40862), .Z(n40861) );
  XOR U44399 ( .A(ein[589]), .B(ein[588]), .Z(n40862) );
  XOR U44400 ( .A(ein[587]), .B(n40863), .Z(ereg_next[588]) );
  AND U44401 ( .A(mul_pow), .B(n40864), .Z(n40863) );
  XOR U44402 ( .A(ein[588]), .B(ein[587]), .Z(n40864) );
  XOR U44403 ( .A(ein[586]), .B(n40865), .Z(ereg_next[587]) );
  AND U44404 ( .A(mul_pow), .B(n40866), .Z(n40865) );
  XOR U44405 ( .A(ein[587]), .B(ein[586]), .Z(n40866) );
  XOR U44406 ( .A(ein[585]), .B(n40867), .Z(ereg_next[586]) );
  AND U44407 ( .A(mul_pow), .B(n40868), .Z(n40867) );
  XOR U44408 ( .A(ein[586]), .B(ein[585]), .Z(n40868) );
  XOR U44409 ( .A(ein[584]), .B(n40869), .Z(ereg_next[585]) );
  AND U44410 ( .A(mul_pow), .B(n40870), .Z(n40869) );
  XOR U44411 ( .A(ein[585]), .B(ein[584]), .Z(n40870) );
  XOR U44412 ( .A(ein[583]), .B(n40871), .Z(ereg_next[584]) );
  AND U44413 ( .A(mul_pow), .B(n40872), .Z(n40871) );
  XOR U44414 ( .A(ein[584]), .B(ein[583]), .Z(n40872) );
  XOR U44415 ( .A(ein[582]), .B(n40873), .Z(ereg_next[583]) );
  AND U44416 ( .A(mul_pow), .B(n40874), .Z(n40873) );
  XOR U44417 ( .A(ein[583]), .B(ein[582]), .Z(n40874) );
  XOR U44418 ( .A(ein[581]), .B(n40875), .Z(ereg_next[582]) );
  AND U44419 ( .A(mul_pow), .B(n40876), .Z(n40875) );
  XOR U44420 ( .A(ein[582]), .B(ein[581]), .Z(n40876) );
  XOR U44421 ( .A(ein[580]), .B(n40877), .Z(ereg_next[581]) );
  AND U44422 ( .A(mul_pow), .B(n40878), .Z(n40877) );
  XOR U44423 ( .A(ein[581]), .B(ein[580]), .Z(n40878) );
  XOR U44424 ( .A(ein[579]), .B(n40879), .Z(ereg_next[580]) );
  AND U44425 ( .A(mul_pow), .B(n40880), .Z(n40879) );
  XOR U44426 ( .A(ein[580]), .B(ein[579]), .Z(n40880) );
  XOR U44427 ( .A(ein[56]), .B(n40881), .Z(ereg_next[57]) );
  AND U44428 ( .A(mul_pow), .B(n40882), .Z(n40881) );
  XOR U44429 ( .A(ein[57]), .B(ein[56]), .Z(n40882) );
  XOR U44430 ( .A(ein[578]), .B(n40883), .Z(ereg_next[579]) );
  AND U44431 ( .A(mul_pow), .B(n40884), .Z(n40883) );
  XOR U44432 ( .A(ein[579]), .B(ein[578]), .Z(n40884) );
  XOR U44433 ( .A(ein[577]), .B(n40885), .Z(ereg_next[578]) );
  AND U44434 ( .A(mul_pow), .B(n40886), .Z(n40885) );
  XOR U44435 ( .A(ein[578]), .B(ein[577]), .Z(n40886) );
  XOR U44436 ( .A(ein[576]), .B(n40887), .Z(ereg_next[577]) );
  AND U44437 ( .A(mul_pow), .B(n40888), .Z(n40887) );
  XOR U44438 ( .A(ein[577]), .B(ein[576]), .Z(n40888) );
  XOR U44439 ( .A(ein[575]), .B(n40889), .Z(ereg_next[576]) );
  AND U44440 ( .A(mul_pow), .B(n40890), .Z(n40889) );
  XOR U44441 ( .A(ein[576]), .B(ein[575]), .Z(n40890) );
  XOR U44442 ( .A(ein[574]), .B(n40891), .Z(ereg_next[575]) );
  AND U44443 ( .A(mul_pow), .B(n40892), .Z(n40891) );
  XOR U44444 ( .A(ein[575]), .B(ein[574]), .Z(n40892) );
  XOR U44445 ( .A(ein[573]), .B(n40893), .Z(ereg_next[574]) );
  AND U44446 ( .A(mul_pow), .B(n40894), .Z(n40893) );
  XOR U44447 ( .A(ein[574]), .B(ein[573]), .Z(n40894) );
  XOR U44448 ( .A(ein[572]), .B(n40895), .Z(ereg_next[573]) );
  AND U44449 ( .A(mul_pow), .B(n40896), .Z(n40895) );
  XOR U44450 ( .A(ein[573]), .B(ein[572]), .Z(n40896) );
  XOR U44451 ( .A(ein[571]), .B(n40897), .Z(ereg_next[572]) );
  AND U44452 ( .A(mul_pow), .B(n40898), .Z(n40897) );
  XOR U44453 ( .A(ein[572]), .B(ein[571]), .Z(n40898) );
  XOR U44454 ( .A(ein[570]), .B(n40899), .Z(ereg_next[571]) );
  AND U44455 ( .A(mul_pow), .B(n40900), .Z(n40899) );
  XOR U44456 ( .A(ein[571]), .B(ein[570]), .Z(n40900) );
  XOR U44457 ( .A(ein[569]), .B(n40901), .Z(ereg_next[570]) );
  AND U44458 ( .A(mul_pow), .B(n40902), .Z(n40901) );
  XOR U44459 ( .A(ein[570]), .B(ein[569]), .Z(n40902) );
  XOR U44460 ( .A(ein[55]), .B(n40903), .Z(ereg_next[56]) );
  AND U44461 ( .A(mul_pow), .B(n40904), .Z(n40903) );
  XOR U44462 ( .A(ein[56]), .B(ein[55]), .Z(n40904) );
  XOR U44463 ( .A(ein[568]), .B(n40905), .Z(ereg_next[569]) );
  AND U44464 ( .A(mul_pow), .B(n40906), .Z(n40905) );
  XOR U44465 ( .A(ein[569]), .B(ein[568]), .Z(n40906) );
  XOR U44466 ( .A(ein[567]), .B(n40907), .Z(ereg_next[568]) );
  AND U44467 ( .A(mul_pow), .B(n40908), .Z(n40907) );
  XOR U44468 ( .A(ein[568]), .B(ein[567]), .Z(n40908) );
  XOR U44469 ( .A(ein[566]), .B(n40909), .Z(ereg_next[567]) );
  AND U44470 ( .A(mul_pow), .B(n40910), .Z(n40909) );
  XOR U44471 ( .A(ein[567]), .B(ein[566]), .Z(n40910) );
  XOR U44472 ( .A(ein[565]), .B(n40911), .Z(ereg_next[566]) );
  AND U44473 ( .A(mul_pow), .B(n40912), .Z(n40911) );
  XOR U44474 ( .A(ein[566]), .B(ein[565]), .Z(n40912) );
  XOR U44475 ( .A(ein[564]), .B(n40913), .Z(ereg_next[565]) );
  AND U44476 ( .A(mul_pow), .B(n40914), .Z(n40913) );
  XOR U44477 ( .A(ein[565]), .B(ein[564]), .Z(n40914) );
  XOR U44478 ( .A(ein[563]), .B(n40915), .Z(ereg_next[564]) );
  AND U44479 ( .A(mul_pow), .B(n40916), .Z(n40915) );
  XOR U44480 ( .A(ein[564]), .B(ein[563]), .Z(n40916) );
  XOR U44481 ( .A(ein[562]), .B(n40917), .Z(ereg_next[563]) );
  AND U44482 ( .A(mul_pow), .B(n40918), .Z(n40917) );
  XOR U44483 ( .A(ein[563]), .B(ein[562]), .Z(n40918) );
  XOR U44484 ( .A(ein[561]), .B(n40919), .Z(ereg_next[562]) );
  AND U44485 ( .A(mul_pow), .B(n40920), .Z(n40919) );
  XOR U44486 ( .A(ein[562]), .B(ein[561]), .Z(n40920) );
  XOR U44487 ( .A(ein[560]), .B(n40921), .Z(ereg_next[561]) );
  AND U44488 ( .A(mul_pow), .B(n40922), .Z(n40921) );
  XOR U44489 ( .A(ein[561]), .B(ein[560]), .Z(n40922) );
  XOR U44490 ( .A(ein[559]), .B(n40923), .Z(ereg_next[560]) );
  AND U44491 ( .A(mul_pow), .B(n40924), .Z(n40923) );
  XOR U44492 ( .A(ein[560]), .B(ein[559]), .Z(n40924) );
  XOR U44493 ( .A(ein[54]), .B(n40925), .Z(ereg_next[55]) );
  AND U44494 ( .A(mul_pow), .B(n40926), .Z(n40925) );
  XOR U44495 ( .A(ein[55]), .B(ein[54]), .Z(n40926) );
  XOR U44496 ( .A(ein[558]), .B(n40927), .Z(ereg_next[559]) );
  AND U44497 ( .A(mul_pow), .B(n40928), .Z(n40927) );
  XOR U44498 ( .A(ein[559]), .B(ein[558]), .Z(n40928) );
  XOR U44499 ( .A(ein[557]), .B(n40929), .Z(ereg_next[558]) );
  AND U44500 ( .A(mul_pow), .B(n40930), .Z(n40929) );
  XOR U44501 ( .A(ein[558]), .B(ein[557]), .Z(n40930) );
  XOR U44502 ( .A(ein[556]), .B(n40931), .Z(ereg_next[557]) );
  AND U44503 ( .A(mul_pow), .B(n40932), .Z(n40931) );
  XOR U44504 ( .A(ein[557]), .B(ein[556]), .Z(n40932) );
  XOR U44505 ( .A(ein[555]), .B(n40933), .Z(ereg_next[556]) );
  AND U44506 ( .A(mul_pow), .B(n40934), .Z(n40933) );
  XOR U44507 ( .A(ein[556]), .B(ein[555]), .Z(n40934) );
  XOR U44508 ( .A(ein[554]), .B(n40935), .Z(ereg_next[555]) );
  AND U44509 ( .A(mul_pow), .B(n40936), .Z(n40935) );
  XOR U44510 ( .A(ein[555]), .B(ein[554]), .Z(n40936) );
  XOR U44511 ( .A(ein[553]), .B(n40937), .Z(ereg_next[554]) );
  AND U44512 ( .A(mul_pow), .B(n40938), .Z(n40937) );
  XOR U44513 ( .A(ein[554]), .B(ein[553]), .Z(n40938) );
  XOR U44514 ( .A(ein[552]), .B(n40939), .Z(ereg_next[553]) );
  AND U44515 ( .A(mul_pow), .B(n40940), .Z(n40939) );
  XOR U44516 ( .A(ein[553]), .B(ein[552]), .Z(n40940) );
  XOR U44517 ( .A(ein[551]), .B(n40941), .Z(ereg_next[552]) );
  AND U44518 ( .A(mul_pow), .B(n40942), .Z(n40941) );
  XOR U44519 ( .A(ein[552]), .B(ein[551]), .Z(n40942) );
  XOR U44520 ( .A(ein[550]), .B(n40943), .Z(ereg_next[551]) );
  AND U44521 ( .A(mul_pow), .B(n40944), .Z(n40943) );
  XOR U44522 ( .A(ein[551]), .B(ein[550]), .Z(n40944) );
  XOR U44523 ( .A(ein[549]), .B(n40945), .Z(ereg_next[550]) );
  AND U44524 ( .A(mul_pow), .B(n40946), .Z(n40945) );
  XOR U44525 ( .A(ein[550]), .B(ein[549]), .Z(n40946) );
  XOR U44526 ( .A(ein[53]), .B(n40947), .Z(ereg_next[54]) );
  AND U44527 ( .A(mul_pow), .B(n40948), .Z(n40947) );
  XOR U44528 ( .A(ein[54]), .B(ein[53]), .Z(n40948) );
  XOR U44529 ( .A(ein[548]), .B(n40949), .Z(ereg_next[549]) );
  AND U44530 ( .A(mul_pow), .B(n40950), .Z(n40949) );
  XOR U44531 ( .A(ein[549]), .B(ein[548]), .Z(n40950) );
  XOR U44532 ( .A(ein[547]), .B(n40951), .Z(ereg_next[548]) );
  AND U44533 ( .A(mul_pow), .B(n40952), .Z(n40951) );
  XOR U44534 ( .A(ein[548]), .B(ein[547]), .Z(n40952) );
  XOR U44535 ( .A(ein[546]), .B(n40953), .Z(ereg_next[547]) );
  AND U44536 ( .A(mul_pow), .B(n40954), .Z(n40953) );
  XOR U44537 ( .A(ein[547]), .B(ein[546]), .Z(n40954) );
  XOR U44538 ( .A(ein[545]), .B(n40955), .Z(ereg_next[546]) );
  AND U44539 ( .A(mul_pow), .B(n40956), .Z(n40955) );
  XOR U44540 ( .A(ein[546]), .B(ein[545]), .Z(n40956) );
  XOR U44541 ( .A(ein[544]), .B(n40957), .Z(ereg_next[545]) );
  AND U44542 ( .A(mul_pow), .B(n40958), .Z(n40957) );
  XOR U44543 ( .A(ein[545]), .B(ein[544]), .Z(n40958) );
  XOR U44544 ( .A(ein[543]), .B(n40959), .Z(ereg_next[544]) );
  AND U44545 ( .A(mul_pow), .B(n40960), .Z(n40959) );
  XOR U44546 ( .A(ein[544]), .B(ein[543]), .Z(n40960) );
  XOR U44547 ( .A(ein[542]), .B(n40961), .Z(ereg_next[543]) );
  AND U44548 ( .A(mul_pow), .B(n40962), .Z(n40961) );
  XOR U44549 ( .A(ein[543]), .B(ein[542]), .Z(n40962) );
  XOR U44550 ( .A(ein[541]), .B(n40963), .Z(ereg_next[542]) );
  AND U44551 ( .A(mul_pow), .B(n40964), .Z(n40963) );
  XOR U44552 ( .A(ein[542]), .B(ein[541]), .Z(n40964) );
  XOR U44553 ( .A(ein[540]), .B(n40965), .Z(ereg_next[541]) );
  AND U44554 ( .A(mul_pow), .B(n40966), .Z(n40965) );
  XOR U44555 ( .A(ein[541]), .B(ein[540]), .Z(n40966) );
  XOR U44556 ( .A(ein[539]), .B(n40967), .Z(ereg_next[540]) );
  AND U44557 ( .A(mul_pow), .B(n40968), .Z(n40967) );
  XOR U44558 ( .A(ein[540]), .B(ein[539]), .Z(n40968) );
  XOR U44559 ( .A(ein[52]), .B(n40969), .Z(ereg_next[53]) );
  AND U44560 ( .A(mul_pow), .B(n40970), .Z(n40969) );
  XOR U44561 ( .A(ein[53]), .B(ein[52]), .Z(n40970) );
  XOR U44562 ( .A(ein[538]), .B(n40971), .Z(ereg_next[539]) );
  AND U44563 ( .A(mul_pow), .B(n40972), .Z(n40971) );
  XOR U44564 ( .A(ein[539]), .B(ein[538]), .Z(n40972) );
  XOR U44565 ( .A(ein[537]), .B(n40973), .Z(ereg_next[538]) );
  AND U44566 ( .A(mul_pow), .B(n40974), .Z(n40973) );
  XOR U44567 ( .A(ein[538]), .B(ein[537]), .Z(n40974) );
  XOR U44568 ( .A(ein[536]), .B(n40975), .Z(ereg_next[537]) );
  AND U44569 ( .A(mul_pow), .B(n40976), .Z(n40975) );
  XOR U44570 ( .A(ein[537]), .B(ein[536]), .Z(n40976) );
  XOR U44571 ( .A(ein[535]), .B(n40977), .Z(ereg_next[536]) );
  AND U44572 ( .A(mul_pow), .B(n40978), .Z(n40977) );
  XOR U44573 ( .A(ein[536]), .B(ein[535]), .Z(n40978) );
  XOR U44574 ( .A(ein[534]), .B(n40979), .Z(ereg_next[535]) );
  AND U44575 ( .A(mul_pow), .B(n40980), .Z(n40979) );
  XOR U44576 ( .A(ein[535]), .B(ein[534]), .Z(n40980) );
  XOR U44577 ( .A(ein[533]), .B(n40981), .Z(ereg_next[534]) );
  AND U44578 ( .A(mul_pow), .B(n40982), .Z(n40981) );
  XOR U44579 ( .A(ein[534]), .B(ein[533]), .Z(n40982) );
  XOR U44580 ( .A(ein[532]), .B(n40983), .Z(ereg_next[533]) );
  AND U44581 ( .A(mul_pow), .B(n40984), .Z(n40983) );
  XOR U44582 ( .A(ein[533]), .B(ein[532]), .Z(n40984) );
  XOR U44583 ( .A(ein[531]), .B(n40985), .Z(ereg_next[532]) );
  AND U44584 ( .A(mul_pow), .B(n40986), .Z(n40985) );
  XOR U44585 ( .A(ein[532]), .B(ein[531]), .Z(n40986) );
  XOR U44586 ( .A(ein[530]), .B(n40987), .Z(ereg_next[531]) );
  AND U44587 ( .A(mul_pow), .B(n40988), .Z(n40987) );
  XOR U44588 ( .A(ein[531]), .B(ein[530]), .Z(n40988) );
  XOR U44589 ( .A(ein[529]), .B(n40989), .Z(ereg_next[530]) );
  AND U44590 ( .A(mul_pow), .B(n40990), .Z(n40989) );
  XOR U44591 ( .A(ein[530]), .B(ein[529]), .Z(n40990) );
  XOR U44592 ( .A(ein[51]), .B(n40991), .Z(ereg_next[52]) );
  AND U44593 ( .A(mul_pow), .B(n40992), .Z(n40991) );
  XOR U44594 ( .A(ein[52]), .B(ein[51]), .Z(n40992) );
  XOR U44595 ( .A(ein[528]), .B(n40993), .Z(ereg_next[529]) );
  AND U44596 ( .A(mul_pow), .B(n40994), .Z(n40993) );
  XOR U44597 ( .A(ein[529]), .B(ein[528]), .Z(n40994) );
  XOR U44598 ( .A(ein[527]), .B(n40995), .Z(ereg_next[528]) );
  AND U44599 ( .A(mul_pow), .B(n40996), .Z(n40995) );
  XOR U44600 ( .A(ein[528]), .B(ein[527]), .Z(n40996) );
  XOR U44601 ( .A(ein[526]), .B(n40997), .Z(ereg_next[527]) );
  AND U44602 ( .A(mul_pow), .B(n40998), .Z(n40997) );
  XOR U44603 ( .A(ein[527]), .B(ein[526]), .Z(n40998) );
  XOR U44604 ( .A(ein[525]), .B(n40999), .Z(ereg_next[526]) );
  AND U44605 ( .A(mul_pow), .B(n41000), .Z(n40999) );
  XOR U44606 ( .A(ein[526]), .B(ein[525]), .Z(n41000) );
  XOR U44607 ( .A(ein[524]), .B(n41001), .Z(ereg_next[525]) );
  AND U44608 ( .A(mul_pow), .B(n41002), .Z(n41001) );
  XOR U44609 ( .A(ein[525]), .B(ein[524]), .Z(n41002) );
  XOR U44610 ( .A(ein[523]), .B(n41003), .Z(ereg_next[524]) );
  AND U44611 ( .A(mul_pow), .B(n41004), .Z(n41003) );
  XOR U44612 ( .A(ein[524]), .B(ein[523]), .Z(n41004) );
  XOR U44613 ( .A(ein[522]), .B(n41005), .Z(ereg_next[523]) );
  AND U44614 ( .A(mul_pow), .B(n41006), .Z(n41005) );
  XOR U44615 ( .A(ein[523]), .B(ein[522]), .Z(n41006) );
  XOR U44616 ( .A(ein[521]), .B(n41007), .Z(ereg_next[522]) );
  AND U44617 ( .A(mul_pow), .B(n41008), .Z(n41007) );
  XOR U44618 ( .A(ein[522]), .B(ein[521]), .Z(n41008) );
  XOR U44619 ( .A(ein[520]), .B(n41009), .Z(ereg_next[521]) );
  AND U44620 ( .A(mul_pow), .B(n41010), .Z(n41009) );
  XOR U44621 ( .A(ein[521]), .B(ein[520]), .Z(n41010) );
  XOR U44622 ( .A(ein[519]), .B(n41011), .Z(ereg_next[520]) );
  AND U44623 ( .A(mul_pow), .B(n41012), .Z(n41011) );
  XOR U44624 ( .A(ein[520]), .B(ein[519]), .Z(n41012) );
  XOR U44625 ( .A(ein[50]), .B(n41013), .Z(ereg_next[51]) );
  AND U44626 ( .A(mul_pow), .B(n41014), .Z(n41013) );
  XOR U44627 ( .A(ein[51]), .B(ein[50]), .Z(n41014) );
  XOR U44628 ( .A(ein[518]), .B(n41015), .Z(ereg_next[519]) );
  AND U44629 ( .A(mul_pow), .B(n41016), .Z(n41015) );
  XOR U44630 ( .A(ein[519]), .B(ein[518]), .Z(n41016) );
  XOR U44631 ( .A(ein[517]), .B(n41017), .Z(ereg_next[518]) );
  AND U44632 ( .A(mul_pow), .B(n41018), .Z(n41017) );
  XOR U44633 ( .A(ein[518]), .B(ein[517]), .Z(n41018) );
  XOR U44634 ( .A(ein[516]), .B(n41019), .Z(ereg_next[517]) );
  AND U44635 ( .A(mul_pow), .B(n41020), .Z(n41019) );
  XOR U44636 ( .A(ein[517]), .B(ein[516]), .Z(n41020) );
  XOR U44637 ( .A(ein[515]), .B(n41021), .Z(ereg_next[516]) );
  AND U44638 ( .A(mul_pow), .B(n41022), .Z(n41021) );
  XOR U44639 ( .A(ein[516]), .B(ein[515]), .Z(n41022) );
  XOR U44640 ( .A(ein[514]), .B(n41023), .Z(ereg_next[515]) );
  AND U44641 ( .A(mul_pow), .B(n41024), .Z(n41023) );
  XOR U44642 ( .A(ein[515]), .B(ein[514]), .Z(n41024) );
  XOR U44643 ( .A(ein[513]), .B(n41025), .Z(ereg_next[514]) );
  AND U44644 ( .A(mul_pow), .B(n41026), .Z(n41025) );
  XOR U44645 ( .A(ein[514]), .B(ein[513]), .Z(n41026) );
  XOR U44646 ( .A(ein[512]), .B(n41027), .Z(ereg_next[513]) );
  AND U44647 ( .A(mul_pow), .B(n41028), .Z(n41027) );
  XOR U44648 ( .A(ein[513]), .B(ein[512]), .Z(n41028) );
  XOR U44649 ( .A(ein[511]), .B(n41029), .Z(ereg_next[512]) );
  AND U44650 ( .A(mul_pow), .B(n41030), .Z(n41029) );
  XOR U44651 ( .A(ein[512]), .B(ein[511]), .Z(n41030) );
  XOR U44652 ( .A(ein[510]), .B(n41031), .Z(ereg_next[511]) );
  AND U44653 ( .A(mul_pow), .B(n41032), .Z(n41031) );
  XOR U44654 ( .A(ein[511]), .B(ein[510]), .Z(n41032) );
  XOR U44655 ( .A(ein[509]), .B(n41033), .Z(ereg_next[510]) );
  AND U44656 ( .A(mul_pow), .B(n41034), .Z(n41033) );
  XOR U44657 ( .A(ein[510]), .B(ein[509]), .Z(n41034) );
  XOR U44658 ( .A(ein[49]), .B(n41035), .Z(ereg_next[50]) );
  AND U44659 ( .A(mul_pow), .B(n41036), .Z(n41035) );
  XOR U44660 ( .A(ein[50]), .B(ein[49]), .Z(n41036) );
  XOR U44661 ( .A(ein[508]), .B(n41037), .Z(ereg_next[509]) );
  AND U44662 ( .A(mul_pow), .B(n41038), .Z(n41037) );
  XOR U44663 ( .A(ein[509]), .B(ein[508]), .Z(n41038) );
  XOR U44664 ( .A(ein[507]), .B(n41039), .Z(ereg_next[508]) );
  AND U44665 ( .A(mul_pow), .B(n41040), .Z(n41039) );
  XOR U44666 ( .A(ein[508]), .B(ein[507]), .Z(n41040) );
  XOR U44667 ( .A(ein[506]), .B(n41041), .Z(ereg_next[507]) );
  AND U44668 ( .A(mul_pow), .B(n41042), .Z(n41041) );
  XOR U44669 ( .A(ein[507]), .B(ein[506]), .Z(n41042) );
  XOR U44670 ( .A(ein[505]), .B(n41043), .Z(ereg_next[506]) );
  AND U44671 ( .A(mul_pow), .B(n41044), .Z(n41043) );
  XOR U44672 ( .A(ein[506]), .B(ein[505]), .Z(n41044) );
  XOR U44673 ( .A(ein[504]), .B(n41045), .Z(ereg_next[505]) );
  AND U44674 ( .A(mul_pow), .B(n41046), .Z(n41045) );
  XOR U44675 ( .A(ein[505]), .B(ein[504]), .Z(n41046) );
  XOR U44676 ( .A(ein[503]), .B(n41047), .Z(ereg_next[504]) );
  AND U44677 ( .A(mul_pow), .B(n41048), .Z(n41047) );
  XOR U44678 ( .A(ein[504]), .B(ein[503]), .Z(n41048) );
  XOR U44679 ( .A(ein[502]), .B(n41049), .Z(ereg_next[503]) );
  AND U44680 ( .A(mul_pow), .B(n41050), .Z(n41049) );
  XOR U44681 ( .A(ein[503]), .B(ein[502]), .Z(n41050) );
  XOR U44682 ( .A(ein[501]), .B(n41051), .Z(ereg_next[502]) );
  AND U44683 ( .A(mul_pow), .B(n41052), .Z(n41051) );
  XOR U44684 ( .A(ein[502]), .B(ein[501]), .Z(n41052) );
  XOR U44685 ( .A(ein[500]), .B(n41053), .Z(ereg_next[501]) );
  AND U44686 ( .A(mul_pow), .B(n41054), .Z(n41053) );
  XOR U44687 ( .A(ein[501]), .B(ein[500]), .Z(n41054) );
  XOR U44688 ( .A(ein[499]), .B(n41055), .Z(ereg_next[500]) );
  AND U44689 ( .A(mul_pow), .B(n41056), .Z(n41055) );
  XOR U44690 ( .A(ein[500]), .B(ein[499]), .Z(n41056) );
  XOR U44691 ( .A(ein[3]), .B(n41057), .Z(ereg_next[4]) );
  AND U44692 ( .A(mul_pow), .B(n41058), .Z(n41057) );
  XOR U44693 ( .A(ein[4]), .B(ein[3]), .Z(n41058) );
  XOR U44694 ( .A(ein[48]), .B(n41059), .Z(ereg_next[49]) );
  AND U44695 ( .A(mul_pow), .B(n41060), .Z(n41059) );
  XOR U44696 ( .A(ein[49]), .B(ein[48]), .Z(n41060) );
  XOR U44697 ( .A(ein[498]), .B(n41061), .Z(ereg_next[499]) );
  AND U44698 ( .A(mul_pow), .B(n41062), .Z(n41061) );
  XOR U44699 ( .A(ein[499]), .B(ein[498]), .Z(n41062) );
  XOR U44700 ( .A(ein[497]), .B(n41063), .Z(ereg_next[498]) );
  AND U44701 ( .A(mul_pow), .B(n41064), .Z(n41063) );
  XOR U44702 ( .A(ein[498]), .B(ein[497]), .Z(n41064) );
  XOR U44703 ( .A(ein[496]), .B(n41065), .Z(ereg_next[497]) );
  AND U44704 ( .A(mul_pow), .B(n41066), .Z(n41065) );
  XOR U44705 ( .A(ein[497]), .B(ein[496]), .Z(n41066) );
  XOR U44706 ( .A(ein[495]), .B(n41067), .Z(ereg_next[496]) );
  AND U44707 ( .A(mul_pow), .B(n41068), .Z(n41067) );
  XOR U44708 ( .A(ein[496]), .B(ein[495]), .Z(n41068) );
  XOR U44709 ( .A(ein[494]), .B(n41069), .Z(ereg_next[495]) );
  AND U44710 ( .A(mul_pow), .B(n41070), .Z(n41069) );
  XOR U44711 ( .A(ein[495]), .B(ein[494]), .Z(n41070) );
  XOR U44712 ( .A(ein[493]), .B(n41071), .Z(ereg_next[494]) );
  AND U44713 ( .A(mul_pow), .B(n41072), .Z(n41071) );
  XOR U44714 ( .A(ein[494]), .B(ein[493]), .Z(n41072) );
  XOR U44715 ( .A(ein[492]), .B(n41073), .Z(ereg_next[493]) );
  AND U44716 ( .A(mul_pow), .B(n41074), .Z(n41073) );
  XOR U44717 ( .A(ein[493]), .B(ein[492]), .Z(n41074) );
  XOR U44718 ( .A(ein[491]), .B(n41075), .Z(ereg_next[492]) );
  AND U44719 ( .A(mul_pow), .B(n41076), .Z(n41075) );
  XOR U44720 ( .A(ein[492]), .B(ein[491]), .Z(n41076) );
  XOR U44721 ( .A(ein[490]), .B(n41077), .Z(ereg_next[491]) );
  AND U44722 ( .A(mul_pow), .B(n41078), .Z(n41077) );
  XOR U44723 ( .A(ein[491]), .B(ein[490]), .Z(n41078) );
  XOR U44724 ( .A(ein[489]), .B(n41079), .Z(ereg_next[490]) );
  AND U44725 ( .A(mul_pow), .B(n41080), .Z(n41079) );
  XOR U44726 ( .A(ein[490]), .B(ein[489]), .Z(n41080) );
  XOR U44727 ( .A(ein[47]), .B(n41081), .Z(ereg_next[48]) );
  AND U44728 ( .A(mul_pow), .B(n41082), .Z(n41081) );
  XOR U44729 ( .A(ein[48]), .B(ein[47]), .Z(n41082) );
  XOR U44730 ( .A(ein[488]), .B(n41083), .Z(ereg_next[489]) );
  AND U44731 ( .A(mul_pow), .B(n41084), .Z(n41083) );
  XOR U44732 ( .A(ein[489]), .B(ein[488]), .Z(n41084) );
  XOR U44733 ( .A(ein[487]), .B(n41085), .Z(ereg_next[488]) );
  AND U44734 ( .A(mul_pow), .B(n41086), .Z(n41085) );
  XOR U44735 ( .A(ein[488]), .B(ein[487]), .Z(n41086) );
  XOR U44736 ( .A(ein[486]), .B(n41087), .Z(ereg_next[487]) );
  AND U44737 ( .A(mul_pow), .B(n41088), .Z(n41087) );
  XOR U44738 ( .A(ein[487]), .B(ein[486]), .Z(n41088) );
  XOR U44739 ( .A(ein[485]), .B(n41089), .Z(ereg_next[486]) );
  AND U44740 ( .A(mul_pow), .B(n41090), .Z(n41089) );
  XOR U44741 ( .A(ein[486]), .B(ein[485]), .Z(n41090) );
  XOR U44742 ( .A(ein[484]), .B(n41091), .Z(ereg_next[485]) );
  AND U44743 ( .A(mul_pow), .B(n41092), .Z(n41091) );
  XOR U44744 ( .A(ein[485]), .B(ein[484]), .Z(n41092) );
  XOR U44745 ( .A(ein[483]), .B(n41093), .Z(ereg_next[484]) );
  AND U44746 ( .A(mul_pow), .B(n41094), .Z(n41093) );
  XOR U44747 ( .A(ein[484]), .B(ein[483]), .Z(n41094) );
  XOR U44748 ( .A(ein[482]), .B(n41095), .Z(ereg_next[483]) );
  AND U44749 ( .A(mul_pow), .B(n41096), .Z(n41095) );
  XOR U44750 ( .A(ein[483]), .B(ein[482]), .Z(n41096) );
  XOR U44751 ( .A(ein[481]), .B(n41097), .Z(ereg_next[482]) );
  AND U44752 ( .A(mul_pow), .B(n41098), .Z(n41097) );
  XOR U44753 ( .A(ein[482]), .B(ein[481]), .Z(n41098) );
  XOR U44754 ( .A(ein[480]), .B(n41099), .Z(ereg_next[481]) );
  AND U44755 ( .A(mul_pow), .B(n41100), .Z(n41099) );
  XOR U44756 ( .A(ein[481]), .B(ein[480]), .Z(n41100) );
  XOR U44757 ( .A(ein[479]), .B(n41101), .Z(ereg_next[480]) );
  AND U44758 ( .A(mul_pow), .B(n41102), .Z(n41101) );
  XOR U44759 ( .A(ein[480]), .B(ein[479]), .Z(n41102) );
  XOR U44760 ( .A(ein[46]), .B(n41103), .Z(ereg_next[47]) );
  AND U44761 ( .A(mul_pow), .B(n41104), .Z(n41103) );
  XOR U44762 ( .A(ein[47]), .B(ein[46]), .Z(n41104) );
  XOR U44763 ( .A(ein[478]), .B(n41105), .Z(ereg_next[479]) );
  AND U44764 ( .A(mul_pow), .B(n41106), .Z(n41105) );
  XOR U44765 ( .A(ein[479]), .B(ein[478]), .Z(n41106) );
  XOR U44766 ( .A(ein[477]), .B(n41107), .Z(ereg_next[478]) );
  AND U44767 ( .A(mul_pow), .B(n41108), .Z(n41107) );
  XOR U44768 ( .A(ein[478]), .B(ein[477]), .Z(n41108) );
  XOR U44769 ( .A(ein[476]), .B(n41109), .Z(ereg_next[477]) );
  AND U44770 ( .A(mul_pow), .B(n41110), .Z(n41109) );
  XOR U44771 ( .A(ein[477]), .B(ein[476]), .Z(n41110) );
  XOR U44772 ( .A(ein[475]), .B(n41111), .Z(ereg_next[476]) );
  AND U44773 ( .A(mul_pow), .B(n41112), .Z(n41111) );
  XOR U44774 ( .A(ein[476]), .B(ein[475]), .Z(n41112) );
  XOR U44775 ( .A(ein[474]), .B(n41113), .Z(ereg_next[475]) );
  AND U44776 ( .A(mul_pow), .B(n41114), .Z(n41113) );
  XOR U44777 ( .A(ein[475]), .B(ein[474]), .Z(n41114) );
  XOR U44778 ( .A(ein[473]), .B(n41115), .Z(ereg_next[474]) );
  AND U44779 ( .A(mul_pow), .B(n41116), .Z(n41115) );
  XOR U44780 ( .A(ein[474]), .B(ein[473]), .Z(n41116) );
  XOR U44781 ( .A(ein[472]), .B(n41117), .Z(ereg_next[473]) );
  AND U44782 ( .A(mul_pow), .B(n41118), .Z(n41117) );
  XOR U44783 ( .A(ein[473]), .B(ein[472]), .Z(n41118) );
  XOR U44784 ( .A(ein[471]), .B(n41119), .Z(ereg_next[472]) );
  AND U44785 ( .A(mul_pow), .B(n41120), .Z(n41119) );
  XOR U44786 ( .A(ein[472]), .B(ein[471]), .Z(n41120) );
  XOR U44787 ( .A(ein[470]), .B(n41121), .Z(ereg_next[471]) );
  AND U44788 ( .A(mul_pow), .B(n41122), .Z(n41121) );
  XOR U44789 ( .A(ein[471]), .B(ein[470]), .Z(n41122) );
  XOR U44790 ( .A(ein[469]), .B(n41123), .Z(ereg_next[470]) );
  AND U44791 ( .A(mul_pow), .B(n41124), .Z(n41123) );
  XOR U44792 ( .A(ein[470]), .B(ein[469]), .Z(n41124) );
  XOR U44793 ( .A(ein[45]), .B(n41125), .Z(ereg_next[46]) );
  AND U44794 ( .A(mul_pow), .B(n41126), .Z(n41125) );
  XOR U44795 ( .A(ein[46]), .B(ein[45]), .Z(n41126) );
  XOR U44796 ( .A(ein[468]), .B(n41127), .Z(ereg_next[469]) );
  AND U44797 ( .A(mul_pow), .B(n41128), .Z(n41127) );
  XOR U44798 ( .A(ein[469]), .B(ein[468]), .Z(n41128) );
  XOR U44799 ( .A(ein[467]), .B(n41129), .Z(ereg_next[468]) );
  AND U44800 ( .A(mul_pow), .B(n41130), .Z(n41129) );
  XOR U44801 ( .A(ein[468]), .B(ein[467]), .Z(n41130) );
  XOR U44802 ( .A(ein[466]), .B(n41131), .Z(ereg_next[467]) );
  AND U44803 ( .A(mul_pow), .B(n41132), .Z(n41131) );
  XOR U44804 ( .A(ein[467]), .B(ein[466]), .Z(n41132) );
  XOR U44805 ( .A(ein[465]), .B(n41133), .Z(ereg_next[466]) );
  AND U44806 ( .A(mul_pow), .B(n41134), .Z(n41133) );
  XOR U44807 ( .A(ein[466]), .B(ein[465]), .Z(n41134) );
  XOR U44808 ( .A(ein[464]), .B(n41135), .Z(ereg_next[465]) );
  AND U44809 ( .A(mul_pow), .B(n41136), .Z(n41135) );
  XOR U44810 ( .A(ein[465]), .B(ein[464]), .Z(n41136) );
  XOR U44811 ( .A(ein[463]), .B(n41137), .Z(ereg_next[464]) );
  AND U44812 ( .A(mul_pow), .B(n41138), .Z(n41137) );
  XOR U44813 ( .A(ein[464]), .B(ein[463]), .Z(n41138) );
  XOR U44814 ( .A(ein[462]), .B(n41139), .Z(ereg_next[463]) );
  AND U44815 ( .A(mul_pow), .B(n41140), .Z(n41139) );
  XOR U44816 ( .A(ein[463]), .B(ein[462]), .Z(n41140) );
  XOR U44817 ( .A(ein[461]), .B(n41141), .Z(ereg_next[462]) );
  AND U44818 ( .A(mul_pow), .B(n41142), .Z(n41141) );
  XOR U44819 ( .A(ein[462]), .B(ein[461]), .Z(n41142) );
  XOR U44820 ( .A(ein[460]), .B(n41143), .Z(ereg_next[461]) );
  AND U44821 ( .A(mul_pow), .B(n41144), .Z(n41143) );
  XOR U44822 ( .A(ein[461]), .B(ein[460]), .Z(n41144) );
  XOR U44823 ( .A(ein[459]), .B(n41145), .Z(ereg_next[460]) );
  AND U44824 ( .A(mul_pow), .B(n41146), .Z(n41145) );
  XOR U44825 ( .A(ein[460]), .B(ein[459]), .Z(n41146) );
  XOR U44826 ( .A(ein[44]), .B(n41147), .Z(ereg_next[45]) );
  AND U44827 ( .A(mul_pow), .B(n41148), .Z(n41147) );
  XOR U44828 ( .A(ein[45]), .B(ein[44]), .Z(n41148) );
  XOR U44829 ( .A(ein[458]), .B(n41149), .Z(ereg_next[459]) );
  AND U44830 ( .A(mul_pow), .B(n41150), .Z(n41149) );
  XOR U44831 ( .A(ein[459]), .B(ein[458]), .Z(n41150) );
  XOR U44832 ( .A(ein[457]), .B(n41151), .Z(ereg_next[458]) );
  AND U44833 ( .A(mul_pow), .B(n41152), .Z(n41151) );
  XOR U44834 ( .A(ein[458]), .B(ein[457]), .Z(n41152) );
  XOR U44835 ( .A(ein[456]), .B(n41153), .Z(ereg_next[457]) );
  AND U44836 ( .A(mul_pow), .B(n41154), .Z(n41153) );
  XOR U44837 ( .A(ein[457]), .B(ein[456]), .Z(n41154) );
  XOR U44838 ( .A(ein[455]), .B(n41155), .Z(ereg_next[456]) );
  AND U44839 ( .A(mul_pow), .B(n41156), .Z(n41155) );
  XOR U44840 ( .A(ein[456]), .B(ein[455]), .Z(n41156) );
  XOR U44841 ( .A(ein[454]), .B(n41157), .Z(ereg_next[455]) );
  AND U44842 ( .A(mul_pow), .B(n41158), .Z(n41157) );
  XOR U44843 ( .A(ein[455]), .B(ein[454]), .Z(n41158) );
  XOR U44844 ( .A(ein[453]), .B(n41159), .Z(ereg_next[454]) );
  AND U44845 ( .A(mul_pow), .B(n41160), .Z(n41159) );
  XOR U44846 ( .A(ein[454]), .B(ein[453]), .Z(n41160) );
  XOR U44847 ( .A(ein[452]), .B(n41161), .Z(ereg_next[453]) );
  AND U44848 ( .A(mul_pow), .B(n41162), .Z(n41161) );
  XOR U44849 ( .A(ein[453]), .B(ein[452]), .Z(n41162) );
  XOR U44850 ( .A(ein[451]), .B(n41163), .Z(ereg_next[452]) );
  AND U44851 ( .A(mul_pow), .B(n41164), .Z(n41163) );
  XOR U44852 ( .A(ein[452]), .B(ein[451]), .Z(n41164) );
  XOR U44853 ( .A(ein[450]), .B(n41165), .Z(ereg_next[451]) );
  AND U44854 ( .A(mul_pow), .B(n41166), .Z(n41165) );
  XOR U44855 ( .A(ein[451]), .B(ein[450]), .Z(n41166) );
  XOR U44856 ( .A(ein[449]), .B(n41167), .Z(ereg_next[450]) );
  AND U44857 ( .A(mul_pow), .B(n41168), .Z(n41167) );
  XOR U44858 ( .A(ein[450]), .B(ein[449]), .Z(n41168) );
  XOR U44859 ( .A(ein[43]), .B(n41169), .Z(ereg_next[44]) );
  AND U44860 ( .A(mul_pow), .B(n41170), .Z(n41169) );
  XOR U44861 ( .A(ein[44]), .B(ein[43]), .Z(n41170) );
  XOR U44862 ( .A(ein[448]), .B(n41171), .Z(ereg_next[449]) );
  AND U44863 ( .A(mul_pow), .B(n41172), .Z(n41171) );
  XOR U44864 ( .A(ein[449]), .B(ein[448]), .Z(n41172) );
  XOR U44865 ( .A(ein[447]), .B(n41173), .Z(ereg_next[448]) );
  AND U44866 ( .A(mul_pow), .B(n41174), .Z(n41173) );
  XOR U44867 ( .A(ein[448]), .B(ein[447]), .Z(n41174) );
  XOR U44868 ( .A(ein[446]), .B(n41175), .Z(ereg_next[447]) );
  AND U44869 ( .A(mul_pow), .B(n41176), .Z(n41175) );
  XOR U44870 ( .A(ein[447]), .B(ein[446]), .Z(n41176) );
  XOR U44871 ( .A(ein[445]), .B(n41177), .Z(ereg_next[446]) );
  AND U44872 ( .A(mul_pow), .B(n41178), .Z(n41177) );
  XOR U44873 ( .A(ein[446]), .B(ein[445]), .Z(n41178) );
  XOR U44874 ( .A(ein[444]), .B(n41179), .Z(ereg_next[445]) );
  AND U44875 ( .A(mul_pow), .B(n41180), .Z(n41179) );
  XOR U44876 ( .A(ein[445]), .B(ein[444]), .Z(n41180) );
  XOR U44877 ( .A(ein[443]), .B(n41181), .Z(ereg_next[444]) );
  AND U44878 ( .A(mul_pow), .B(n41182), .Z(n41181) );
  XOR U44879 ( .A(ein[444]), .B(ein[443]), .Z(n41182) );
  XOR U44880 ( .A(ein[442]), .B(n41183), .Z(ereg_next[443]) );
  AND U44881 ( .A(mul_pow), .B(n41184), .Z(n41183) );
  XOR U44882 ( .A(ein[443]), .B(ein[442]), .Z(n41184) );
  XOR U44883 ( .A(ein[441]), .B(n41185), .Z(ereg_next[442]) );
  AND U44884 ( .A(mul_pow), .B(n41186), .Z(n41185) );
  XOR U44885 ( .A(ein[442]), .B(ein[441]), .Z(n41186) );
  XOR U44886 ( .A(ein[440]), .B(n41187), .Z(ereg_next[441]) );
  AND U44887 ( .A(mul_pow), .B(n41188), .Z(n41187) );
  XOR U44888 ( .A(ein[441]), .B(ein[440]), .Z(n41188) );
  XOR U44889 ( .A(ein[439]), .B(n41189), .Z(ereg_next[440]) );
  AND U44890 ( .A(mul_pow), .B(n41190), .Z(n41189) );
  XOR U44891 ( .A(ein[440]), .B(ein[439]), .Z(n41190) );
  XOR U44892 ( .A(ein[42]), .B(n41191), .Z(ereg_next[43]) );
  AND U44893 ( .A(mul_pow), .B(n41192), .Z(n41191) );
  XOR U44894 ( .A(ein[43]), .B(ein[42]), .Z(n41192) );
  XOR U44895 ( .A(ein[438]), .B(n41193), .Z(ereg_next[439]) );
  AND U44896 ( .A(mul_pow), .B(n41194), .Z(n41193) );
  XOR U44897 ( .A(ein[439]), .B(ein[438]), .Z(n41194) );
  XOR U44898 ( .A(ein[437]), .B(n41195), .Z(ereg_next[438]) );
  AND U44899 ( .A(mul_pow), .B(n41196), .Z(n41195) );
  XOR U44900 ( .A(ein[438]), .B(ein[437]), .Z(n41196) );
  XOR U44901 ( .A(ein[436]), .B(n41197), .Z(ereg_next[437]) );
  AND U44902 ( .A(mul_pow), .B(n41198), .Z(n41197) );
  XOR U44903 ( .A(ein[437]), .B(ein[436]), .Z(n41198) );
  XOR U44904 ( .A(ein[435]), .B(n41199), .Z(ereg_next[436]) );
  AND U44905 ( .A(mul_pow), .B(n41200), .Z(n41199) );
  XOR U44906 ( .A(ein[436]), .B(ein[435]), .Z(n41200) );
  XOR U44907 ( .A(ein[434]), .B(n41201), .Z(ereg_next[435]) );
  AND U44908 ( .A(mul_pow), .B(n41202), .Z(n41201) );
  XOR U44909 ( .A(ein[435]), .B(ein[434]), .Z(n41202) );
  XOR U44910 ( .A(ein[433]), .B(n41203), .Z(ereg_next[434]) );
  AND U44911 ( .A(mul_pow), .B(n41204), .Z(n41203) );
  XOR U44912 ( .A(ein[434]), .B(ein[433]), .Z(n41204) );
  XOR U44913 ( .A(ein[432]), .B(n41205), .Z(ereg_next[433]) );
  AND U44914 ( .A(mul_pow), .B(n41206), .Z(n41205) );
  XOR U44915 ( .A(ein[433]), .B(ein[432]), .Z(n41206) );
  XOR U44916 ( .A(ein[431]), .B(n41207), .Z(ereg_next[432]) );
  AND U44917 ( .A(mul_pow), .B(n41208), .Z(n41207) );
  XOR U44918 ( .A(ein[432]), .B(ein[431]), .Z(n41208) );
  XOR U44919 ( .A(ein[430]), .B(n41209), .Z(ereg_next[431]) );
  AND U44920 ( .A(mul_pow), .B(n41210), .Z(n41209) );
  XOR U44921 ( .A(ein[431]), .B(ein[430]), .Z(n41210) );
  XOR U44922 ( .A(ein[429]), .B(n41211), .Z(ereg_next[430]) );
  AND U44923 ( .A(mul_pow), .B(n41212), .Z(n41211) );
  XOR U44924 ( .A(ein[430]), .B(ein[429]), .Z(n41212) );
  XOR U44925 ( .A(ein[41]), .B(n41213), .Z(ereg_next[42]) );
  AND U44926 ( .A(mul_pow), .B(n41214), .Z(n41213) );
  XOR U44927 ( .A(ein[42]), .B(ein[41]), .Z(n41214) );
  XOR U44928 ( .A(ein[428]), .B(n41215), .Z(ereg_next[429]) );
  AND U44929 ( .A(mul_pow), .B(n41216), .Z(n41215) );
  XOR U44930 ( .A(ein[429]), .B(ein[428]), .Z(n41216) );
  XOR U44931 ( .A(ein[427]), .B(n41217), .Z(ereg_next[428]) );
  AND U44932 ( .A(mul_pow), .B(n41218), .Z(n41217) );
  XOR U44933 ( .A(ein[428]), .B(ein[427]), .Z(n41218) );
  XOR U44934 ( .A(ein[426]), .B(n41219), .Z(ereg_next[427]) );
  AND U44935 ( .A(mul_pow), .B(n41220), .Z(n41219) );
  XOR U44936 ( .A(ein[427]), .B(ein[426]), .Z(n41220) );
  XOR U44937 ( .A(ein[425]), .B(n41221), .Z(ereg_next[426]) );
  AND U44938 ( .A(mul_pow), .B(n41222), .Z(n41221) );
  XOR U44939 ( .A(ein[426]), .B(ein[425]), .Z(n41222) );
  XOR U44940 ( .A(ein[424]), .B(n41223), .Z(ereg_next[425]) );
  AND U44941 ( .A(mul_pow), .B(n41224), .Z(n41223) );
  XOR U44942 ( .A(ein[425]), .B(ein[424]), .Z(n41224) );
  XOR U44943 ( .A(ein[423]), .B(n41225), .Z(ereg_next[424]) );
  AND U44944 ( .A(mul_pow), .B(n41226), .Z(n41225) );
  XOR U44945 ( .A(ein[424]), .B(ein[423]), .Z(n41226) );
  XOR U44946 ( .A(ein[422]), .B(n41227), .Z(ereg_next[423]) );
  AND U44947 ( .A(mul_pow), .B(n41228), .Z(n41227) );
  XOR U44948 ( .A(ein[423]), .B(ein[422]), .Z(n41228) );
  XOR U44949 ( .A(ein[421]), .B(n41229), .Z(ereg_next[422]) );
  AND U44950 ( .A(mul_pow), .B(n41230), .Z(n41229) );
  XOR U44951 ( .A(ein[422]), .B(ein[421]), .Z(n41230) );
  XOR U44952 ( .A(ein[420]), .B(n41231), .Z(ereg_next[421]) );
  AND U44953 ( .A(mul_pow), .B(n41232), .Z(n41231) );
  XOR U44954 ( .A(ein[421]), .B(ein[420]), .Z(n41232) );
  XOR U44955 ( .A(ein[419]), .B(n41233), .Z(ereg_next[420]) );
  AND U44956 ( .A(mul_pow), .B(n41234), .Z(n41233) );
  XOR U44957 ( .A(ein[420]), .B(ein[419]), .Z(n41234) );
  XOR U44958 ( .A(ein[40]), .B(n41235), .Z(ereg_next[41]) );
  AND U44959 ( .A(mul_pow), .B(n41236), .Z(n41235) );
  XOR U44960 ( .A(ein[41]), .B(ein[40]), .Z(n41236) );
  XOR U44961 ( .A(ein[418]), .B(n41237), .Z(ereg_next[419]) );
  AND U44962 ( .A(mul_pow), .B(n41238), .Z(n41237) );
  XOR U44963 ( .A(ein[419]), .B(ein[418]), .Z(n41238) );
  XOR U44964 ( .A(ein[417]), .B(n41239), .Z(ereg_next[418]) );
  AND U44965 ( .A(mul_pow), .B(n41240), .Z(n41239) );
  XOR U44966 ( .A(ein[418]), .B(ein[417]), .Z(n41240) );
  XOR U44967 ( .A(ein[416]), .B(n41241), .Z(ereg_next[417]) );
  AND U44968 ( .A(mul_pow), .B(n41242), .Z(n41241) );
  XOR U44969 ( .A(ein[417]), .B(ein[416]), .Z(n41242) );
  XOR U44970 ( .A(ein[415]), .B(n41243), .Z(ereg_next[416]) );
  AND U44971 ( .A(mul_pow), .B(n41244), .Z(n41243) );
  XOR U44972 ( .A(ein[416]), .B(ein[415]), .Z(n41244) );
  XOR U44973 ( .A(ein[414]), .B(n41245), .Z(ereg_next[415]) );
  AND U44974 ( .A(mul_pow), .B(n41246), .Z(n41245) );
  XOR U44975 ( .A(ein[415]), .B(ein[414]), .Z(n41246) );
  XOR U44976 ( .A(ein[413]), .B(n41247), .Z(ereg_next[414]) );
  AND U44977 ( .A(mul_pow), .B(n41248), .Z(n41247) );
  XOR U44978 ( .A(ein[414]), .B(ein[413]), .Z(n41248) );
  XOR U44979 ( .A(ein[412]), .B(n41249), .Z(ereg_next[413]) );
  AND U44980 ( .A(mul_pow), .B(n41250), .Z(n41249) );
  XOR U44981 ( .A(ein[413]), .B(ein[412]), .Z(n41250) );
  XOR U44982 ( .A(ein[411]), .B(n41251), .Z(ereg_next[412]) );
  AND U44983 ( .A(mul_pow), .B(n41252), .Z(n41251) );
  XOR U44984 ( .A(ein[412]), .B(ein[411]), .Z(n41252) );
  XOR U44985 ( .A(ein[410]), .B(n41253), .Z(ereg_next[411]) );
  AND U44986 ( .A(mul_pow), .B(n41254), .Z(n41253) );
  XOR U44987 ( .A(ein[411]), .B(ein[410]), .Z(n41254) );
  XOR U44988 ( .A(ein[409]), .B(n41255), .Z(ereg_next[410]) );
  AND U44989 ( .A(mul_pow), .B(n41256), .Z(n41255) );
  XOR U44990 ( .A(ein[410]), .B(ein[409]), .Z(n41256) );
  XOR U44991 ( .A(ein[39]), .B(n41257), .Z(ereg_next[40]) );
  AND U44992 ( .A(mul_pow), .B(n41258), .Z(n41257) );
  XOR U44993 ( .A(ein[40]), .B(ein[39]), .Z(n41258) );
  XOR U44994 ( .A(ein[408]), .B(n41259), .Z(ereg_next[409]) );
  AND U44995 ( .A(mul_pow), .B(n41260), .Z(n41259) );
  XOR U44996 ( .A(ein[409]), .B(ein[408]), .Z(n41260) );
  XOR U44997 ( .A(ein[407]), .B(n41261), .Z(ereg_next[408]) );
  AND U44998 ( .A(mul_pow), .B(n41262), .Z(n41261) );
  XOR U44999 ( .A(ein[408]), .B(ein[407]), .Z(n41262) );
  XOR U45000 ( .A(ein[406]), .B(n41263), .Z(ereg_next[407]) );
  AND U45001 ( .A(mul_pow), .B(n41264), .Z(n41263) );
  XOR U45002 ( .A(ein[407]), .B(ein[406]), .Z(n41264) );
  XOR U45003 ( .A(ein[405]), .B(n41265), .Z(ereg_next[406]) );
  AND U45004 ( .A(mul_pow), .B(n41266), .Z(n41265) );
  XOR U45005 ( .A(ein[406]), .B(ein[405]), .Z(n41266) );
  XOR U45006 ( .A(ein[404]), .B(n41267), .Z(ereg_next[405]) );
  AND U45007 ( .A(mul_pow), .B(n41268), .Z(n41267) );
  XOR U45008 ( .A(ein[405]), .B(ein[404]), .Z(n41268) );
  XOR U45009 ( .A(ein[403]), .B(n41269), .Z(ereg_next[404]) );
  AND U45010 ( .A(mul_pow), .B(n41270), .Z(n41269) );
  XOR U45011 ( .A(ein[404]), .B(ein[403]), .Z(n41270) );
  XOR U45012 ( .A(ein[402]), .B(n41271), .Z(ereg_next[403]) );
  AND U45013 ( .A(mul_pow), .B(n41272), .Z(n41271) );
  XOR U45014 ( .A(ein[403]), .B(ein[402]), .Z(n41272) );
  XOR U45015 ( .A(ein[401]), .B(n41273), .Z(ereg_next[402]) );
  AND U45016 ( .A(mul_pow), .B(n41274), .Z(n41273) );
  XOR U45017 ( .A(ein[402]), .B(ein[401]), .Z(n41274) );
  XOR U45018 ( .A(ein[400]), .B(n41275), .Z(ereg_next[401]) );
  AND U45019 ( .A(mul_pow), .B(n41276), .Z(n41275) );
  XOR U45020 ( .A(ein[401]), .B(ein[400]), .Z(n41276) );
  XOR U45021 ( .A(ein[399]), .B(n41277), .Z(ereg_next[400]) );
  AND U45022 ( .A(mul_pow), .B(n41278), .Z(n41277) );
  XOR U45023 ( .A(ein[400]), .B(ein[399]), .Z(n41278) );
  XOR U45024 ( .A(ein[2]), .B(n41279), .Z(ereg_next[3]) );
  AND U45025 ( .A(mul_pow), .B(n41280), .Z(n41279) );
  XOR U45026 ( .A(ein[3]), .B(ein[2]), .Z(n41280) );
  XOR U45027 ( .A(ein[38]), .B(n41281), .Z(ereg_next[39]) );
  AND U45028 ( .A(mul_pow), .B(n41282), .Z(n41281) );
  XOR U45029 ( .A(ein[39]), .B(ein[38]), .Z(n41282) );
  XOR U45030 ( .A(ein[398]), .B(n41283), .Z(ereg_next[399]) );
  AND U45031 ( .A(mul_pow), .B(n41284), .Z(n41283) );
  XOR U45032 ( .A(ein[399]), .B(ein[398]), .Z(n41284) );
  XOR U45033 ( .A(ein[397]), .B(n41285), .Z(ereg_next[398]) );
  AND U45034 ( .A(mul_pow), .B(n41286), .Z(n41285) );
  XOR U45035 ( .A(ein[398]), .B(ein[397]), .Z(n41286) );
  XOR U45036 ( .A(ein[396]), .B(n41287), .Z(ereg_next[397]) );
  AND U45037 ( .A(mul_pow), .B(n41288), .Z(n41287) );
  XOR U45038 ( .A(ein[397]), .B(ein[396]), .Z(n41288) );
  XOR U45039 ( .A(ein[395]), .B(n41289), .Z(ereg_next[396]) );
  AND U45040 ( .A(mul_pow), .B(n41290), .Z(n41289) );
  XOR U45041 ( .A(ein[396]), .B(ein[395]), .Z(n41290) );
  XOR U45042 ( .A(ein[394]), .B(n41291), .Z(ereg_next[395]) );
  AND U45043 ( .A(mul_pow), .B(n41292), .Z(n41291) );
  XOR U45044 ( .A(ein[395]), .B(ein[394]), .Z(n41292) );
  XOR U45045 ( .A(ein[393]), .B(n41293), .Z(ereg_next[394]) );
  AND U45046 ( .A(mul_pow), .B(n41294), .Z(n41293) );
  XOR U45047 ( .A(ein[394]), .B(ein[393]), .Z(n41294) );
  XOR U45048 ( .A(ein[392]), .B(n41295), .Z(ereg_next[393]) );
  AND U45049 ( .A(mul_pow), .B(n41296), .Z(n41295) );
  XOR U45050 ( .A(ein[393]), .B(ein[392]), .Z(n41296) );
  XOR U45051 ( .A(ein[391]), .B(n41297), .Z(ereg_next[392]) );
  AND U45052 ( .A(mul_pow), .B(n41298), .Z(n41297) );
  XOR U45053 ( .A(ein[392]), .B(ein[391]), .Z(n41298) );
  XOR U45054 ( .A(ein[390]), .B(n41299), .Z(ereg_next[391]) );
  AND U45055 ( .A(mul_pow), .B(n41300), .Z(n41299) );
  XOR U45056 ( .A(ein[391]), .B(ein[390]), .Z(n41300) );
  XOR U45057 ( .A(ein[389]), .B(n41301), .Z(ereg_next[390]) );
  AND U45058 ( .A(mul_pow), .B(n41302), .Z(n41301) );
  XOR U45059 ( .A(ein[390]), .B(ein[389]), .Z(n41302) );
  XOR U45060 ( .A(ein[37]), .B(n41303), .Z(ereg_next[38]) );
  AND U45061 ( .A(mul_pow), .B(n41304), .Z(n41303) );
  XOR U45062 ( .A(ein[38]), .B(ein[37]), .Z(n41304) );
  XOR U45063 ( .A(ein[388]), .B(n41305), .Z(ereg_next[389]) );
  AND U45064 ( .A(mul_pow), .B(n41306), .Z(n41305) );
  XOR U45065 ( .A(ein[389]), .B(ein[388]), .Z(n41306) );
  XOR U45066 ( .A(ein[387]), .B(n41307), .Z(ereg_next[388]) );
  AND U45067 ( .A(mul_pow), .B(n41308), .Z(n41307) );
  XOR U45068 ( .A(ein[388]), .B(ein[387]), .Z(n41308) );
  XOR U45069 ( .A(ein[386]), .B(n41309), .Z(ereg_next[387]) );
  AND U45070 ( .A(mul_pow), .B(n41310), .Z(n41309) );
  XOR U45071 ( .A(ein[387]), .B(ein[386]), .Z(n41310) );
  XOR U45072 ( .A(ein[385]), .B(n41311), .Z(ereg_next[386]) );
  AND U45073 ( .A(mul_pow), .B(n41312), .Z(n41311) );
  XOR U45074 ( .A(ein[386]), .B(ein[385]), .Z(n41312) );
  XOR U45075 ( .A(ein[384]), .B(n41313), .Z(ereg_next[385]) );
  AND U45076 ( .A(mul_pow), .B(n41314), .Z(n41313) );
  XOR U45077 ( .A(ein[385]), .B(ein[384]), .Z(n41314) );
  XOR U45078 ( .A(ein[383]), .B(n41315), .Z(ereg_next[384]) );
  AND U45079 ( .A(mul_pow), .B(n41316), .Z(n41315) );
  XOR U45080 ( .A(ein[384]), .B(ein[383]), .Z(n41316) );
  XOR U45081 ( .A(ein[382]), .B(n41317), .Z(ereg_next[383]) );
  AND U45082 ( .A(mul_pow), .B(n41318), .Z(n41317) );
  XOR U45083 ( .A(ein[383]), .B(ein[382]), .Z(n41318) );
  XOR U45084 ( .A(ein[381]), .B(n41319), .Z(ereg_next[382]) );
  AND U45085 ( .A(mul_pow), .B(n41320), .Z(n41319) );
  XOR U45086 ( .A(ein[382]), .B(ein[381]), .Z(n41320) );
  XOR U45087 ( .A(ein[380]), .B(n41321), .Z(ereg_next[381]) );
  AND U45088 ( .A(mul_pow), .B(n41322), .Z(n41321) );
  XOR U45089 ( .A(ein[381]), .B(ein[380]), .Z(n41322) );
  XOR U45090 ( .A(ein[379]), .B(n41323), .Z(ereg_next[380]) );
  AND U45091 ( .A(mul_pow), .B(n41324), .Z(n41323) );
  XOR U45092 ( .A(ein[380]), .B(ein[379]), .Z(n41324) );
  XOR U45093 ( .A(ein[36]), .B(n41325), .Z(ereg_next[37]) );
  AND U45094 ( .A(mul_pow), .B(n41326), .Z(n41325) );
  XOR U45095 ( .A(ein[37]), .B(ein[36]), .Z(n41326) );
  XOR U45096 ( .A(ein[378]), .B(n41327), .Z(ereg_next[379]) );
  AND U45097 ( .A(mul_pow), .B(n41328), .Z(n41327) );
  XOR U45098 ( .A(ein[379]), .B(ein[378]), .Z(n41328) );
  XOR U45099 ( .A(ein[377]), .B(n41329), .Z(ereg_next[378]) );
  AND U45100 ( .A(mul_pow), .B(n41330), .Z(n41329) );
  XOR U45101 ( .A(ein[378]), .B(ein[377]), .Z(n41330) );
  XOR U45102 ( .A(ein[376]), .B(n41331), .Z(ereg_next[377]) );
  AND U45103 ( .A(mul_pow), .B(n41332), .Z(n41331) );
  XOR U45104 ( .A(ein[377]), .B(ein[376]), .Z(n41332) );
  XOR U45105 ( .A(ein[375]), .B(n41333), .Z(ereg_next[376]) );
  AND U45106 ( .A(mul_pow), .B(n41334), .Z(n41333) );
  XOR U45107 ( .A(ein[376]), .B(ein[375]), .Z(n41334) );
  XOR U45108 ( .A(ein[374]), .B(n41335), .Z(ereg_next[375]) );
  AND U45109 ( .A(mul_pow), .B(n41336), .Z(n41335) );
  XOR U45110 ( .A(ein[375]), .B(ein[374]), .Z(n41336) );
  XOR U45111 ( .A(ein[373]), .B(n41337), .Z(ereg_next[374]) );
  AND U45112 ( .A(mul_pow), .B(n41338), .Z(n41337) );
  XOR U45113 ( .A(ein[374]), .B(ein[373]), .Z(n41338) );
  XOR U45114 ( .A(ein[372]), .B(n41339), .Z(ereg_next[373]) );
  AND U45115 ( .A(mul_pow), .B(n41340), .Z(n41339) );
  XOR U45116 ( .A(ein[373]), .B(ein[372]), .Z(n41340) );
  XOR U45117 ( .A(ein[371]), .B(n41341), .Z(ereg_next[372]) );
  AND U45118 ( .A(mul_pow), .B(n41342), .Z(n41341) );
  XOR U45119 ( .A(ein[372]), .B(ein[371]), .Z(n41342) );
  XOR U45120 ( .A(ein[370]), .B(n41343), .Z(ereg_next[371]) );
  AND U45121 ( .A(mul_pow), .B(n41344), .Z(n41343) );
  XOR U45122 ( .A(ein[371]), .B(ein[370]), .Z(n41344) );
  XOR U45123 ( .A(ein[369]), .B(n41345), .Z(ereg_next[370]) );
  AND U45124 ( .A(mul_pow), .B(n41346), .Z(n41345) );
  XOR U45125 ( .A(ein[370]), .B(ein[369]), .Z(n41346) );
  XOR U45126 ( .A(ein[35]), .B(n41347), .Z(ereg_next[36]) );
  AND U45127 ( .A(mul_pow), .B(n41348), .Z(n41347) );
  XOR U45128 ( .A(ein[36]), .B(ein[35]), .Z(n41348) );
  XOR U45129 ( .A(ein[368]), .B(n41349), .Z(ereg_next[369]) );
  AND U45130 ( .A(mul_pow), .B(n41350), .Z(n41349) );
  XOR U45131 ( .A(ein[369]), .B(ein[368]), .Z(n41350) );
  XOR U45132 ( .A(ein[367]), .B(n41351), .Z(ereg_next[368]) );
  AND U45133 ( .A(mul_pow), .B(n41352), .Z(n41351) );
  XOR U45134 ( .A(ein[368]), .B(ein[367]), .Z(n41352) );
  XOR U45135 ( .A(ein[366]), .B(n41353), .Z(ereg_next[367]) );
  AND U45136 ( .A(mul_pow), .B(n41354), .Z(n41353) );
  XOR U45137 ( .A(ein[367]), .B(ein[366]), .Z(n41354) );
  XOR U45138 ( .A(ein[365]), .B(n41355), .Z(ereg_next[366]) );
  AND U45139 ( .A(mul_pow), .B(n41356), .Z(n41355) );
  XOR U45140 ( .A(ein[366]), .B(ein[365]), .Z(n41356) );
  XOR U45141 ( .A(ein[364]), .B(n41357), .Z(ereg_next[365]) );
  AND U45142 ( .A(mul_pow), .B(n41358), .Z(n41357) );
  XOR U45143 ( .A(ein[365]), .B(ein[364]), .Z(n41358) );
  XOR U45144 ( .A(ein[363]), .B(n41359), .Z(ereg_next[364]) );
  AND U45145 ( .A(mul_pow), .B(n41360), .Z(n41359) );
  XOR U45146 ( .A(ein[364]), .B(ein[363]), .Z(n41360) );
  XOR U45147 ( .A(ein[362]), .B(n41361), .Z(ereg_next[363]) );
  AND U45148 ( .A(mul_pow), .B(n41362), .Z(n41361) );
  XOR U45149 ( .A(ein[363]), .B(ein[362]), .Z(n41362) );
  XOR U45150 ( .A(ein[361]), .B(n41363), .Z(ereg_next[362]) );
  AND U45151 ( .A(mul_pow), .B(n41364), .Z(n41363) );
  XOR U45152 ( .A(ein[362]), .B(ein[361]), .Z(n41364) );
  XOR U45153 ( .A(ein[360]), .B(n41365), .Z(ereg_next[361]) );
  AND U45154 ( .A(mul_pow), .B(n41366), .Z(n41365) );
  XOR U45155 ( .A(ein[361]), .B(ein[360]), .Z(n41366) );
  XOR U45156 ( .A(ein[359]), .B(n41367), .Z(ereg_next[360]) );
  AND U45157 ( .A(mul_pow), .B(n41368), .Z(n41367) );
  XOR U45158 ( .A(ein[360]), .B(ein[359]), .Z(n41368) );
  XOR U45159 ( .A(ein[34]), .B(n41369), .Z(ereg_next[35]) );
  AND U45160 ( .A(mul_pow), .B(n41370), .Z(n41369) );
  XOR U45161 ( .A(ein[35]), .B(ein[34]), .Z(n41370) );
  XOR U45162 ( .A(ein[358]), .B(n41371), .Z(ereg_next[359]) );
  AND U45163 ( .A(mul_pow), .B(n41372), .Z(n41371) );
  XOR U45164 ( .A(ein[359]), .B(ein[358]), .Z(n41372) );
  XOR U45165 ( .A(ein[357]), .B(n41373), .Z(ereg_next[358]) );
  AND U45166 ( .A(mul_pow), .B(n41374), .Z(n41373) );
  XOR U45167 ( .A(ein[358]), .B(ein[357]), .Z(n41374) );
  XOR U45168 ( .A(ein[356]), .B(n41375), .Z(ereg_next[357]) );
  AND U45169 ( .A(mul_pow), .B(n41376), .Z(n41375) );
  XOR U45170 ( .A(ein[357]), .B(ein[356]), .Z(n41376) );
  XOR U45171 ( .A(ein[355]), .B(n41377), .Z(ereg_next[356]) );
  AND U45172 ( .A(mul_pow), .B(n41378), .Z(n41377) );
  XOR U45173 ( .A(ein[356]), .B(ein[355]), .Z(n41378) );
  XOR U45174 ( .A(ein[354]), .B(n41379), .Z(ereg_next[355]) );
  AND U45175 ( .A(mul_pow), .B(n41380), .Z(n41379) );
  XOR U45176 ( .A(ein[355]), .B(ein[354]), .Z(n41380) );
  XOR U45177 ( .A(ein[353]), .B(n41381), .Z(ereg_next[354]) );
  AND U45178 ( .A(mul_pow), .B(n41382), .Z(n41381) );
  XOR U45179 ( .A(ein[354]), .B(ein[353]), .Z(n41382) );
  XOR U45180 ( .A(ein[352]), .B(n41383), .Z(ereg_next[353]) );
  AND U45181 ( .A(mul_pow), .B(n41384), .Z(n41383) );
  XOR U45182 ( .A(ein[353]), .B(ein[352]), .Z(n41384) );
  XOR U45183 ( .A(ein[351]), .B(n41385), .Z(ereg_next[352]) );
  AND U45184 ( .A(mul_pow), .B(n41386), .Z(n41385) );
  XOR U45185 ( .A(ein[352]), .B(ein[351]), .Z(n41386) );
  XOR U45186 ( .A(ein[350]), .B(n41387), .Z(ereg_next[351]) );
  AND U45187 ( .A(mul_pow), .B(n41388), .Z(n41387) );
  XOR U45188 ( .A(ein[351]), .B(ein[350]), .Z(n41388) );
  XOR U45189 ( .A(ein[349]), .B(n41389), .Z(ereg_next[350]) );
  AND U45190 ( .A(mul_pow), .B(n41390), .Z(n41389) );
  XOR U45191 ( .A(ein[350]), .B(ein[349]), .Z(n41390) );
  XOR U45192 ( .A(ein[33]), .B(n41391), .Z(ereg_next[34]) );
  AND U45193 ( .A(mul_pow), .B(n41392), .Z(n41391) );
  XOR U45194 ( .A(ein[34]), .B(ein[33]), .Z(n41392) );
  XOR U45195 ( .A(ein[348]), .B(n41393), .Z(ereg_next[349]) );
  AND U45196 ( .A(mul_pow), .B(n41394), .Z(n41393) );
  XOR U45197 ( .A(ein[349]), .B(ein[348]), .Z(n41394) );
  XOR U45198 ( .A(ein[347]), .B(n41395), .Z(ereg_next[348]) );
  AND U45199 ( .A(mul_pow), .B(n41396), .Z(n41395) );
  XOR U45200 ( .A(ein[348]), .B(ein[347]), .Z(n41396) );
  XOR U45201 ( .A(ein[346]), .B(n41397), .Z(ereg_next[347]) );
  AND U45202 ( .A(mul_pow), .B(n41398), .Z(n41397) );
  XOR U45203 ( .A(ein[347]), .B(ein[346]), .Z(n41398) );
  XOR U45204 ( .A(ein[345]), .B(n41399), .Z(ereg_next[346]) );
  AND U45205 ( .A(mul_pow), .B(n41400), .Z(n41399) );
  XOR U45206 ( .A(ein[346]), .B(ein[345]), .Z(n41400) );
  XOR U45207 ( .A(ein[344]), .B(n41401), .Z(ereg_next[345]) );
  AND U45208 ( .A(mul_pow), .B(n41402), .Z(n41401) );
  XOR U45209 ( .A(ein[345]), .B(ein[344]), .Z(n41402) );
  XOR U45210 ( .A(ein[343]), .B(n41403), .Z(ereg_next[344]) );
  AND U45211 ( .A(mul_pow), .B(n41404), .Z(n41403) );
  XOR U45212 ( .A(ein[344]), .B(ein[343]), .Z(n41404) );
  XOR U45213 ( .A(ein[342]), .B(n41405), .Z(ereg_next[343]) );
  AND U45214 ( .A(mul_pow), .B(n41406), .Z(n41405) );
  XOR U45215 ( .A(ein[343]), .B(ein[342]), .Z(n41406) );
  XOR U45216 ( .A(ein[341]), .B(n41407), .Z(ereg_next[342]) );
  AND U45217 ( .A(mul_pow), .B(n41408), .Z(n41407) );
  XOR U45218 ( .A(ein[342]), .B(ein[341]), .Z(n41408) );
  XOR U45219 ( .A(ein[340]), .B(n41409), .Z(ereg_next[341]) );
  AND U45220 ( .A(mul_pow), .B(n41410), .Z(n41409) );
  XOR U45221 ( .A(ein[341]), .B(ein[340]), .Z(n41410) );
  XOR U45222 ( .A(ein[339]), .B(n41411), .Z(ereg_next[340]) );
  AND U45223 ( .A(mul_pow), .B(n41412), .Z(n41411) );
  XOR U45224 ( .A(ein[340]), .B(ein[339]), .Z(n41412) );
  XOR U45225 ( .A(ein[32]), .B(n41413), .Z(ereg_next[33]) );
  AND U45226 ( .A(mul_pow), .B(n41414), .Z(n41413) );
  XOR U45227 ( .A(ein[33]), .B(ein[32]), .Z(n41414) );
  XOR U45228 ( .A(ein[338]), .B(n41415), .Z(ereg_next[339]) );
  AND U45229 ( .A(mul_pow), .B(n41416), .Z(n41415) );
  XOR U45230 ( .A(ein[339]), .B(ein[338]), .Z(n41416) );
  XOR U45231 ( .A(ein[337]), .B(n41417), .Z(ereg_next[338]) );
  AND U45232 ( .A(mul_pow), .B(n41418), .Z(n41417) );
  XOR U45233 ( .A(ein[338]), .B(ein[337]), .Z(n41418) );
  XOR U45234 ( .A(ein[336]), .B(n41419), .Z(ereg_next[337]) );
  AND U45235 ( .A(mul_pow), .B(n41420), .Z(n41419) );
  XOR U45236 ( .A(ein[337]), .B(ein[336]), .Z(n41420) );
  XOR U45237 ( .A(ein[335]), .B(n41421), .Z(ereg_next[336]) );
  AND U45238 ( .A(mul_pow), .B(n41422), .Z(n41421) );
  XOR U45239 ( .A(ein[336]), .B(ein[335]), .Z(n41422) );
  XOR U45240 ( .A(ein[334]), .B(n41423), .Z(ereg_next[335]) );
  AND U45241 ( .A(mul_pow), .B(n41424), .Z(n41423) );
  XOR U45242 ( .A(ein[335]), .B(ein[334]), .Z(n41424) );
  XOR U45243 ( .A(ein[333]), .B(n41425), .Z(ereg_next[334]) );
  AND U45244 ( .A(mul_pow), .B(n41426), .Z(n41425) );
  XOR U45245 ( .A(ein[334]), .B(ein[333]), .Z(n41426) );
  XOR U45246 ( .A(ein[332]), .B(n41427), .Z(ereg_next[333]) );
  AND U45247 ( .A(mul_pow), .B(n41428), .Z(n41427) );
  XOR U45248 ( .A(ein[333]), .B(ein[332]), .Z(n41428) );
  XOR U45249 ( .A(ein[331]), .B(n41429), .Z(ereg_next[332]) );
  AND U45250 ( .A(mul_pow), .B(n41430), .Z(n41429) );
  XOR U45251 ( .A(ein[332]), .B(ein[331]), .Z(n41430) );
  XOR U45252 ( .A(ein[330]), .B(n41431), .Z(ereg_next[331]) );
  AND U45253 ( .A(mul_pow), .B(n41432), .Z(n41431) );
  XOR U45254 ( .A(ein[331]), .B(ein[330]), .Z(n41432) );
  XOR U45255 ( .A(ein[329]), .B(n41433), .Z(ereg_next[330]) );
  AND U45256 ( .A(mul_pow), .B(n41434), .Z(n41433) );
  XOR U45257 ( .A(ein[330]), .B(ein[329]), .Z(n41434) );
  XOR U45258 ( .A(ein[31]), .B(n41435), .Z(ereg_next[32]) );
  AND U45259 ( .A(mul_pow), .B(n41436), .Z(n41435) );
  XOR U45260 ( .A(ein[32]), .B(ein[31]), .Z(n41436) );
  XOR U45261 ( .A(ein[328]), .B(n41437), .Z(ereg_next[329]) );
  AND U45262 ( .A(mul_pow), .B(n41438), .Z(n41437) );
  XOR U45263 ( .A(ein[329]), .B(ein[328]), .Z(n41438) );
  XOR U45264 ( .A(ein[327]), .B(n41439), .Z(ereg_next[328]) );
  AND U45265 ( .A(mul_pow), .B(n41440), .Z(n41439) );
  XOR U45266 ( .A(ein[328]), .B(ein[327]), .Z(n41440) );
  XOR U45267 ( .A(ein[326]), .B(n41441), .Z(ereg_next[327]) );
  AND U45268 ( .A(mul_pow), .B(n41442), .Z(n41441) );
  XOR U45269 ( .A(ein[327]), .B(ein[326]), .Z(n41442) );
  XOR U45270 ( .A(ein[325]), .B(n41443), .Z(ereg_next[326]) );
  AND U45271 ( .A(mul_pow), .B(n41444), .Z(n41443) );
  XOR U45272 ( .A(ein[326]), .B(ein[325]), .Z(n41444) );
  XOR U45273 ( .A(ein[324]), .B(n41445), .Z(ereg_next[325]) );
  AND U45274 ( .A(mul_pow), .B(n41446), .Z(n41445) );
  XOR U45275 ( .A(ein[325]), .B(ein[324]), .Z(n41446) );
  XOR U45276 ( .A(ein[323]), .B(n41447), .Z(ereg_next[324]) );
  AND U45277 ( .A(mul_pow), .B(n41448), .Z(n41447) );
  XOR U45278 ( .A(ein[324]), .B(ein[323]), .Z(n41448) );
  XOR U45279 ( .A(ein[322]), .B(n41449), .Z(ereg_next[323]) );
  AND U45280 ( .A(mul_pow), .B(n41450), .Z(n41449) );
  XOR U45281 ( .A(ein[323]), .B(ein[322]), .Z(n41450) );
  XOR U45282 ( .A(ein[321]), .B(n41451), .Z(ereg_next[322]) );
  AND U45283 ( .A(mul_pow), .B(n41452), .Z(n41451) );
  XOR U45284 ( .A(ein[322]), .B(ein[321]), .Z(n41452) );
  XOR U45285 ( .A(ein[320]), .B(n41453), .Z(ereg_next[321]) );
  AND U45286 ( .A(mul_pow), .B(n41454), .Z(n41453) );
  XOR U45287 ( .A(ein[321]), .B(ein[320]), .Z(n41454) );
  XOR U45288 ( .A(ein[319]), .B(n41455), .Z(ereg_next[320]) );
  AND U45289 ( .A(mul_pow), .B(n41456), .Z(n41455) );
  XOR U45290 ( .A(ein[320]), .B(ein[319]), .Z(n41456) );
  XOR U45291 ( .A(ein[30]), .B(n41457), .Z(ereg_next[31]) );
  AND U45292 ( .A(mul_pow), .B(n41458), .Z(n41457) );
  XOR U45293 ( .A(ein[31]), .B(ein[30]), .Z(n41458) );
  XOR U45294 ( .A(ein[318]), .B(n41459), .Z(ereg_next[319]) );
  AND U45295 ( .A(mul_pow), .B(n41460), .Z(n41459) );
  XOR U45296 ( .A(ein[319]), .B(ein[318]), .Z(n41460) );
  XOR U45297 ( .A(ein[317]), .B(n41461), .Z(ereg_next[318]) );
  AND U45298 ( .A(mul_pow), .B(n41462), .Z(n41461) );
  XOR U45299 ( .A(ein[318]), .B(ein[317]), .Z(n41462) );
  XOR U45300 ( .A(ein[316]), .B(n41463), .Z(ereg_next[317]) );
  AND U45301 ( .A(mul_pow), .B(n41464), .Z(n41463) );
  XOR U45302 ( .A(ein[317]), .B(ein[316]), .Z(n41464) );
  XOR U45303 ( .A(ein[315]), .B(n41465), .Z(ereg_next[316]) );
  AND U45304 ( .A(mul_pow), .B(n41466), .Z(n41465) );
  XOR U45305 ( .A(ein[316]), .B(ein[315]), .Z(n41466) );
  XOR U45306 ( .A(ein[314]), .B(n41467), .Z(ereg_next[315]) );
  AND U45307 ( .A(mul_pow), .B(n41468), .Z(n41467) );
  XOR U45308 ( .A(ein[315]), .B(ein[314]), .Z(n41468) );
  XOR U45309 ( .A(ein[313]), .B(n41469), .Z(ereg_next[314]) );
  AND U45310 ( .A(mul_pow), .B(n41470), .Z(n41469) );
  XOR U45311 ( .A(ein[314]), .B(ein[313]), .Z(n41470) );
  XOR U45312 ( .A(ein[312]), .B(n41471), .Z(ereg_next[313]) );
  AND U45313 ( .A(mul_pow), .B(n41472), .Z(n41471) );
  XOR U45314 ( .A(ein[313]), .B(ein[312]), .Z(n41472) );
  XOR U45315 ( .A(ein[311]), .B(n41473), .Z(ereg_next[312]) );
  AND U45316 ( .A(mul_pow), .B(n41474), .Z(n41473) );
  XOR U45317 ( .A(ein[312]), .B(ein[311]), .Z(n41474) );
  XOR U45318 ( .A(ein[310]), .B(n41475), .Z(ereg_next[311]) );
  AND U45319 ( .A(mul_pow), .B(n41476), .Z(n41475) );
  XOR U45320 ( .A(ein[311]), .B(ein[310]), .Z(n41476) );
  XOR U45321 ( .A(ein[309]), .B(n41477), .Z(ereg_next[310]) );
  AND U45322 ( .A(mul_pow), .B(n41478), .Z(n41477) );
  XOR U45323 ( .A(ein[310]), .B(ein[309]), .Z(n41478) );
  XOR U45324 ( .A(ein[29]), .B(n41479), .Z(ereg_next[30]) );
  AND U45325 ( .A(mul_pow), .B(n41480), .Z(n41479) );
  XOR U45326 ( .A(ein[30]), .B(ein[29]), .Z(n41480) );
  XOR U45327 ( .A(ein[308]), .B(n41481), .Z(ereg_next[309]) );
  AND U45328 ( .A(mul_pow), .B(n41482), .Z(n41481) );
  XOR U45329 ( .A(ein[309]), .B(ein[308]), .Z(n41482) );
  XOR U45330 ( .A(ein[307]), .B(n41483), .Z(ereg_next[308]) );
  AND U45331 ( .A(mul_pow), .B(n41484), .Z(n41483) );
  XOR U45332 ( .A(ein[308]), .B(ein[307]), .Z(n41484) );
  XOR U45333 ( .A(ein[306]), .B(n41485), .Z(ereg_next[307]) );
  AND U45334 ( .A(mul_pow), .B(n41486), .Z(n41485) );
  XOR U45335 ( .A(ein[307]), .B(ein[306]), .Z(n41486) );
  XOR U45336 ( .A(ein[305]), .B(n41487), .Z(ereg_next[306]) );
  AND U45337 ( .A(mul_pow), .B(n41488), .Z(n41487) );
  XOR U45338 ( .A(ein[306]), .B(ein[305]), .Z(n41488) );
  XOR U45339 ( .A(ein[304]), .B(n41489), .Z(ereg_next[305]) );
  AND U45340 ( .A(mul_pow), .B(n41490), .Z(n41489) );
  XOR U45341 ( .A(ein[305]), .B(ein[304]), .Z(n41490) );
  XOR U45342 ( .A(ein[303]), .B(n41491), .Z(ereg_next[304]) );
  AND U45343 ( .A(mul_pow), .B(n41492), .Z(n41491) );
  XOR U45344 ( .A(ein[304]), .B(ein[303]), .Z(n41492) );
  XOR U45345 ( .A(ein[302]), .B(n41493), .Z(ereg_next[303]) );
  AND U45346 ( .A(mul_pow), .B(n41494), .Z(n41493) );
  XOR U45347 ( .A(ein[303]), .B(ein[302]), .Z(n41494) );
  XOR U45348 ( .A(ein[301]), .B(n41495), .Z(ereg_next[302]) );
  AND U45349 ( .A(mul_pow), .B(n41496), .Z(n41495) );
  XOR U45350 ( .A(ein[302]), .B(ein[301]), .Z(n41496) );
  XOR U45351 ( .A(ein[300]), .B(n41497), .Z(ereg_next[301]) );
  AND U45352 ( .A(mul_pow), .B(n41498), .Z(n41497) );
  XOR U45353 ( .A(ein[301]), .B(ein[300]), .Z(n41498) );
  XOR U45354 ( .A(ein[299]), .B(n41499), .Z(ereg_next[300]) );
  AND U45355 ( .A(mul_pow), .B(n41500), .Z(n41499) );
  XOR U45356 ( .A(ein[300]), .B(ein[299]), .Z(n41500) );
  XOR U45357 ( .A(ein[1]), .B(n41501), .Z(ereg_next[2]) );
  AND U45358 ( .A(mul_pow), .B(n41502), .Z(n41501) );
  XOR U45359 ( .A(ein[2]), .B(ein[1]), .Z(n41502) );
  XOR U45360 ( .A(ein[28]), .B(n41503), .Z(ereg_next[29]) );
  AND U45361 ( .A(mul_pow), .B(n41504), .Z(n41503) );
  XOR U45362 ( .A(ein[29]), .B(ein[28]), .Z(n41504) );
  XOR U45363 ( .A(ein[298]), .B(n41505), .Z(ereg_next[299]) );
  AND U45364 ( .A(mul_pow), .B(n41506), .Z(n41505) );
  XOR U45365 ( .A(ein[299]), .B(ein[298]), .Z(n41506) );
  XOR U45366 ( .A(ein[297]), .B(n41507), .Z(ereg_next[298]) );
  AND U45367 ( .A(mul_pow), .B(n41508), .Z(n41507) );
  XOR U45368 ( .A(ein[298]), .B(ein[297]), .Z(n41508) );
  XOR U45369 ( .A(ein[296]), .B(n41509), .Z(ereg_next[297]) );
  AND U45370 ( .A(mul_pow), .B(n41510), .Z(n41509) );
  XOR U45371 ( .A(ein[297]), .B(ein[296]), .Z(n41510) );
  XOR U45372 ( .A(ein[295]), .B(n41511), .Z(ereg_next[296]) );
  AND U45373 ( .A(mul_pow), .B(n41512), .Z(n41511) );
  XOR U45374 ( .A(ein[296]), .B(ein[295]), .Z(n41512) );
  XOR U45375 ( .A(ein[294]), .B(n41513), .Z(ereg_next[295]) );
  AND U45376 ( .A(mul_pow), .B(n41514), .Z(n41513) );
  XOR U45377 ( .A(ein[295]), .B(ein[294]), .Z(n41514) );
  XOR U45378 ( .A(ein[293]), .B(n41515), .Z(ereg_next[294]) );
  AND U45379 ( .A(mul_pow), .B(n41516), .Z(n41515) );
  XOR U45380 ( .A(ein[294]), .B(ein[293]), .Z(n41516) );
  XOR U45381 ( .A(ein[292]), .B(n41517), .Z(ereg_next[293]) );
  AND U45382 ( .A(mul_pow), .B(n41518), .Z(n41517) );
  XOR U45383 ( .A(ein[293]), .B(ein[292]), .Z(n41518) );
  XOR U45384 ( .A(ein[291]), .B(n41519), .Z(ereg_next[292]) );
  AND U45385 ( .A(mul_pow), .B(n41520), .Z(n41519) );
  XOR U45386 ( .A(ein[292]), .B(ein[291]), .Z(n41520) );
  XOR U45387 ( .A(ein[290]), .B(n41521), .Z(ereg_next[291]) );
  AND U45388 ( .A(mul_pow), .B(n41522), .Z(n41521) );
  XOR U45389 ( .A(ein[291]), .B(ein[290]), .Z(n41522) );
  XOR U45390 ( .A(ein[289]), .B(n41523), .Z(ereg_next[290]) );
  AND U45391 ( .A(mul_pow), .B(n41524), .Z(n41523) );
  XOR U45392 ( .A(ein[290]), .B(ein[289]), .Z(n41524) );
  XOR U45393 ( .A(ein[27]), .B(n41525), .Z(ereg_next[28]) );
  AND U45394 ( .A(mul_pow), .B(n41526), .Z(n41525) );
  XOR U45395 ( .A(ein[28]), .B(ein[27]), .Z(n41526) );
  XOR U45396 ( .A(ein[288]), .B(n41527), .Z(ereg_next[289]) );
  AND U45397 ( .A(mul_pow), .B(n41528), .Z(n41527) );
  XOR U45398 ( .A(ein[289]), .B(ein[288]), .Z(n41528) );
  XOR U45399 ( .A(ein[287]), .B(n41529), .Z(ereg_next[288]) );
  AND U45400 ( .A(mul_pow), .B(n41530), .Z(n41529) );
  XOR U45401 ( .A(ein[288]), .B(ein[287]), .Z(n41530) );
  XOR U45402 ( .A(ein[286]), .B(n41531), .Z(ereg_next[287]) );
  AND U45403 ( .A(mul_pow), .B(n41532), .Z(n41531) );
  XOR U45404 ( .A(ein[287]), .B(ein[286]), .Z(n41532) );
  XOR U45405 ( .A(ein[285]), .B(n41533), .Z(ereg_next[286]) );
  AND U45406 ( .A(mul_pow), .B(n41534), .Z(n41533) );
  XOR U45407 ( .A(ein[286]), .B(ein[285]), .Z(n41534) );
  XOR U45408 ( .A(ein[284]), .B(n41535), .Z(ereg_next[285]) );
  AND U45409 ( .A(mul_pow), .B(n41536), .Z(n41535) );
  XOR U45410 ( .A(ein[285]), .B(ein[284]), .Z(n41536) );
  XOR U45411 ( .A(ein[283]), .B(n41537), .Z(ereg_next[284]) );
  AND U45412 ( .A(mul_pow), .B(n41538), .Z(n41537) );
  XOR U45413 ( .A(ein[284]), .B(ein[283]), .Z(n41538) );
  XOR U45414 ( .A(ein[282]), .B(n41539), .Z(ereg_next[283]) );
  AND U45415 ( .A(mul_pow), .B(n41540), .Z(n41539) );
  XOR U45416 ( .A(ein[283]), .B(ein[282]), .Z(n41540) );
  XOR U45417 ( .A(ein[281]), .B(n41541), .Z(ereg_next[282]) );
  AND U45418 ( .A(mul_pow), .B(n41542), .Z(n41541) );
  XOR U45419 ( .A(ein[282]), .B(ein[281]), .Z(n41542) );
  XOR U45420 ( .A(ein[280]), .B(n41543), .Z(ereg_next[281]) );
  AND U45421 ( .A(mul_pow), .B(n41544), .Z(n41543) );
  XOR U45422 ( .A(ein[281]), .B(ein[280]), .Z(n41544) );
  XOR U45423 ( .A(ein[279]), .B(n41545), .Z(ereg_next[280]) );
  AND U45424 ( .A(mul_pow), .B(n41546), .Z(n41545) );
  XOR U45425 ( .A(ein[280]), .B(ein[279]), .Z(n41546) );
  XOR U45426 ( .A(ein[26]), .B(n41547), .Z(ereg_next[27]) );
  AND U45427 ( .A(mul_pow), .B(n41548), .Z(n41547) );
  XOR U45428 ( .A(ein[27]), .B(ein[26]), .Z(n41548) );
  XOR U45429 ( .A(ein[278]), .B(n41549), .Z(ereg_next[279]) );
  AND U45430 ( .A(mul_pow), .B(n41550), .Z(n41549) );
  XOR U45431 ( .A(ein[279]), .B(ein[278]), .Z(n41550) );
  XOR U45432 ( .A(ein[277]), .B(n41551), .Z(ereg_next[278]) );
  AND U45433 ( .A(mul_pow), .B(n41552), .Z(n41551) );
  XOR U45434 ( .A(ein[278]), .B(ein[277]), .Z(n41552) );
  XOR U45435 ( .A(ein[276]), .B(n41553), .Z(ereg_next[277]) );
  AND U45436 ( .A(mul_pow), .B(n41554), .Z(n41553) );
  XOR U45437 ( .A(ein[277]), .B(ein[276]), .Z(n41554) );
  XOR U45438 ( .A(ein[275]), .B(n41555), .Z(ereg_next[276]) );
  AND U45439 ( .A(mul_pow), .B(n41556), .Z(n41555) );
  XOR U45440 ( .A(ein[276]), .B(ein[275]), .Z(n41556) );
  XOR U45441 ( .A(ein[274]), .B(n41557), .Z(ereg_next[275]) );
  AND U45442 ( .A(mul_pow), .B(n41558), .Z(n41557) );
  XOR U45443 ( .A(ein[275]), .B(ein[274]), .Z(n41558) );
  XOR U45444 ( .A(ein[273]), .B(n41559), .Z(ereg_next[274]) );
  AND U45445 ( .A(mul_pow), .B(n41560), .Z(n41559) );
  XOR U45446 ( .A(ein[274]), .B(ein[273]), .Z(n41560) );
  XOR U45447 ( .A(ein[272]), .B(n41561), .Z(ereg_next[273]) );
  AND U45448 ( .A(mul_pow), .B(n41562), .Z(n41561) );
  XOR U45449 ( .A(ein[273]), .B(ein[272]), .Z(n41562) );
  XOR U45450 ( .A(ein[271]), .B(n41563), .Z(ereg_next[272]) );
  AND U45451 ( .A(mul_pow), .B(n41564), .Z(n41563) );
  XOR U45452 ( .A(ein[272]), .B(ein[271]), .Z(n41564) );
  XOR U45453 ( .A(ein[270]), .B(n41565), .Z(ereg_next[271]) );
  AND U45454 ( .A(mul_pow), .B(n41566), .Z(n41565) );
  XOR U45455 ( .A(ein[271]), .B(ein[270]), .Z(n41566) );
  XOR U45456 ( .A(ein[269]), .B(n41567), .Z(ereg_next[270]) );
  AND U45457 ( .A(mul_pow), .B(n41568), .Z(n41567) );
  XOR U45458 ( .A(ein[270]), .B(ein[269]), .Z(n41568) );
  XOR U45459 ( .A(ein[25]), .B(n41569), .Z(ereg_next[26]) );
  AND U45460 ( .A(mul_pow), .B(n41570), .Z(n41569) );
  XOR U45461 ( .A(ein[26]), .B(ein[25]), .Z(n41570) );
  XOR U45462 ( .A(ein[268]), .B(n41571), .Z(ereg_next[269]) );
  AND U45463 ( .A(mul_pow), .B(n41572), .Z(n41571) );
  XOR U45464 ( .A(ein[269]), .B(ein[268]), .Z(n41572) );
  XOR U45465 ( .A(ein[267]), .B(n41573), .Z(ereg_next[268]) );
  AND U45466 ( .A(mul_pow), .B(n41574), .Z(n41573) );
  XOR U45467 ( .A(ein[268]), .B(ein[267]), .Z(n41574) );
  XOR U45468 ( .A(ein[266]), .B(n41575), .Z(ereg_next[267]) );
  AND U45469 ( .A(mul_pow), .B(n41576), .Z(n41575) );
  XOR U45470 ( .A(ein[267]), .B(ein[266]), .Z(n41576) );
  XOR U45471 ( .A(ein[265]), .B(n41577), .Z(ereg_next[266]) );
  AND U45472 ( .A(mul_pow), .B(n41578), .Z(n41577) );
  XOR U45473 ( .A(ein[266]), .B(ein[265]), .Z(n41578) );
  XOR U45474 ( .A(ein[264]), .B(n41579), .Z(ereg_next[265]) );
  AND U45475 ( .A(mul_pow), .B(n41580), .Z(n41579) );
  XOR U45476 ( .A(ein[265]), .B(ein[264]), .Z(n41580) );
  XOR U45477 ( .A(ein[263]), .B(n41581), .Z(ereg_next[264]) );
  AND U45478 ( .A(mul_pow), .B(n41582), .Z(n41581) );
  XOR U45479 ( .A(ein[264]), .B(ein[263]), .Z(n41582) );
  XOR U45480 ( .A(ein[262]), .B(n41583), .Z(ereg_next[263]) );
  AND U45481 ( .A(mul_pow), .B(n41584), .Z(n41583) );
  XOR U45482 ( .A(ein[263]), .B(ein[262]), .Z(n41584) );
  XOR U45483 ( .A(ein[261]), .B(n41585), .Z(ereg_next[262]) );
  AND U45484 ( .A(mul_pow), .B(n41586), .Z(n41585) );
  XOR U45485 ( .A(ein[262]), .B(ein[261]), .Z(n41586) );
  XOR U45486 ( .A(ein[260]), .B(n41587), .Z(ereg_next[261]) );
  AND U45487 ( .A(mul_pow), .B(n41588), .Z(n41587) );
  XOR U45488 ( .A(ein[261]), .B(ein[260]), .Z(n41588) );
  XOR U45489 ( .A(ein[259]), .B(n41589), .Z(ereg_next[260]) );
  AND U45490 ( .A(mul_pow), .B(n41590), .Z(n41589) );
  XOR U45491 ( .A(ein[260]), .B(ein[259]), .Z(n41590) );
  XOR U45492 ( .A(ein[24]), .B(n41591), .Z(ereg_next[25]) );
  AND U45493 ( .A(mul_pow), .B(n41592), .Z(n41591) );
  XOR U45494 ( .A(ein[25]), .B(ein[24]), .Z(n41592) );
  XOR U45495 ( .A(ein[258]), .B(n41593), .Z(ereg_next[259]) );
  AND U45496 ( .A(mul_pow), .B(n41594), .Z(n41593) );
  XOR U45497 ( .A(ein[259]), .B(ein[258]), .Z(n41594) );
  XOR U45498 ( .A(ein[257]), .B(n41595), .Z(ereg_next[258]) );
  AND U45499 ( .A(mul_pow), .B(n41596), .Z(n41595) );
  XOR U45500 ( .A(ein[258]), .B(ein[257]), .Z(n41596) );
  XOR U45501 ( .A(ein[256]), .B(n41597), .Z(ereg_next[257]) );
  AND U45502 ( .A(mul_pow), .B(n41598), .Z(n41597) );
  XOR U45503 ( .A(ein[257]), .B(ein[256]), .Z(n41598) );
  XOR U45504 ( .A(ein[255]), .B(n41599), .Z(ereg_next[256]) );
  AND U45505 ( .A(mul_pow), .B(n41600), .Z(n41599) );
  XOR U45506 ( .A(ein[256]), .B(ein[255]), .Z(n41600) );
  XOR U45507 ( .A(ein[254]), .B(n41601), .Z(ereg_next[255]) );
  AND U45508 ( .A(mul_pow), .B(n41602), .Z(n41601) );
  XOR U45509 ( .A(ein[255]), .B(ein[254]), .Z(n41602) );
  XOR U45510 ( .A(ein[253]), .B(n41603), .Z(ereg_next[254]) );
  AND U45511 ( .A(mul_pow), .B(n41604), .Z(n41603) );
  XOR U45512 ( .A(ein[254]), .B(ein[253]), .Z(n41604) );
  XOR U45513 ( .A(ein[252]), .B(n41605), .Z(ereg_next[253]) );
  AND U45514 ( .A(mul_pow), .B(n41606), .Z(n41605) );
  XOR U45515 ( .A(ein[253]), .B(ein[252]), .Z(n41606) );
  XOR U45516 ( .A(ein[251]), .B(n41607), .Z(ereg_next[252]) );
  AND U45517 ( .A(mul_pow), .B(n41608), .Z(n41607) );
  XOR U45518 ( .A(ein[252]), .B(ein[251]), .Z(n41608) );
  XOR U45519 ( .A(ein[250]), .B(n41609), .Z(ereg_next[251]) );
  AND U45520 ( .A(mul_pow), .B(n41610), .Z(n41609) );
  XOR U45521 ( .A(ein[251]), .B(ein[250]), .Z(n41610) );
  XOR U45522 ( .A(ein[249]), .B(n41611), .Z(ereg_next[250]) );
  AND U45523 ( .A(mul_pow), .B(n41612), .Z(n41611) );
  XOR U45524 ( .A(ein[250]), .B(ein[249]), .Z(n41612) );
  XOR U45525 ( .A(ein[23]), .B(n41613), .Z(ereg_next[24]) );
  AND U45526 ( .A(mul_pow), .B(n41614), .Z(n41613) );
  XOR U45527 ( .A(ein[24]), .B(ein[23]), .Z(n41614) );
  XOR U45528 ( .A(ein[248]), .B(n41615), .Z(ereg_next[249]) );
  AND U45529 ( .A(mul_pow), .B(n41616), .Z(n41615) );
  XOR U45530 ( .A(ein[249]), .B(ein[248]), .Z(n41616) );
  XOR U45531 ( .A(ein[247]), .B(n41617), .Z(ereg_next[248]) );
  AND U45532 ( .A(mul_pow), .B(n41618), .Z(n41617) );
  XOR U45533 ( .A(ein[248]), .B(ein[247]), .Z(n41618) );
  XOR U45534 ( .A(ein[246]), .B(n41619), .Z(ereg_next[247]) );
  AND U45535 ( .A(mul_pow), .B(n41620), .Z(n41619) );
  XOR U45536 ( .A(ein[247]), .B(ein[246]), .Z(n41620) );
  XOR U45537 ( .A(ein[245]), .B(n41621), .Z(ereg_next[246]) );
  AND U45538 ( .A(mul_pow), .B(n41622), .Z(n41621) );
  XOR U45539 ( .A(ein[246]), .B(ein[245]), .Z(n41622) );
  XOR U45540 ( .A(ein[244]), .B(n41623), .Z(ereg_next[245]) );
  AND U45541 ( .A(mul_pow), .B(n41624), .Z(n41623) );
  XOR U45542 ( .A(ein[245]), .B(ein[244]), .Z(n41624) );
  XOR U45543 ( .A(ein[243]), .B(n41625), .Z(ereg_next[244]) );
  AND U45544 ( .A(mul_pow), .B(n41626), .Z(n41625) );
  XOR U45545 ( .A(ein[244]), .B(ein[243]), .Z(n41626) );
  XOR U45546 ( .A(ein[242]), .B(n41627), .Z(ereg_next[243]) );
  AND U45547 ( .A(mul_pow), .B(n41628), .Z(n41627) );
  XOR U45548 ( .A(ein[243]), .B(ein[242]), .Z(n41628) );
  XOR U45549 ( .A(ein[241]), .B(n41629), .Z(ereg_next[242]) );
  AND U45550 ( .A(mul_pow), .B(n41630), .Z(n41629) );
  XOR U45551 ( .A(ein[242]), .B(ein[241]), .Z(n41630) );
  XOR U45552 ( .A(ein[240]), .B(n41631), .Z(ereg_next[241]) );
  AND U45553 ( .A(mul_pow), .B(n41632), .Z(n41631) );
  XOR U45554 ( .A(ein[241]), .B(ein[240]), .Z(n41632) );
  XOR U45555 ( .A(ein[239]), .B(n41633), .Z(ereg_next[240]) );
  AND U45556 ( .A(mul_pow), .B(n41634), .Z(n41633) );
  XOR U45557 ( .A(ein[240]), .B(ein[239]), .Z(n41634) );
  XOR U45558 ( .A(ein[22]), .B(n41635), .Z(ereg_next[23]) );
  AND U45559 ( .A(mul_pow), .B(n41636), .Z(n41635) );
  XOR U45560 ( .A(ein[23]), .B(ein[22]), .Z(n41636) );
  XOR U45561 ( .A(ein[238]), .B(n41637), .Z(ereg_next[239]) );
  AND U45562 ( .A(mul_pow), .B(n41638), .Z(n41637) );
  XOR U45563 ( .A(ein[239]), .B(ein[238]), .Z(n41638) );
  XOR U45564 ( .A(ein[237]), .B(n41639), .Z(ereg_next[238]) );
  AND U45565 ( .A(mul_pow), .B(n41640), .Z(n41639) );
  XOR U45566 ( .A(ein[238]), .B(ein[237]), .Z(n41640) );
  XOR U45567 ( .A(ein[236]), .B(n41641), .Z(ereg_next[237]) );
  AND U45568 ( .A(mul_pow), .B(n41642), .Z(n41641) );
  XOR U45569 ( .A(ein[237]), .B(ein[236]), .Z(n41642) );
  XOR U45570 ( .A(ein[235]), .B(n41643), .Z(ereg_next[236]) );
  AND U45571 ( .A(mul_pow), .B(n41644), .Z(n41643) );
  XOR U45572 ( .A(ein[236]), .B(ein[235]), .Z(n41644) );
  XOR U45573 ( .A(ein[234]), .B(n41645), .Z(ereg_next[235]) );
  AND U45574 ( .A(mul_pow), .B(n41646), .Z(n41645) );
  XOR U45575 ( .A(ein[235]), .B(ein[234]), .Z(n41646) );
  XOR U45576 ( .A(ein[233]), .B(n41647), .Z(ereg_next[234]) );
  AND U45577 ( .A(mul_pow), .B(n41648), .Z(n41647) );
  XOR U45578 ( .A(ein[234]), .B(ein[233]), .Z(n41648) );
  XOR U45579 ( .A(ein[232]), .B(n41649), .Z(ereg_next[233]) );
  AND U45580 ( .A(mul_pow), .B(n41650), .Z(n41649) );
  XOR U45581 ( .A(ein[233]), .B(ein[232]), .Z(n41650) );
  XOR U45582 ( .A(ein[231]), .B(n41651), .Z(ereg_next[232]) );
  AND U45583 ( .A(mul_pow), .B(n41652), .Z(n41651) );
  XOR U45584 ( .A(ein[232]), .B(ein[231]), .Z(n41652) );
  XOR U45585 ( .A(ein[230]), .B(n41653), .Z(ereg_next[231]) );
  AND U45586 ( .A(mul_pow), .B(n41654), .Z(n41653) );
  XOR U45587 ( .A(ein[231]), .B(ein[230]), .Z(n41654) );
  XOR U45588 ( .A(ein[229]), .B(n41655), .Z(ereg_next[230]) );
  AND U45589 ( .A(mul_pow), .B(n41656), .Z(n41655) );
  XOR U45590 ( .A(ein[230]), .B(ein[229]), .Z(n41656) );
  XOR U45591 ( .A(ein[21]), .B(n41657), .Z(ereg_next[22]) );
  AND U45592 ( .A(mul_pow), .B(n41658), .Z(n41657) );
  XOR U45593 ( .A(ein[22]), .B(ein[21]), .Z(n41658) );
  XOR U45594 ( .A(ein[228]), .B(n41659), .Z(ereg_next[229]) );
  AND U45595 ( .A(mul_pow), .B(n41660), .Z(n41659) );
  XOR U45596 ( .A(ein[229]), .B(ein[228]), .Z(n41660) );
  XOR U45597 ( .A(ein[227]), .B(n41661), .Z(ereg_next[228]) );
  AND U45598 ( .A(mul_pow), .B(n41662), .Z(n41661) );
  XOR U45599 ( .A(ein[228]), .B(ein[227]), .Z(n41662) );
  XOR U45600 ( .A(ein[226]), .B(n41663), .Z(ereg_next[227]) );
  AND U45601 ( .A(mul_pow), .B(n41664), .Z(n41663) );
  XOR U45602 ( .A(ein[227]), .B(ein[226]), .Z(n41664) );
  XOR U45603 ( .A(ein[225]), .B(n41665), .Z(ereg_next[226]) );
  AND U45604 ( .A(mul_pow), .B(n41666), .Z(n41665) );
  XOR U45605 ( .A(ein[226]), .B(ein[225]), .Z(n41666) );
  XOR U45606 ( .A(ein[224]), .B(n41667), .Z(ereg_next[225]) );
  AND U45607 ( .A(mul_pow), .B(n41668), .Z(n41667) );
  XOR U45608 ( .A(ein[225]), .B(ein[224]), .Z(n41668) );
  XOR U45609 ( .A(ein[223]), .B(n41669), .Z(ereg_next[224]) );
  AND U45610 ( .A(mul_pow), .B(n41670), .Z(n41669) );
  XOR U45611 ( .A(ein[224]), .B(ein[223]), .Z(n41670) );
  XOR U45612 ( .A(ein[222]), .B(n41671), .Z(ereg_next[223]) );
  AND U45613 ( .A(mul_pow), .B(n41672), .Z(n41671) );
  XOR U45614 ( .A(ein[223]), .B(ein[222]), .Z(n41672) );
  XOR U45615 ( .A(ein[221]), .B(n41673), .Z(ereg_next[222]) );
  AND U45616 ( .A(mul_pow), .B(n41674), .Z(n41673) );
  XOR U45617 ( .A(ein[222]), .B(ein[221]), .Z(n41674) );
  XOR U45618 ( .A(ein[220]), .B(n41675), .Z(ereg_next[221]) );
  AND U45619 ( .A(mul_pow), .B(n41676), .Z(n41675) );
  XOR U45620 ( .A(ein[221]), .B(ein[220]), .Z(n41676) );
  XOR U45621 ( .A(ein[219]), .B(n41677), .Z(ereg_next[220]) );
  AND U45622 ( .A(mul_pow), .B(n41678), .Z(n41677) );
  XOR U45623 ( .A(ein[220]), .B(ein[219]), .Z(n41678) );
  XOR U45624 ( .A(ein[20]), .B(n41679), .Z(ereg_next[21]) );
  AND U45625 ( .A(mul_pow), .B(n41680), .Z(n41679) );
  XOR U45626 ( .A(ein[21]), .B(ein[20]), .Z(n41680) );
  XOR U45627 ( .A(ein[218]), .B(n41681), .Z(ereg_next[219]) );
  AND U45628 ( .A(mul_pow), .B(n41682), .Z(n41681) );
  XOR U45629 ( .A(ein[219]), .B(ein[218]), .Z(n41682) );
  XOR U45630 ( .A(ein[217]), .B(n41683), .Z(ereg_next[218]) );
  AND U45631 ( .A(mul_pow), .B(n41684), .Z(n41683) );
  XOR U45632 ( .A(ein[218]), .B(ein[217]), .Z(n41684) );
  XOR U45633 ( .A(ein[216]), .B(n41685), .Z(ereg_next[217]) );
  AND U45634 ( .A(mul_pow), .B(n41686), .Z(n41685) );
  XOR U45635 ( .A(ein[217]), .B(ein[216]), .Z(n41686) );
  XOR U45636 ( .A(ein[215]), .B(n41687), .Z(ereg_next[216]) );
  AND U45637 ( .A(mul_pow), .B(n41688), .Z(n41687) );
  XOR U45638 ( .A(ein[216]), .B(ein[215]), .Z(n41688) );
  XOR U45639 ( .A(ein[214]), .B(n41689), .Z(ereg_next[215]) );
  AND U45640 ( .A(mul_pow), .B(n41690), .Z(n41689) );
  XOR U45641 ( .A(ein[215]), .B(ein[214]), .Z(n41690) );
  XOR U45642 ( .A(ein[213]), .B(n41691), .Z(ereg_next[214]) );
  AND U45643 ( .A(mul_pow), .B(n41692), .Z(n41691) );
  XOR U45644 ( .A(ein[214]), .B(ein[213]), .Z(n41692) );
  XOR U45645 ( .A(ein[212]), .B(n41693), .Z(ereg_next[213]) );
  AND U45646 ( .A(mul_pow), .B(n41694), .Z(n41693) );
  XOR U45647 ( .A(ein[213]), .B(ein[212]), .Z(n41694) );
  XOR U45648 ( .A(ein[211]), .B(n41695), .Z(ereg_next[212]) );
  AND U45649 ( .A(mul_pow), .B(n41696), .Z(n41695) );
  XOR U45650 ( .A(ein[212]), .B(ein[211]), .Z(n41696) );
  XOR U45651 ( .A(ein[210]), .B(n41697), .Z(ereg_next[211]) );
  AND U45652 ( .A(mul_pow), .B(n41698), .Z(n41697) );
  XOR U45653 ( .A(ein[211]), .B(ein[210]), .Z(n41698) );
  XOR U45654 ( .A(ein[209]), .B(n41699), .Z(ereg_next[210]) );
  AND U45655 ( .A(mul_pow), .B(n41700), .Z(n41699) );
  XOR U45656 ( .A(ein[210]), .B(ein[209]), .Z(n41700) );
  XOR U45657 ( .A(ein[19]), .B(n41701), .Z(ereg_next[20]) );
  AND U45658 ( .A(mul_pow), .B(n41702), .Z(n41701) );
  XOR U45659 ( .A(ein[20]), .B(ein[19]), .Z(n41702) );
  XOR U45660 ( .A(ein[208]), .B(n41703), .Z(ereg_next[209]) );
  AND U45661 ( .A(mul_pow), .B(n41704), .Z(n41703) );
  XOR U45662 ( .A(ein[209]), .B(ein[208]), .Z(n41704) );
  XOR U45663 ( .A(ein[207]), .B(n41705), .Z(ereg_next[208]) );
  AND U45664 ( .A(mul_pow), .B(n41706), .Z(n41705) );
  XOR U45665 ( .A(ein[208]), .B(ein[207]), .Z(n41706) );
  XOR U45666 ( .A(ein[206]), .B(n41707), .Z(ereg_next[207]) );
  AND U45667 ( .A(mul_pow), .B(n41708), .Z(n41707) );
  XOR U45668 ( .A(ein[207]), .B(ein[206]), .Z(n41708) );
  XOR U45669 ( .A(ein[205]), .B(n41709), .Z(ereg_next[206]) );
  AND U45670 ( .A(mul_pow), .B(n41710), .Z(n41709) );
  XOR U45671 ( .A(ein[206]), .B(ein[205]), .Z(n41710) );
  XOR U45672 ( .A(ein[204]), .B(n41711), .Z(ereg_next[205]) );
  AND U45673 ( .A(mul_pow), .B(n41712), .Z(n41711) );
  XOR U45674 ( .A(ein[205]), .B(ein[204]), .Z(n41712) );
  XOR U45675 ( .A(ein[203]), .B(n41713), .Z(ereg_next[204]) );
  AND U45676 ( .A(mul_pow), .B(n41714), .Z(n41713) );
  XOR U45677 ( .A(ein[204]), .B(ein[203]), .Z(n41714) );
  XOR U45678 ( .A(ein[202]), .B(n41715), .Z(ereg_next[203]) );
  AND U45679 ( .A(mul_pow), .B(n41716), .Z(n41715) );
  XOR U45680 ( .A(ein[203]), .B(ein[202]), .Z(n41716) );
  XOR U45681 ( .A(ein[201]), .B(n41717), .Z(ereg_next[202]) );
  AND U45682 ( .A(mul_pow), .B(n41718), .Z(n41717) );
  XOR U45683 ( .A(ein[202]), .B(ein[201]), .Z(n41718) );
  XOR U45684 ( .A(ein[200]), .B(n41719), .Z(ereg_next[201]) );
  AND U45685 ( .A(mul_pow), .B(n41720), .Z(n41719) );
  XOR U45686 ( .A(ein[201]), .B(ein[200]), .Z(n41720) );
  XOR U45687 ( .A(ein[199]), .B(n41721), .Z(ereg_next[200]) );
  AND U45688 ( .A(mul_pow), .B(n41722), .Z(n41721) );
  XOR U45689 ( .A(ein[200]), .B(ein[199]), .Z(n41722) );
  XOR U45690 ( .A(ein[0]), .B(n41723), .Z(ereg_next[1]) );
  AND U45691 ( .A(mul_pow), .B(n41724), .Z(n41723) );
  XOR U45692 ( .A(ein[1]), .B(ein[0]), .Z(n41724) );
  XOR U45693 ( .A(ein[18]), .B(n41725), .Z(ereg_next[19]) );
  AND U45694 ( .A(mul_pow), .B(n41726), .Z(n41725) );
  XOR U45695 ( .A(ein[19]), .B(ein[18]), .Z(n41726) );
  XOR U45696 ( .A(ein[198]), .B(n41727), .Z(ereg_next[199]) );
  AND U45697 ( .A(mul_pow), .B(n41728), .Z(n41727) );
  XOR U45698 ( .A(ein[199]), .B(ein[198]), .Z(n41728) );
  XOR U45699 ( .A(ein[197]), .B(n41729), .Z(ereg_next[198]) );
  AND U45700 ( .A(mul_pow), .B(n41730), .Z(n41729) );
  XOR U45701 ( .A(ein[198]), .B(ein[197]), .Z(n41730) );
  XOR U45702 ( .A(ein[196]), .B(n41731), .Z(ereg_next[197]) );
  AND U45703 ( .A(mul_pow), .B(n41732), .Z(n41731) );
  XOR U45704 ( .A(ein[197]), .B(ein[196]), .Z(n41732) );
  XOR U45705 ( .A(ein[195]), .B(n41733), .Z(ereg_next[196]) );
  AND U45706 ( .A(mul_pow), .B(n41734), .Z(n41733) );
  XOR U45707 ( .A(ein[196]), .B(ein[195]), .Z(n41734) );
  XOR U45708 ( .A(ein[194]), .B(n41735), .Z(ereg_next[195]) );
  AND U45709 ( .A(mul_pow), .B(n41736), .Z(n41735) );
  XOR U45710 ( .A(ein[195]), .B(ein[194]), .Z(n41736) );
  XOR U45711 ( .A(ein[193]), .B(n41737), .Z(ereg_next[194]) );
  AND U45712 ( .A(mul_pow), .B(n41738), .Z(n41737) );
  XOR U45713 ( .A(ein[194]), .B(ein[193]), .Z(n41738) );
  XOR U45714 ( .A(ein[192]), .B(n41739), .Z(ereg_next[193]) );
  AND U45715 ( .A(mul_pow), .B(n41740), .Z(n41739) );
  XOR U45716 ( .A(ein[193]), .B(ein[192]), .Z(n41740) );
  XOR U45717 ( .A(ein[191]), .B(n41741), .Z(ereg_next[192]) );
  AND U45718 ( .A(mul_pow), .B(n41742), .Z(n41741) );
  XOR U45719 ( .A(ein[192]), .B(ein[191]), .Z(n41742) );
  XOR U45720 ( .A(ein[190]), .B(n41743), .Z(ereg_next[191]) );
  AND U45721 ( .A(mul_pow), .B(n41744), .Z(n41743) );
  XOR U45722 ( .A(ein[191]), .B(ein[190]), .Z(n41744) );
  XOR U45723 ( .A(ein[189]), .B(n41745), .Z(ereg_next[190]) );
  AND U45724 ( .A(mul_pow), .B(n41746), .Z(n41745) );
  XOR U45725 ( .A(ein[190]), .B(ein[189]), .Z(n41746) );
  XOR U45726 ( .A(ein[17]), .B(n41747), .Z(ereg_next[18]) );
  AND U45727 ( .A(mul_pow), .B(n41748), .Z(n41747) );
  XOR U45728 ( .A(ein[18]), .B(ein[17]), .Z(n41748) );
  XOR U45729 ( .A(ein[188]), .B(n41749), .Z(ereg_next[189]) );
  AND U45730 ( .A(mul_pow), .B(n41750), .Z(n41749) );
  XOR U45731 ( .A(ein[189]), .B(ein[188]), .Z(n41750) );
  XOR U45732 ( .A(ein[187]), .B(n41751), .Z(ereg_next[188]) );
  AND U45733 ( .A(mul_pow), .B(n41752), .Z(n41751) );
  XOR U45734 ( .A(ein[188]), .B(ein[187]), .Z(n41752) );
  XOR U45735 ( .A(ein[186]), .B(n41753), .Z(ereg_next[187]) );
  AND U45736 ( .A(mul_pow), .B(n41754), .Z(n41753) );
  XOR U45737 ( .A(ein[187]), .B(ein[186]), .Z(n41754) );
  XOR U45738 ( .A(ein[185]), .B(n41755), .Z(ereg_next[186]) );
  AND U45739 ( .A(mul_pow), .B(n41756), .Z(n41755) );
  XOR U45740 ( .A(ein[186]), .B(ein[185]), .Z(n41756) );
  XOR U45741 ( .A(ein[184]), .B(n41757), .Z(ereg_next[185]) );
  AND U45742 ( .A(mul_pow), .B(n41758), .Z(n41757) );
  XOR U45743 ( .A(ein[185]), .B(ein[184]), .Z(n41758) );
  XOR U45744 ( .A(ein[183]), .B(n41759), .Z(ereg_next[184]) );
  AND U45745 ( .A(mul_pow), .B(n41760), .Z(n41759) );
  XOR U45746 ( .A(ein[184]), .B(ein[183]), .Z(n41760) );
  XOR U45747 ( .A(ein[182]), .B(n41761), .Z(ereg_next[183]) );
  AND U45748 ( .A(mul_pow), .B(n41762), .Z(n41761) );
  XOR U45749 ( .A(ein[183]), .B(ein[182]), .Z(n41762) );
  XOR U45750 ( .A(ein[181]), .B(n41763), .Z(ereg_next[182]) );
  AND U45751 ( .A(mul_pow), .B(n41764), .Z(n41763) );
  XOR U45752 ( .A(ein[182]), .B(ein[181]), .Z(n41764) );
  XOR U45753 ( .A(ein[180]), .B(n41765), .Z(ereg_next[181]) );
  AND U45754 ( .A(mul_pow), .B(n41766), .Z(n41765) );
  XOR U45755 ( .A(ein[181]), .B(ein[180]), .Z(n41766) );
  XOR U45756 ( .A(ein[179]), .B(n41767), .Z(ereg_next[180]) );
  AND U45757 ( .A(mul_pow), .B(n41768), .Z(n41767) );
  XOR U45758 ( .A(ein[180]), .B(ein[179]), .Z(n41768) );
  XOR U45759 ( .A(ein[16]), .B(n41769), .Z(ereg_next[17]) );
  AND U45760 ( .A(mul_pow), .B(n41770), .Z(n41769) );
  XOR U45761 ( .A(ein[17]), .B(ein[16]), .Z(n41770) );
  XOR U45762 ( .A(ein[178]), .B(n41771), .Z(ereg_next[179]) );
  AND U45763 ( .A(mul_pow), .B(n41772), .Z(n41771) );
  XOR U45764 ( .A(ein[179]), .B(ein[178]), .Z(n41772) );
  XOR U45765 ( .A(ein[177]), .B(n41773), .Z(ereg_next[178]) );
  AND U45766 ( .A(mul_pow), .B(n41774), .Z(n41773) );
  XOR U45767 ( .A(ein[178]), .B(ein[177]), .Z(n41774) );
  XOR U45768 ( .A(ein[176]), .B(n41775), .Z(ereg_next[177]) );
  AND U45769 ( .A(mul_pow), .B(n41776), .Z(n41775) );
  XOR U45770 ( .A(ein[177]), .B(ein[176]), .Z(n41776) );
  XOR U45771 ( .A(ein[175]), .B(n41777), .Z(ereg_next[176]) );
  AND U45772 ( .A(mul_pow), .B(n41778), .Z(n41777) );
  XOR U45773 ( .A(ein[176]), .B(ein[175]), .Z(n41778) );
  XOR U45774 ( .A(ein[174]), .B(n41779), .Z(ereg_next[175]) );
  AND U45775 ( .A(mul_pow), .B(n41780), .Z(n41779) );
  XOR U45776 ( .A(ein[175]), .B(ein[174]), .Z(n41780) );
  XOR U45777 ( .A(ein[173]), .B(n41781), .Z(ereg_next[174]) );
  AND U45778 ( .A(mul_pow), .B(n41782), .Z(n41781) );
  XOR U45779 ( .A(ein[174]), .B(ein[173]), .Z(n41782) );
  XOR U45780 ( .A(ein[172]), .B(n41783), .Z(ereg_next[173]) );
  AND U45781 ( .A(mul_pow), .B(n41784), .Z(n41783) );
  XOR U45782 ( .A(ein[173]), .B(ein[172]), .Z(n41784) );
  XOR U45783 ( .A(ein[171]), .B(n41785), .Z(ereg_next[172]) );
  AND U45784 ( .A(mul_pow), .B(n41786), .Z(n41785) );
  XOR U45785 ( .A(ein[172]), .B(ein[171]), .Z(n41786) );
  XOR U45786 ( .A(ein[170]), .B(n41787), .Z(ereg_next[171]) );
  AND U45787 ( .A(mul_pow), .B(n41788), .Z(n41787) );
  XOR U45788 ( .A(ein[171]), .B(ein[170]), .Z(n41788) );
  XOR U45789 ( .A(ein[169]), .B(n41789), .Z(ereg_next[170]) );
  AND U45790 ( .A(mul_pow), .B(n41790), .Z(n41789) );
  XOR U45791 ( .A(ein[170]), .B(ein[169]), .Z(n41790) );
  XOR U45792 ( .A(ein[15]), .B(n41791), .Z(ereg_next[16]) );
  AND U45793 ( .A(mul_pow), .B(n41792), .Z(n41791) );
  XOR U45794 ( .A(ein[16]), .B(ein[15]), .Z(n41792) );
  XOR U45795 ( .A(ein[168]), .B(n41793), .Z(ereg_next[169]) );
  AND U45796 ( .A(mul_pow), .B(n41794), .Z(n41793) );
  XOR U45797 ( .A(ein[169]), .B(ein[168]), .Z(n41794) );
  XOR U45798 ( .A(ein[167]), .B(n41795), .Z(ereg_next[168]) );
  AND U45799 ( .A(mul_pow), .B(n41796), .Z(n41795) );
  XOR U45800 ( .A(ein[168]), .B(ein[167]), .Z(n41796) );
  XOR U45801 ( .A(ein[166]), .B(n41797), .Z(ereg_next[167]) );
  AND U45802 ( .A(mul_pow), .B(n41798), .Z(n41797) );
  XOR U45803 ( .A(ein[167]), .B(ein[166]), .Z(n41798) );
  XOR U45804 ( .A(ein[165]), .B(n41799), .Z(ereg_next[166]) );
  AND U45805 ( .A(mul_pow), .B(n41800), .Z(n41799) );
  XOR U45806 ( .A(ein[166]), .B(ein[165]), .Z(n41800) );
  XOR U45807 ( .A(ein[164]), .B(n41801), .Z(ereg_next[165]) );
  AND U45808 ( .A(mul_pow), .B(n41802), .Z(n41801) );
  XOR U45809 ( .A(ein[165]), .B(ein[164]), .Z(n41802) );
  XOR U45810 ( .A(ein[163]), .B(n41803), .Z(ereg_next[164]) );
  AND U45811 ( .A(mul_pow), .B(n41804), .Z(n41803) );
  XOR U45812 ( .A(ein[164]), .B(ein[163]), .Z(n41804) );
  XOR U45813 ( .A(ein[162]), .B(n41805), .Z(ereg_next[163]) );
  AND U45814 ( .A(mul_pow), .B(n41806), .Z(n41805) );
  XOR U45815 ( .A(ein[163]), .B(ein[162]), .Z(n41806) );
  XOR U45816 ( .A(ein[161]), .B(n41807), .Z(ereg_next[162]) );
  AND U45817 ( .A(mul_pow), .B(n41808), .Z(n41807) );
  XOR U45818 ( .A(ein[162]), .B(ein[161]), .Z(n41808) );
  XOR U45819 ( .A(ein[160]), .B(n41809), .Z(ereg_next[161]) );
  AND U45820 ( .A(mul_pow), .B(n41810), .Z(n41809) );
  XOR U45821 ( .A(ein[161]), .B(ein[160]), .Z(n41810) );
  XOR U45822 ( .A(ein[159]), .B(n41811), .Z(ereg_next[160]) );
  AND U45823 ( .A(mul_pow), .B(n41812), .Z(n41811) );
  XOR U45824 ( .A(ein[160]), .B(ein[159]), .Z(n41812) );
  XOR U45825 ( .A(ein[14]), .B(n41813), .Z(ereg_next[15]) );
  AND U45826 ( .A(mul_pow), .B(n41814), .Z(n41813) );
  XOR U45827 ( .A(ein[15]), .B(ein[14]), .Z(n41814) );
  XOR U45828 ( .A(ein[158]), .B(n41815), .Z(ereg_next[159]) );
  AND U45829 ( .A(mul_pow), .B(n41816), .Z(n41815) );
  XOR U45830 ( .A(ein[159]), .B(ein[158]), .Z(n41816) );
  XOR U45831 ( .A(ein[157]), .B(n41817), .Z(ereg_next[158]) );
  AND U45832 ( .A(mul_pow), .B(n41818), .Z(n41817) );
  XOR U45833 ( .A(ein[158]), .B(ein[157]), .Z(n41818) );
  XOR U45834 ( .A(ein[156]), .B(n41819), .Z(ereg_next[157]) );
  AND U45835 ( .A(mul_pow), .B(n41820), .Z(n41819) );
  XOR U45836 ( .A(ein[157]), .B(ein[156]), .Z(n41820) );
  XOR U45837 ( .A(ein[155]), .B(n41821), .Z(ereg_next[156]) );
  AND U45838 ( .A(mul_pow), .B(n41822), .Z(n41821) );
  XOR U45839 ( .A(ein[156]), .B(ein[155]), .Z(n41822) );
  XOR U45840 ( .A(ein[154]), .B(n41823), .Z(ereg_next[155]) );
  AND U45841 ( .A(mul_pow), .B(n41824), .Z(n41823) );
  XOR U45842 ( .A(ein[155]), .B(ein[154]), .Z(n41824) );
  XOR U45843 ( .A(ein[153]), .B(n41825), .Z(ereg_next[154]) );
  AND U45844 ( .A(mul_pow), .B(n41826), .Z(n41825) );
  XOR U45845 ( .A(ein[154]), .B(ein[153]), .Z(n41826) );
  XOR U45846 ( .A(ein[152]), .B(n41827), .Z(ereg_next[153]) );
  AND U45847 ( .A(mul_pow), .B(n41828), .Z(n41827) );
  XOR U45848 ( .A(ein[153]), .B(ein[152]), .Z(n41828) );
  XOR U45849 ( .A(ein[151]), .B(n41829), .Z(ereg_next[152]) );
  AND U45850 ( .A(mul_pow), .B(n41830), .Z(n41829) );
  XOR U45851 ( .A(ein[152]), .B(ein[151]), .Z(n41830) );
  XOR U45852 ( .A(ein[150]), .B(n41831), .Z(ereg_next[151]) );
  AND U45853 ( .A(mul_pow), .B(n41832), .Z(n41831) );
  XOR U45854 ( .A(ein[151]), .B(ein[150]), .Z(n41832) );
  XOR U45855 ( .A(ein[149]), .B(n41833), .Z(ereg_next[150]) );
  AND U45856 ( .A(mul_pow), .B(n41834), .Z(n41833) );
  XOR U45857 ( .A(ein[150]), .B(ein[149]), .Z(n41834) );
  XOR U45858 ( .A(ein[13]), .B(n41835), .Z(ereg_next[14]) );
  AND U45859 ( .A(mul_pow), .B(n41836), .Z(n41835) );
  XOR U45860 ( .A(ein[14]), .B(ein[13]), .Z(n41836) );
  XOR U45861 ( .A(ein[148]), .B(n41837), .Z(ereg_next[149]) );
  AND U45862 ( .A(mul_pow), .B(n41838), .Z(n41837) );
  XOR U45863 ( .A(ein[149]), .B(ein[148]), .Z(n41838) );
  XOR U45864 ( .A(ein[147]), .B(n41839), .Z(ereg_next[148]) );
  AND U45865 ( .A(mul_pow), .B(n41840), .Z(n41839) );
  XOR U45866 ( .A(ein[148]), .B(ein[147]), .Z(n41840) );
  XOR U45867 ( .A(ein[146]), .B(n41841), .Z(ereg_next[147]) );
  AND U45868 ( .A(mul_pow), .B(n41842), .Z(n41841) );
  XOR U45869 ( .A(ein[147]), .B(ein[146]), .Z(n41842) );
  XOR U45870 ( .A(ein[145]), .B(n41843), .Z(ereg_next[146]) );
  AND U45871 ( .A(mul_pow), .B(n41844), .Z(n41843) );
  XOR U45872 ( .A(ein[146]), .B(ein[145]), .Z(n41844) );
  XOR U45873 ( .A(ein[144]), .B(n41845), .Z(ereg_next[145]) );
  AND U45874 ( .A(mul_pow), .B(n41846), .Z(n41845) );
  XOR U45875 ( .A(ein[145]), .B(ein[144]), .Z(n41846) );
  XOR U45876 ( .A(ein[143]), .B(n41847), .Z(ereg_next[144]) );
  AND U45877 ( .A(mul_pow), .B(n41848), .Z(n41847) );
  XOR U45878 ( .A(ein[144]), .B(ein[143]), .Z(n41848) );
  XOR U45879 ( .A(ein[142]), .B(n41849), .Z(ereg_next[143]) );
  AND U45880 ( .A(mul_pow), .B(n41850), .Z(n41849) );
  XOR U45881 ( .A(ein[143]), .B(ein[142]), .Z(n41850) );
  XOR U45882 ( .A(ein[141]), .B(n41851), .Z(ereg_next[142]) );
  AND U45883 ( .A(mul_pow), .B(n41852), .Z(n41851) );
  XOR U45884 ( .A(ein[142]), .B(ein[141]), .Z(n41852) );
  XOR U45885 ( .A(ein[140]), .B(n41853), .Z(ereg_next[141]) );
  AND U45886 ( .A(mul_pow), .B(n41854), .Z(n41853) );
  XOR U45887 ( .A(ein[141]), .B(ein[140]), .Z(n41854) );
  XOR U45888 ( .A(ein[139]), .B(n41855), .Z(ereg_next[140]) );
  AND U45889 ( .A(mul_pow), .B(n41856), .Z(n41855) );
  XOR U45890 ( .A(ein[140]), .B(ein[139]), .Z(n41856) );
  XOR U45891 ( .A(ein[12]), .B(n41857), .Z(ereg_next[13]) );
  AND U45892 ( .A(mul_pow), .B(n41858), .Z(n41857) );
  XOR U45893 ( .A(ein[13]), .B(ein[12]), .Z(n41858) );
  XOR U45894 ( .A(ein[138]), .B(n41859), .Z(ereg_next[139]) );
  AND U45895 ( .A(mul_pow), .B(n41860), .Z(n41859) );
  XOR U45896 ( .A(ein[139]), .B(ein[138]), .Z(n41860) );
  XOR U45897 ( .A(ein[137]), .B(n41861), .Z(ereg_next[138]) );
  AND U45898 ( .A(mul_pow), .B(n41862), .Z(n41861) );
  XOR U45899 ( .A(ein[138]), .B(ein[137]), .Z(n41862) );
  XOR U45900 ( .A(ein[136]), .B(n41863), .Z(ereg_next[137]) );
  AND U45901 ( .A(mul_pow), .B(n41864), .Z(n41863) );
  XOR U45902 ( .A(ein[137]), .B(ein[136]), .Z(n41864) );
  XOR U45903 ( .A(ein[135]), .B(n41865), .Z(ereg_next[136]) );
  AND U45904 ( .A(mul_pow), .B(n41866), .Z(n41865) );
  XOR U45905 ( .A(ein[136]), .B(ein[135]), .Z(n41866) );
  XOR U45906 ( .A(ein[134]), .B(n41867), .Z(ereg_next[135]) );
  AND U45907 ( .A(mul_pow), .B(n41868), .Z(n41867) );
  XOR U45908 ( .A(ein[135]), .B(ein[134]), .Z(n41868) );
  XOR U45909 ( .A(ein[133]), .B(n41869), .Z(ereg_next[134]) );
  AND U45910 ( .A(mul_pow), .B(n41870), .Z(n41869) );
  XOR U45911 ( .A(ein[134]), .B(ein[133]), .Z(n41870) );
  XOR U45912 ( .A(ein[132]), .B(n41871), .Z(ereg_next[133]) );
  AND U45913 ( .A(mul_pow), .B(n41872), .Z(n41871) );
  XOR U45914 ( .A(ein[133]), .B(ein[132]), .Z(n41872) );
  XOR U45915 ( .A(ein[131]), .B(n41873), .Z(ereg_next[132]) );
  AND U45916 ( .A(mul_pow), .B(n41874), .Z(n41873) );
  XOR U45917 ( .A(ein[132]), .B(ein[131]), .Z(n41874) );
  XOR U45918 ( .A(ein[130]), .B(n41875), .Z(ereg_next[131]) );
  AND U45919 ( .A(mul_pow), .B(n41876), .Z(n41875) );
  XOR U45920 ( .A(ein[131]), .B(ein[130]), .Z(n41876) );
  XOR U45921 ( .A(ein[129]), .B(n41877), .Z(ereg_next[130]) );
  AND U45922 ( .A(mul_pow), .B(n41878), .Z(n41877) );
  XOR U45923 ( .A(ein[130]), .B(ein[129]), .Z(n41878) );
  XOR U45924 ( .A(ein[11]), .B(n41879), .Z(ereg_next[12]) );
  AND U45925 ( .A(mul_pow), .B(n41880), .Z(n41879) );
  XOR U45926 ( .A(ein[12]), .B(ein[11]), .Z(n41880) );
  XOR U45927 ( .A(ein[128]), .B(n41881), .Z(ereg_next[129]) );
  AND U45928 ( .A(mul_pow), .B(n41882), .Z(n41881) );
  XOR U45929 ( .A(ein[129]), .B(ein[128]), .Z(n41882) );
  XOR U45930 ( .A(ein[127]), .B(n41883), .Z(ereg_next[128]) );
  AND U45931 ( .A(mul_pow), .B(n41884), .Z(n41883) );
  XOR U45932 ( .A(ein[128]), .B(ein[127]), .Z(n41884) );
  XOR U45933 ( .A(ein[126]), .B(n41885), .Z(ereg_next[127]) );
  AND U45934 ( .A(mul_pow), .B(n41886), .Z(n41885) );
  XOR U45935 ( .A(ein[127]), .B(ein[126]), .Z(n41886) );
  XOR U45936 ( .A(ein[125]), .B(n41887), .Z(ereg_next[126]) );
  AND U45937 ( .A(mul_pow), .B(n41888), .Z(n41887) );
  XOR U45938 ( .A(ein[126]), .B(ein[125]), .Z(n41888) );
  XOR U45939 ( .A(ein[124]), .B(n41889), .Z(ereg_next[125]) );
  AND U45940 ( .A(mul_pow), .B(n41890), .Z(n41889) );
  XOR U45941 ( .A(ein[125]), .B(ein[124]), .Z(n41890) );
  XOR U45942 ( .A(ein[123]), .B(n41891), .Z(ereg_next[124]) );
  AND U45943 ( .A(mul_pow), .B(n41892), .Z(n41891) );
  XOR U45944 ( .A(ein[124]), .B(ein[123]), .Z(n41892) );
  XOR U45945 ( .A(ein[122]), .B(n41893), .Z(ereg_next[123]) );
  AND U45946 ( .A(mul_pow), .B(n41894), .Z(n41893) );
  XOR U45947 ( .A(ein[123]), .B(ein[122]), .Z(n41894) );
  XOR U45948 ( .A(ein[121]), .B(n41895), .Z(ereg_next[122]) );
  AND U45949 ( .A(mul_pow), .B(n41896), .Z(n41895) );
  XOR U45950 ( .A(ein[122]), .B(ein[121]), .Z(n41896) );
  XOR U45951 ( .A(ein[120]), .B(n41897), .Z(ereg_next[121]) );
  AND U45952 ( .A(mul_pow), .B(n41898), .Z(n41897) );
  XOR U45953 ( .A(ein[121]), .B(ein[120]), .Z(n41898) );
  XOR U45954 ( .A(ein[119]), .B(n41899), .Z(ereg_next[120]) );
  AND U45955 ( .A(mul_pow), .B(n41900), .Z(n41899) );
  XOR U45956 ( .A(ein[120]), .B(ein[119]), .Z(n41900) );
  XOR U45957 ( .A(ein[10]), .B(n41901), .Z(ereg_next[11]) );
  AND U45958 ( .A(mul_pow), .B(n41902), .Z(n41901) );
  XOR U45959 ( .A(ein[11]), .B(ein[10]), .Z(n41902) );
  XOR U45960 ( .A(ein[118]), .B(n41903), .Z(ereg_next[119]) );
  AND U45961 ( .A(mul_pow), .B(n41904), .Z(n41903) );
  XOR U45962 ( .A(ein[119]), .B(ein[118]), .Z(n41904) );
  XOR U45963 ( .A(ein[117]), .B(n41905), .Z(ereg_next[118]) );
  AND U45964 ( .A(mul_pow), .B(n41906), .Z(n41905) );
  XOR U45965 ( .A(ein[118]), .B(ein[117]), .Z(n41906) );
  XOR U45966 ( .A(ein[116]), .B(n41907), .Z(ereg_next[117]) );
  AND U45967 ( .A(mul_pow), .B(n41908), .Z(n41907) );
  XOR U45968 ( .A(ein[117]), .B(ein[116]), .Z(n41908) );
  XOR U45969 ( .A(ein[115]), .B(n41909), .Z(ereg_next[116]) );
  AND U45970 ( .A(mul_pow), .B(n41910), .Z(n41909) );
  XOR U45971 ( .A(ein[116]), .B(ein[115]), .Z(n41910) );
  XOR U45972 ( .A(ein[114]), .B(n41911), .Z(ereg_next[115]) );
  AND U45973 ( .A(mul_pow), .B(n41912), .Z(n41911) );
  XOR U45974 ( .A(ein[115]), .B(ein[114]), .Z(n41912) );
  XOR U45975 ( .A(ein[113]), .B(n41913), .Z(ereg_next[114]) );
  AND U45976 ( .A(mul_pow), .B(n41914), .Z(n41913) );
  XOR U45977 ( .A(ein[114]), .B(ein[113]), .Z(n41914) );
  XOR U45978 ( .A(ein[112]), .B(n41915), .Z(ereg_next[113]) );
  AND U45979 ( .A(mul_pow), .B(n41916), .Z(n41915) );
  XOR U45980 ( .A(ein[113]), .B(ein[112]), .Z(n41916) );
  XOR U45981 ( .A(ein[111]), .B(n41917), .Z(ereg_next[112]) );
  AND U45982 ( .A(mul_pow), .B(n41918), .Z(n41917) );
  XOR U45983 ( .A(ein[112]), .B(ein[111]), .Z(n41918) );
  XOR U45984 ( .A(ein[110]), .B(n41919), .Z(ereg_next[111]) );
  AND U45985 ( .A(mul_pow), .B(n41920), .Z(n41919) );
  XOR U45986 ( .A(ein[111]), .B(ein[110]), .Z(n41920) );
  XOR U45987 ( .A(ein[109]), .B(n41921), .Z(ereg_next[110]) );
  AND U45988 ( .A(mul_pow), .B(n41922), .Z(n41921) );
  XOR U45989 ( .A(ein[110]), .B(ein[109]), .Z(n41922) );
  XOR U45990 ( .A(ein[9]), .B(n41923), .Z(ereg_next[10]) );
  AND U45991 ( .A(mul_pow), .B(n41924), .Z(n41923) );
  XOR U45992 ( .A(ein[9]), .B(ein[10]), .Z(n41924) );
  XOR U45993 ( .A(ein[108]), .B(n41925), .Z(ereg_next[109]) );
  AND U45994 ( .A(mul_pow), .B(n41926), .Z(n41925) );
  XOR U45995 ( .A(ein[109]), .B(ein[108]), .Z(n41926) );
  XOR U45996 ( .A(ein[107]), .B(n41927), .Z(ereg_next[108]) );
  AND U45997 ( .A(mul_pow), .B(n41928), .Z(n41927) );
  XOR U45998 ( .A(ein[108]), .B(ein[107]), .Z(n41928) );
  XOR U45999 ( .A(ein[106]), .B(n41929), .Z(ereg_next[107]) );
  AND U46000 ( .A(mul_pow), .B(n41930), .Z(n41929) );
  XOR U46001 ( .A(ein[107]), .B(ein[106]), .Z(n41930) );
  XOR U46002 ( .A(ein[105]), .B(n41931), .Z(ereg_next[106]) );
  AND U46003 ( .A(mul_pow), .B(n41932), .Z(n41931) );
  XOR U46004 ( .A(ein[106]), .B(ein[105]), .Z(n41932) );
  XOR U46005 ( .A(ein[104]), .B(n41933), .Z(ereg_next[105]) );
  AND U46006 ( .A(mul_pow), .B(n41934), .Z(n41933) );
  XOR U46007 ( .A(ein[105]), .B(ein[104]), .Z(n41934) );
  XOR U46008 ( .A(ein[103]), .B(n41935), .Z(ereg_next[104]) );
  AND U46009 ( .A(mul_pow), .B(n41936), .Z(n41935) );
  XOR U46010 ( .A(ein[104]), .B(ein[103]), .Z(n41936) );
  XOR U46011 ( .A(ein[102]), .B(n41937), .Z(ereg_next[103]) );
  AND U46012 ( .A(mul_pow), .B(n41938), .Z(n41937) );
  XOR U46013 ( .A(ein[103]), .B(ein[102]), .Z(n41938) );
  XOR U46014 ( .A(ein[101]), .B(n41939), .Z(ereg_next[102]) );
  AND U46015 ( .A(mul_pow), .B(n41940), .Z(n41939) );
  XOR U46016 ( .A(ein[102]), .B(ein[101]), .Z(n41940) );
  XOR U46017 ( .A(ein[1022]), .B(n41941), .Z(ereg_next[1023]) );
  AND U46018 ( .A(mul_pow), .B(n41942), .Z(n41941) );
  XOR U46019 ( .A(ein[1023]), .B(ein[1022]), .Z(n41942) );
  XOR U46020 ( .A(ein[1021]), .B(n41943), .Z(ereg_next[1022]) );
  AND U46021 ( .A(mul_pow), .B(n41944), .Z(n41943) );
  XOR U46022 ( .A(ein[1022]), .B(ein[1021]), .Z(n41944) );
  XOR U46023 ( .A(ein[1020]), .B(n41945), .Z(ereg_next[1021]) );
  AND U46024 ( .A(mul_pow), .B(n41946), .Z(n41945) );
  XOR U46025 ( .A(ein[1021]), .B(ein[1020]), .Z(n41946) );
  XOR U46026 ( .A(ein[1019]), .B(n41947), .Z(ereg_next[1020]) );
  AND U46027 ( .A(mul_pow), .B(n41948), .Z(n41947) );
  XOR U46028 ( .A(ein[1020]), .B(ein[1019]), .Z(n41948) );
  XOR U46029 ( .A(ein[100]), .B(n41949), .Z(ereg_next[101]) );
  AND U46030 ( .A(mul_pow), .B(n41950), .Z(n41949) );
  XOR U46031 ( .A(ein[101]), .B(ein[100]), .Z(n41950) );
  XOR U46032 ( .A(ein[1018]), .B(n41951), .Z(ereg_next[1019]) );
  AND U46033 ( .A(mul_pow), .B(n41952), .Z(n41951) );
  XOR U46034 ( .A(ein[1019]), .B(ein[1018]), .Z(n41952) );
  XOR U46035 ( .A(ein[1017]), .B(n41953), .Z(ereg_next[1018]) );
  AND U46036 ( .A(mul_pow), .B(n41954), .Z(n41953) );
  XOR U46037 ( .A(ein[1018]), .B(ein[1017]), .Z(n41954) );
  XOR U46038 ( .A(ein[1016]), .B(n41955), .Z(ereg_next[1017]) );
  AND U46039 ( .A(mul_pow), .B(n41956), .Z(n41955) );
  XOR U46040 ( .A(ein[1017]), .B(ein[1016]), .Z(n41956) );
  XOR U46041 ( .A(ein[1015]), .B(n41957), .Z(ereg_next[1016]) );
  AND U46042 ( .A(mul_pow), .B(n41958), .Z(n41957) );
  XOR U46043 ( .A(ein[1016]), .B(ein[1015]), .Z(n41958) );
  XOR U46044 ( .A(ein[1014]), .B(n41959), .Z(ereg_next[1015]) );
  AND U46045 ( .A(mul_pow), .B(n41960), .Z(n41959) );
  XOR U46046 ( .A(ein[1015]), .B(ein[1014]), .Z(n41960) );
  XOR U46047 ( .A(ein[1013]), .B(n41961), .Z(ereg_next[1014]) );
  AND U46048 ( .A(mul_pow), .B(n41962), .Z(n41961) );
  XOR U46049 ( .A(ein[1014]), .B(ein[1013]), .Z(n41962) );
  XOR U46050 ( .A(ein[1012]), .B(n41963), .Z(ereg_next[1013]) );
  AND U46051 ( .A(mul_pow), .B(n41964), .Z(n41963) );
  XOR U46052 ( .A(ein[1013]), .B(ein[1012]), .Z(n41964) );
  XOR U46053 ( .A(ein[1011]), .B(n41965), .Z(ereg_next[1012]) );
  AND U46054 ( .A(mul_pow), .B(n41966), .Z(n41965) );
  XOR U46055 ( .A(ein[1012]), .B(ein[1011]), .Z(n41966) );
  XOR U46056 ( .A(ein[1010]), .B(n41967), .Z(ereg_next[1011]) );
  AND U46057 ( .A(mul_pow), .B(n41968), .Z(n41967) );
  XOR U46058 ( .A(ein[1011]), .B(ein[1010]), .Z(n41968) );
  XOR U46059 ( .A(ein[1009]), .B(n41969), .Z(ereg_next[1010]) );
  AND U46060 ( .A(mul_pow), .B(n41970), .Z(n41969) );
  XOR U46061 ( .A(ein[1010]), .B(ein[1009]), .Z(n41970) );
  XOR U46062 ( .A(ein[99]), .B(n41971), .Z(ereg_next[100]) );
  AND U46063 ( .A(mul_pow), .B(n41972), .Z(n41971) );
  XOR U46064 ( .A(ein[99]), .B(ein[100]), .Z(n41972) );
  XOR U46065 ( .A(ein[1008]), .B(n41973), .Z(ereg_next[1009]) );
  AND U46066 ( .A(mul_pow), .B(n41974), .Z(n41973) );
  XOR U46067 ( .A(ein[1009]), .B(ein[1008]), .Z(n41974) );
  XOR U46068 ( .A(ein[1007]), .B(n41975), .Z(ereg_next[1008]) );
  AND U46069 ( .A(mul_pow), .B(n41976), .Z(n41975) );
  XOR U46070 ( .A(ein[1008]), .B(ein[1007]), .Z(n41976) );
  XOR U46071 ( .A(ein[1006]), .B(n41977), .Z(ereg_next[1007]) );
  AND U46072 ( .A(mul_pow), .B(n41978), .Z(n41977) );
  XOR U46073 ( .A(ein[1007]), .B(ein[1006]), .Z(n41978) );
  XOR U46074 ( .A(ein[1005]), .B(n41979), .Z(ereg_next[1006]) );
  AND U46075 ( .A(mul_pow), .B(n41980), .Z(n41979) );
  XOR U46076 ( .A(ein[1006]), .B(ein[1005]), .Z(n41980) );
  XOR U46077 ( .A(ein[1004]), .B(n41981), .Z(ereg_next[1005]) );
  AND U46078 ( .A(mul_pow), .B(n41982), .Z(n41981) );
  XOR U46079 ( .A(ein[1005]), .B(ein[1004]), .Z(n41982) );
  XOR U46080 ( .A(ein[1003]), .B(n41983), .Z(ereg_next[1004]) );
  AND U46081 ( .A(mul_pow), .B(n41984), .Z(n41983) );
  XOR U46082 ( .A(ein[1004]), .B(ein[1003]), .Z(n41984) );
  XOR U46083 ( .A(ein[1002]), .B(n41985), .Z(ereg_next[1003]) );
  AND U46084 ( .A(mul_pow), .B(n41986), .Z(n41985) );
  XOR U46085 ( .A(ein[1003]), .B(ein[1002]), .Z(n41986) );
  XOR U46086 ( .A(ein[1001]), .B(n41987), .Z(ereg_next[1002]) );
  AND U46087 ( .A(mul_pow), .B(n41988), .Z(n41987) );
  XOR U46088 ( .A(ein[1002]), .B(ein[1001]), .Z(n41988) );
  XOR U46089 ( .A(ein[1000]), .B(n41989), .Z(ereg_next[1001]) );
  AND U46090 ( .A(mul_pow), .B(n41990), .Z(n41989) );
  XOR U46091 ( .A(ein[1001]), .B(ein[1000]), .Z(n41990) );
  XOR U46092 ( .A(ein[999]), .B(n41991), .Z(ereg_next[1000]) );
  AND U46093 ( .A(mul_pow), .B(n41992), .Z(n41991) );
  XOR U46094 ( .A(ein[999]), .B(ein[1000]), .Z(n41992) );
  AND U46095 ( .A(ein[0]), .B(mul_pow), .Z(ereg_next[0]) );
endmodule

