
module compare_N16384_CC256 ( clk, rst, x, y, g, e );
  input [63:0] x;
  input [63:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  IV U10 ( .A(ebreg), .Z(e) );
  XNOR U11 ( .A(y[45]), .B(x[45]), .Z(n9) );
  NANDN U12 ( .A(x[44]), .B(y[44]), .Z(n8) );
  NAND U13 ( .A(n9), .B(n8), .Z(n269) );
  XNOR U14 ( .A(y[41]), .B(x[41]), .Z(n11) );
  NANDN U15 ( .A(x[40]), .B(y[40]), .Z(n10) );
  NAND U16 ( .A(n11), .B(n10), .Z(n257) );
  XNOR U17 ( .A(y[43]), .B(x[43]), .Z(n13) );
  NANDN U18 ( .A(x[42]), .B(y[42]), .Z(n12) );
  NAND U19 ( .A(n13), .B(n12), .Z(n263) );
  NOR U20 ( .A(n257), .B(n263), .Z(n16) );
  XNOR U21 ( .A(y[47]), .B(x[47]), .Z(n15) );
  NANDN U22 ( .A(x[46]), .B(y[46]), .Z(n14) );
  NAND U23 ( .A(n15), .B(n14), .Z(n275) );
  ANDN U24 ( .B(n16), .A(n275), .Z(n17) );
  NANDN U25 ( .A(n269), .B(n17), .Z(n29) );
  XNOR U26 ( .A(y[37]), .B(x[37]), .Z(n19) );
  NANDN U27 ( .A(x[36]), .B(y[36]), .Z(n18) );
  NAND U28 ( .A(n19), .B(n18), .Z(n245) );
  XNOR U29 ( .A(y[33]), .B(x[33]), .Z(n21) );
  NANDN U30 ( .A(x[32]), .B(y[32]), .Z(n20) );
  NAND U31 ( .A(n21), .B(n20), .Z(n233) );
  XNOR U32 ( .A(y[35]), .B(x[35]), .Z(n23) );
  NANDN U33 ( .A(x[34]), .B(y[34]), .Z(n22) );
  NAND U34 ( .A(n23), .B(n22), .Z(n239) );
  NOR U35 ( .A(n233), .B(n239), .Z(n26) );
  XNOR U36 ( .A(y[39]), .B(x[39]), .Z(n25) );
  NANDN U37 ( .A(x[38]), .B(y[38]), .Z(n24) );
  NAND U38 ( .A(n25), .B(n24), .Z(n251) );
  ANDN U39 ( .B(n26), .A(n251), .Z(n27) );
  NANDN U40 ( .A(n245), .B(n27), .Z(n28) );
  NOR U41 ( .A(n29), .B(n28), .Z(n85) );
  ANDN U42 ( .B(x[60]), .A(y[60]), .Z(n313) );
  ANDN U43 ( .B(x[56]), .A(y[56]), .Z(n301) );
  ANDN U44 ( .B(x[58]), .A(y[58]), .Z(n307) );
  NOR U45 ( .A(n301), .B(n307), .Z(n30) );
  ANDN U46 ( .B(x[62]), .A(y[62]), .Z(n319) );
  ANDN U47 ( .B(n30), .A(n319), .Z(n31) );
  NANDN U48 ( .A(n313), .B(n31), .Z(n43) );
  ANDN U49 ( .B(x[44]), .A(y[44]), .Z(n265) );
  ANDN U50 ( .B(x[40]), .A(y[40]), .Z(n253) );
  ANDN U51 ( .B(x[42]), .A(y[42]), .Z(n259) );
  NOR U52 ( .A(n253), .B(n259), .Z(n32) );
  ANDN U53 ( .B(x[46]), .A(y[46]), .Z(n271) );
  ANDN U54 ( .B(n32), .A(n271), .Z(n33) );
  NANDN U55 ( .A(n265), .B(n33), .Z(n37) );
  ANDN U56 ( .B(x[36]), .A(y[36]), .Z(n241) );
  ANDN U57 ( .B(x[32]), .A(y[32]), .Z(n231) );
  ANDN U58 ( .B(x[34]), .A(y[34]), .Z(n235) );
  NOR U59 ( .A(n231), .B(n235), .Z(n34) );
  ANDN U60 ( .B(x[38]), .A(y[38]), .Z(n247) );
  ANDN U61 ( .B(n34), .A(n247), .Z(n35) );
  NANDN U62 ( .A(n241), .B(n35), .Z(n36) );
  NOR U63 ( .A(n37), .B(n36), .Z(n41) );
  ANDN U64 ( .B(x[52]), .A(y[52]), .Z(n289) );
  ANDN U65 ( .B(x[48]), .A(y[48]), .Z(n277) );
  ANDN U66 ( .B(x[50]), .A(y[50]), .Z(n283) );
  NOR U67 ( .A(n277), .B(n283), .Z(n38) );
  ANDN U68 ( .B(x[54]), .A(y[54]), .Z(n295) );
  ANDN U69 ( .B(n38), .A(n295), .Z(n39) );
  NANDN U70 ( .A(n289), .B(n39), .Z(n40) );
  ANDN U71 ( .B(n41), .A(n40), .Z(n42) );
  NANDN U72 ( .A(n43), .B(n42), .Z(n83) );
  XNOR U73 ( .A(y[61]), .B(x[61]), .Z(n45) );
  NANDN U74 ( .A(x[60]), .B(y[60]), .Z(n44) );
  NAND U75 ( .A(n45), .B(n44), .Z(n317) );
  XNOR U76 ( .A(y[57]), .B(x[57]), .Z(n47) );
  NANDN U77 ( .A(x[56]), .B(y[56]), .Z(n46) );
  NAND U78 ( .A(n47), .B(n46), .Z(n305) );
  XNOR U79 ( .A(y[59]), .B(x[59]), .Z(n49) );
  NANDN U80 ( .A(x[58]), .B(y[58]), .Z(n48) );
  NAND U81 ( .A(n49), .B(n48), .Z(n311) );
  NOR U82 ( .A(n305), .B(n311), .Z(n52) );
  XNOR U83 ( .A(y[63]), .B(x[63]), .Z(n51) );
  NANDN U84 ( .A(x[62]), .B(y[62]), .Z(n50) );
  NAND U85 ( .A(n51), .B(n50), .Z(n323) );
  ANDN U86 ( .B(n52), .A(n323), .Z(n53) );
  NANDN U87 ( .A(n317), .B(n53), .Z(n65) );
  XNOR U88 ( .A(y[53]), .B(x[53]), .Z(n55) );
  NANDN U89 ( .A(x[52]), .B(y[52]), .Z(n54) );
  NAND U90 ( .A(n55), .B(n54), .Z(n293) );
  XNOR U91 ( .A(y[49]), .B(x[49]), .Z(n57) );
  NANDN U92 ( .A(x[48]), .B(y[48]), .Z(n56) );
  NAND U93 ( .A(n57), .B(n56), .Z(n281) );
  XNOR U94 ( .A(y[51]), .B(x[51]), .Z(n59) );
  NANDN U95 ( .A(x[50]), .B(y[50]), .Z(n58) );
  NAND U96 ( .A(n59), .B(n58), .Z(n287) );
  NOR U97 ( .A(n281), .B(n287), .Z(n62) );
  XNOR U98 ( .A(y[55]), .B(x[55]), .Z(n61) );
  NANDN U99 ( .A(x[54]), .B(y[54]), .Z(n60) );
  NAND U100 ( .A(n61), .B(n60), .Z(n299) );
  ANDN U101 ( .B(n62), .A(n299), .Z(n63) );
  NANDN U102 ( .A(n293), .B(n63), .Z(n64) );
  NOR U103 ( .A(n65), .B(n64), .Z(n81) );
  ANDN U104 ( .B(x[28]), .A(y[28]), .Z(n219) );
  ANDN U105 ( .B(x[24]), .A(y[24]), .Z(n207) );
  ANDN U106 ( .B(x[26]), .A(y[26]), .Z(n213) );
  NOR U107 ( .A(n207), .B(n213), .Z(n66) );
  ANDN U108 ( .B(x[30]), .A(y[30]), .Z(n225) );
  ANDN U109 ( .B(n66), .A(n225), .Z(n67) );
  NANDN U110 ( .A(n219), .B(n67), .Z(n79) );
  NANDN U111 ( .A(y[8]), .B(x[8]), .Z(n141) );
  ANDN U112 ( .B(x[10]), .A(y[10]), .Z(n138) );
  ANDN U113 ( .B(n141), .A(n138), .Z(n68) );
  ANDN U114 ( .B(x[14]), .A(y[14]), .Z(n177) );
  ANDN U115 ( .B(n68), .A(n177), .Z(n69) );
  NANDN U116 ( .A(y[12]), .B(x[12]), .Z(n137) );
  NAND U117 ( .A(n69), .B(n137), .Z(n73) );
  NANDN U118 ( .A(y[6]), .B(x[6]), .Z(n143) );
  NANDN U119 ( .A(y[0]), .B(x[0]), .Z(n146) );
  NANDN U120 ( .A(y[4]), .B(x[4]), .Z(n145) );
  AND U121 ( .A(n146), .B(n145), .Z(n70) );
  AND U122 ( .A(n143), .B(n70), .Z(n71) );
  NANDN U123 ( .A(y[2]), .B(x[2]), .Z(n151) );
  NAND U124 ( .A(n71), .B(n151), .Z(n72) );
  NOR U125 ( .A(n73), .B(n72), .Z(n77) );
  ANDN U126 ( .B(x[20]), .A(y[20]), .Z(n195) );
  ANDN U127 ( .B(x[16]), .A(y[16]), .Z(n183) );
  ANDN U128 ( .B(x[18]), .A(y[18]), .Z(n189) );
  NOR U129 ( .A(n183), .B(n189), .Z(n74) );
  ANDN U130 ( .B(x[22]), .A(y[22]), .Z(n201) );
  ANDN U131 ( .B(n74), .A(n201), .Z(n75) );
  NANDN U132 ( .A(n195), .B(n75), .Z(n76) );
  ANDN U133 ( .B(n77), .A(n76), .Z(n78) );
  NANDN U134 ( .A(n79), .B(n78), .Z(n80) );
  ANDN U135 ( .B(n81), .A(n80), .Z(n82) );
  NANDN U136 ( .A(n83), .B(n82), .Z(n84) );
  ANDN U137 ( .B(n85), .A(n84), .Z(n134) );
  XNOR U138 ( .A(y[21]), .B(x[21]), .Z(n87) );
  NANDN U139 ( .A(x[20]), .B(y[20]), .Z(n86) );
  NAND U140 ( .A(n87), .B(n86), .Z(n197) );
  XNOR U141 ( .A(y[17]), .B(x[17]), .Z(n89) );
  NANDN U142 ( .A(x[16]), .B(y[16]), .Z(n88) );
  NAND U143 ( .A(n89), .B(n88), .Z(n185) );
  XNOR U144 ( .A(y[19]), .B(x[19]), .Z(n91) );
  NANDN U145 ( .A(x[18]), .B(y[18]), .Z(n90) );
  NAND U146 ( .A(n91), .B(n90), .Z(n191) );
  NOR U147 ( .A(n185), .B(n191), .Z(n94) );
  XNOR U148 ( .A(y[23]), .B(x[23]), .Z(n93) );
  NANDN U149 ( .A(x[22]), .B(y[22]), .Z(n92) );
  NAND U150 ( .A(n93), .B(n92), .Z(n203) );
  ANDN U151 ( .B(n94), .A(n203), .Z(n95) );
  NANDN U152 ( .A(n197), .B(n95), .Z(n132) );
  XNOR U153 ( .A(y[7]), .B(x[7]), .Z(n97) );
  NANDN U154 ( .A(x[6]), .B(y[6]), .Z(n96) );
  NAND U155 ( .A(n97), .B(n96), .Z(n161) );
  XNOR U156 ( .A(y[3]), .B(x[3]), .Z(n99) );
  NANDN U157 ( .A(x[2]), .B(y[2]), .Z(n98) );
  NAND U158 ( .A(n99), .B(n98), .Z(n153) );
  XNOR U159 ( .A(y[5]), .B(x[5]), .Z(n101) );
  NANDN U160 ( .A(x[4]), .B(y[4]), .Z(n100) );
  NAND U161 ( .A(n101), .B(n100), .Z(n157) );
  NOR U162 ( .A(n153), .B(n157), .Z(n105) );
  XNOR U163 ( .A(y[1]), .B(x[1]), .Z(n103) );
  NANDN U164 ( .A(x[0]), .B(y[0]), .Z(n102) );
  NAND U165 ( .A(n103), .B(n102), .Z(n104) );
  ANDN U166 ( .B(n105), .A(n104), .Z(n106) );
  NANDN U167 ( .A(n161), .B(n106), .Z(n118) );
  XNOR U168 ( .A(y[13]), .B(x[13]), .Z(n108) );
  NANDN U169 ( .A(x[12]), .B(y[12]), .Z(n107) );
  NAND U170 ( .A(n108), .B(n107), .Z(n173) );
  XNOR U171 ( .A(y[9]), .B(x[9]), .Z(n110) );
  NANDN U172 ( .A(x[8]), .B(y[8]), .Z(n109) );
  NAND U173 ( .A(n110), .B(n109), .Z(n165) );
  XNOR U174 ( .A(y[11]), .B(x[11]), .Z(n112) );
  NANDN U175 ( .A(x[10]), .B(y[10]), .Z(n111) );
  NAND U176 ( .A(n112), .B(n111), .Z(n169) );
  NOR U177 ( .A(n165), .B(n169), .Z(n115) );
  XNOR U178 ( .A(y[15]), .B(x[15]), .Z(n114) );
  NANDN U179 ( .A(x[14]), .B(y[14]), .Z(n113) );
  NAND U180 ( .A(n114), .B(n113), .Z(n179) );
  ANDN U181 ( .B(n115), .A(n179), .Z(n116) );
  NANDN U182 ( .A(n173), .B(n116), .Z(n117) );
  NOR U183 ( .A(n118), .B(n117), .Z(n130) );
  XNOR U184 ( .A(y[29]), .B(x[29]), .Z(n120) );
  NANDN U185 ( .A(x[28]), .B(y[28]), .Z(n119) );
  NAND U186 ( .A(n120), .B(n119), .Z(n221) );
  XNOR U187 ( .A(y[25]), .B(x[25]), .Z(n122) );
  NANDN U188 ( .A(x[24]), .B(y[24]), .Z(n121) );
  NAND U189 ( .A(n122), .B(n121), .Z(n209) );
  XNOR U190 ( .A(y[27]), .B(x[27]), .Z(n124) );
  NANDN U191 ( .A(x[26]), .B(y[26]), .Z(n123) );
  NAND U192 ( .A(n124), .B(n123), .Z(n215) );
  NOR U193 ( .A(n209), .B(n215), .Z(n127) );
  XNOR U194 ( .A(y[31]), .B(x[31]), .Z(n126) );
  NANDN U195 ( .A(x[30]), .B(y[30]), .Z(n125) );
  NAND U196 ( .A(n126), .B(n125), .Z(n227) );
  ANDN U197 ( .B(n127), .A(n227), .Z(n128) );
  NANDN U198 ( .A(n221), .B(n128), .Z(n129) );
  ANDN U199 ( .B(n130), .A(n129), .Z(n131) );
  NANDN U200 ( .A(n132), .B(n131), .Z(n133) );
  ANDN U201 ( .B(n134), .A(n133), .Z(n135) );
  NAND U202 ( .A(e), .B(n135), .Z(n5) );
  NANDN U203 ( .A(n135), .B(e), .Z(n327) );
  ANDN U204 ( .B(x[63]), .A(y[63]), .Z(n325) );
  ANDN U205 ( .B(x[31]), .A(y[31]), .Z(n229) );
  ANDN U206 ( .B(x[29]), .A(y[29]), .Z(n223) );
  ANDN U207 ( .B(x[27]), .A(y[27]), .Z(n217) );
  ANDN U208 ( .B(x[25]), .A(y[25]), .Z(n211) );
  ANDN U209 ( .B(x[23]), .A(y[23]), .Z(n205) );
  ANDN U210 ( .B(x[21]), .A(y[21]), .Z(n199) );
  ANDN U211 ( .B(x[19]), .A(y[19]), .Z(n193) );
  ANDN U212 ( .B(x[17]), .A(y[17]), .Z(n187) );
  ANDN U213 ( .B(x[15]), .A(y[15]), .Z(n181) );
  NANDN U214 ( .A(y[13]), .B(x[13]), .Z(n175) );
  NANDN U215 ( .A(y[11]), .B(x[11]), .Z(n136) );
  AND U216 ( .A(n137), .B(n136), .Z(n171) );
  NANDN U217 ( .A(y[9]), .B(x[9]), .Z(n139) );
  ANDN U218 ( .B(n139), .A(n138), .Z(n167) );
  NANDN U219 ( .A(y[7]), .B(x[7]), .Z(n140) );
  AND U220 ( .A(n141), .B(n140), .Z(n163) );
  NANDN U221 ( .A(y[5]), .B(x[5]), .Z(n142) );
  AND U222 ( .A(n143), .B(n142), .Z(n159) );
  NANDN U223 ( .A(y[3]), .B(x[3]), .Z(n144) );
  AND U224 ( .A(n145), .B(n144), .Z(n155) );
  NANDN U225 ( .A(x[1]), .B(n146), .Z(n149) );
  XNOR U226 ( .A(n146), .B(x[1]), .Z(n147) );
  NAND U227 ( .A(n147), .B(y[1]), .Z(n148) );
  NAND U228 ( .A(n149), .B(n148), .Z(n150) );
  AND U229 ( .A(n151), .B(n150), .Z(n152) );
  OR U230 ( .A(n153), .B(n152), .Z(n154) );
  AND U231 ( .A(n155), .B(n154), .Z(n156) );
  OR U232 ( .A(n157), .B(n156), .Z(n158) );
  AND U233 ( .A(n159), .B(n158), .Z(n160) );
  OR U234 ( .A(n161), .B(n160), .Z(n162) );
  AND U235 ( .A(n163), .B(n162), .Z(n164) );
  OR U236 ( .A(n165), .B(n164), .Z(n166) );
  AND U237 ( .A(n167), .B(n166), .Z(n168) );
  OR U238 ( .A(n169), .B(n168), .Z(n170) );
  AND U239 ( .A(n171), .B(n170), .Z(n172) );
  OR U240 ( .A(n173), .B(n172), .Z(n174) );
  AND U241 ( .A(n175), .B(n174), .Z(n176) );
  NANDN U242 ( .A(n177), .B(n176), .Z(n178) );
  NANDN U243 ( .A(n179), .B(n178), .Z(n180) );
  NANDN U244 ( .A(n181), .B(n180), .Z(n182) );
  OR U245 ( .A(n183), .B(n182), .Z(n184) );
  NANDN U246 ( .A(n185), .B(n184), .Z(n186) );
  NANDN U247 ( .A(n187), .B(n186), .Z(n188) );
  OR U248 ( .A(n189), .B(n188), .Z(n190) );
  NANDN U249 ( .A(n191), .B(n190), .Z(n192) );
  NANDN U250 ( .A(n193), .B(n192), .Z(n194) );
  OR U251 ( .A(n195), .B(n194), .Z(n196) );
  NANDN U252 ( .A(n197), .B(n196), .Z(n198) );
  NANDN U253 ( .A(n199), .B(n198), .Z(n200) );
  OR U254 ( .A(n201), .B(n200), .Z(n202) );
  NANDN U255 ( .A(n203), .B(n202), .Z(n204) );
  NANDN U256 ( .A(n205), .B(n204), .Z(n206) );
  OR U257 ( .A(n207), .B(n206), .Z(n208) );
  NANDN U258 ( .A(n209), .B(n208), .Z(n210) );
  NANDN U259 ( .A(n211), .B(n210), .Z(n212) );
  OR U260 ( .A(n213), .B(n212), .Z(n214) );
  NANDN U261 ( .A(n215), .B(n214), .Z(n216) );
  NANDN U262 ( .A(n217), .B(n216), .Z(n218) );
  OR U263 ( .A(n219), .B(n218), .Z(n220) );
  NANDN U264 ( .A(n221), .B(n220), .Z(n222) );
  NANDN U265 ( .A(n223), .B(n222), .Z(n224) );
  OR U266 ( .A(n225), .B(n224), .Z(n226) );
  NANDN U267 ( .A(n227), .B(n226), .Z(n228) );
  NANDN U268 ( .A(n229), .B(n228), .Z(n230) );
  OR U269 ( .A(n231), .B(n230), .Z(n232) );
  NANDN U270 ( .A(n233), .B(n232), .Z(n234) );
  NANDN U271 ( .A(n235), .B(n234), .Z(n237) );
  ANDN U272 ( .B(x[33]), .A(y[33]), .Z(n236) );
  OR U273 ( .A(n237), .B(n236), .Z(n238) );
  NANDN U274 ( .A(n239), .B(n238), .Z(n240) );
  NANDN U275 ( .A(n241), .B(n240), .Z(n243) );
  ANDN U276 ( .B(x[35]), .A(y[35]), .Z(n242) );
  OR U277 ( .A(n243), .B(n242), .Z(n244) );
  NANDN U278 ( .A(n245), .B(n244), .Z(n246) );
  NANDN U279 ( .A(n247), .B(n246), .Z(n249) );
  ANDN U280 ( .B(x[37]), .A(y[37]), .Z(n248) );
  OR U281 ( .A(n249), .B(n248), .Z(n250) );
  NANDN U282 ( .A(n251), .B(n250), .Z(n252) );
  NANDN U283 ( .A(n253), .B(n252), .Z(n255) );
  ANDN U284 ( .B(x[39]), .A(y[39]), .Z(n254) );
  OR U285 ( .A(n255), .B(n254), .Z(n256) );
  NANDN U286 ( .A(n257), .B(n256), .Z(n258) );
  NANDN U287 ( .A(n259), .B(n258), .Z(n261) );
  ANDN U288 ( .B(x[41]), .A(y[41]), .Z(n260) );
  OR U289 ( .A(n261), .B(n260), .Z(n262) );
  NANDN U290 ( .A(n263), .B(n262), .Z(n264) );
  NANDN U291 ( .A(n265), .B(n264), .Z(n267) );
  ANDN U292 ( .B(x[43]), .A(y[43]), .Z(n266) );
  OR U293 ( .A(n267), .B(n266), .Z(n268) );
  NANDN U294 ( .A(n269), .B(n268), .Z(n270) );
  NANDN U295 ( .A(n271), .B(n270), .Z(n273) );
  ANDN U296 ( .B(x[45]), .A(y[45]), .Z(n272) );
  OR U297 ( .A(n273), .B(n272), .Z(n274) );
  NANDN U298 ( .A(n275), .B(n274), .Z(n276) );
  NANDN U299 ( .A(n277), .B(n276), .Z(n279) );
  ANDN U300 ( .B(x[47]), .A(y[47]), .Z(n278) );
  OR U301 ( .A(n279), .B(n278), .Z(n280) );
  NANDN U302 ( .A(n281), .B(n280), .Z(n282) );
  NANDN U303 ( .A(n283), .B(n282), .Z(n285) );
  ANDN U304 ( .B(x[49]), .A(y[49]), .Z(n284) );
  OR U305 ( .A(n285), .B(n284), .Z(n286) );
  NANDN U306 ( .A(n287), .B(n286), .Z(n288) );
  NANDN U307 ( .A(n289), .B(n288), .Z(n291) );
  ANDN U308 ( .B(x[51]), .A(y[51]), .Z(n290) );
  OR U309 ( .A(n291), .B(n290), .Z(n292) );
  NANDN U310 ( .A(n293), .B(n292), .Z(n294) );
  NANDN U311 ( .A(n295), .B(n294), .Z(n297) );
  ANDN U312 ( .B(x[53]), .A(y[53]), .Z(n296) );
  OR U313 ( .A(n297), .B(n296), .Z(n298) );
  NANDN U314 ( .A(n299), .B(n298), .Z(n300) );
  NANDN U315 ( .A(n301), .B(n300), .Z(n303) );
  ANDN U316 ( .B(x[55]), .A(y[55]), .Z(n302) );
  OR U317 ( .A(n303), .B(n302), .Z(n304) );
  NANDN U318 ( .A(n305), .B(n304), .Z(n306) );
  NANDN U319 ( .A(n307), .B(n306), .Z(n309) );
  ANDN U320 ( .B(x[57]), .A(y[57]), .Z(n308) );
  OR U321 ( .A(n309), .B(n308), .Z(n310) );
  NANDN U322 ( .A(n311), .B(n310), .Z(n312) );
  NANDN U323 ( .A(n313), .B(n312), .Z(n315) );
  ANDN U324 ( .B(x[59]), .A(y[59]), .Z(n314) );
  OR U325 ( .A(n315), .B(n314), .Z(n316) );
  NANDN U326 ( .A(n317), .B(n316), .Z(n318) );
  NANDN U327 ( .A(n319), .B(n318), .Z(n321) );
  ANDN U328 ( .B(x[61]), .A(y[61]), .Z(n320) );
  OR U329 ( .A(n321), .B(n320), .Z(n322) );
  NANDN U330 ( .A(n323), .B(n322), .Z(n324) );
  NANDN U331 ( .A(n325), .B(n324), .Z(n326) );
  NANDN U332 ( .A(n327), .B(n326), .Z(n329) );
  NAND U333 ( .A(n327), .B(g), .Z(n328) );
  NAND U334 ( .A(n329), .B(n328), .Z(n4) );
endmodule

