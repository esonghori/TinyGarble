
module FA_0 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(A), .B(B), .Z(CO) );
  XOR U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_99 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_98 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_97 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_96 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_95 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_94 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_93 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_92 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_91 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_90 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_89 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_88 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_87 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_86 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_85 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_84 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_83 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_82 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_81 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_80 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_79 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_78 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_77 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_76 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_75 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_74 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_73 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_72 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_71 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_70 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_69 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_68 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_67 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_66 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_65 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_64 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_63 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_62 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_61 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_60 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_59 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_58 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_57 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_56 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_55 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_54 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_53 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_52 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_51 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_50 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_49 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_48 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_47 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_46 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_45 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_44 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_43 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_42 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_41 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_40 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_39 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_38 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_37 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_36 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_35 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_34 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_33 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_32 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_31 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_30 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_29 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_28 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_27 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_26 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_25 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_24 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_23 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_22 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_21 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_20 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_19 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_18 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_17 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_16 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_15 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_14 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_13 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_12 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_11 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_10 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_9 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_8 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_7 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_6 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_5 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_4 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XNOR U2 ( .A(A), .B(CI), .Z(n1) );
  XOR U3 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_1 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N1024 ( A, B, CI, S, CO );
  input [1023:0] A;
  input [1023:0] B;
  output [1023:0] S;
  input CI;
  output CO;

  wire   [1023:1] C;

  FA_0 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(B[0]), .CI(1'b0), .S(
        S[0]), .CO(C[1]) );
  FA_1023 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(B[1]), .CI(C[1]), .S(
        S[1]), .CO(C[2]) );
  FA_1022 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(
        S[2]), .CO(C[3]) );
  FA_1021 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(
        S[3]), .CO(C[4]) );
  FA_1020 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(
        S[4]), .CO(C[5]) );
  FA_1019 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(
        S[5]), .CO(C[6]) );
  FA_1018 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(
        S[6]), .CO(C[7]) );
  FA_1017 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(
        S[7]), .CO(C[8]) );
  FA_1016 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(
        S[8]), .CO(C[9]) );
  FA_1015 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(
        S[9]), .CO(C[10]) );
  FA_1014 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_1013 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_1012 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_1011 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_1010 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_1009 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_1008 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_1007 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_1006 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_1005 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_1004 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_1003 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_1002 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_1001 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_1000 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_999 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_998 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_997 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_996 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_995 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_994 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_993 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_992 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_991 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_990 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_989 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_988 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_987 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_986 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_985 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_984 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_983 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_982 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_981 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_980 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_979 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_978 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_977 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_976 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_975 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_974 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_973 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_972 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_971 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_970 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_969 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_968 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_967 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_966 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_965 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_964 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_963 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_962 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_961 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_960 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_959 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_958 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_957 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_956 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_955 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_954 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_953 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_952 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_951 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_950 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_949 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_948 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_947 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_946 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_945 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_944 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_943 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_942 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_941 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_940 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_939 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_938 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_937 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_936 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_935 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_934 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_933 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_932 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_931 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_930 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_929 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_928 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_927 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_926 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_925 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_924 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(B[100]), .CI(
        C[100]), .S(S[100]), .CO(C[101]) );
  FA_923 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(B[101]), .CI(
        C[101]), .S(S[101]), .CO(C[102]) );
  FA_922 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(B[102]), .CI(
        C[102]), .S(S[102]), .CO(C[103]) );
  FA_921 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(B[103]), .CI(
        C[103]), .S(S[103]), .CO(C[104]) );
  FA_920 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(B[104]), .CI(
        C[104]), .S(S[104]), .CO(C[105]) );
  FA_919 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(B[105]), .CI(
        C[105]), .S(S[105]), .CO(C[106]) );
  FA_918 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(B[106]), .CI(
        C[106]), .S(S[106]), .CO(C[107]) );
  FA_917 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(B[107]), .CI(
        C[107]), .S(S[107]), .CO(C[108]) );
  FA_916 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(B[108]), .CI(
        C[108]), .S(S[108]), .CO(C[109]) );
  FA_915 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(B[109]), .CI(
        C[109]), .S(S[109]), .CO(C[110]) );
  FA_914 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(B[110]), .CI(
        C[110]), .S(S[110]), .CO(C[111]) );
  FA_913 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(B[111]), .CI(
        C[111]), .S(S[111]), .CO(C[112]) );
  FA_912 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(B[112]), .CI(
        C[112]), .S(S[112]), .CO(C[113]) );
  FA_911 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(B[113]), .CI(
        C[113]), .S(S[113]), .CO(C[114]) );
  FA_910 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(B[114]), .CI(
        C[114]), .S(S[114]), .CO(C[115]) );
  FA_909 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(B[115]), .CI(
        C[115]), .S(S[115]), .CO(C[116]) );
  FA_908 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(B[116]), .CI(
        C[116]), .S(S[116]), .CO(C[117]) );
  FA_907 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(B[117]), .CI(
        C[117]), .S(S[117]), .CO(C[118]) );
  FA_906 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(B[118]), .CI(
        C[118]), .S(S[118]), .CO(C[119]) );
  FA_905 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(B[119]), .CI(
        C[119]), .S(S[119]), .CO(C[120]) );
  FA_904 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(B[120]), .CI(
        C[120]), .S(S[120]), .CO(C[121]) );
  FA_903 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(B[121]), .CI(
        C[121]), .S(S[121]), .CO(C[122]) );
  FA_902 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(B[122]), .CI(
        C[122]), .S(S[122]), .CO(C[123]) );
  FA_901 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(B[123]), .CI(
        C[123]), .S(S[123]), .CO(C[124]) );
  FA_900 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(B[124]), .CI(
        C[124]), .S(S[124]), .CO(C[125]) );
  FA_899 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(B[125]), .CI(
        C[125]), .S(S[125]), .CO(C[126]) );
  FA_898 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(B[126]), .CI(
        C[126]), .S(S[126]), .CO(C[127]) );
  FA_897 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(B[127]), .CI(
        C[127]), .S(S[127]), .CO(C[128]) );
  FA_896 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(B[128]), .CI(
        C[128]), .S(S[128]), .CO(C[129]) );
  FA_895 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(B[129]), .CI(
        C[129]), .S(S[129]), .CO(C[130]) );
  FA_894 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(B[130]), .CI(
        C[130]), .S(S[130]), .CO(C[131]) );
  FA_893 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(B[131]), .CI(
        C[131]), .S(S[131]), .CO(C[132]) );
  FA_892 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(B[132]), .CI(
        C[132]), .S(S[132]), .CO(C[133]) );
  FA_891 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(B[133]), .CI(
        C[133]), .S(S[133]), .CO(C[134]) );
  FA_890 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(B[134]), .CI(
        C[134]), .S(S[134]), .CO(C[135]) );
  FA_889 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(B[135]), .CI(
        C[135]), .S(S[135]), .CO(C[136]) );
  FA_888 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(B[136]), .CI(
        C[136]), .S(S[136]), .CO(C[137]) );
  FA_887 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(B[137]), .CI(
        C[137]), .S(S[137]), .CO(C[138]) );
  FA_886 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(B[138]), .CI(
        C[138]), .S(S[138]), .CO(C[139]) );
  FA_885 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(B[139]), .CI(
        C[139]), .S(S[139]), .CO(C[140]) );
  FA_884 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(B[140]), .CI(
        C[140]), .S(S[140]), .CO(C[141]) );
  FA_883 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(B[141]), .CI(
        C[141]), .S(S[141]), .CO(C[142]) );
  FA_882 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(B[142]), .CI(
        C[142]), .S(S[142]), .CO(C[143]) );
  FA_881 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(B[143]), .CI(
        C[143]), .S(S[143]), .CO(C[144]) );
  FA_880 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(B[144]), .CI(
        C[144]), .S(S[144]), .CO(C[145]) );
  FA_879 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(B[145]), .CI(
        C[145]), .S(S[145]), .CO(C[146]) );
  FA_878 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(B[146]), .CI(
        C[146]), .S(S[146]), .CO(C[147]) );
  FA_877 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(B[147]), .CI(
        C[147]), .S(S[147]), .CO(C[148]) );
  FA_876 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(B[148]), .CI(
        C[148]), .S(S[148]), .CO(C[149]) );
  FA_875 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(B[149]), .CI(
        C[149]), .S(S[149]), .CO(C[150]) );
  FA_874 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(B[150]), .CI(
        C[150]), .S(S[150]), .CO(C[151]) );
  FA_873 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(B[151]), .CI(
        C[151]), .S(S[151]), .CO(C[152]) );
  FA_872 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(B[152]), .CI(
        C[152]), .S(S[152]), .CO(C[153]) );
  FA_871 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(B[153]), .CI(
        C[153]), .S(S[153]), .CO(C[154]) );
  FA_870 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(B[154]), .CI(
        C[154]), .S(S[154]), .CO(C[155]) );
  FA_869 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(B[155]), .CI(
        C[155]), .S(S[155]), .CO(C[156]) );
  FA_868 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(B[156]), .CI(
        C[156]), .S(S[156]), .CO(C[157]) );
  FA_867 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(B[157]), .CI(
        C[157]), .S(S[157]), .CO(C[158]) );
  FA_866 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(B[158]), .CI(
        C[158]), .S(S[158]), .CO(C[159]) );
  FA_865 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(B[159]), .CI(
        C[159]), .S(S[159]), .CO(C[160]) );
  FA_864 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(B[160]), .CI(
        C[160]), .S(S[160]), .CO(C[161]) );
  FA_863 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(B[161]), .CI(
        C[161]), .S(S[161]), .CO(C[162]) );
  FA_862 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(B[162]), .CI(
        C[162]), .S(S[162]), .CO(C[163]) );
  FA_861 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(B[163]), .CI(
        C[163]), .S(S[163]), .CO(C[164]) );
  FA_860 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(B[164]), .CI(
        C[164]), .S(S[164]), .CO(C[165]) );
  FA_859 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(B[165]), .CI(
        C[165]), .S(S[165]), .CO(C[166]) );
  FA_858 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(B[166]), .CI(
        C[166]), .S(S[166]), .CO(C[167]) );
  FA_857 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(B[167]), .CI(
        C[167]), .S(S[167]), .CO(C[168]) );
  FA_856 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(B[168]), .CI(
        C[168]), .S(S[168]), .CO(C[169]) );
  FA_855 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(B[169]), .CI(
        C[169]), .S(S[169]), .CO(C[170]) );
  FA_854 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(B[170]), .CI(
        C[170]), .S(S[170]), .CO(C[171]) );
  FA_853 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(B[171]), .CI(
        C[171]), .S(S[171]), .CO(C[172]) );
  FA_852 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(B[172]), .CI(
        C[172]), .S(S[172]), .CO(C[173]) );
  FA_851 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(B[173]), .CI(
        C[173]), .S(S[173]), .CO(C[174]) );
  FA_850 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(B[174]), .CI(
        C[174]), .S(S[174]), .CO(C[175]) );
  FA_849 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(B[175]), .CI(
        C[175]), .S(S[175]), .CO(C[176]) );
  FA_848 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(B[176]), .CI(
        C[176]), .S(S[176]), .CO(C[177]) );
  FA_847 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(B[177]), .CI(
        C[177]), .S(S[177]), .CO(C[178]) );
  FA_846 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(B[178]), .CI(
        C[178]), .S(S[178]), .CO(C[179]) );
  FA_845 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(B[179]), .CI(
        C[179]), .S(S[179]), .CO(C[180]) );
  FA_844 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(B[180]), .CI(
        C[180]), .S(S[180]), .CO(C[181]) );
  FA_843 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(B[181]), .CI(
        C[181]), .S(S[181]), .CO(C[182]) );
  FA_842 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(B[182]), .CI(
        C[182]), .S(S[182]), .CO(C[183]) );
  FA_841 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(B[183]), .CI(
        C[183]), .S(S[183]), .CO(C[184]) );
  FA_840 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(B[184]), .CI(
        C[184]), .S(S[184]), .CO(C[185]) );
  FA_839 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(B[185]), .CI(
        C[185]), .S(S[185]), .CO(C[186]) );
  FA_838 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(B[186]), .CI(
        C[186]), .S(S[186]), .CO(C[187]) );
  FA_837 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(B[187]), .CI(
        C[187]), .S(S[187]), .CO(C[188]) );
  FA_836 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(B[188]), .CI(
        C[188]), .S(S[188]), .CO(C[189]) );
  FA_835 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(B[189]), .CI(
        C[189]), .S(S[189]), .CO(C[190]) );
  FA_834 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(B[190]), .CI(
        C[190]), .S(S[190]), .CO(C[191]) );
  FA_833 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(B[191]), .CI(
        C[191]), .S(S[191]), .CO(C[192]) );
  FA_832 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(B[192]), .CI(
        C[192]), .S(S[192]), .CO(C[193]) );
  FA_831 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(B[193]), .CI(
        C[193]), .S(S[193]), .CO(C[194]) );
  FA_830 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(B[194]), .CI(
        C[194]), .S(S[194]), .CO(C[195]) );
  FA_829 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(B[195]), .CI(
        C[195]), .S(S[195]), .CO(C[196]) );
  FA_828 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(B[196]), .CI(
        C[196]), .S(S[196]), .CO(C[197]) );
  FA_827 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(B[197]), .CI(
        C[197]), .S(S[197]), .CO(C[198]) );
  FA_826 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(B[198]), .CI(
        C[198]), .S(S[198]), .CO(C[199]) );
  FA_825 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(B[199]), .CI(
        C[199]), .S(S[199]), .CO(C[200]) );
  FA_824 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(B[200]), .CI(
        C[200]), .S(S[200]), .CO(C[201]) );
  FA_823 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(B[201]), .CI(
        C[201]), .S(S[201]), .CO(C[202]) );
  FA_822 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(B[202]), .CI(
        C[202]), .S(S[202]), .CO(C[203]) );
  FA_821 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(B[203]), .CI(
        C[203]), .S(S[203]), .CO(C[204]) );
  FA_820 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(B[204]), .CI(
        C[204]), .S(S[204]), .CO(C[205]) );
  FA_819 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(B[205]), .CI(
        C[205]), .S(S[205]), .CO(C[206]) );
  FA_818 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(B[206]), .CI(
        C[206]), .S(S[206]), .CO(C[207]) );
  FA_817 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(B[207]), .CI(
        C[207]), .S(S[207]), .CO(C[208]) );
  FA_816 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(B[208]), .CI(
        C[208]), .S(S[208]), .CO(C[209]) );
  FA_815 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(B[209]), .CI(
        C[209]), .S(S[209]), .CO(C[210]) );
  FA_814 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(B[210]), .CI(
        C[210]), .S(S[210]), .CO(C[211]) );
  FA_813 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(B[211]), .CI(
        C[211]), .S(S[211]), .CO(C[212]) );
  FA_812 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(B[212]), .CI(
        C[212]), .S(S[212]), .CO(C[213]) );
  FA_811 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(B[213]), .CI(
        C[213]), .S(S[213]), .CO(C[214]) );
  FA_810 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(B[214]), .CI(
        C[214]), .S(S[214]), .CO(C[215]) );
  FA_809 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(B[215]), .CI(
        C[215]), .S(S[215]), .CO(C[216]) );
  FA_808 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(B[216]), .CI(
        C[216]), .S(S[216]), .CO(C[217]) );
  FA_807 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(B[217]), .CI(
        C[217]), .S(S[217]), .CO(C[218]) );
  FA_806 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(B[218]), .CI(
        C[218]), .S(S[218]), .CO(C[219]) );
  FA_805 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(B[219]), .CI(
        C[219]), .S(S[219]), .CO(C[220]) );
  FA_804 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(B[220]), .CI(
        C[220]), .S(S[220]), .CO(C[221]) );
  FA_803 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(B[221]), .CI(
        C[221]), .S(S[221]), .CO(C[222]) );
  FA_802 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(B[222]), .CI(
        C[222]), .S(S[222]), .CO(C[223]) );
  FA_801 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(B[223]), .CI(
        C[223]), .S(S[223]), .CO(C[224]) );
  FA_800 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(B[224]), .CI(
        C[224]), .S(S[224]), .CO(C[225]) );
  FA_799 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(B[225]), .CI(
        C[225]), .S(S[225]), .CO(C[226]) );
  FA_798 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(B[226]), .CI(
        C[226]), .S(S[226]), .CO(C[227]) );
  FA_797 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(B[227]), .CI(
        C[227]), .S(S[227]), .CO(C[228]) );
  FA_796 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(B[228]), .CI(
        C[228]), .S(S[228]), .CO(C[229]) );
  FA_795 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(B[229]), .CI(
        C[229]), .S(S[229]), .CO(C[230]) );
  FA_794 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(B[230]), .CI(
        C[230]), .S(S[230]), .CO(C[231]) );
  FA_793 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(B[231]), .CI(
        C[231]), .S(S[231]), .CO(C[232]) );
  FA_792 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(B[232]), .CI(
        C[232]), .S(S[232]), .CO(C[233]) );
  FA_791 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(B[233]), .CI(
        C[233]), .S(S[233]), .CO(C[234]) );
  FA_790 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(B[234]), .CI(
        C[234]), .S(S[234]), .CO(C[235]) );
  FA_789 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(B[235]), .CI(
        C[235]), .S(S[235]), .CO(C[236]) );
  FA_788 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(B[236]), .CI(
        C[236]), .S(S[236]), .CO(C[237]) );
  FA_787 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(B[237]), .CI(
        C[237]), .S(S[237]), .CO(C[238]) );
  FA_786 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(B[238]), .CI(
        C[238]), .S(S[238]), .CO(C[239]) );
  FA_785 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(B[239]), .CI(
        C[239]), .S(S[239]), .CO(C[240]) );
  FA_784 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(B[240]), .CI(
        C[240]), .S(S[240]), .CO(C[241]) );
  FA_783 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(B[241]), .CI(
        C[241]), .S(S[241]), .CO(C[242]) );
  FA_782 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(B[242]), .CI(
        C[242]), .S(S[242]), .CO(C[243]) );
  FA_781 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(B[243]), .CI(
        C[243]), .S(S[243]), .CO(C[244]) );
  FA_780 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(B[244]), .CI(
        C[244]), .S(S[244]), .CO(C[245]) );
  FA_779 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(B[245]), .CI(
        C[245]), .S(S[245]), .CO(C[246]) );
  FA_778 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(B[246]), .CI(
        C[246]), .S(S[246]), .CO(C[247]) );
  FA_777 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(B[247]), .CI(
        C[247]), .S(S[247]), .CO(C[248]) );
  FA_776 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(B[248]), .CI(
        C[248]), .S(S[248]), .CO(C[249]) );
  FA_775 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(B[249]), .CI(
        C[249]), .S(S[249]), .CO(C[250]) );
  FA_774 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(B[250]), .CI(
        C[250]), .S(S[250]), .CO(C[251]) );
  FA_773 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(B[251]), .CI(
        C[251]), .S(S[251]), .CO(C[252]) );
  FA_772 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(B[252]), .CI(
        C[252]), .S(S[252]), .CO(C[253]) );
  FA_771 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(B[253]), .CI(
        C[253]), .S(S[253]), .CO(C[254]) );
  FA_770 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(B[254]), .CI(
        C[254]), .S(S[254]), .CO(C[255]) );
  FA_769 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(B[255]), .CI(
        C[255]), .S(S[255]), .CO(C[256]) );
  FA_768 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(B[256]), .CI(
        C[256]), .S(S[256]), .CO(C[257]) );
  FA_767 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(B[257]), .CI(
        C[257]), .S(S[257]), .CO(C[258]) );
  FA_766 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(B[258]), .CI(
        C[258]), .S(S[258]), .CO(C[259]) );
  FA_765 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(B[259]), .CI(
        C[259]), .S(S[259]), .CO(C[260]) );
  FA_764 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(B[260]), .CI(
        C[260]), .S(S[260]), .CO(C[261]) );
  FA_763 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(B[261]), .CI(
        C[261]), .S(S[261]), .CO(C[262]) );
  FA_762 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(B[262]), .CI(
        C[262]), .S(S[262]), .CO(C[263]) );
  FA_761 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(B[263]), .CI(
        C[263]), .S(S[263]), .CO(C[264]) );
  FA_760 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(B[264]), .CI(
        C[264]), .S(S[264]), .CO(C[265]) );
  FA_759 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(B[265]), .CI(
        C[265]), .S(S[265]), .CO(C[266]) );
  FA_758 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(B[266]), .CI(
        C[266]), .S(S[266]), .CO(C[267]) );
  FA_757 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(B[267]), .CI(
        C[267]), .S(S[267]), .CO(C[268]) );
  FA_756 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(B[268]), .CI(
        C[268]), .S(S[268]), .CO(C[269]) );
  FA_755 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(B[269]), .CI(
        C[269]), .S(S[269]), .CO(C[270]) );
  FA_754 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(B[270]), .CI(
        C[270]), .S(S[270]), .CO(C[271]) );
  FA_753 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(B[271]), .CI(
        C[271]), .S(S[271]), .CO(C[272]) );
  FA_752 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(B[272]), .CI(
        C[272]), .S(S[272]), .CO(C[273]) );
  FA_751 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(B[273]), .CI(
        C[273]), .S(S[273]), .CO(C[274]) );
  FA_750 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(B[274]), .CI(
        C[274]), .S(S[274]), .CO(C[275]) );
  FA_749 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(B[275]), .CI(
        C[275]), .S(S[275]), .CO(C[276]) );
  FA_748 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(B[276]), .CI(
        C[276]), .S(S[276]), .CO(C[277]) );
  FA_747 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(B[277]), .CI(
        C[277]), .S(S[277]), .CO(C[278]) );
  FA_746 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(B[278]), .CI(
        C[278]), .S(S[278]), .CO(C[279]) );
  FA_745 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(B[279]), .CI(
        C[279]), .S(S[279]), .CO(C[280]) );
  FA_744 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(B[280]), .CI(
        C[280]), .S(S[280]), .CO(C[281]) );
  FA_743 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(B[281]), .CI(
        C[281]), .S(S[281]), .CO(C[282]) );
  FA_742 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(B[282]), .CI(
        C[282]), .S(S[282]), .CO(C[283]) );
  FA_741 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(B[283]), .CI(
        C[283]), .S(S[283]), .CO(C[284]) );
  FA_740 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(B[284]), .CI(
        C[284]), .S(S[284]), .CO(C[285]) );
  FA_739 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(B[285]), .CI(
        C[285]), .S(S[285]), .CO(C[286]) );
  FA_738 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(B[286]), .CI(
        C[286]), .S(S[286]), .CO(C[287]) );
  FA_737 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(B[287]), .CI(
        C[287]), .S(S[287]), .CO(C[288]) );
  FA_736 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(B[288]), .CI(
        C[288]), .S(S[288]), .CO(C[289]) );
  FA_735 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(B[289]), .CI(
        C[289]), .S(S[289]), .CO(C[290]) );
  FA_734 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(B[290]), .CI(
        C[290]), .S(S[290]), .CO(C[291]) );
  FA_733 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(B[291]), .CI(
        C[291]), .S(S[291]), .CO(C[292]) );
  FA_732 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(B[292]), .CI(
        C[292]), .S(S[292]), .CO(C[293]) );
  FA_731 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(B[293]), .CI(
        C[293]), .S(S[293]), .CO(C[294]) );
  FA_730 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(B[294]), .CI(
        C[294]), .S(S[294]), .CO(C[295]) );
  FA_729 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(B[295]), .CI(
        C[295]), .S(S[295]), .CO(C[296]) );
  FA_728 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(B[296]), .CI(
        C[296]), .S(S[296]), .CO(C[297]) );
  FA_727 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(B[297]), .CI(
        C[297]), .S(S[297]), .CO(C[298]) );
  FA_726 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(B[298]), .CI(
        C[298]), .S(S[298]), .CO(C[299]) );
  FA_725 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(B[299]), .CI(
        C[299]), .S(S[299]), .CO(C[300]) );
  FA_724 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(B[300]), .CI(
        C[300]), .S(S[300]), .CO(C[301]) );
  FA_723 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(B[301]), .CI(
        C[301]), .S(S[301]), .CO(C[302]) );
  FA_722 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(B[302]), .CI(
        C[302]), .S(S[302]), .CO(C[303]) );
  FA_721 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(B[303]), .CI(
        C[303]), .S(S[303]), .CO(C[304]) );
  FA_720 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(B[304]), .CI(
        C[304]), .S(S[304]), .CO(C[305]) );
  FA_719 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(B[305]), .CI(
        C[305]), .S(S[305]), .CO(C[306]) );
  FA_718 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(B[306]), .CI(
        C[306]), .S(S[306]), .CO(C[307]) );
  FA_717 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(B[307]), .CI(
        C[307]), .S(S[307]), .CO(C[308]) );
  FA_716 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(B[308]), .CI(
        C[308]), .S(S[308]), .CO(C[309]) );
  FA_715 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(B[309]), .CI(
        C[309]), .S(S[309]), .CO(C[310]) );
  FA_714 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(B[310]), .CI(
        C[310]), .S(S[310]), .CO(C[311]) );
  FA_713 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(B[311]), .CI(
        C[311]), .S(S[311]), .CO(C[312]) );
  FA_712 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(B[312]), .CI(
        C[312]), .S(S[312]), .CO(C[313]) );
  FA_711 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(B[313]), .CI(
        C[313]), .S(S[313]), .CO(C[314]) );
  FA_710 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(B[314]), .CI(
        C[314]), .S(S[314]), .CO(C[315]) );
  FA_709 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(B[315]), .CI(
        C[315]), .S(S[315]), .CO(C[316]) );
  FA_708 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(B[316]), .CI(
        C[316]), .S(S[316]), .CO(C[317]) );
  FA_707 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(B[317]), .CI(
        C[317]), .S(S[317]), .CO(C[318]) );
  FA_706 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(B[318]), .CI(
        C[318]), .S(S[318]), .CO(C[319]) );
  FA_705 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(B[319]), .CI(
        C[319]), .S(S[319]), .CO(C[320]) );
  FA_704 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(B[320]), .CI(
        C[320]), .S(S[320]), .CO(C[321]) );
  FA_703 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(B[321]), .CI(
        C[321]), .S(S[321]), .CO(C[322]) );
  FA_702 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(B[322]), .CI(
        C[322]), .S(S[322]), .CO(C[323]) );
  FA_701 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(B[323]), .CI(
        C[323]), .S(S[323]), .CO(C[324]) );
  FA_700 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(B[324]), .CI(
        C[324]), .S(S[324]), .CO(C[325]) );
  FA_699 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(B[325]), .CI(
        C[325]), .S(S[325]), .CO(C[326]) );
  FA_698 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(B[326]), .CI(
        C[326]), .S(S[326]), .CO(C[327]) );
  FA_697 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(B[327]), .CI(
        C[327]), .S(S[327]), .CO(C[328]) );
  FA_696 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(B[328]), .CI(
        C[328]), .S(S[328]), .CO(C[329]) );
  FA_695 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(B[329]), .CI(
        C[329]), .S(S[329]), .CO(C[330]) );
  FA_694 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(B[330]), .CI(
        C[330]), .S(S[330]), .CO(C[331]) );
  FA_693 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(B[331]), .CI(
        C[331]), .S(S[331]), .CO(C[332]) );
  FA_692 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(B[332]), .CI(
        C[332]), .S(S[332]), .CO(C[333]) );
  FA_691 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(B[333]), .CI(
        C[333]), .S(S[333]), .CO(C[334]) );
  FA_690 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(B[334]), .CI(
        C[334]), .S(S[334]), .CO(C[335]) );
  FA_689 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(B[335]), .CI(
        C[335]), .S(S[335]), .CO(C[336]) );
  FA_688 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(B[336]), .CI(
        C[336]), .S(S[336]), .CO(C[337]) );
  FA_687 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(B[337]), .CI(
        C[337]), .S(S[337]), .CO(C[338]) );
  FA_686 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(B[338]), .CI(
        C[338]), .S(S[338]), .CO(C[339]) );
  FA_685 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(B[339]), .CI(
        C[339]), .S(S[339]), .CO(C[340]) );
  FA_684 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(B[340]), .CI(
        C[340]), .S(S[340]), .CO(C[341]) );
  FA_683 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(B[341]), .CI(
        C[341]), .S(S[341]), .CO(C[342]) );
  FA_682 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(B[342]), .CI(
        C[342]), .S(S[342]), .CO(C[343]) );
  FA_681 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(B[343]), .CI(
        C[343]), .S(S[343]), .CO(C[344]) );
  FA_680 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(B[344]), .CI(
        C[344]), .S(S[344]), .CO(C[345]) );
  FA_679 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(B[345]), .CI(
        C[345]), .S(S[345]), .CO(C[346]) );
  FA_678 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(B[346]), .CI(
        C[346]), .S(S[346]), .CO(C[347]) );
  FA_677 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(B[347]), .CI(
        C[347]), .S(S[347]), .CO(C[348]) );
  FA_676 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(B[348]), .CI(
        C[348]), .S(S[348]), .CO(C[349]) );
  FA_675 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(B[349]), .CI(
        C[349]), .S(S[349]), .CO(C[350]) );
  FA_674 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(B[350]), .CI(
        C[350]), .S(S[350]), .CO(C[351]) );
  FA_673 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(B[351]), .CI(
        C[351]), .S(S[351]), .CO(C[352]) );
  FA_672 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(B[352]), .CI(
        C[352]), .S(S[352]), .CO(C[353]) );
  FA_671 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(B[353]), .CI(
        C[353]), .S(S[353]), .CO(C[354]) );
  FA_670 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(B[354]), .CI(
        C[354]), .S(S[354]), .CO(C[355]) );
  FA_669 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(B[355]), .CI(
        C[355]), .S(S[355]), .CO(C[356]) );
  FA_668 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(B[356]), .CI(
        C[356]), .S(S[356]), .CO(C[357]) );
  FA_667 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(B[357]), .CI(
        C[357]), .S(S[357]), .CO(C[358]) );
  FA_666 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(B[358]), .CI(
        C[358]), .S(S[358]), .CO(C[359]) );
  FA_665 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(B[359]), .CI(
        C[359]), .S(S[359]), .CO(C[360]) );
  FA_664 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(B[360]), .CI(
        C[360]), .S(S[360]), .CO(C[361]) );
  FA_663 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(B[361]), .CI(
        C[361]), .S(S[361]), .CO(C[362]) );
  FA_662 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(B[362]), .CI(
        C[362]), .S(S[362]), .CO(C[363]) );
  FA_661 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(B[363]), .CI(
        C[363]), .S(S[363]), .CO(C[364]) );
  FA_660 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(B[364]), .CI(
        C[364]), .S(S[364]), .CO(C[365]) );
  FA_659 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(B[365]), .CI(
        C[365]), .S(S[365]), .CO(C[366]) );
  FA_658 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(B[366]), .CI(
        C[366]), .S(S[366]), .CO(C[367]) );
  FA_657 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(B[367]), .CI(
        C[367]), .S(S[367]), .CO(C[368]) );
  FA_656 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(B[368]), .CI(
        C[368]), .S(S[368]), .CO(C[369]) );
  FA_655 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(B[369]), .CI(
        C[369]), .S(S[369]), .CO(C[370]) );
  FA_654 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(B[370]), .CI(
        C[370]), .S(S[370]), .CO(C[371]) );
  FA_653 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(B[371]), .CI(
        C[371]), .S(S[371]), .CO(C[372]) );
  FA_652 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(B[372]), .CI(
        C[372]), .S(S[372]), .CO(C[373]) );
  FA_651 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(B[373]), .CI(
        C[373]), .S(S[373]), .CO(C[374]) );
  FA_650 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(B[374]), .CI(
        C[374]), .S(S[374]), .CO(C[375]) );
  FA_649 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(B[375]), .CI(
        C[375]), .S(S[375]), .CO(C[376]) );
  FA_648 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(B[376]), .CI(
        C[376]), .S(S[376]), .CO(C[377]) );
  FA_647 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(B[377]), .CI(
        C[377]), .S(S[377]), .CO(C[378]) );
  FA_646 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(B[378]), .CI(
        C[378]), .S(S[378]), .CO(C[379]) );
  FA_645 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(B[379]), .CI(
        C[379]), .S(S[379]), .CO(C[380]) );
  FA_644 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(B[380]), .CI(
        C[380]), .S(S[380]), .CO(C[381]) );
  FA_643 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(B[381]), .CI(
        C[381]), .S(S[381]), .CO(C[382]) );
  FA_642 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(B[382]), .CI(
        C[382]), .S(S[382]), .CO(C[383]) );
  FA_641 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(B[383]), .CI(
        C[383]), .S(S[383]), .CO(C[384]) );
  FA_640 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(B[384]), .CI(
        C[384]), .S(S[384]), .CO(C[385]) );
  FA_639 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(B[385]), .CI(
        C[385]), .S(S[385]), .CO(C[386]) );
  FA_638 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(B[386]), .CI(
        C[386]), .S(S[386]), .CO(C[387]) );
  FA_637 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(B[387]), .CI(
        C[387]), .S(S[387]), .CO(C[388]) );
  FA_636 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(B[388]), .CI(
        C[388]), .S(S[388]), .CO(C[389]) );
  FA_635 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(B[389]), .CI(
        C[389]), .S(S[389]), .CO(C[390]) );
  FA_634 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(B[390]), .CI(
        C[390]), .S(S[390]), .CO(C[391]) );
  FA_633 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(B[391]), .CI(
        C[391]), .S(S[391]), .CO(C[392]) );
  FA_632 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(B[392]), .CI(
        C[392]), .S(S[392]), .CO(C[393]) );
  FA_631 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(B[393]), .CI(
        C[393]), .S(S[393]), .CO(C[394]) );
  FA_630 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(B[394]), .CI(
        C[394]), .S(S[394]), .CO(C[395]) );
  FA_629 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(B[395]), .CI(
        C[395]), .S(S[395]), .CO(C[396]) );
  FA_628 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(B[396]), .CI(
        C[396]), .S(S[396]), .CO(C[397]) );
  FA_627 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(B[397]), .CI(
        C[397]), .S(S[397]), .CO(C[398]) );
  FA_626 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(B[398]), .CI(
        C[398]), .S(S[398]), .CO(C[399]) );
  FA_625 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(B[399]), .CI(
        C[399]), .S(S[399]), .CO(C[400]) );
  FA_624 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(B[400]), .CI(
        C[400]), .S(S[400]), .CO(C[401]) );
  FA_623 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(B[401]), .CI(
        C[401]), .S(S[401]), .CO(C[402]) );
  FA_622 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(B[402]), .CI(
        C[402]), .S(S[402]), .CO(C[403]) );
  FA_621 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(B[403]), .CI(
        C[403]), .S(S[403]), .CO(C[404]) );
  FA_620 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(B[404]), .CI(
        C[404]), .S(S[404]), .CO(C[405]) );
  FA_619 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(B[405]), .CI(
        C[405]), .S(S[405]), .CO(C[406]) );
  FA_618 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(B[406]), .CI(
        C[406]), .S(S[406]), .CO(C[407]) );
  FA_617 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(B[407]), .CI(
        C[407]), .S(S[407]), .CO(C[408]) );
  FA_616 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(B[408]), .CI(
        C[408]), .S(S[408]), .CO(C[409]) );
  FA_615 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(B[409]), .CI(
        C[409]), .S(S[409]), .CO(C[410]) );
  FA_614 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(B[410]), .CI(
        C[410]), .S(S[410]), .CO(C[411]) );
  FA_613 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(B[411]), .CI(
        C[411]), .S(S[411]), .CO(C[412]) );
  FA_612 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(B[412]), .CI(
        C[412]), .S(S[412]), .CO(C[413]) );
  FA_611 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(B[413]), .CI(
        C[413]), .S(S[413]), .CO(C[414]) );
  FA_610 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(B[414]), .CI(
        C[414]), .S(S[414]), .CO(C[415]) );
  FA_609 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(B[415]), .CI(
        C[415]), .S(S[415]), .CO(C[416]) );
  FA_608 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(B[416]), .CI(
        C[416]), .S(S[416]), .CO(C[417]) );
  FA_607 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(B[417]), .CI(
        C[417]), .S(S[417]), .CO(C[418]) );
  FA_606 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(B[418]), .CI(
        C[418]), .S(S[418]), .CO(C[419]) );
  FA_605 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(B[419]), .CI(
        C[419]), .S(S[419]), .CO(C[420]) );
  FA_604 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(B[420]), .CI(
        C[420]), .S(S[420]), .CO(C[421]) );
  FA_603 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(B[421]), .CI(
        C[421]), .S(S[421]), .CO(C[422]) );
  FA_602 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(B[422]), .CI(
        C[422]), .S(S[422]), .CO(C[423]) );
  FA_601 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(B[423]), .CI(
        C[423]), .S(S[423]), .CO(C[424]) );
  FA_600 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(B[424]), .CI(
        C[424]), .S(S[424]), .CO(C[425]) );
  FA_599 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(B[425]), .CI(
        C[425]), .S(S[425]), .CO(C[426]) );
  FA_598 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(B[426]), .CI(
        C[426]), .S(S[426]), .CO(C[427]) );
  FA_597 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(B[427]), .CI(
        C[427]), .S(S[427]), .CO(C[428]) );
  FA_596 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(B[428]), .CI(
        C[428]), .S(S[428]), .CO(C[429]) );
  FA_595 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(B[429]), .CI(
        C[429]), .S(S[429]), .CO(C[430]) );
  FA_594 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(B[430]), .CI(
        C[430]), .S(S[430]), .CO(C[431]) );
  FA_593 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(B[431]), .CI(
        C[431]), .S(S[431]), .CO(C[432]) );
  FA_592 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(B[432]), .CI(
        C[432]), .S(S[432]), .CO(C[433]) );
  FA_591 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(B[433]), .CI(
        C[433]), .S(S[433]), .CO(C[434]) );
  FA_590 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(B[434]), .CI(
        C[434]), .S(S[434]), .CO(C[435]) );
  FA_589 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(B[435]), .CI(
        C[435]), .S(S[435]), .CO(C[436]) );
  FA_588 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(B[436]), .CI(
        C[436]), .S(S[436]), .CO(C[437]) );
  FA_587 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(B[437]), .CI(
        C[437]), .S(S[437]), .CO(C[438]) );
  FA_586 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(B[438]), .CI(
        C[438]), .S(S[438]), .CO(C[439]) );
  FA_585 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(B[439]), .CI(
        C[439]), .S(S[439]), .CO(C[440]) );
  FA_584 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(B[440]), .CI(
        C[440]), .S(S[440]), .CO(C[441]) );
  FA_583 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(B[441]), .CI(
        C[441]), .S(S[441]), .CO(C[442]) );
  FA_582 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(B[442]), .CI(
        C[442]), .S(S[442]), .CO(C[443]) );
  FA_581 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(B[443]), .CI(
        C[443]), .S(S[443]), .CO(C[444]) );
  FA_580 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(B[444]), .CI(
        C[444]), .S(S[444]), .CO(C[445]) );
  FA_579 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(B[445]), .CI(
        C[445]), .S(S[445]), .CO(C[446]) );
  FA_578 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(B[446]), .CI(
        C[446]), .S(S[446]), .CO(C[447]) );
  FA_577 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(B[447]), .CI(
        C[447]), .S(S[447]), .CO(C[448]) );
  FA_576 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(B[448]), .CI(
        C[448]), .S(S[448]), .CO(C[449]) );
  FA_575 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(B[449]), .CI(
        C[449]), .S(S[449]), .CO(C[450]) );
  FA_574 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(B[450]), .CI(
        C[450]), .S(S[450]), .CO(C[451]) );
  FA_573 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(B[451]), .CI(
        C[451]), .S(S[451]), .CO(C[452]) );
  FA_572 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(B[452]), .CI(
        C[452]), .S(S[452]), .CO(C[453]) );
  FA_571 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(B[453]), .CI(
        C[453]), .S(S[453]), .CO(C[454]) );
  FA_570 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(B[454]), .CI(
        C[454]), .S(S[454]), .CO(C[455]) );
  FA_569 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(B[455]), .CI(
        C[455]), .S(S[455]), .CO(C[456]) );
  FA_568 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(B[456]), .CI(
        C[456]), .S(S[456]), .CO(C[457]) );
  FA_567 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(B[457]), .CI(
        C[457]), .S(S[457]), .CO(C[458]) );
  FA_566 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(B[458]), .CI(
        C[458]), .S(S[458]), .CO(C[459]) );
  FA_565 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(B[459]), .CI(
        C[459]), .S(S[459]), .CO(C[460]) );
  FA_564 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(B[460]), .CI(
        C[460]), .S(S[460]), .CO(C[461]) );
  FA_563 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(B[461]), .CI(
        C[461]), .S(S[461]), .CO(C[462]) );
  FA_562 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(B[462]), .CI(
        C[462]), .S(S[462]), .CO(C[463]) );
  FA_561 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(B[463]), .CI(
        C[463]), .S(S[463]), .CO(C[464]) );
  FA_560 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(B[464]), .CI(
        C[464]), .S(S[464]), .CO(C[465]) );
  FA_559 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(B[465]), .CI(
        C[465]), .S(S[465]), .CO(C[466]) );
  FA_558 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(B[466]), .CI(
        C[466]), .S(S[466]), .CO(C[467]) );
  FA_557 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(B[467]), .CI(
        C[467]), .S(S[467]), .CO(C[468]) );
  FA_556 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(B[468]), .CI(
        C[468]), .S(S[468]), .CO(C[469]) );
  FA_555 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(B[469]), .CI(
        C[469]), .S(S[469]), .CO(C[470]) );
  FA_554 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(B[470]), .CI(
        C[470]), .S(S[470]), .CO(C[471]) );
  FA_553 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(B[471]), .CI(
        C[471]), .S(S[471]), .CO(C[472]) );
  FA_552 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(B[472]), .CI(
        C[472]), .S(S[472]), .CO(C[473]) );
  FA_551 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(B[473]), .CI(
        C[473]), .S(S[473]), .CO(C[474]) );
  FA_550 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(B[474]), .CI(
        C[474]), .S(S[474]), .CO(C[475]) );
  FA_549 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(B[475]), .CI(
        C[475]), .S(S[475]), .CO(C[476]) );
  FA_548 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(B[476]), .CI(
        C[476]), .S(S[476]), .CO(C[477]) );
  FA_547 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(B[477]), .CI(
        C[477]), .S(S[477]), .CO(C[478]) );
  FA_546 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(B[478]), .CI(
        C[478]), .S(S[478]), .CO(C[479]) );
  FA_545 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(B[479]), .CI(
        C[479]), .S(S[479]), .CO(C[480]) );
  FA_544 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(B[480]), .CI(
        C[480]), .S(S[480]), .CO(C[481]) );
  FA_543 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(B[481]), .CI(
        C[481]), .S(S[481]), .CO(C[482]) );
  FA_542 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(B[482]), .CI(
        C[482]), .S(S[482]), .CO(C[483]) );
  FA_541 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(B[483]), .CI(
        C[483]), .S(S[483]), .CO(C[484]) );
  FA_540 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(B[484]), .CI(
        C[484]), .S(S[484]), .CO(C[485]) );
  FA_539 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(B[485]), .CI(
        C[485]), .S(S[485]), .CO(C[486]) );
  FA_538 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(B[486]), .CI(
        C[486]), .S(S[486]), .CO(C[487]) );
  FA_537 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(B[487]), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_536 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(B[488]), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_535 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(B[489]), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_534 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(B[490]), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_533 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(B[491]), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_532 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(B[492]), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_531 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(B[493]), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_530 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(B[494]), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_529 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(B[495]), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_528 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(B[496]), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_527 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(B[497]), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_526 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(B[498]), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_525 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(B[499]), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_524 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(B[500]), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_523 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(B[501]), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_522 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(B[502]), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_521 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(B[503]), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_520 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(B[504]), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_519 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(B[505]), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_518 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(B[506]), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_517 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(B[507]), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_516 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(B[508]), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_515 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(B[509]), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_514 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(B[510]), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_513 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(B[511]), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_512 \FA_INST_0[1].FA_INST_1[0].FA_  ( .A(A[512]), .B(B[512]), .CI(C[512]), 
        .S(S[512]), .CO(C[513]) );
  FA_511 \FA_INST_0[1].FA_INST_1[1].FA_  ( .A(A[513]), .B(B[513]), .CI(C[513]), 
        .S(S[513]), .CO(C[514]) );
  FA_510 \FA_INST_0[1].FA_INST_1[2].FA_  ( .A(A[514]), .B(B[514]), .CI(C[514]), 
        .S(S[514]), .CO(C[515]) );
  FA_509 \FA_INST_0[1].FA_INST_1[3].FA_  ( .A(A[515]), .B(B[515]), .CI(C[515]), 
        .S(S[515]), .CO(C[516]) );
  FA_508 \FA_INST_0[1].FA_INST_1[4].FA_  ( .A(A[516]), .B(B[516]), .CI(C[516]), 
        .S(S[516]), .CO(C[517]) );
  FA_507 \FA_INST_0[1].FA_INST_1[5].FA_  ( .A(A[517]), .B(B[517]), .CI(C[517]), 
        .S(S[517]), .CO(C[518]) );
  FA_506 \FA_INST_0[1].FA_INST_1[6].FA_  ( .A(A[518]), .B(B[518]), .CI(C[518]), 
        .S(S[518]), .CO(C[519]) );
  FA_505 \FA_INST_0[1].FA_INST_1[7].FA_  ( .A(A[519]), .B(B[519]), .CI(C[519]), 
        .S(S[519]), .CO(C[520]) );
  FA_504 \FA_INST_0[1].FA_INST_1[8].FA_  ( .A(A[520]), .B(B[520]), .CI(C[520]), 
        .S(S[520]), .CO(C[521]) );
  FA_503 \FA_INST_0[1].FA_INST_1[9].FA_  ( .A(A[521]), .B(B[521]), .CI(C[521]), 
        .S(S[521]), .CO(C[522]) );
  FA_502 \FA_INST_0[1].FA_INST_1[10].FA_  ( .A(A[522]), .B(B[522]), .CI(C[522]), .S(S[522]), .CO(C[523]) );
  FA_501 \FA_INST_0[1].FA_INST_1[11].FA_  ( .A(A[523]), .B(B[523]), .CI(C[523]), .S(S[523]), .CO(C[524]) );
  FA_500 \FA_INST_0[1].FA_INST_1[12].FA_  ( .A(A[524]), .B(B[524]), .CI(C[524]), .S(S[524]), .CO(C[525]) );
  FA_499 \FA_INST_0[1].FA_INST_1[13].FA_  ( .A(A[525]), .B(B[525]), .CI(C[525]), .S(S[525]), .CO(C[526]) );
  FA_498 \FA_INST_0[1].FA_INST_1[14].FA_  ( .A(A[526]), .B(B[526]), .CI(C[526]), .S(S[526]), .CO(C[527]) );
  FA_497 \FA_INST_0[1].FA_INST_1[15].FA_  ( .A(A[527]), .B(B[527]), .CI(C[527]), .S(S[527]), .CO(C[528]) );
  FA_496 \FA_INST_0[1].FA_INST_1[16].FA_  ( .A(A[528]), .B(B[528]), .CI(C[528]), .S(S[528]), .CO(C[529]) );
  FA_495 \FA_INST_0[1].FA_INST_1[17].FA_  ( .A(A[529]), .B(B[529]), .CI(C[529]), .S(S[529]), .CO(C[530]) );
  FA_494 \FA_INST_0[1].FA_INST_1[18].FA_  ( .A(A[530]), .B(B[530]), .CI(C[530]), .S(S[530]), .CO(C[531]) );
  FA_493 \FA_INST_0[1].FA_INST_1[19].FA_  ( .A(A[531]), .B(B[531]), .CI(C[531]), .S(S[531]), .CO(C[532]) );
  FA_492 \FA_INST_0[1].FA_INST_1[20].FA_  ( .A(A[532]), .B(B[532]), .CI(C[532]), .S(S[532]), .CO(C[533]) );
  FA_491 \FA_INST_0[1].FA_INST_1[21].FA_  ( .A(A[533]), .B(B[533]), .CI(C[533]), .S(S[533]), .CO(C[534]) );
  FA_490 \FA_INST_0[1].FA_INST_1[22].FA_  ( .A(A[534]), .B(B[534]), .CI(C[534]), .S(S[534]), .CO(C[535]) );
  FA_489 \FA_INST_0[1].FA_INST_1[23].FA_  ( .A(A[535]), .B(B[535]), .CI(C[535]), .S(S[535]), .CO(C[536]) );
  FA_488 \FA_INST_0[1].FA_INST_1[24].FA_  ( .A(A[536]), .B(B[536]), .CI(C[536]), .S(S[536]), .CO(C[537]) );
  FA_487 \FA_INST_0[1].FA_INST_1[25].FA_  ( .A(A[537]), .B(B[537]), .CI(C[537]), .S(S[537]), .CO(C[538]) );
  FA_486 \FA_INST_0[1].FA_INST_1[26].FA_  ( .A(A[538]), .B(B[538]), .CI(C[538]), .S(S[538]), .CO(C[539]) );
  FA_485 \FA_INST_0[1].FA_INST_1[27].FA_  ( .A(A[539]), .B(B[539]), .CI(C[539]), .S(S[539]), .CO(C[540]) );
  FA_484 \FA_INST_0[1].FA_INST_1[28].FA_  ( .A(A[540]), .B(B[540]), .CI(C[540]), .S(S[540]), .CO(C[541]) );
  FA_483 \FA_INST_0[1].FA_INST_1[29].FA_  ( .A(A[541]), .B(B[541]), .CI(C[541]), .S(S[541]), .CO(C[542]) );
  FA_482 \FA_INST_0[1].FA_INST_1[30].FA_  ( .A(A[542]), .B(B[542]), .CI(C[542]), .S(S[542]), .CO(C[543]) );
  FA_481 \FA_INST_0[1].FA_INST_1[31].FA_  ( .A(A[543]), .B(B[543]), .CI(C[543]), .S(S[543]), .CO(C[544]) );
  FA_480 \FA_INST_0[1].FA_INST_1[32].FA_  ( .A(A[544]), .B(B[544]), .CI(C[544]), .S(S[544]), .CO(C[545]) );
  FA_479 \FA_INST_0[1].FA_INST_1[33].FA_  ( .A(A[545]), .B(B[545]), .CI(C[545]), .S(S[545]), .CO(C[546]) );
  FA_478 \FA_INST_0[1].FA_INST_1[34].FA_  ( .A(A[546]), .B(B[546]), .CI(C[546]), .S(S[546]), .CO(C[547]) );
  FA_477 \FA_INST_0[1].FA_INST_1[35].FA_  ( .A(A[547]), .B(B[547]), .CI(C[547]), .S(S[547]), .CO(C[548]) );
  FA_476 \FA_INST_0[1].FA_INST_1[36].FA_  ( .A(A[548]), .B(B[548]), .CI(C[548]), .S(S[548]), .CO(C[549]) );
  FA_475 \FA_INST_0[1].FA_INST_1[37].FA_  ( .A(A[549]), .B(B[549]), .CI(C[549]), .S(S[549]), .CO(C[550]) );
  FA_474 \FA_INST_0[1].FA_INST_1[38].FA_  ( .A(A[550]), .B(B[550]), .CI(C[550]), .S(S[550]), .CO(C[551]) );
  FA_473 \FA_INST_0[1].FA_INST_1[39].FA_  ( .A(A[551]), .B(B[551]), .CI(C[551]), .S(S[551]), .CO(C[552]) );
  FA_472 \FA_INST_0[1].FA_INST_1[40].FA_  ( .A(A[552]), .B(B[552]), .CI(C[552]), .S(S[552]), .CO(C[553]) );
  FA_471 \FA_INST_0[1].FA_INST_1[41].FA_  ( .A(A[553]), .B(B[553]), .CI(C[553]), .S(S[553]), .CO(C[554]) );
  FA_470 \FA_INST_0[1].FA_INST_1[42].FA_  ( .A(A[554]), .B(B[554]), .CI(C[554]), .S(S[554]), .CO(C[555]) );
  FA_469 \FA_INST_0[1].FA_INST_1[43].FA_  ( .A(A[555]), .B(B[555]), .CI(C[555]), .S(S[555]), .CO(C[556]) );
  FA_468 \FA_INST_0[1].FA_INST_1[44].FA_  ( .A(A[556]), .B(B[556]), .CI(C[556]), .S(S[556]), .CO(C[557]) );
  FA_467 \FA_INST_0[1].FA_INST_1[45].FA_  ( .A(A[557]), .B(B[557]), .CI(C[557]), .S(S[557]), .CO(C[558]) );
  FA_466 \FA_INST_0[1].FA_INST_1[46].FA_  ( .A(A[558]), .B(B[558]), .CI(C[558]), .S(S[558]), .CO(C[559]) );
  FA_465 \FA_INST_0[1].FA_INST_1[47].FA_  ( .A(A[559]), .B(B[559]), .CI(C[559]), .S(S[559]), .CO(C[560]) );
  FA_464 \FA_INST_0[1].FA_INST_1[48].FA_  ( .A(A[560]), .B(B[560]), .CI(C[560]), .S(S[560]), .CO(C[561]) );
  FA_463 \FA_INST_0[1].FA_INST_1[49].FA_  ( .A(A[561]), .B(B[561]), .CI(C[561]), .S(S[561]), .CO(C[562]) );
  FA_462 \FA_INST_0[1].FA_INST_1[50].FA_  ( .A(A[562]), .B(B[562]), .CI(C[562]), .S(S[562]), .CO(C[563]) );
  FA_461 \FA_INST_0[1].FA_INST_1[51].FA_  ( .A(A[563]), .B(B[563]), .CI(C[563]), .S(S[563]), .CO(C[564]) );
  FA_460 \FA_INST_0[1].FA_INST_1[52].FA_  ( .A(A[564]), .B(B[564]), .CI(C[564]), .S(S[564]), .CO(C[565]) );
  FA_459 \FA_INST_0[1].FA_INST_1[53].FA_  ( .A(A[565]), .B(B[565]), .CI(C[565]), .S(S[565]), .CO(C[566]) );
  FA_458 \FA_INST_0[1].FA_INST_1[54].FA_  ( .A(A[566]), .B(B[566]), .CI(C[566]), .S(S[566]), .CO(C[567]) );
  FA_457 \FA_INST_0[1].FA_INST_1[55].FA_  ( .A(A[567]), .B(B[567]), .CI(C[567]), .S(S[567]), .CO(C[568]) );
  FA_456 \FA_INST_0[1].FA_INST_1[56].FA_  ( .A(A[568]), .B(B[568]), .CI(C[568]), .S(S[568]), .CO(C[569]) );
  FA_455 \FA_INST_0[1].FA_INST_1[57].FA_  ( .A(A[569]), .B(B[569]), .CI(C[569]), .S(S[569]), .CO(C[570]) );
  FA_454 \FA_INST_0[1].FA_INST_1[58].FA_  ( .A(A[570]), .B(B[570]), .CI(C[570]), .S(S[570]), .CO(C[571]) );
  FA_453 \FA_INST_0[1].FA_INST_1[59].FA_  ( .A(A[571]), .B(B[571]), .CI(C[571]), .S(S[571]), .CO(C[572]) );
  FA_452 \FA_INST_0[1].FA_INST_1[60].FA_  ( .A(A[572]), .B(B[572]), .CI(C[572]), .S(S[572]), .CO(C[573]) );
  FA_451 \FA_INST_0[1].FA_INST_1[61].FA_  ( .A(A[573]), .B(B[573]), .CI(C[573]), .S(S[573]), .CO(C[574]) );
  FA_450 \FA_INST_0[1].FA_INST_1[62].FA_  ( .A(A[574]), .B(B[574]), .CI(C[574]), .S(S[574]), .CO(C[575]) );
  FA_449 \FA_INST_0[1].FA_INST_1[63].FA_  ( .A(A[575]), .B(B[575]), .CI(C[575]), .S(S[575]), .CO(C[576]) );
  FA_448 \FA_INST_0[1].FA_INST_1[64].FA_  ( .A(A[576]), .B(B[576]), .CI(C[576]), .S(S[576]), .CO(C[577]) );
  FA_447 \FA_INST_0[1].FA_INST_1[65].FA_  ( .A(A[577]), .B(B[577]), .CI(C[577]), .S(S[577]), .CO(C[578]) );
  FA_446 \FA_INST_0[1].FA_INST_1[66].FA_  ( .A(A[578]), .B(B[578]), .CI(C[578]), .S(S[578]), .CO(C[579]) );
  FA_445 \FA_INST_0[1].FA_INST_1[67].FA_  ( .A(A[579]), .B(B[579]), .CI(C[579]), .S(S[579]), .CO(C[580]) );
  FA_444 \FA_INST_0[1].FA_INST_1[68].FA_  ( .A(A[580]), .B(B[580]), .CI(C[580]), .S(S[580]), .CO(C[581]) );
  FA_443 \FA_INST_0[1].FA_INST_1[69].FA_  ( .A(A[581]), .B(B[581]), .CI(C[581]), .S(S[581]), .CO(C[582]) );
  FA_442 \FA_INST_0[1].FA_INST_1[70].FA_  ( .A(A[582]), .B(B[582]), .CI(C[582]), .S(S[582]), .CO(C[583]) );
  FA_441 \FA_INST_0[1].FA_INST_1[71].FA_  ( .A(A[583]), .B(B[583]), .CI(C[583]), .S(S[583]), .CO(C[584]) );
  FA_440 \FA_INST_0[1].FA_INST_1[72].FA_  ( .A(A[584]), .B(B[584]), .CI(C[584]), .S(S[584]), .CO(C[585]) );
  FA_439 \FA_INST_0[1].FA_INST_1[73].FA_  ( .A(A[585]), .B(B[585]), .CI(C[585]), .S(S[585]), .CO(C[586]) );
  FA_438 \FA_INST_0[1].FA_INST_1[74].FA_  ( .A(A[586]), .B(B[586]), .CI(C[586]), .S(S[586]), .CO(C[587]) );
  FA_437 \FA_INST_0[1].FA_INST_1[75].FA_  ( .A(A[587]), .B(B[587]), .CI(C[587]), .S(S[587]), .CO(C[588]) );
  FA_436 \FA_INST_0[1].FA_INST_1[76].FA_  ( .A(A[588]), .B(B[588]), .CI(C[588]), .S(S[588]), .CO(C[589]) );
  FA_435 \FA_INST_0[1].FA_INST_1[77].FA_  ( .A(A[589]), .B(B[589]), .CI(C[589]), .S(S[589]), .CO(C[590]) );
  FA_434 \FA_INST_0[1].FA_INST_1[78].FA_  ( .A(A[590]), .B(B[590]), .CI(C[590]), .S(S[590]), .CO(C[591]) );
  FA_433 \FA_INST_0[1].FA_INST_1[79].FA_  ( .A(A[591]), .B(B[591]), .CI(C[591]), .S(S[591]), .CO(C[592]) );
  FA_432 \FA_INST_0[1].FA_INST_1[80].FA_  ( .A(A[592]), .B(B[592]), .CI(C[592]), .S(S[592]), .CO(C[593]) );
  FA_431 \FA_INST_0[1].FA_INST_1[81].FA_  ( .A(A[593]), .B(B[593]), .CI(C[593]), .S(S[593]), .CO(C[594]) );
  FA_430 \FA_INST_0[1].FA_INST_1[82].FA_  ( .A(A[594]), .B(B[594]), .CI(C[594]), .S(S[594]), .CO(C[595]) );
  FA_429 \FA_INST_0[1].FA_INST_1[83].FA_  ( .A(A[595]), .B(B[595]), .CI(C[595]), .S(S[595]), .CO(C[596]) );
  FA_428 \FA_INST_0[1].FA_INST_1[84].FA_  ( .A(A[596]), .B(B[596]), .CI(C[596]), .S(S[596]), .CO(C[597]) );
  FA_427 \FA_INST_0[1].FA_INST_1[85].FA_  ( .A(A[597]), .B(B[597]), .CI(C[597]), .S(S[597]), .CO(C[598]) );
  FA_426 \FA_INST_0[1].FA_INST_1[86].FA_  ( .A(A[598]), .B(B[598]), .CI(C[598]), .S(S[598]), .CO(C[599]) );
  FA_425 \FA_INST_0[1].FA_INST_1[87].FA_  ( .A(A[599]), .B(B[599]), .CI(C[599]), .S(S[599]), .CO(C[600]) );
  FA_424 \FA_INST_0[1].FA_INST_1[88].FA_  ( .A(A[600]), .B(B[600]), .CI(C[600]), .S(S[600]), .CO(C[601]) );
  FA_423 \FA_INST_0[1].FA_INST_1[89].FA_  ( .A(A[601]), .B(B[601]), .CI(C[601]), .S(S[601]), .CO(C[602]) );
  FA_422 \FA_INST_0[1].FA_INST_1[90].FA_  ( .A(A[602]), .B(B[602]), .CI(C[602]), .S(S[602]), .CO(C[603]) );
  FA_421 \FA_INST_0[1].FA_INST_1[91].FA_  ( .A(A[603]), .B(B[603]), .CI(C[603]), .S(S[603]), .CO(C[604]) );
  FA_420 \FA_INST_0[1].FA_INST_1[92].FA_  ( .A(A[604]), .B(B[604]), .CI(C[604]), .S(S[604]), .CO(C[605]) );
  FA_419 \FA_INST_0[1].FA_INST_1[93].FA_  ( .A(A[605]), .B(B[605]), .CI(C[605]), .S(S[605]), .CO(C[606]) );
  FA_418 \FA_INST_0[1].FA_INST_1[94].FA_  ( .A(A[606]), .B(B[606]), .CI(C[606]), .S(S[606]), .CO(C[607]) );
  FA_417 \FA_INST_0[1].FA_INST_1[95].FA_  ( .A(A[607]), .B(B[607]), .CI(C[607]), .S(S[607]), .CO(C[608]) );
  FA_416 \FA_INST_0[1].FA_INST_1[96].FA_  ( .A(A[608]), .B(B[608]), .CI(C[608]), .S(S[608]), .CO(C[609]) );
  FA_415 \FA_INST_0[1].FA_INST_1[97].FA_  ( .A(A[609]), .B(B[609]), .CI(C[609]), .S(S[609]), .CO(C[610]) );
  FA_414 \FA_INST_0[1].FA_INST_1[98].FA_  ( .A(A[610]), .B(B[610]), .CI(C[610]), .S(S[610]), .CO(C[611]) );
  FA_413 \FA_INST_0[1].FA_INST_1[99].FA_  ( .A(A[611]), .B(B[611]), .CI(C[611]), .S(S[611]), .CO(C[612]) );
  FA_412 \FA_INST_0[1].FA_INST_1[100].FA_  ( .A(A[612]), .B(B[612]), .CI(
        C[612]), .S(S[612]), .CO(C[613]) );
  FA_411 \FA_INST_0[1].FA_INST_1[101].FA_  ( .A(A[613]), .B(B[613]), .CI(
        C[613]), .S(S[613]), .CO(C[614]) );
  FA_410 \FA_INST_0[1].FA_INST_1[102].FA_  ( .A(A[614]), .B(B[614]), .CI(
        C[614]), .S(S[614]), .CO(C[615]) );
  FA_409 \FA_INST_0[1].FA_INST_1[103].FA_  ( .A(A[615]), .B(B[615]), .CI(
        C[615]), .S(S[615]), .CO(C[616]) );
  FA_408 \FA_INST_0[1].FA_INST_1[104].FA_  ( .A(A[616]), .B(B[616]), .CI(
        C[616]), .S(S[616]), .CO(C[617]) );
  FA_407 \FA_INST_0[1].FA_INST_1[105].FA_  ( .A(A[617]), .B(B[617]), .CI(
        C[617]), .S(S[617]), .CO(C[618]) );
  FA_406 \FA_INST_0[1].FA_INST_1[106].FA_  ( .A(A[618]), .B(B[618]), .CI(
        C[618]), .S(S[618]), .CO(C[619]) );
  FA_405 \FA_INST_0[1].FA_INST_1[107].FA_  ( .A(A[619]), .B(B[619]), .CI(
        C[619]), .S(S[619]), .CO(C[620]) );
  FA_404 \FA_INST_0[1].FA_INST_1[108].FA_  ( .A(A[620]), .B(B[620]), .CI(
        C[620]), .S(S[620]), .CO(C[621]) );
  FA_403 \FA_INST_0[1].FA_INST_1[109].FA_  ( .A(A[621]), .B(B[621]), .CI(
        C[621]), .S(S[621]), .CO(C[622]) );
  FA_402 \FA_INST_0[1].FA_INST_1[110].FA_  ( .A(A[622]), .B(B[622]), .CI(
        C[622]), .S(S[622]), .CO(C[623]) );
  FA_401 \FA_INST_0[1].FA_INST_1[111].FA_  ( .A(A[623]), .B(B[623]), .CI(
        C[623]), .S(S[623]), .CO(C[624]) );
  FA_400 \FA_INST_0[1].FA_INST_1[112].FA_  ( .A(A[624]), .B(B[624]), .CI(
        C[624]), .S(S[624]), .CO(C[625]) );
  FA_399 \FA_INST_0[1].FA_INST_1[113].FA_  ( .A(A[625]), .B(B[625]), .CI(
        C[625]), .S(S[625]), .CO(C[626]) );
  FA_398 \FA_INST_0[1].FA_INST_1[114].FA_  ( .A(A[626]), .B(B[626]), .CI(
        C[626]), .S(S[626]), .CO(C[627]) );
  FA_397 \FA_INST_0[1].FA_INST_1[115].FA_  ( .A(A[627]), .B(B[627]), .CI(
        C[627]), .S(S[627]), .CO(C[628]) );
  FA_396 \FA_INST_0[1].FA_INST_1[116].FA_  ( .A(A[628]), .B(B[628]), .CI(
        C[628]), .S(S[628]), .CO(C[629]) );
  FA_395 \FA_INST_0[1].FA_INST_1[117].FA_  ( .A(A[629]), .B(B[629]), .CI(
        C[629]), .S(S[629]), .CO(C[630]) );
  FA_394 \FA_INST_0[1].FA_INST_1[118].FA_  ( .A(A[630]), .B(B[630]), .CI(
        C[630]), .S(S[630]), .CO(C[631]) );
  FA_393 \FA_INST_0[1].FA_INST_1[119].FA_  ( .A(A[631]), .B(B[631]), .CI(
        C[631]), .S(S[631]), .CO(C[632]) );
  FA_392 \FA_INST_0[1].FA_INST_1[120].FA_  ( .A(A[632]), .B(B[632]), .CI(
        C[632]), .S(S[632]), .CO(C[633]) );
  FA_391 \FA_INST_0[1].FA_INST_1[121].FA_  ( .A(A[633]), .B(B[633]), .CI(
        C[633]), .S(S[633]), .CO(C[634]) );
  FA_390 \FA_INST_0[1].FA_INST_1[122].FA_  ( .A(A[634]), .B(B[634]), .CI(
        C[634]), .S(S[634]), .CO(C[635]) );
  FA_389 \FA_INST_0[1].FA_INST_1[123].FA_  ( .A(A[635]), .B(B[635]), .CI(
        C[635]), .S(S[635]), .CO(C[636]) );
  FA_388 \FA_INST_0[1].FA_INST_1[124].FA_  ( .A(A[636]), .B(B[636]), .CI(
        C[636]), .S(S[636]), .CO(C[637]) );
  FA_387 \FA_INST_0[1].FA_INST_1[125].FA_  ( .A(A[637]), .B(B[637]), .CI(
        C[637]), .S(S[637]), .CO(C[638]) );
  FA_386 \FA_INST_0[1].FA_INST_1[126].FA_  ( .A(A[638]), .B(B[638]), .CI(
        C[638]), .S(S[638]), .CO(C[639]) );
  FA_385 \FA_INST_0[1].FA_INST_1[127].FA_  ( .A(A[639]), .B(B[639]), .CI(
        C[639]), .S(S[639]), .CO(C[640]) );
  FA_384 \FA_INST_0[1].FA_INST_1[128].FA_  ( .A(A[640]), .B(B[640]), .CI(
        C[640]), .S(S[640]), .CO(C[641]) );
  FA_383 \FA_INST_0[1].FA_INST_1[129].FA_  ( .A(A[641]), .B(B[641]), .CI(
        C[641]), .S(S[641]), .CO(C[642]) );
  FA_382 \FA_INST_0[1].FA_INST_1[130].FA_  ( .A(A[642]), .B(B[642]), .CI(
        C[642]), .S(S[642]), .CO(C[643]) );
  FA_381 \FA_INST_0[1].FA_INST_1[131].FA_  ( .A(A[643]), .B(B[643]), .CI(
        C[643]), .S(S[643]), .CO(C[644]) );
  FA_380 \FA_INST_0[1].FA_INST_1[132].FA_  ( .A(A[644]), .B(B[644]), .CI(
        C[644]), .S(S[644]), .CO(C[645]) );
  FA_379 \FA_INST_0[1].FA_INST_1[133].FA_  ( .A(A[645]), .B(B[645]), .CI(
        C[645]), .S(S[645]), .CO(C[646]) );
  FA_378 \FA_INST_0[1].FA_INST_1[134].FA_  ( .A(A[646]), .B(B[646]), .CI(
        C[646]), .S(S[646]), .CO(C[647]) );
  FA_377 \FA_INST_0[1].FA_INST_1[135].FA_  ( .A(A[647]), .B(B[647]), .CI(
        C[647]), .S(S[647]), .CO(C[648]) );
  FA_376 \FA_INST_0[1].FA_INST_1[136].FA_  ( .A(A[648]), .B(B[648]), .CI(
        C[648]), .S(S[648]), .CO(C[649]) );
  FA_375 \FA_INST_0[1].FA_INST_1[137].FA_  ( .A(A[649]), .B(B[649]), .CI(
        C[649]), .S(S[649]), .CO(C[650]) );
  FA_374 \FA_INST_0[1].FA_INST_1[138].FA_  ( .A(A[650]), .B(B[650]), .CI(
        C[650]), .S(S[650]), .CO(C[651]) );
  FA_373 \FA_INST_0[1].FA_INST_1[139].FA_  ( .A(A[651]), .B(B[651]), .CI(
        C[651]), .S(S[651]), .CO(C[652]) );
  FA_372 \FA_INST_0[1].FA_INST_1[140].FA_  ( .A(A[652]), .B(B[652]), .CI(
        C[652]), .S(S[652]), .CO(C[653]) );
  FA_371 \FA_INST_0[1].FA_INST_1[141].FA_  ( .A(A[653]), .B(B[653]), .CI(
        C[653]), .S(S[653]), .CO(C[654]) );
  FA_370 \FA_INST_0[1].FA_INST_1[142].FA_  ( .A(A[654]), .B(B[654]), .CI(
        C[654]), .S(S[654]), .CO(C[655]) );
  FA_369 \FA_INST_0[1].FA_INST_1[143].FA_  ( .A(A[655]), .B(B[655]), .CI(
        C[655]), .S(S[655]), .CO(C[656]) );
  FA_368 \FA_INST_0[1].FA_INST_1[144].FA_  ( .A(A[656]), .B(B[656]), .CI(
        C[656]), .S(S[656]), .CO(C[657]) );
  FA_367 \FA_INST_0[1].FA_INST_1[145].FA_  ( .A(A[657]), .B(B[657]), .CI(
        C[657]), .S(S[657]), .CO(C[658]) );
  FA_366 \FA_INST_0[1].FA_INST_1[146].FA_  ( .A(A[658]), .B(B[658]), .CI(
        C[658]), .S(S[658]), .CO(C[659]) );
  FA_365 \FA_INST_0[1].FA_INST_1[147].FA_  ( .A(A[659]), .B(B[659]), .CI(
        C[659]), .S(S[659]), .CO(C[660]) );
  FA_364 \FA_INST_0[1].FA_INST_1[148].FA_  ( .A(A[660]), .B(B[660]), .CI(
        C[660]), .S(S[660]), .CO(C[661]) );
  FA_363 \FA_INST_0[1].FA_INST_1[149].FA_  ( .A(A[661]), .B(B[661]), .CI(
        C[661]), .S(S[661]), .CO(C[662]) );
  FA_362 \FA_INST_0[1].FA_INST_1[150].FA_  ( .A(A[662]), .B(B[662]), .CI(
        C[662]), .S(S[662]), .CO(C[663]) );
  FA_361 \FA_INST_0[1].FA_INST_1[151].FA_  ( .A(A[663]), .B(B[663]), .CI(
        C[663]), .S(S[663]), .CO(C[664]) );
  FA_360 \FA_INST_0[1].FA_INST_1[152].FA_  ( .A(A[664]), .B(B[664]), .CI(
        C[664]), .S(S[664]), .CO(C[665]) );
  FA_359 \FA_INST_0[1].FA_INST_1[153].FA_  ( .A(A[665]), .B(B[665]), .CI(
        C[665]), .S(S[665]), .CO(C[666]) );
  FA_358 \FA_INST_0[1].FA_INST_1[154].FA_  ( .A(A[666]), .B(B[666]), .CI(
        C[666]), .S(S[666]), .CO(C[667]) );
  FA_357 \FA_INST_0[1].FA_INST_1[155].FA_  ( .A(A[667]), .B(B[667]), .CI(
        C[667]), .S(S[667]), .CO(C[668]) );
  FA_356 \FA_INST_0[1].FA_INST_1[156].FA_  ( .A(A[668]), .B(B[668]), .CI(
        C[668]), .S(S[668]), .CO(C[669]) );
  FA_355 \FA_INST_0[1].FA_INST_1[157].FA_  ( .A(A[669]), .B(B[669]), .CI(
        C[669]), .S(S[669]), .CO(C[670]) );
  FA_354 \FA_INST_0[1].FA_INST_1[158].FA_  ( .A(A[670]), .B(B[670]), .CI(
        C[670]), .S(S[670]), .CO(C[671]) );
  FA_353 \FA_INST_0[1].FA_INST_1[159].FA_  ( .A(A[671]), .B(B[671]), .CI(
        C[671]), .S(S[671]), .CO(C[672]) );
  FA_352 \FA_INST_0[1].FA_INST_1[160].FA_  ( .A(A[672]), .B(B[672]), .CI(
        C[672]), .S(S[672]), .CO(C[673]) );
  FA_351 \FA_INST_0[1].FA_INST_1[161].FA_  ( .A(A[673]), .B(B[673]), .CI(
        C[673]), .S(S[673]), .CO(C[674]) );
  FA_350 \FA_INST_0[1].FA_INST_1[162].FA_  ( .A(A[674]), .B(B[674]), .CI(
        C[674]), .S(S[674]), .CO(C[675]) );
  FA_349 \FA_INST_0[1].FA_INST_1[163].FA_  ( .A(A[675]), .B(B[675]), .CI(
        C[675]), .S(S[675]), .CO(C[676]) );
  FA_348 \FA_INST_0[1].FA_INST_1[164].FA_  ( .A(A[676]), .B(B[676]), .CI(
        C[676]), .S(S[676]), .CO(C[677]) );
  FA_347 \FA_INST_0[1].FA_INST_1[165].FA_  ( .A(A[677]), .B(B[677]), .CI(
        C[677]), .S(S[677]), .CO(C[678]) );
  FA_346 \FA_INST_0[1].FA_INST_1[166].FA_  ( .A(A[678]), .B(B[678]), .CI(
        C[678]), .S(S[678]), .CO(C[679]) );
  FA_345 \FA_INST_0[1].FA_INST_1[167].FA_  ( .A(A[679]), .B(B[679]), .CI(
        C[679]), .S(S[679]), .CO(C[680]) );
  FA_344 \FA_INST_0[1].FA_INST_1[168].FA_  ( .A(A[680]), .B(B[680]), .CI(
        C[680]), .S(S[680]), .CO(C[681]) );
  FA_343 \FA_INST_0[1].FA_INST_1[169].FA_  ( .A(A[681]), .B(B[681]), .CI(
        C[681]), .S(S[681]), .CO(C[682]) );
  FA_342 \FA_INST_0[1].FA_INST_1[170].FA_  ( .A(A[682]), .B(B[682]), .CI(
        C[682]), .S(S[682]), .CO(C[683]) );
  FA_341 \FA_INST_0[1].FA_INST_1[171].FA_  ( .A(A[683]), .B(B[683]), .CI(
        C[683]), .S(S[683]), .CO(C[684]) );
  FA_340 \FA_INST_0[1].FA_INST_1[172].FA_  ( .A(A[684]), .B(B[684]), .CI(
        C[684]), .S(S[684]), .CO(C[685]) );
  FA_339 \FA_INST_0[1].FA_INST_1[173].FA_  ( .A(A[685]), .B(B[685]), .CI(
        C[685]), .S(S[685]), .CO(C[686]) );
  FA_338 \FA_INST_0[1].FA_INST_1[174].FA_  ( .A(A[686]), .B(B[686]), .CI(
        C[686]), .S(S[686]), .CO(C[687]) );
  FA_337 \FA_INST_0[1].FA_INST_1[175].FA_  ( .A(A[687]), .B(B[687]), .CI(
        C[687]), .S(S[687]), .CO(C[688]) );
  FA_336 \FA_INST_0[1].FA_INST_1[176].FA_  ( .A(A[688]), .B(B[688]), .CI(
        C[688]), .S(S[688]), .CO(C[689]) );
  FA_335 \FA_INST_0[1].FA_INST_1[177].FA_  ( .A(A[689]), .B(B[689]), .CI(
        C[689]), .S(S[689]), .CO(C[690]) );
  FA_334 \FA_INST_0[1].FA_INST_1[178].FA_  ( .A(A[690]), .B(B[690]), .CI(
        C[690]), .S(S[690]), .CO(C[691]) );
  FA_333 \FA_INST_0[1].FA_INST_1[179].FA_  ( .A(A[691]), .B(B[691]), .CI(
        C[691]), .S(S[691]), .CO(C[692]) );
  FA_332 \FA_INST_0[1].FA_INST_1[180].FA_  ( .A(A[692]), .B(B[692]), .CI(
        C[692]), .S(S[692]), .CO(C[693]) );
  FA_331 \FA_INST_0[1].FA_INST_1[181].FA_  ( .A(A[693]), .B(B[693]), .CI(
        C[693]), .S(S[693]), .CO(C[694]) );
  FA_330 \FA_INST_0[1].FA_INST_1[182].FA_  ( .A(A[694]), .B(B[694]), .CI(
        C[694]), .S(S[694]), .CO(C[695]) );
  FA_329 \FA_INST_0[1].FA_INST_1[183].FA_  ( .A(A[695]), .B(B[695]), .CI(
        C[695]), .S(S[695]), .CO(C[696]) );
  FA_328 \FA_INST_0[1].FA_INST_1[184].FA_  ( .A(A[696]), .B(B[696]), .CI(
        C[696]), .S(S[696]), .CO(C[697]) );
  FA_327 \FA_INST_0[1].FA_INST_1[185].FA_  ( .A(A[697]), .B(B[697]), .CI(
        C[697]), .S(S[697]), .CO(C[698]) );
  FA_326 \FA_INST_0[1].FA_INST_1[186].FA_  ( .A(A[698]), .B(B[698]), .CI(
        C[698]), .S(S[698]), .CO(C[699]) );
  FA_325 \FA_INST_0[1].FA_INST_1[187].FA_  ( .A(A[699]), .B(B[699]), .CI(
        C[699]), .S(S[699]), .CO(C[700]) );
  FA_324 \FA_INST_0[1].FA_INST_1[188].FA_  ( .A(A[700]), .B(B[700]), .CI(
        C[700]), .S(S[700]), .CO(C[701]) );
  FA_323 \FA_INST_0[1].FA_INST_1[189].FA_  ( .A(A[701]), .B(B[701]), .CI(
        C[701]), .S(S[701]), .CO(C[702]) );
  FA_322 \FA_INST_0[1].FA_INST_1[190].FA_  ( .A(A[702]), .B(B[702]), .CI(
        C[702]), .S(S[702]), .CO(C[703]) );
  FA_321 \FA_INST_0[1].FA_INST_1[191].FA_  ( .A(A[703]), .B(B[703]), .CI(
        C[703]), .S(S[703]), .CO(C[704]) );
  FA_320 \FA_INST_0[1].FA_INST_1[192].FA_  ( .A(A[704]), .B(B[704]), .CI(
        C[704]), .S(S[704]), .CO(C[705]) );
  FA_319 \FA_INST_0[1].FA_INST_1[193].FA_  ( .A(A[705]), .B(B[705]), .CI(
        C[705]), .S(S[705]), .CO(C[706]) );
  FA_318 \FA_INST_0[1].FA_INST_1[194].FA_  ( .A(A[706]), .B(B[706]), .CI(
        C[706]), .S(S[706]), .CO(C[707]) );
  FA_317 \FA_INST_0[1].FA_INST_1[195].FA_  ( .A(A[707]), .B(B[707]), .CI(
        C[707]), .S(S[707]), .CO(C[708]) );
  FA_316 \FA_INST_0[1].FA_INST_1[196].FA_  ( .A(A[708]), .B(B[708]), .CI(
        C[708]), .S(S[708]), .CO(C[709]) );
  FA_315 \FA_INST_0[1].FA_INST_1[197].FA_  ( .A(A[709]), .B(B[709]), .CI(
        C[709]), .S(S[709]), .CO(C[710]) );
  FA_314 \FA_INST_0[1].FA_INST_1[198].FA_  ( .A(A[710]), .B(B[710]), .CI(
        C[710]), .S(S[710]), .CO(C[711]) );
  FA_313 \FA_INST_0[1].FA_INST_1[199].FA_  ( .A(A[711]), .B(B[711]), .CI(
        C[711]), .S(S[711]), .CO(C[712]) );
  FA_312 \FA_INST_0[1].FA_INST_1[200].FA_  ( .A(A[712]), .B(B[712]), .CI(
        C[712]), .S(S[712]), .CO(C[713]) );
  FA_311 \FA_INST_0[1].FA_INST_1[201].FA_  ( .A(A[713]), .B(B[713]), .CI(
        C[713]), .S(S[713]), .CO(C[714]) );
  FA_310 \FA_INST_0[1].FA_INST_1[202].FA_  ( .A(A[714]), .B(B[714]), .CI(
        C[714]), .S(S[714]), .CO(C[715]) );
  FA_309 \FA_INST_0[1].FA_INST_1[203].FA_  ( .A(A[715]), .B(B[715]), .CI(
        C[715]), .S(S[715]), .CO(C[716]) );
  FA_308 \FA_INST_0[1].FA_INST_1[204].FA_  ( .A(A[716]), .B(B[716]), .CI(
        C[716]), .S(S[716]), .CO(C[717]) );
  FA_307 \FA_INST_0[1].FA_INST_1[205].FA_  ( .A(A[717]), .B(B[717]), .CI(
        C[717]), .S(S[717]), .CO(C[718]) );
  FA_306 \FA_INST_0[1].FA_INST_1[206].FA_  ( .A(A[718]), .B(B[718]), .CI(
        C[718]), .S(S[718]), .CO(C[719]) );
  FA_305 \FA_INST_0[1].FA_INST_1[207].FA_  ( .A(A[719]), .B(B[719]), .CI(
        C[719]), .S(S[719]), .CO(C[720]) );
  FA_304 \FA_INST_0[1].FA_INST_1[208].FA_  ( .A(A[720]), .B(B[720]), .CI(
        C[720]), .S(S[720]), .CO(C[721]) );
  FA_303 \FA_INST_0[1].FA_INST_1[209].FA_  ( .A(A[721]), .B(B[721]), .CI(
        C[721]), .S(S[721]), .CO(C[722]) );
  FA_302 \FA_INST_0[1].FA_INST_1[210].FA_  ( .A(A[722]), .B(B[722]), .CI(
        C[722]), .S(S[722]), .CO(C[723]) );
  FA_301 \FA_INST_0[1].FA_INST_1[211].FA_  ( .A(A[723]), .B(B[723]), .CI(
        C[723]), .S(S[723]), .CO(C[724]) );
  FA_300 \FA_INST_0[1].FA_INST_1[212].FA_  ( .A(A[724]), .B(B[724]), .CI(
        C[724]), .S(S[724]), .CO(C[725]) );
  FA_299 \FA_INST_0[1].FA_INST_1[213].FA_  ( .A(A[725]), .B(B[725]), .CI(
        C[725]), .S(S[725]), .CO(C[726]) );
  FA_298 \FA_INST_0[1].FA_INST_1[214].FA_  ( .A(A[726]), .B(B[726]), .CI(
        C[726]), .S(S[726]), .CO(C[727]) );
  FA_297 \FA_INST_0[1].FA_INST_1[215].FA_  ( .A(A[727]), .B(B[727]), .CI(
        C[727]), .S(S[727]), .CO(C[728]) );
  FA_296 \FA_INST_0[1].FA_INST_1[216].FA_  ( .A(A[728]), .B(B[728]), .CI(
        C[728]), .S(S[728]), .CO(C[729]) );
  FA_295 \FA_INST_0[1].FA_INST_1[217].FA_  ( .A(A[729]), .B(B[729]), .CI(
        C[729]), .S(S[729]), .CO(C[730]) );
  FA_294 \FA_INST_0[1].FA_INST_1[218].FA_  ( .A(A[730]), .B(B[730]), .CI(
        C[730]), .S(S[730]), .CO(C[731]) );
  FA_293 \FA_INST_0[1].FA_INST_1[219].FA_  ( .A(A[731]), .B(B[731]), .CI(
        C[731]), .S(S[731]), .CO(C[732]) );
  FA_292 \FA_INST_0[1].FA_INST_1[220].FA_  ( .A(A[732]), .B(B[732]), .CI(
        C[732]), .S(S[732]), .CO(C[733]) );
  FA_291 \FA_INST_0[1].FA_INST_1[221].FA_  ( .A(A[733]), .B(B[733]), .CI(
        C[733]), .S(S[733]), .CO(C[734]) );
  FA_290 \FA_INST_0[1].FA_INST_1[222].FA_  ( .A(A[734]), .B(B[734]), .CI(
        C[734]), .S(S[734]), .CO(C[735]) );
  FA_289 \FA_INST_0[1].FA_INST_1[223].FA_  ( .A(A[735]), .B(B[735]), .CI(
        C[735]), .S(S[735]), .CO(C[736]) );
  FA_288 \FA_INST_0[1].FA_INST_1[224].FA_  ( .A(A[736]), .B(B[736]), .CI(
        C[736]), .S(S[736]), .CO(C[737]) );
  FA_287 \FA_INST_0[1].FA_INST_1[225].FA_  ( .A(A[737]), .B(B[737]), .CI(
        C[737]), .S(S[737]), .CO(C[738]) );
  FA_286 \FA_INST_0[1].FA_INST_1[226].FA_  ( .A(A[738]), .B(B[738]), .CI(
        C[738]), .S(S[738]), .CO(C[739]) );
  FA_285 \FA_INST_0[1].FA_INST_1[227].FA_  ( .A(A[739]), .B(B[739]), .CI(
        C[739]), .S(S[739]), .CO(C[740]) );
  FA_284 \FA_INST_0[1].FA_INST_1[228].FA_  ( .A(A[740]), .B(B[740]), .CI(
        C[740]), .S(S[740]), .CO(C[741]) );
  FA_283 \FA_INST_0[1].FA_INST_1[229].FA_  ( .A(A[741]), .B(B[741]), .CI(
        C[741]), .S(S[741]), .CO(C[742]) );
  FA_282 \FA_INST_0[1].FA_INST_1[230].FA_  ( .A(A[742]), .B(B[742]), .CI(
        C[742]), .S(S[742]), .CO(C[743]) );
  FA_281 \FA_INST_0[1].FA_INST_1[231].FA_  ( .A(A[743]), .B(B[743]), .CI(
        C[743]), .S(S[743]), .CO(C[744]) );
  FA_280 \FA_INST_0[1].FA_INST_1[232].FA_  ( .A(A[744]), .B(B[744]), .CI(
        C[744]), .S(S[744]), .CO(C[745]) );
  FA_279 \FA_INST_0[1].FA_INST_1[233].FA_  ( .A(A[745]), .B(B[745]), .CI(
        C[745]), .S(S[745]), .CO(C[746]) );
  FA_278 \FA_INST_0[1].FA_INST_1[234].FA_  ( .A(A[746]), .B(B[746]), .CI(
        C[746]), .S(S[746]), .CO(C[747]) );
  FA_277 \FA_INST_0[1].FA_INST_1[235].FA_  ( .A(A[747]), .B(B[747]), .CI(
        C[747]), .S(S[747]), .CO(C[748]) );
  FA_276 \FA_INST_0[1].FA_INST_1[236].FA_  ( .A(A[748]), .B(B[748]), .CI(
        C[748]), .S(S[748]), .CO(C[749]) );
  FA_275 \FA_INST_0[1].FA_INST_1[237].FA_  ( .A(A[749]), .B(B[749]), .CI(
        C[749]), .S(S[749]), .CO(C[750]) );
  FA_274 \FA_INST_0[1].FA_INST_1[238].FA_  ( .A(A[750]), .B(B[750]), .CI(
        C[750]), .S(S[750]), .CO(C[751]) );
  FA_273 \FA_INST_0[1].FA_INST_1[239].FA_  ( .A(A[751]), .B(B[751]), .CI(
        C[751]), .S(S[751]), .CO(C[752]) );
  FA_272 \FA_INST_0[1].FA_INST_1[240].FA_  ( .A(A[752]), .B(B[752]), .CI(
        C[752]), .S(S[752]), .CO(C[753]) );
  FA_271 \FA_INST_0[1].FA_INST_1[241].FA_  ( .A(A[753]), .B(B[753]), .CI(
        C[753]), .S(S[753]), .CO(C[754]) );
  FA_270 \FA_INST_0[1].FA_INST_1[242].FA_  ( .A(A[754]), .B(B[754]), .CI(
        C[754]), .S(S[754]), .CO(C[755]) );
  FA_269 \FA_INST_0[1].FA_INST_1[243].FA_  ( .A(A[755]), .B(B[755]), .CI(
        C[755]), .S(S[755]), .CO(C[756]) );
  FA_268 \FA_INST_0[1].FA_INST_1[244].FA_  ( .A(A[756]), .B(B[756]), .CI(
        C[756]), .S(S[756]), .CO(C[757]) );
  FA_267 \FA_INST_0[1].FA_INST_1[245].FA_  ( .A(A[757]), .B(B[757]), .CI(
        C[757]), .S(S[757]), .CO(C[758]) );
  FA_266 \FA_INST_0[1].FA_INST_1[246].FA_  ( .A(A[758]), .B(B[758]), .CI(
        C[758]), .S(S[758]), .CO(C[759]) );
  FA_265 \FA_INST_0[1].FA_INST_1[247].FA_  ( .A(A[759]), .B(B[759]), .CI(
        C[759]), .S(S[759]), .CO(C[760]) );
  FA_264 \FA_INST_0[1].FA_INST_1[248].FA_  ( .A(A[760]), .B(B[760]), .CI(
        C[760]), .S(S[760]), .CO(C[761]) );
  FA_263 \FA_INST_0[1].FA_INST_1[249].FA_  ( .A(A[761]), .B(B[761]), .CI(
        C[761]), .S(S[761]), .CO(C[762]) );
  FA_262 \FA_INST_0[1].FA_INST_1[250].FA_  ( .A(A[762]), .B(B[762]), .CI(
        C[762]), .S(S[762]), .CO(C[763]) );
  FA_261 \FA_INST_0[1].FA_INST_1[251].FA_  ( .A(A[763]), .B(B[763]), .CI(
        C[763]), .S(S[763]), .CO(C[764]) );
  FA_260 \FA_INST_0[1].FA_INST_1[252].FA_  ( .A(A[764]), .B(B[764]), .CI(
        C[764]), .S(S[764]), .CO(C[765]) );
  FA_259 \FA_INST_0[1].FA_INST_1[253].FA_  ( .A(A[765]), .B(B[765]), .CI(
        C[765]), .S(S[765]), .CO(C[766]) );
  FA_258 \FA_INST_0[1].FA_INST_1[254].FA_  ( .A(A[766]), .B(B[766]), .CI(
        C[766]), .S(S[766]), .CO(C[767]) );
  FA_257 \FA_INST_0[1].FA_INST_1[255].FA_  ( .A(A[767]), .B(B[767]), .CI(
        C[767]), .S(S[767]), .CO(C[768]) );
  FA_256 \FA_INST_0[1].FA_INST_1[256].FA_  ( .A(A[768]), .B(B[768]), .CI(
        C[768]), .S(S[768]), .CO(C[769]) );
  FA_255 \FA_INST_0[1].FA_INST_1[257].FA_  ( .A(A[769]), .B(B[769]), .CI(
        C[769]), .S(S[769]), .CO(C[770]) );
  FA_254 \FA_INST_0[1].FA_INST_1[258].FA_  ( .A(A[770]), .B(B[770]), .CI(
        C[770]), .S(S[770]), .CO(C[771]) );
  FA_253 \FA_INST_0[1].FA_INST_1[259].FA_  ( .A(A[771]), .B(B[771]), .CI(
        C[771]), .S(S[771]), .CO(C[772]) );
  FA_252 \FA_INST_0[1].FA_INST_1[260].FA_  ( .A(A[772]), .B(B[772]), .CI(
        C[772]), .S(S[772]), .CO(C[773]) );
  FA_251 \FA_INST_0[1].FA_INST_1[261].FA_  ( .A(A[773]), .B(B[773]), .CI(
        C[773]), .S(S[773]), .CO(C[774]) );
  FA_250 \FA_INST_0[1].FA_INST_1[262].FA_  ( .A(A[774]), .B(B[774]), .CI(
        C[774]), .S(S[774]), .CO(C[775]) );
  FA_249 \FA_INST_0[1].FA_INST_1[263].FA_  ( .A(A[775]), .B(B[775]), .CI(
        C[775]), .S(S[775]), .CO(C[776]) );
  FA_248 \FA_INST_0[1].FA_INST_1[264].FA_  ( .A(A[776]), .B(B[776]), .CI(
        C[776]), .S(S[776]), .CO(C[777]) );
  FA_247 \FA_INST_0[1].FA_INST_1[265].FA_  ( .A(A[777]), .B(B[777]), .CI(
        C[777]), .S(S[777]), .CO(C[778]) );
  FA_246 \FA_INST_0[1].FA_INST_1[266].FA_  ( .A(A[778]), .B(B[778]), .CI(
        C[778]), .S(S[778]), .CO(C[779]) );
  FA_245 \FA_INST_0[1].FA_INST_1[267].FA_  ( .A(A[779]), .B(B[779]), .CI(
        C[779]), .S(S[779]), .CO(C[780]) );
  FA_244 \FA_INST_0[1].FA_INST_1[268].FA_  ( .A(A[780]), .B(B[780]), .CI(
        C[780]), .S(S[780]), .CO(C[781]) );
  FA_243 \FA_INST_0[1].FA_INST_1[269].FA_  ( .A(A[781]), .B(B[781]), .CI(
        C[781]), .S(S[781]), .CO(C[782]) );
  FA_242 \FA_INST_0[1].FA_INST_1[270].FA_  ( .A(A[782]), .B(B[782]), .CI(
        C[782]), .S(S[782]), .CO(C[783]) );
  FA_241 \FA_INST_0[1].FA_INST_1[271].FA_  ( .A(A[783]), .B(B[783]), .CI(
        C[783]), .S(S[783]), .CO(C[784]) );
  FA_240 \FA_INST_0[1].FA_INST_1[272].FA_  ( .A(A[784]), .B(B[784]), .CI(
        C[784]), .S(S[784]), .CO(C[785]) );
  FA_239 \FA_INST_0[1].FA_INST_1[273].FA_  ( .A(A[785]), .B(B[785]), .CI(
        C[785]), .S(S[785]), .CO(C[786]) );
  FA_238 \FA_INST_0[1].FA_INST_1[274].FA_  ( .A(A[786]), .B(B[786]), .CI(
        C[786]), .S(S[786]), .CO(C[787]) );
  FA_237 \FA_INST_0[1].FA_INST_1[275].FA_  ( .A(A[787]), .B(B[787]), .CI(
        C[787]), .S(S[787]), .CO(C[788]) );
  FA_236 \FA_INST_0[1].FA_INST_1[276].FA_  ( .A(A[788]), .B(B[788]), .CI(
        C[788]), .S(S[788]), .CO(C[789]) );
  FA_235 \FA_INST_0[1].FA_INST_1[277].FA_  ( .A(A[789]), .B(B[789]), .CI(
        C[789]), .S(S[789]), .CO(C[790]) );
  FA_234 \FA_INST_0[1].FA_INST_1[278].FA_  ( .A(A[790]), .B(B[790]), .CI(
        C[790]), .S(S[790]), .CO(C[791]) );
  FA_233 \FA_INST_0[1].FA_INST_1[279].FA_  ( .A(A[791]), .B(B[791]), .CI(
        C[791]), .S(S[791]), .CO(C[792]) );
  FA_232 \FA_INST_0[1].FA_INST_1[280].FA_  ( .A(A[792]), .B(B[792]), .CI(
        C[792]), .S(S[792]), .CO(C[793]) );
  FA_231 \FA_INST_0[1].FA_INST_1[281].FA_  ( .A(A[793]), .B(B[793]), .CI(
        C[793]), .S(S[793]), .CO(C[794]) );
  FA_230 \FA_INST_0[1].FA_INST_1[282].FA_  ( .A(A[794]), .B(B[794]), .CI(
        C[794]), .S(S[794]), .CO(C[795]) );
  FA_229 \FA_INST_0[1].FA_INST_1[283].FA_  ( .A(A[795]), .B(B[795]), .CI(
        C[795]), .S(S[795]), .CO(C[796]) );
  FA_228 \FA_INST_0[1].FA_INST_1[284].FA_  ( .A(A[796]), .B(B[796]), .CI(
        C[796]), .S(S[796]), .CO(C[797]) );
  FA_227 \FA_INST_0[1].FA_INST_1[285].FA_  ( .A(A[797]), .B(B[797]), .CI(
        C[797]), .S(S[797]), .CO(C[798]) );
  FA_226 \FA_INST_0[1].FA_INST_1[286].FA_  ( .A(A[798]), .B(B[798]), .CI(
        C[798]), .S(S[798]), .CO(C[799]) );
  FA_225 \FA_INST_0[1].FA_INST_1[287].FA_  ( .A(A[799]), .B(B[799]), .CI(
        C[799]), .S(S[799]), .CO(C[800]) );
  FA_224 \FA_INST_0[1].FA_INST_1[288].FA_  ( .A(A[800]), .B(B[800]), .CI(
        C[800]), .S(S[800]), .CO(C[801]) );
  FA_223 \FA_INST_0[1].FA_INST_1[289].FA_  ( .A(A[801]), .B(B[801]), .CI(
        C[801]), .S(S[801]), .CO(C[802]) );
  FA_222 \FA_INST_0[1].FA_INST_1[290].FA_  ( .A(A[802]), .B(B[802]), .CI(
        C[802]), .S(S[802]), .CO(C[803]) );
  FA_221 \FA_INST_0[1].FA_INST_1[291].FA_  ( .A(A[803]), .B(B[803]), .CI(
        C[803]), .S(S[803]), .CO(C[804]) );
  FA_220 \FA_INST_0[1].FA_INST_1[292].FA_  ( .A(A[804]), .B(B[804]), .CI(
        C[804]), .S(S[804]), .CO(C[805]) );
  FA_219 \FA_INST_0[1].FA_INST_1[293].FA_  ( .A(A[805]), .B(B[805]), .CI(
        C[805]), .S(S[805]), .CO(C[806]) );
  FA_218 \FA_INST_0[1].FA_INST_1[294].FA_  ( .A(A[806]), .B(B[806]), .CI(
        C[806]), .S(S[806]), .CO(C[807]) );
  FA_217 \FA_INST_0[1].FA_INST_1[295].FA_  ( .A(A[807]), .B(B[807]), .CI(
        C[807]), .S(S[807]), .CO(C[808]) );
  FA_216 \FA_INST_0[1].FA_INST_1[296].FA_  ( .A(A[808]), .B(B[808]), .CI(
        C[808]), .S(S[808]), .CO(C[809]) );
  FA_215 \FA_INST_0[1].FA_INST_1[297].FA_  ( .A(A[809]), .B(B[809]), .CI(
        C[809]), .S(S[809]), .CO(C[810]) );
  FA_214 \FA_INST_0[1].FA_INST_1[298].FA_  ( .A(A[810]), .B(B[810]), .CI(
        C[810]), .S(S[810]), .CO(C[811]) );
  FA_213 \FA_INST_0[1].FA_INST_1[299].FA_  ( .A(A[811]), .B(B[811]), .CI(
        C[811]), .S(S[811]), .CO(C[812]) );
  FA_212 \FA_INST_0[1].FA_INST_1[300].FA_  ( .A(A[812]), .B(B[812]), .CI(
        C[812]), .S(S[812]), .CO(C[813]) );
  FA_211 \FA_INST_0[1].FA_INST_1[301].FA_  ( .A(A[813]), .B(B[813]), .CI(
        C[813]), .S(S[813]), .CO(C[814]) );
  FA_210 \FA_INST_0[1].FA_INST_1[302].FA_  ( .A(A[814]), .B(B[814]), .CI(
        C[814]), .S(S[814]), .CO(C[815]) );
  FA_209 \FA_INST_0[1].FA_INST_1[303].FA_  ( .A(A[815]), .B(B[815]), .CI(
        C[815]), .S(S[815]), .CO(C[816]) );
  FA_208 \FA_INST_0[1].FA_INST_1[304].FA_  ( .A(A[816]), .B(B[816]), .CI(
        C[816]), .S(S[816]), .CO(C[817]) );
  FA_207 \FA_INST_0[1].FA_INST_1[305].FA_  ( .A(A[817]), .B(B[817]), .CI(
        C[817]), .S(S[817]), .CO(C[818]) );
  FA_206 \FA_INST_0[1].FA_INST_1[306].FA_  ( .A(A[818]), .B(B[818]), .CI(
        C[818]), .S(S[818]), .CO(C[819]) );
  FA_205 \FA_INST_0[1].FA_INST_1[307].FA_  ( .A(A[819]), .B(B[819]), .CI(
        C[819]), .S(S[819]), .CO(C[820]) );
  FA_204 \FA_INST_0[1].FA_INST_1[308].FA_  ( .A(A[820]), .B(B[820]), .CI(
        C[820]), .S(S[820]), .CO(C[821]) );
  FA_203 \FA_INST_0[1].FA_INST_1[309].FA_  ( .A(A[821]), .B(B[821]), .CI(
        C[821]), .S(S[821]), .CO(C[822]) );
  FA_202 \FA_INST_0[1].FA_INST_1[310].FA_  ( .A(A[822]), .B(B[822]), .CI(
        C[822]), .S(S[822]), .CO(C[823]) );
  FA_201 \FA_INST_0[1].FA_INST_1[311].FA_  ( .A(A[823]), .B(B[823]), .CI(
        C[823]), .S(S[823]), .CO(C[824]) );
  FA_200 \FA_INST_0[1].FA_INST_1[312].FA_  ( .A(A[824]), .B(B[824]), .CI(
        C[824]), .S(S[824]), .CO(C[825]) );
  FA_199 \FA_INST_0[1].FA_INST_1[313].FA_  ( .A(A[825]), .B(B[825]), .CI(
        C[825]), .S(S[825]), .CO(C[826]) );
  FA_198 \FA_INST_0[1].FA_INST_1[314].FA_  ( .A(A[826]), .B(B[826]), .CI(
        C[826]), .S(S[826]), .CO(C[827]) );
  FA_197 \FA_INST_0[1].FA_INST_1[315].FA_  ( .A(A[827]), .B(B[827]), .CI(
        C[827]), .S(S[827]), .CO(C[828]) );
  FA_196 \FA_INST_0[1].FA_INST_1[316].FA_  ( .A(A[828]), .B(B[828]), .CI(
        C[828]), .S(S[828]), .CO(C[829]) );
  FA_195 \FA_INST_0[1].FA_INST_1[317].FA_  ( .A(A[829]), .B(B[829]), .CI(
        C[829]), .S(S[829]), .CO(C[830]) );
  FA_194 \FA_INST_0[1].FA_INST_1[318].FA_  ( .A(A[830]), .B(B[830]), .CI(
        C[830]), .S(S[830]), .CO(C[831]) );
  FA_193 \FA_INST_0[1].FA_INST_1[319].FA_  ( .A(A[831]), .B(B[831]), .CI(
        C[831]), .S(S[831]), .CO(C[832]) );
  FA_192 \FA_INST_0[1].FA_INST_1[320].FA_  ( .A(A[832]), .B(B[832]), .CI(
        C[832]), .S(S[832]), .CO(C[833]) );
  FA_191 \FA_INST_0[1].FA_INST_1[321].FA_  ( .A(A[833]), .B(B[833]), .CI(
        C[833]), .S(S[833]), .CO(C[834]) );
  FA_190 \FA_INST_0[1].FA_INST_1[322].FA_  ( .A(A[834]), .B(B[834]), .CI(
        C[834]), .S(S[834]), .CO(C[835]) );
  FA_189 \FA_INST_0[1].FA_INST_1[323].FA_  ( .A(A[835]), .B(B[835]), .CI(
        C[835]), .S(S[835]), .CO(C[836]) );
  FA_188 \FA_INST_0[1].FA_INST_1[324].FA_  ( .A(A[836]), .B(B[836]), .CI(
        C[836]), .S(S[836]), .CO(C[837]) );
  FA_187 \FA_INST_0[1].FA_INST_1[325].FA_  ( .A(A[837]), .B(B[837]), .CI(
        C[837]), .S(S[837]), .CO(C[838]) );
  FA_186 \FA_INST_0[1].FA_INST_1[326].FA_  ( .A(A[838]), .B(B[838]), .CI(
        C[838]), .S(S[838]), .CO(C[839]) );
  FA_185 \FA_INST_0[1].FA_INST_1[327].FA_  ( .A(A[839]), .B(B[839]), .CI(
        C[839]), .S(S[839]), .CO(C[840]) );
  FA_184 \FA_INST_0[1].FA_INST_1[328].FA_  ( .A(A[840]), .B(B[840]), .CI(
        C[840]), .S(S[840]), .CO(C[841]) );
  FA_183 \FA_INST_0[1].FA_INST_1[329].FA_  ( .A(A[841]), .B(B[841]), .CI(
        C[841]), .S(S[841]), .CO(C[842]) );
  FA_182 \FA_INST_0[1].FA_INST_1[330].FA_  ( .A(A[842]), .B(B[842]), .CI(
        C[842]), .S(S[842]), .CO(C[843]) );
  FA_181 \FA_INST_0[1].FA_INST_1[331].FA_  ( .A(A[843]), .B(B[843]), .CI(
        C[843]), .S(S[843]), .CO(C[844]) );
  FA_180 \FA_INST_0[1].FA_INST_1[332].FA_  ( .A(A[844]), .B(B[844]), .CI(
        C[844]), .S(S[844]), .CO(C[845]) );
  FA_179 \FA_INST_0[1].FA_INST_1[333].FA_  ( .A(A[845]), .B(B[845]), .CI(
        C[845]), .S(S[845]), .CO(C[846]) );
  FA_178 \FA_INST_0[1].FA_INST_1[334].FA_  ( .A(A[846]), .B(B[846]), .CI(
        C[846]), .S(S[846]), .CO(C[847]) );
  FA_177 \FA_INST_0[1].FA_INST_1[335].FA_  ( .A(A[847]), .B(B[847]), .CI(
        C[847]), .S(S[847]), .CO(C[848]) );
  FA_176 \FA_INST_0[1].FA_INST_1[336].FA_  ( .A(A[848]), .B(B[848]), .CI(
        C[848]), .S(S[848]), .CO(C[849]) );
  FA_175 \FA_INST_0[1].FA_INST_1[337].FA_  ( .A(A[849]), .B(B[849]), .CI(
        C[849]), .S(S[849]), .CO(C[850]) );
  FA_174 \FA_INST_0[1].FA_INST_1[338].FA_  ( .A(A[850]), .B(B[850]), .CI(
        C[850]), .S(S[850]), .CO(C[851]) );
  FA_173 \FA_INST_0[1].FA_INST_1[339].FA_  ( .A(A[851]), .B(B[851]), .CI(
        C[851]), .S(S[851]), .CO(C[852]) );
  FA_172 \FA_INST_0[1].FA_INST_1[340].FA_  ( .A(A[852]), .B(B[852]), .CI(
        C[852]), .S(S[852]), .CO(C[853]) );
  FA_171 \FA_INST_0[1].FA_INST_1[341].FA_  ( .A(A[853]), .B(B[853]), .CI(
        C[853]), .S(S[853]), .CO(C[854]) );
  FA_170 \FA_INST_0[1].FA_INST_1[342].FA_  ( .A(A[854]), .B(B[854]), .CI(
        C[854]), .S(S[854]), .CO(C[855]) );
  FA_169 \FA_INST_0[1].FA_INST_1[343].FA_  ( .A(A[855]), .B(B[855]), .CI(
        C[855]), .S(S[855]), .CO(C[856]) );
  FA_168 \FA_INST_0[1].FA_INST_1[344].FA_  ( .A(A[856]), .B(B[856]), .CI(
        C[856]), .S(S[856]), .CO(C[857]) );
  FA_167 \FA_INST_0[1].FA_INST_1[345].FA_  ( .A(A[857]), .B(B[857]), .CI(
        C[857]), .S(S[857]), .CO(C[858]) );
  FA_166 \FA_INST_0[1].FA_INST_1[346].FA_  ( .A(A[858]), .B(B[858]), .CI(
        C[858]), .S(S[858]), .CO(C[859]) );
  FA_165 \FA_INST_0[1].FA_INST_1[347].FA_  ( .A(A[859]), .B(B[859]), .CI(
        C[859]), .S(S[859]), .CO(C[860]) );
  FA_164 \FA_INST_0[1].FA_INST_1[348].FA_  ( .A(A[860]), .B(B[860]), .CI(
        C[860]), .S(S[860]), .CO(C[861]) );
  FA_163 \FA_INST_0[1].FA_INST_1[349].FA_  ( .A(A[861]), .B(B[861]), .CI(
        C[861]), .S(S[861]), .CO(C[862]) );
  FA_162 \FA_INST_0[1].FA_INST_1[350].FA_  ( .A(A[862]), .B(B[862]), .CI(
        C[862]), .S(S[862]), .CO(C[863]) );
  FA_161 \FA_INST_0[1].FA_INST_1[351].FA_  ( .A(A[863]), .B(B[863]), .CI(
        C[863]), .S(S[863]), .CO(C[864]) );
  FA_160 \FA_INST_0[1].FA_INST_1[352].FA_  ( .A(A[864]), .B(B[864]), .CI(
        C[864]), .S(S[864]), .CO(C[865]) );
  FA_159 \FA_INST_0[1].FA_INST_1[353].FA_  ( .A(A[865]), .B(B[865]), .CI(
        C[865]), .S(S[865]), .CO(C[866]) );
  FA_158 \FA_INST_0[1].FA_INST_1[354].FA_  ( .A(A[866]), .B(B[866]), .CI(
        C[866]), .S(S[866]), .CO(C[867]) );
  FA_157 \FA_INST_0[1].FA_INST_1[355].FA_  ( .A(A[867]), .B(B[867]), .CI(
        C[867]), .S(S[867]), .CO(C[868]) );
  FA_156 \FA_INST_0[1].FA_INST_1[356].FA_  ( .A(A[868]), .B(B[868]), .CI(
        C[868]), .S(S[868]), .CO(C[869]) );
  FA_155 \FA_INST_0[1].FA_INST_1[357].FA_  ( .A(A[869]), .B(B[869]), .CI(
        C[869]), .S(S[869]), .CO(C[870]) );
  FA_154 \FA_INST_0[1].FA_INST_1[358].FA_  ( .A(A[870]), .B(B[870]), .CI(
        C[870]), .S(S[870]), .CO(C[871]) );
  FA_153 \FA_INST_0[1].FA_INST_1[359].FA_  ( .A(A[871]), .B(B[871]), .CI(
        C[871]), .S(S[871]), .CO(C[872]) );
  FA_152 \FA_INST_0[1].FA_INST_1[360].FA_  ( .A(A[872]), .B(B[872]), .CI(
        C[872]), .S(S[872]), .CO(C[873]) );
  FA_151 \FA_INST_0[1].FA_INST_1[361].FA_  ( .A(A[873]), .B(B[873]), .CI(
        C[873]), .S(S[873]), .CO(C[874]) );
  FA_150 \FA_INST_0[1].FA_INST_1[362].FA_  ( .A(A[874]), .B(B[874]), .CI(
        C[874]), .S(S[874]), .CO(C[875]) );
  FA_149 \FA_INST_0[1].FA_INST_1[363].FA_  ( .A(A[875]), .B(B[875]), .CI(
        C[875]), .S(S[875]), .CO(C[876]) );
  FA_148 \FA_INST_0[1].FA_INST_1[364].FA_  ( .A(A[876]), .B(B[876]), .CI(
        C[876]), .S(S[876]), .CO(C[877]) );
  FA_147 \FA_INST_0[1].FA_INST_1[365].FA_  ( .A(A[877]), .B(B[877]), .CI(
        C[877]), .S(S[877]), .CO(C[878]) );
  FA_146 \FA_INST_0[1].FA_INST_1[366].FA_  ( .A(A[878]), .B(B[878]), .CI(
        C[878]), .S(S[878]), .CO(C[879]) );
  FA_145 \FA_INST_0[1].FA_INST_1[367].FA_  ( .A(A[879]), .B(B[879]), .CI(
        C[879]), .S(S[879]), .CO(C[880]) );
  FA_144 \FA_INST_0[1].FA_INST_1[368].FA_  ( .A(A[880]), .B(B[880]), .CI(
        C[880]), .S(S[880]), .CO(C[881]) );
  FA_143 \FA_INST_0[1].FA_INST_1[369].FA_  ( .A(A[881]), .B(B[881]), .CI(
        C[881]), .S(S[881]), .CO(C[882]) );
  FA_142 \FA_INST_0[1].FA_INST_1[370].FA_  ( .A(A[882]), .B(B[882]), .CI(
        C[882]), .S(S[882]), .CO(C[883]) );
  FA_141 \FA_INST_0[1].FA_INST_1[371].FA_  ( .A(A[883]), .B(B[883]), .CI(
        C[883]), .S(S[883]), .CO(C[884]) );
  FA_140 \FA_INST_0[1].FA_INST_1[372].FA_  ( .A(A[884]), .B(B[884]), .CI(
        C[884]), .S(S[884]), .CO(C[885]) );
  FA_139 \FA_INST_0[1].FA_INST_1[373].FA_  ( .A(A[885]), .B(B[885]), .CI(
        C[885]), .S(S[885]), .CO(C[886]) );
  FA_138 \FA_INST_0[1].FA_INST_1[374].FA_  ( .A(A[886]), .B(B[886]), .CI(
        C[886]), .S(S[886]), .CO(C[887]) );
  FA_137 \FA_INST_0[1].FA_INST_1[375].FA_  ( .A(A[887]), .B(B[887]), .CI(
        C[887]), .S(S[887]), .CO(C[888]) );
  FA_136 \FA_INST_0[1].FA_INST_1[376].FA_  ( .A(A[888]), .B(B[888]), .CI(
        C[888]), .S(S[888]), .CO(C[889]) );
  FA_135 \FA_INST_0[1].FA_INST_1[377].FA_  ( .A(A[889]), .B(B[889]), .CI(
        C[889]), .S(S[889]), .CO(C[890]) );
  FA_134 \FA_INST_0[1].FA_INST_1[378].FA_  ( .A(A[890]), .B(B[890]), .CI(
        C[890]), .S(S[890]), .CO(C[891]) );
  FA_133 \FA_INST_0[1].FA_INST_1[379].FA_  ( .A(A[891]), .B(B[891]), .CI(
        C[891]), .S(S[891]), .CO(C[892]) );
  FA_132 \FA_INST_0[1].FA_INST_1[380].FA_  ( .A(A[892]), .B(B[892]), .CI(
        C[892]), .S(S[892]), .CO(C[893]) );
  FA_131 \FA_INST_0[1].FA_INST_1[381].FA_  ( .A(A[893]), .B(B[893]), .CI(
        C[893]), .S(S[893]), .CO(C[894]) );
  FA_130 \FA_INST_0[1].FA_INST_1[382].FA_  ( .A(A[894]), .B(B[894]), .CI(
        C[894]), .S(S[894]), .CO(C[895]) );
  FA_129 \FA_INST_0[1].FA_INST_1[383].FA_  ( .A(A[895]), .B(B[895]), .CI(
        C[895]), .S(S[895]), .CO(C[896]) );
  FA_128 \FA_INST_0[1].FA_INST_1[384].FA_  ( .A(A[896]), .B(B[896]), .CI(
        C[896]), .S(S[896]), .CO(C[897]) );
  FA_127 \FA_INST_0[1].FA_INST_1[385].FA_  ( .A(A[897]), .B(B[897]), .CI(
        C[897]), .S(S[897]), .CO(C[898]) );
  FA_126 \FA_INST_0[1].FA_INST_1[386].FA_  ( .A(A[898]), .B(B[898]), .CI(
        C[898]), .S(S[898]), .CO(C[899]) );
  FA_125 \FA_INST_0[1].FA_INST_1[387].FA_  ( .A(A[899]), .B(B[899]), .CI(
        C[899]), .S(S[899]), .CO(C[900]) );
  FA_124 \FA_INST_0[1].FA_INST_1[388].FA_  ( .A(A[900]), .B(B[900]), .CI(
        C[900]), .S(S[900]), .CO(C[901]) );
  FA_123 \FA_INST_0[1].FA_INST_1[389].FA_  ( .A(A[901]), .B(B[901]), .CI(
        C[901]), .S(S[901]), .CO(C[902]) );
  FA_122 \FA_INST_0[1].FA_INST_1[390].FA_  ( .A(A[902]), .B(B[902]), .CI(
        C[902]), .S(S[902]), .CO(C[903]) );
  FA_121 \FA_INST_0[1].FA_INST_1[391].FA_  ( .A(A[903]), .B(B[903]), .CI(
        C[903]), .S(S[903]), .CO(C[904]) );
  FA_120 \FA_INST_0[1].FA_INST_1[392].FA_  ( .A(A[904]), .B(B[904]), .CI(
        C[904]), .S(S[904]), .CO(C[905]) );
  FA_119 \FA_INST_0[1].FA_INST_1[393].FA_  ( .A(A[905]), .B(B[905]), .CI(
        C[905]), .S(S[905]), .CO(C[906]) );
  FA_118 \FA_INST_0[1].FA_INST_1[394].FA_  ( .A(A[906]), .B(B[906]), .CI(
        C[906]), .S(S[906]), .CO(C[907]) );
  FA_117 \FA_INST_0[1].FA_INST_1[395].FA_  ( .A(A[907]), .B(B[907]), .CI(
        C[907]), .S(S[907]), .CO(C[908]) );
  FA_116 \FA_INST_0[1].FA_INST_1[396].FA_  ( .A(A[908]), .B(B[908]), .CI(
        C[908]), .S(S[908]), .CO(C[909]) );
  FA_115 \FA_INST_0[1].FA_INST_1[397].FA_  ( .A(A[909]), .B(B[909]), .CI(
        C[909]), .S(S[909]), .CO(C[910]) );
  FA_114 \FA_INST_0[1].FA_INST_1[398].FA_  ( .A(A[910]), .B(B[910]), .CI(
        C[910]), .S(S[910]), .CO(C[911]) );
  FA_113 \FA_INST_0[1].FA_INST_1[399].FA_  ( .A(A[911]), .B(B[911]), .CI(
        C[911]), .S(S[911]), .CO(C[912]) );
  FA_112 \FA_INST_0[1].FA_INST_1[400].FA_  ( .A(A[912]), .B(B[912]), .CI(
        C[912]), .S(S[912]), .CO(C[913]) );
  FA_111 \FA_INST_0[1].FA_INST_1[401].FA_  ( .A(A[913]), .B(B[913]), .CI(
        C[913]), .S(S[913]), .CO(C[914]) );
  FA_110 \FA_INST_0[1].FA_INST_1[402].FA_  ( .A(A[914]), .B(B[914]), .CI(
        C[914]), .S(S[914]), .CO(C[915]) );
  FA_109 \FA_INST_0[1].FA_INST_1[403].FA_  ( .A(A[915]), .B(B[915]), .CI(
        C[915]), .S(S[915]), .CO(C[916]) );
  FA_108 \FA_INST_0[1].FA_INST_1[404].FA_  ( .A(A[916]), .B(B[916]), .CI(
        C[916]), .S(S[916]), .CO(C[917]) );
  FA_107 \FA_INST_0[1].FA_INST_1[405].FA_  ( .A(A[917]), .B(B[917]), .CI(
        C[917]), .S(S[917]), .CO(C[918]) );
  FA_106 \FA_INST_0[1].FA_INST_1[406].FA_  ( .A(A[918]), .B(B[918]), .CI(
        C[918]), .S(S[918]), .CO(C[919]) );
  FA_105 \FA_INST_0[1].FA_INST_1[407].FA_  ( .A(A[919]), .B(B[919]), .CI(
        C[919]), .S(S[919]), .CO(C[920]) );
  FA_104 \FA_INST_0[1].FA_INST_1[408].FA_  ( .A(A[920]), .B(B[920]), .CI(
        C[920]), .S(S[920]), .CO(C[921]) );
  FA_103 \FA_INST_0[1].FA_INST_1[409].FA_  ( .A(A[921]), .B(B[921]), .CI(
        C[921]), .S(S[921]), .CO(C[922]) );
  FA_102 \FA_INST_0[1].FA_INST_1[410].FA_  ( .A(A[922]), .B(B[922]), .CI(
        C[922]), .S(S[922]), .CO(C[923]) );
  FA_101 \FA_INST_0[1].FA_INST_1[411].FA_  ( .A(A[923]), .B(B[923]), .CI(
        C[923]), .S(S[923]), .CO(C[924]) );
  FA_100 \FA_INST_0[1].FA_INST_1[412].FA_  ( .A(A[924]), .B(B[924]), .CI(
        C[924]), .S(S[924]), .CO(C[925]) );
  FA_99 \FA_INST_0[1].FA_INST_1[413].FA_  ( .A(A[925]), .B(B[925]), .CI(C[925]), .S(S[925]), .CO(C[926]) );
  FA_98 \FA_INST_0[1].FA_INST_1[414].FA_  ( .A(A[926]), .B(B[926]), .CI(C[926]), .S(S[926]), .CO(C[927]) );
  FA_97 \FA_INST_0[1].FA_INST_1[415].FA_  ( .A(A[927]), .B(B[927]), .CI(C[927]), .S(S[927]), .CO(C[928]) );
  FA_96 \FA_INST_0[1].FA_INST_1[416].FA_  ( .A(A[928]), .B(B[928]), .CI(C[928]), .S(S[928]), .CO(C[929]) );
  FA_95 \FA_INST_0[1].FA_INST_1[417].FA_  ( .A(A[929]), .B(B[929]), .CI(C[929]), .S(S[929]), .CO(C[930]) );
  FA_94 \FA_INST_0[1].FA_INST_1[418].FA_  ( .A(A[930]), .B(B[930]), .CI(C[930]), .S(S[930]), .CO(C[931]) );
  FA_93 \FA_INST_0[1].FA_INST_1[419].FA_  ( .A(A[931]), .B(B[931]), .CI(C[931]), .S(S[931]), .CO(C[932]) );
  FA_92 \FA_INST_0[1].FA_INST_1[420].FA_  ( .A(A[932]), .B(B[932]), .CI(C[932]), .S(S[932]), .CO(C[933]) );
  FA_91 \FA_INST_0[1].FA_INST_1[421].FA_  ( .A(A[933]), .B(B[933]), .CI(C[933]), .S(S[933]), .CO(C[934]) );
  FA_90 \FA_INST_0[1].FA_INST_1[422].FA_  ( .A(A[934]), .B(B[934]), .CI(C[934]), .S(S[934]), .CO(C[935]) );
  FA_89 \FA_INST_0[1].FA_INST_1[423].FA_  ( .A(A[935]), .B(B[935]), .CI(C[935]), .S(S[935]), .CO(C[936]) );
  FA_88 \FA_INST_0[1].FA_INST_1[424].FA_  ( .A(A[936]), .B(B[936]), .CI(C[936]), .S(S[936]), .CO(C[937]) );
  FA_87 \FA_INST_0[1].FA_INST_1[425].FA_  ( .A(A[937]), .B(B[937]), .CI(C[937]), .S(S[937]), .CO(C[938]) );
  FA_86 \FA_INST_0[1].FA_INST_1[426].FA_  ( .A(A[938]), .B(B[938]), .CI(C[938]), .S(S[938]), .CO(C[939]) );
  FA_85 \FA_INST_0[1].FA_INST_1[427].FA_  ( .A(A[939]), .B(B[939]), .CI(C[939]), .S(S[939]), .CO(C[940]) );
  FA_84 \FA_INST_0[1].FA_INST_1[428].FA_  ( .A(A[940]), .B(B[940]), .CI(C[940]), .S(S[940]), .CO(C[941]) );
  FA_83 \FA_INST_0[1].FA_INST_1[429].FA_  ( .A(A[941]), .B(B[941]), .CI(C[941]), .S(S[941]), .CO(C[942]) );
  FA_82 \FA_INST_0[1].FA_INST_1[430].FA_  ( .A(A[942]), .B(B[942]), .CI(C[942]), .S(S[942]), .CO(C[943]) );
  FA_81 \FA_INST_0[1].FA_INST_1[431].FA_  ( .A(A[943]), .B(B[943]), .CI(C[943]), .S(S[943]), .CO(C[944]) );
  FA_80 \FA_INST_0[1].FA_INST_1[432].FA_  ( .A(A[944]), .B(B[944]), .CI(C[944]), .S(S[944]), .CO(C[945]) );
  FA_79 \FA_INST_0[1].FA_INST_1[433].FA_  ( .A(A[945]), .B(B[945]), .CI(C[945]), .S(S[945]), .CO(C[946]) );
  FA_78 \FA_INST_0[1].FA_INST_1[434].FA_  ( .A(A[946]), .B(B[946]), .CI(C[946]), .S(S[946]), .CO(C[947]) );
  FA_77 \FA_INST_0[1].FA_INST_1[435].FA_  ( .A(A[947]), .B(B[947]), .CI(C[947]), .S(S[947]), .CO(C[948]) );
  FA_76 \FA_INST_0[1].FA_INST_1[436].FA_  ( .A(A[948]), .B(B[948]), .CI(C[948]), .S(S[948]), .CO(C[949]) );
  FA_75 \FA_INST_0[1].FA_INST_1[437].FA_  ( .A(A[949]), .B(B[949]), .CI(C[949]), .S(S[949]), .CO(C[950]) );
  FA_74 \FA_INST_0[1].FA_INST_1[438].FA_  ( .A(A[950]), .B(B[950]), .CI(C[950]), .S(S[950]), .CO(C[951]) );
  FA_73 \FA_INST_0[1].FA_INST_1[439].FA_  ( .A(A[951]), .B(B[951]), .CI(C[951]), .S(S[951]), .CO(C[952]) );
  FA_72 \FA_INST_0[1].FA_INST_1[440].FA_  ( .A(A[952]), .B(B[952]), .CI(C[952]), .S(S[952]), .CO(C[953]) );
  FA_71 \FA_INST_0[1].FA_INST_1[441].FA_  ( .A(A[953]), .B(B[953]), .CI(C[953]), .S(S[953]), .CO(C[954]) );
  FA_70 \FA_INST_0[1].FA_INST_1[442].FA_  ( .A(A[954]), .B(B[954]), .CI(C[954]), .S(S[954]), .CO(C[955]) );
  FA_69 \FA_INST_0[1].FA_INST_1[443].FA_  ( .A(A[955]), .B(B[955]), .CI(C[955]), .S(S[955]), .CO(C[956]) );
  FA_68 \FA_INST_0[1].FA_INST_1[444].FA_  ( .A(A[956]), .B(B[956]), .CI(C[956]), .S(S[956]), .CO(C[957]) );
  FA_67 \FA_INST_0[1].FA_INST_1[445].FA_  ( .A(A[957]), .B(B[957]), .CI(C[957]), .S(S[957]), .CO(C[958]) );
  FA_66 \FA_INST_0[1].FA_INST_1[446].FA_  ( .A(A[958]), .B(B[958]), .CI(C[958]), .S(S[958]), .CO(C[959]) );
  FA_65 \FA_INST_0[1].FA_INST_1[447].FA_  ( .A(A[959]), .B(B[959]), .CI(C[959]), .S(S[959]), .CO(C[960]) );
  FA_64 \FA_INST_0[1].FA_INST_1[448].FA_  ( .A(A[960]), .B(B[960]), .CI(C[960]), .S(S[960]), .CO(C[961]) );
  FA_63 \FA_INST_0[1].FA_INST_1[449].FA_  ( .A(A[961]), .B(B[961]), .CI(C[961]), .S(S[961]), .CO(C[962]) );
  FA_62 \FA_INST_0[1].FA_INST_1[450].FA_  ( .A(A[962]), .B(B[962]), .CI(C[962]), .S(S[962]), .CO(C[963]) );
  FA_61 \FA_INST_0[1].FA_INST_1[451].FA_  ( .A(A[963]), .B(B[963]), .CI(C[963]), .S(S[963]), .CO(C[964]) );
  FA_60 \FA_INST_0[1].FA_INST_1[452].FA_  ( .A(A[964]), .B(B[964]), .CI(C[964]), .S(S[964]), .CO(C[965]) );
  FA_59 \FA_INST_0[1].FA_INST_1[453].FA_  ( .A(A[965]), .B(B[965]), .CI(C[965]), .S(S[965]), .CO(C[966]) );
  FA_58 \FA_INST_0[1].FA_INST_1[454].FA_  ( .A(A[966]), .B(B[966]), .CI(C[966]), .S(S[966]), .CO(C[967]) );
  FA_57 \FA_INST_0[1].FA_INST_1[455].FA_  ( .A(A[967]), .B(B[967]), .CI(C[967]), .S(S[967]), .CO(C[968]) );
  FA_56 \FA_INST_0[1].FA_INST_1[456].FA_  ( .A(A[968]), .B(B[968]), .CI(C[968]), .S(S[968]), .CO(C[969]) );
  FA_55 \FA_INST_0[1].FA_INST_1[457].FA_  ( .A(A[969]), .B(B[969]), .CI(C[969]), .S(S[969]), .CO(C[970]) );
  FA_54 \FA_INST_0[1].FA_INST_1[458].FA_  ( .A(A[970]), .B(B[970]), .CI(C[970]), .S(S[970]), .CO(C[971]) );
  FA_53 \FA_INST_0[1].FA_INST_1[459].FA_  ( .A(A[971]), .B(B[971]), .CI(C[971]), .S(S[971]), .CO(C[972]) );
  FA_52 \FA_INST_0[1].FA_INST_1[460].FA_  ( .A(A[972]), .B(B[972]), .CI(C[972]), .S(S[972]), .CO(C[973]) );
  FA_51 \FA_INST_0[1].FA_INST_1[461].FA_  ( .A(A[973]), .B(B[973]), .CI(C[973]), .S(S[973]), .CO(C[974]) );
  FA_50 \FA_INST_0[1].FA_INST_1[462].FA_  ( .A(A[974]), .B(B[974]), .CI(C[974]), .S(S[974]), .CO(C[975]) );
  FA_49 \FA_INST_0[1].FA_INST_1[463].FA_  ( .A(A[975]), .B(B[975]), .CI(C[975]), .S(S[975]), .CO(C[976]) );
  FA_48 \FA_INST_0[1].FA_INST_1[464].FA_  ( .A(A[976]), .B(B[976]), .CI(C[976]), .S(S[976]), .CO(C[977]) );
  FA_47 \FA_INST_0[1].FA_INST_1[465].FA_  ( .A(A[977]), .B(B[977]), .CI(C[977]), .S(S[977]), .CO(C[978]) );
  FA_46 \FA_INST_0[1].FA_INST_1[466].FA_  ( .A(A[978]), .B(B[978]), .CI(C[978]), .S(S[978]), .CO(C[979]) );
  FA_45 \FA_INST_0[1].FA_INST_1[467].FA_  ( .A(A[979]), .B(B[979]), .CI(C[979]), .S(S[979]), .CO(C[980]) );
  FA_44 \FA_INST_0[1].FA_INST_1[468].FA_  ( .A(A[980]), .B(B[980]), .CI(C[980]), .S(S[980]), .CO(C[981]) );
  FA_43 \FA_INST_0[1].FA_INST_1[469].FA_  ( .A(A[981]), .B(B[981]), .CI(C[981]), .S(S[981]), .CO(C[982]) );
  FA_42 \FA_INST_0[1].FA_INST_1[470].FA_  ( .A(A[982]), .B(B[982]), .CI(C[982]), .S(S[982]), .CO(C[983]) );
  FA_41 \FA_INST_0[1].FA_INST_1[471].FA_  ( .A(A[983]), .B(B[983]), .CI(C[983]), .S(S[983]), .CO(C[984]) );
  FA_40 \FA_INST_0[1].FA_INST_1[472].FA_  ( .A(A[984]), .B(B[984]), .CI(C[984]), .S(S[984]), .CO(C[985]) );
  FA_39 \FA_INST_0[1].FA_INST_1[473].FA_  ( .A(A[985]), .B(B[985]), .CI(C[985]), .S(S[985]), .CO(C[986]) );
  FA_38 \FA_INST_0[1].FA_INST_1[474].FA_  ( .A(A[986]), .B(B[986]), .CI(C[986]), .S(S[986]), .CO(C[987]) );
  FA_37 \FA_INST_0[1].FA_INST_1[475].FA_  ( .A(A[987]), .B(B[987]), .CI(C[987]), .S(S[987]), .CO(C[988]) );
  FA_36 \FA_INST_0[1].FA_INST_1[476].FA_  ( .A(A[988]), .B(B[988]), .CI(C[988]), .S(S[988]), .CO(C[989]) );
  FA_35 \FA_INST_0[1].FA_INST_1[477].FA_  ( .A(A[989]), .B(B[989]), .CI(C[989]), .S(S[989]), .CO(C[990]) );
  FA_34 \FA_INST_0[1].FA_INST_1[478].FA_  ( .A(A[990]), .B(B[990]), .CI(C[990]), .S(S[990]), .CO(C[991]) );
  FA_33 \FA_INST_0[1].FA_INST_1[479].FA_  ( .A(A[991]), .B(B[991]), .CI(C[991]), .S(S[991]), .CO(C[992]) );
  FA_32 \FA_INST_0[1].FA_INST_1[480].FA_  ( .A(A[992]), .B(B[992]), .CI(C[992]), .S(S[992]), .CO(C[993]) );
  FA_31 \FA_INST_0[1].FA_INST_1[481].FA_  ( .A(A[993]), .B(B[993]), .CI(C[993]), .S(S[993]), .CO(C[994]) );
  FA_30 \FA_INST_0[1].FA_INST_1[482].FA_  ( .A(A[994]), .B(B[994]), .CI(C[994]), .S(S[994]), .CO(C[995]) );
  FA_29 \FA_INST_0[1].FA_INST_1[483].FA_  ( .A(A[995]), .B(B[995]), .CI(C[995]), .S(S[995]), .CO(C[996]) );
  FA_28 \FA_INST_0[1].FA_INST_1[484].FA_  ( .A(A[996]), .B(B[996]), .CI(C[996]), .S(S[996]), .CO(C[997]) );
  FA_27 \FA_INST_0[1].FA_INST_1[485].FA_  ( .A(A[997]), .B(B[997]), .CI(C[997]), .S(S[997]), .CO(C[998]) );
  FA_26 \FA_INST_0[1].FA_INST_1[486].FA_  ( .A(A[998]), .B(B[998]), .CI(C[998]), .S(S[998]), .CO(C[999]) );
  FA_25 \FA_INST_0[1].FA_INST_1[487].FA_  ( .A(A[999]), .B(B[999]), .CI(C[999]), .S(S[999]), .CO(C[1000]) );
  FA_24 \FA_INST_0[1].FA_INST_1[488].FA_  ( .A(A[1000]), .B(B[1000]), .CI(
        C[1000]), .S(S[1000]), .CO(C[1001]) );
  FA_23 \FA_INST_0[1].FA_INST_1[489].FA_  ( .A(A[1001]), .B(B[1001]), .CI(
        C[1001]), .S(S[1001]), .CO(C[1002]) );
  FA_22 \FA_INST_0[1].FA_INST_1[490].FA_  ( .A(A[1002]), .B(B[1002]), .CI(
        C[1002]), .S(S[1002]), .CO(C[1003]) );
  FA_21 \FA_INST_0[1].FA_INST_1[491].FA_  ( .A(A[1003]), .B(B[1003]), .CI(
        C[1003]), .S(S[1003]), .CO(C[1004]) );
  FA_20 \FA_INST_0[1].FA_INST_1[492].FA_  ( .A(A[1004]), .B(B[1004]), .CI(
        C[1004]), .S(S[1004]), .CO(C[1005]) );
  FA_19 \FA_INST_0[1].FA_INST_1[493].FA_  ( .A(A[1005]), .B(B[1005]), .CI(
        C[1005]), .S(S[1005]), .CO(C[1006]) );
  FA_18 \FA_INST_0[1].FA_INST_1[494].FA_  ( .A(A[1006]), .B(B[1006]), .CI(
        C[1006]), .S(S[1006]), .CO(C[1007]) );
  FA_17 \FA_INST_0[1].FA_INST_1[495].FA_  ( .A(A[1007]), .B(B[1007]), .CI(
        C[1007]), .S(S[1007]), .CO(C[1008]) );
  FA_16 \FA_INST_0[1].FA_INST_1[496].FA_  ( .A(A[1008]), .B(B[1008]), .CI(
        C[1008]), .S(S[1008]), .CO(C[1009]) );
  FA_15 \FA_INST_0[1].FA_INST_1[497].FA_  ( .A(A[1009]), .B(B[1009]), .CI(
        C[1009]), .S(S[1009]), .CO(C[1010]) );
  FA_14 \FA_INST_0[1].FA_INST_1[498].FA_  ( .A(A[1010]), .B(B[1010]), .CI(
        C[1010]), .S(S[1010]), .CO(C[1011]) );
  FA_13 \FA_INST_0[1].FA_INST_1[499].FA_  ( .A(A[1011]), .B(B[1011]), .CI(
        C[1011]), .S(S[1011]), .CO(C[1012]) );
  FA_12 \FA_INST_0[1].FA_INST_1[500].FA_  ( .A(A[1012]), .B(B[1012]), .CI(
        C[1012]), .S(S[1012]), .CO(C[1013]) );
  FA_11 \FA_INST_0[1].FA_INST_1[501].FA_  ( .A(A[1013]), .B(B[1013]), .CI(
        C[1013]), .S(S[1013]), .CO(C[1014]) );
  FA_10 \FA_INST_0[1].FA_INST_1[502].FA_  ( .A(A[1014]), .B(B[1014]), .CI(
        C[1014]), .S(S[1014]), .CO(C[1015]) );
  FA_9 \FA_INST_0[1].FA_INST_1[503].FA_  ( .A(A[1015]), .B(B[1015]), .CI(
        C[1015]), .S(S[1015]), .CO(C[1016]) );
  FA_8 \FA_INST_0[1].FA_INST_1[504].FA_  ( .A(A[1016]), .B(B[1016]), .CI(
        C[1016]), .S(S[1016]), .CO(C[1017]) );
  FA_7 \FA_INST_0[1].FA_INST_1[505].FA_  ( .A(A[1017]), .B(B[1017]), .CI(
        C[1017]), .S(S[1017]), .CO(C[1018]) );
  FA_6 \FA_INST_0[1].FA_INST_1[506].FA_  ( .A(A[1018]), .B(B[1018]), .CI(
        C[1018]), .S(S[1018]), .CO(C[1019]) );
  FA_5 \FA_INST_0[1].FA_INST_1[507].FA_  ( .A(A[1019]), .B(B[1019]), .CI(
        C[1019]), .S(S[1019]), .CO(C[1020]) );
  FA_4 \FA_INST_0[1].FA_INST_1[508].FA_  ( .A(A[1020]), .B(B[1020]), .CI(
        C[1020]), .S(S[1020]), .CO(C[1021]) );
  FA_3 \FA_INST_0[1].FA_INST_1[509].FA_  ( .A(A[1021]), .B(B[1021]), .CI(
        C[1021]), .S(S[1021]), .CO(C[1022]) );
  FA_2 \FA_INST_0[1].FA_INST_1[510].FA_  ( .A(A[1022]), .B(B[1022]), .CI(
        C[1022]), .S(S[1022]) );
  FA_1 \FA_INST_0[1].FA_INST_1[511].FA_  ( .A(1'b0), .B(B[1023]), .CI(1'b0), 
        .S(S[1023]) );
endmodule


module mult_N1024_CC1024_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [1023:0] A;
  input [0:0] B;
  output [1024:0] PRODUCT;
  input TC;


  AND U2 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  AND U3 ( .A(A[1]), .B(B[0]), .Z(PRODUCT[1]) );
  AND U4 ( .A(A[2]), .B(B[0]), .Z(PRODUCT[2]) );
  AND U5 ( .A(A[3]), .B(B[0]), .Z(PRODUCT[3]) );
  AND U6 ( .A(A[4]), .B(B[0]), .Z(PRODUCT[4]) );
  AND U7 ( .A(A[5]), .B(B[0]), .Z(PRODUCT[5]) );
  AND U8 ( .A(A[6]), .B(B[0]), .Z(PRODUCT[6]) );
  AND U9 ( .A(A[7]), .B(B[0]), .Z(PRODUCT[7]) );
  AND U10 ( .A(A[8]), .B(B[0]), .Z(PRODUCT[8]) );
  AND U11 ( .A(A[9]), .B(B[0]), .Z(PRODUCT[9]) );
  AND U12 ( .A(A[10]), .B(B[0]), .Z(PRODUCT[10]) );
  AND U13 ( .A(A[11]), .B(B[0]), .Z(PRODUCT[11]) );
  AND U14 ( .A(A[12]), .B(B[0]), .Z(PRODUCT[12]) );
  AND U15 ( .A(A[13]), .B(B[0]), .Z(PRODUCT[13]) );
  AND U16 ( .A(A[14]), .B(B[0]), .Z(PRODUCT[14]) );
  AND U17 ( .A(A[15]), .B(B[0]), .Z(PRODUCT[15]) );
  AND U18 ( .A(A[16]), .B(B[0]), .Z(PRODUCT[16]) );
  AND U19 ( .A(A[17]), .B(B[0]), .Z(PRODUCT[17]) );
  AND U20 ( .A(A[18]), .B(B[0]), .Z(PRODUCT[18]) );
  AND U21 ( .A(A[19]), .B(B[0]), .Z(PRODUCT[19]) );
  AND U22 ( .A(A[20]), .B(B[0]), .Z(PRODUCT[20]) );
  AND U23 ( .A(A[21]), .B(B[0]), .Z(PRODUCT[21]) );
  AND U24 ( .A(A[22]), .B(B[0]), .Z(PRODUCT[22]) );
  AND U25 ( .A(A[23]), .B(B[0]), .Z(PRODUCT[23]) );
  AND U26 ( .A(A[24]), .B(B[0]), .Z(PRODUCT[24]) );
  AND U27 ( .A(A[25]), .B(B[0]), .Z(PRODUCT[25]) );
  AND U28 ( .A(A[26]), .B(B[0]), .Z(PRODUCT[26]) );
  AND U29 ( .A(A[27]), .B(B[0]), .Z(PRODUCT[27]) );
  AND U30 ( .A(A[28]), .B(B[0]), .Z(PRODUCT[28]) );
  AND U31 ( .A(A[29]), .B(B[0]), .Z(PRODUCT[29]) );
  AND U32 ( .A(A[30]), .B(B[0]), .Z(PRODUCT[30]) );
  AND U33 ( .A(A[31]), .B(B[0]), .Z(PRODUCT[31]) );
  AND U34 ( .A(A[32]), .B(B[0]), .Z(PRODUCT[32]) );
  AND U35 ( .A(A[33]), .B(B[0]), .Z(PRODUCT[33]) );
  AND U36 ( .A(A[34]), .B(B[0]), .Z(PRODUCT[34]) );
  AND U37 ( .A(A[35]), .B(B[0]), .Z(PRODUCT[35]) );
  AND U38 ( .A(A[36]), .B(B[0]), .Z(PRODUCT[36]) );
  AND U39 ( .A(A[37]), .B(B[0]), .Z(PRODUCT[37]) );
  AND U40 ( .A(A[38]), .B(B[0]), .Z(PRODUCT[38]) );
  AND U41 ( .A(A[39]), .B(B[0]), .Z(PRODUCT[39]) );
  AND U42 ( .A(A[40]), .B(B[0]), .Z(PRODUCT[40]) );
  AND U43 ( .A(A[41]), .B(B[0]), .Z(PRODUCT[41]) );
  AND U44 ( .A(A[42]), .B(B[0]), .Z(PRODUCT[42]) );
  AND U45 ( .A(A[43]), .B(B[0]), .Z(PRODUCT[43]) );
  AND U46 ( .A(A[44]), .B(B[0]), .Z(PRODUCT[44]) );
  AND U47 ( .A(A[45]), .B(B[0]), .Z(PRODUCT[45]) );
  AND U48 ( .A(A[46]), .B(B[0]), .Z(PRODUCT[46]) );
  AND U49 ( .A(A[47]), .B(B[0]), .Z(PRODUCT[47]) );
  AND U50 ( .A(A[48]), .B(B[0]), .Z(PRODUCT[48]) );
  AND U51 ( .A(A[49]), .B(B[0]), .Z(PRODUCT[49]) );
  AND U52 ( .A(A[50]), .B(B[0]), .Z(PRODUCT[50]) );
  AND U53 ( .A(A[51]), .B(B[0]), .Z(PRODUCT[51]) );
  AND U54 ( .A(A[52]), .B(B[0]), .Z(PRODUCT[52]) );
  AND U55 ( .A(A[53]), .B(B[0]), .Z(PRODUCT[53]) );
  AND U56 ( .A(A[54]), .B(B[0]), .Z(PRODUCT[54]) );
  AND U57 ( .A(A[55]), .B(B[0]), .Z(PRODUCT[55]) );
  AND U58 ( .A(A[56]), .B(B[0]), .Z(PRODUCT[56]) );
  AND U59 ( .A(A[57]), .B(B[0]), .Z(PRODUCT[57]) );
  AND U60 ( .A(A[58]), .B(B[0]), .Z(PRODUCT[58]) );
  AND U61 ( .A(A[59]), .B(B[0]), .Z(PRODUCT[59]) );
  AND U62 ( .A(A[60]), .B(B[0]), .Z(PRODUCT[60]) );
  AND U63 ( .A(A[61]), .B(B[0]), .Z(PRODUCT[61]) );
  AND U64 ( .A(A[62]), .B(B[0]), .Z(PRODUCT[62]) );
  AND U65 ( .A(A[63]), .B(B[0]), .Z(PRODUCT[63]) );
  AND U66 ( .A(A[64]), .B(B[0]), .Z(PRODUCT[64]) );
  AND U67 ( .A(A[65]), .B(B[0]), .Z(PRODUCT[65]) );
  AND U68 ( .A(A[66]), .B(B[0]), .Z(PRODUCT[66]) );
  AND U69 ( .A(A[67]), .B(B[0]), .Z(PRODUCT[67]) );
  AND U70 ( .A(A[68]), .B(B[0]), .Z(PRODUCT[68]) );
  AND U71 ( .A(A[69]), .B(B[0]), .Z(PRODUCT[69]) );
  AND U72 ( .A(A[70]), .B(B[0]), .Z(PRODUCT[70]) );
  AND U73 ( .A(A[71]), .B(B[0]), .Z(PRODUCT[71]) );
  AND U74 ( .A(A[72]), .B(B[0]), .Z(PRODUCT[72]) );
  AND U75 ( .A(A[73]), .B(B[0]), .Z(PRODUCT[73]) );
  AND U76 ( .A(A[74]), .B(B[0]), .Z(PRODUCT[74]) );
  AND U77 ( .A(A[75]), .B(B[0]), .Z(PRODUCT[75]) );
  AND U78 ( .A(A[76]), .B(B[0]), .Z(PRODUCT[76]) );
  AND U79 ( .A(A[77]), .B(B[0]), .Z(PRODUCT[77]) );
  AND U80 ( .A(A[78]), .B(B[0]), .Z(PRODUCT[78]) );
  AND U81 ( .A(A[79]), .B(B[0]), .Z(PRODUCT[79]) );
  AND U82 ( .A(A[80]), .B(B[0]), .Z(PRODUCT[80]) );
  AND U83 ( .A(A[81]), .B(B[0]), .Z(PRODUCT[81]) );
  AND U84 ( .A(A[82]), .B(B[0]), .Z(PRODUCT[82]) );
  AND U85 ( .A(A[83]), .B(B[0]), .Z(PRODUCT[83]) );
  AND U86 ( .A(A[84]), .B(B[0]), .Z(PRODUCT[84]) );
  AND U87 ( .A(A[85]), .B(B[0]), .Z(PRODUCT[85]) );
  AND U88 ( .A(A[86]), .B(B[0]), .Z(PRODUCT[86]) );
  AND U89 ( .A(A[87]), .B(B[0]), .Z(PRODUCT[87]) );
  AND U90 ( .A(A[88]), .B(B[0]), .Z(PRODUCT[88]) );
  AND U91 ( .A(A[89]), .B(B[0]), .Z(PRODUCT[89]) );
  AND U92 ( .A(A[90]), .B(B[0]), .Z(PRODUCT[90]) );
  AND U93 ( .A(A[91]), .B(B[0]), .Z(PRODUCT[91]) );
  AND U94 ( .A(A[92]), .B(B[0]), .Z(PRODUCT[92]) );
  AND U95 ( .A(A[93]), .B(B[0]), .Z(PRODUCT[93]) );
  AND U96 ( .A(A[94]), .B(B[0]), .Z(PRODUCT[94]) );
  AND U97 ( .A(A[95]), .B(B[0]), .Z(PRODUCT[95]) );
  AND U98 ( .A(A[96]), .B(B[0]), .Z(PRODUCT[96]) );
  AND U99 ( .A(A[97]), .B(B[0]), .Z(PRODUCT[97]) );
  AND U100 ( .A(A[98]), .B(B[0]), .Z(PRODUCT[98]) );
  AND U101 ( .A(A[99]), .B(B[0]), .Z(PRODUCT[99]) );
  AND U102 ( .A(A[100]), .B(B[0]), .Z(PRODUCT[100]) );
  AND U103 ( .A(A[101]), .B(B[0]), .Z(PRODUCT[101]) );
  AND U104 ( .A(A[102]), .B(B[0]), .Z(PRODUCT[102]) );
  AND U105 ( .A(A[103]), .B(B[0]), .Z(PRODUCT[103]) );
  AND U106 ( .A(A[104]), .B(B[0]), .Z(PRODUCT[104]) );
  AND U107 ( .A(A[105]), .B(B[0]), .Z(PRODUCT[105]) );
  AND U108 ( .A(A[106]), .B(B[0]), .Z(PRODUCT[106]) );
  AND U109 ( .A(A[107]), .B(B[0]), .Z(PRODUCT[107]) );
  AND U110 ( .A(A[108]), .B(B[0]), .Z(PRODUCT[108]) );
  AND U111 ( .A(A[109]), .B(B[0]), .Z(PRODUCT[109]) );
  AND U112 ( .A(A[110]), .B(B[0]), .Z(PRODUCT[110]) );
  AND U113 ( .A(A[111]), .B(B[0]), .Z(PRODUCT[111]) );
  AND U114 ( .A(A[112]), .B(B[0]), .Z(PRODUCT[112]) );
  AND U115 ( .A(A[113]), .B(B[0]), .Z(PRODUCT[113]) );
  AND U116 ( .A(A[114]), .B(B[0]), .Z(PRODUCT[114]) );
  AND U117 ( .A(A[115]), .B(B[0]), .Z(PRODUCT[115]) );
  AND U118 ( .A(A[116]), .B(B[0]), .Z(PRODUCT[116]) );
  AND U119 ( .A(A[117]), .B(B[0]), .Z(PRODUCT[117]) );
  AND U120 ( .A(A[118]), .B(B[0]), .Z(PRODUCT[118]) );
  AND U121 ( .A(A[119]), .B(B[0]), .Z(PRODUCT[119]) );
  AND U122 ( .A(A[120]), .B(B[0]), .Z(PRODUCT[120]) );
  AND U123 ( .A(A[121]), .B(B[0]), .Z(PRODUCT[121]) );
  AND U124 ( .A(A[122]), .B(B[0]), .Z(PRODUCT[122]) );
  AND U125 ( .A(A[123]), .B(B[0]), .Z(PRODUCT[123]) );
  AND U126 ( .A(A[124]), .B(B[0]), .Z(PRODUCT[124]) );
  AND U127 ( .A(A[125]), .B(B[0]), .Z(PRODUCT[125]) );
  AND U128 ( .A(A[126]), .B(B[0]), .Z(PRODUCT[126]) );
  AND U129 ( .A(A[127]), .B(B[0]), .Z(PRODUCT[127]) );
  AND U130 ( .A(A[128]), .B(B[0]), .Z(PRODUCT[128]) );
  AND U131 ( .A(A[129]), .B(B[0]), .Z(PRODUCT[129]) );
  AND U132 ( .A(A[130]), .B(B[0]), .Z(PRODUCT[130]) );
  AND U133 ( .A(A[131]), .B(B[0]), .Z(PRODUCT[131]) );
  AND U134 ( .A(A[132]), .B(B[0]), .Z(PRODUCT[132]) );
  AND U135 ( .A(A[133]), .B(B[0]), .Z(PRODUCT[133]) );
  AND U136 ( .A(A[134]), .B(B[0]), .Z(PRODUCT[134]) );
  AND U137 ( .A(A[135]), .B(B[0]), .Z(PRODUCT[135]) );
  AND U138 ( .A(A[136]), .B(B[0]), .Z(PRODUCT[136]) );
  AND U139 ( .A(A[137]), .B(B[0]), .Z(PRODUCT[137]) );
  AND U140 ( .A(A[138]), .B(B[0]), .Z(PRODUCT[138]) );
  AND U141 ( .A(A[139]), .B(B[0]), .Z(PRODUCT[139]) );
  AND U142 ( .A(A[140]), .B(B[0]), .Z(PRODUCT[140]) );
  AND U143 ( .A(A[141]), .B(B[0]), .Z(PRODUCT[141]) );
  AND U144 ( .A(A[142]), .B(B[0]), .Z(PRODUCT[142]) );
  AND U145 ( .A(A[143]), .B(B[0]), .Z(PRODUCT[143]) );
  AND U146 ( .A(A[144]), .B(B[0]), .Z(PRODUCT[144]) );
  AND U147 ( .A(A[145]), .B(B[0]), .Z(PRODUCT[145]) );
  AND U148 ( .A(A[146]), .B(B[0]), .Z(PRODUCT[146]) );
  AND U149 ( .A(A[147]), .B(B[0]), .Z(PRODUCT[147]) );
  AND U150 ( .A(A[148]), .B(B[0]), .Z(PRODUCT[148]) );
  AND U151 ( .A(A[149]), .B(B[0]), .Z(PRODUCT[149]) );
  AND U152 ( .A(A[150]), .B(B[0]), .Z(PRODUCT[150]) );
  AND U153 ( .A(A[151]), .B(B[0]), .Z(PRODUCT[151]) );
  AND U154 ( .A(A[152]), .B(B[0]), .Z(PRODUCT[152]) );
  AND U155 ( .A(A[153]), .B(B[0]), .Z(PRODUCT[153]) );
  AND U156 ( .A(A[154]), .B(B[0]), .Z(PRODUCT[154]) );
  AND U157 ( .A(A[155]), .B(B[0]), .Z(PRODUCT[155]) );
  AND U158 ( .A(A[156]), .B(B[0]), .Z(PRODUCT[156]) );
  AND U159 ( .A(A[157]), .B(B[0]), .Z(PRODUCT[157]) );
  AND U160 ( .A(A[158]), .B(B[0]), .Z(PRODUCT[158]) );
  AND U161 ( .A(A[159]), .B(B[0]), .Z(PRODUCT[159]) );
  AND U162 ( .A(A[160]), .B(B[0]), .Z(PRODUCT[160]) );
  AND U163 ( .A(A[161]), .B(B[0]), .Z(PRODUCT[161]) );
  AND U164 ( .A(A[162]), .B(B[0]), .Z(PRODUCT[162]) );
  AND U165 ( .A(A[163]), .B(B[0]), .Z(PRODUCT[163]) );
  AND U166 ( .A(A[164]), .B(B[0]), .Z(PRODUCT[164]) );
  AND U167 ( .A(A[165]), .B(B[0]), .Z(PRODUCT[165]) );
  AND U168 ( .A(A[166]), .B(B[0]), .Z(PRODUCT[166]) );
  AND U169 ( .A(A[167]), .B(B[0]), .Z(PRODUCT[167]) );
  AND U170 ( .A(A[168]), .B(B[0]), .Z(PRODUCT[168]) );
  AND U171 ( .A(A[169]), .B(B[0]), .Z(PRODUCT[169]) );
  AND U172 ( .A(A[170]), .B(B[0]), .Z(PRODUCT[170]) );
  AND U173 ( .A(A[171]), .B(B[0]), .Z(PRODUCT[171]) );
  AND U174 ( .A(A[172]), .B(B[0]), .Z(PRODUCT[172]) );
  AND U175 ( .A(A[173]), .B(B[0]), .Z(PRODUCT[173]) );
  AND U176 ( .A(A[174]), .B(B[0]), .Z(PRODUCT[174]) );
  AND U177 ( .A(A[175]), .B(B[0]), .Z(PRODUCT[175]) );
  AND U178 ( .A(A[176]), .B(B[0]), .Z(PRODUCT[176]) );
  AND U179 ( .A(A[177]), .B(B[0]), .Z(PRODUCT[177]) );
  AND U180 ( .A(A[178]), .B(B[0]), .Z(PRODUCT[178]) );
  AND U181 ( .A(A[179]), .B(B[0]), .Z(PRODUCT[179]) );
  AND U182 ( .A(A[180]), .B(B[0]), .Z(PRODUCT[180]) );
  AND U183 ( .A(A[181]), .B(B[0]), .Z(PRODUCT[181]) );
  AND U184 ( .A(A[182]), .B(B[0]), .Z(PRODUCT[182]) );
  AND U185 ( .A(A[183]), .B(B[0]), .Z(PRODUCT[183]) );
  AND U186 ( .A(A[184]), .B(B[0]), .Z(PRODUCT[184]) );
  AND U187 ( .A(A[185]), .B(B[0]), .Z(PRODUCT[185]) );
  AND U188 ( .A(A[186]), .B(B[0]), .Z(PRODUCT[186]) );
  AND U189 ( .A(A[187]), .B(B[0]), .Z(PRODUCT[187]) );
  AND U190 ( .A(A[188]), .B(B[0]), .Z(PRODUCT[188]) );
  AND U191 ( .A(A[189]), .B(B[0]), .Z(PRODUCT[189]) );
  AND U192 ( .A(A[190]), .B(B[0]), .Z(PRODUCT[190]) );
  AND U193 ( .A(A[191]), .B(B[0]), .Z(PRODUCT[191]) );
  AND U194 ( .A(A[192]), .B(B[0]), .Z(PRODUCT[192]) );
  AND U195 ( .A(A[193]), .B(B[0]), .Z(PRODUCT[193]) );
  AND U196 ( .A(A[194]), .B(B[0]), .Z(PRODUCT[194]) );
  AND U197 ( .A(A[195]), .B(B[0]), .Z(PRODUCT[195]) );
  AND U198 ( .A(A[196]), .B(B[0]), .Z(PRODUCT[196]) );
  AND U199 ( .A(A[197]), .B(B[0]), .Z(PRODUCT[197]) );
  AND U200 ( .A(A[198]), .B(B[0]), .Z(PRODUCT[198]) );
  AND U201 ( .A(A[199]), .B(B[0]), .Z(PRODUCT[199]) );
  AND U202 ( .A(A[200]), .B(B[0]), .Z(PRODUCT[200]) );
  AND U203 ( .A(A[201]), .B(B[0]), .Z(PRODUCT[201]) );
  AND U204 ( .A(A[202]), .B(B[0]), .Z(PRODUCT[202]) );
  AND U205 ( .A(A[203]), .B(B[0]), .Z(PRODUCT[203]) );
  AND U206 ( .A(A[204]), .B(B[0]), .Z(PRODUCT[204]) );
  AND U207 ( .A(A[205]), .B(B[0]), .Z(PRODUCT[205]) );
  AND U208 ( .A(A[206]), .B(B[0]), .Z(PRODUCT[206]) );
  AND U209 ( .A(A[207]), .B(B[0]), .Z(PRODUCT[207]) );
  AND U210 ( .A(A[208]), .B(B[0]), .Z(PRODUCT[208]) );
  AND U211 ( .A(A[209]), .B(B[0]), .Z(PRODUCT[209]) );
  AND U212 ( .A(A[210]), .B(B[0]), .Z(PRODUCT[210]) );
  AND U213 ( .A(A[211]), .B(B[0]), .Z(PRODUCT[211]) );
  AND U214 ( .A(A[212]), .B(B[0]), .Z(PRODUCT[212]) );
  AND U215 ( .A(A[213]), .B(B[0]), .Z(PRODUCT[213]) );
  AND U216 ( .A(A[214]), .B(B[0]), .Z(PRODUCT[214]) );
  AND U217 ( .A(A[215]), .B(B[0]), .Z(PRODUCT[215]) );
  AND U218 ( .A(A[216]), .B(B[0]), .Z(PRODUCT[216]) );
  AND U219 ( .A(A[217]), .B(B[0]), .Z(PRODUCT[217]) );
  AND U220 ( .A(A[218]), .B(B[0]), .Z(PRODUCT[218]) );
  AND U221 ( .A(A[219]), .B(B[0]), .Z(PRODUCT[219]) );
  AND U222 ( .A(A[220]), .B(B[0]), .Z(PRODUCT[220]) );
  AND U223 ( .A(A[221]), .B(B[0]), .Z(PRODUCT[221]) );
  AND U224 ( .A(A[222]), .B(B[0]), .Z(PRODUCT[222]) );
  AND U225 ( .A(A[223]), .B(B[0]), .Z(PRODUCT[223]) );
  AND U226 ( .A(A[224]), .B(B[0]), .Z(PRODUCT[224]) );
  AND U227 ( .A(A[225]), .B(B[0]), .Z(PRODUCT[225]) );
  AND U228 ( .A(A[226]), .B(B[0]), .Z(PRODUCT[226]) );
  AND U229 ( .A(A[227]), .B(B[0]), .Z(PRODUCT[227]) );
  AND U230 ( .A(A[228]), .B(B[0]), .Z(PRODUCT[228]) );
  AND U231 ( .A(A[229]), .B(B[0]), .Z(PRODUCT[229]) );
  AND U232 ( .A(A[230]), .B(B[0]), .Z(PRODUCT[230]) );
  AND U233 ( .A(A[231]), .B(B[0]), .Z(PRODUCT[231]) );
  AND U234 ( .A(A[232]), .B(B[0]), .Z(PRODUCT[232]) );
  AND U235 ( .A(A[233]), .B(B[0]), .Z(PRODUCT[233]) );
  AND U236 ( .A(A[234]), .B(B[0]), .Z(PRODUCT[234]) );
  AND U237 ( .A(A[235]), .B(B[0]), .Z(PRODUCT[235]) );
  AND U238 ( .A(A[236]), .B(B[0]), .Z(PRODUCT[236]) );
  AND U239 ( .A(A[237]), .B(B[0]), .Z(PRODUCT[237]) );
  AND U240 ( .A(A[238]), .B(B[0]), .Z(PRODUCT[238]) );
  AND U241 ( .A(A[239]), .B(B[0]), .Z(PRODUCT[239]) );
  AND U242 ( .A(A[240]), .B(B[0]), .Z(PRODUCT[240]) );
  AND U243 ( .A(A[241]), .B(B[0]), .Z(PRODUCT[241]) );
  AND U244 ( .A(A[242]), .B(B[0]), .Z(PRODUCT[242]) );
  AND U245 ( .A(A[243]), .B(B[0]), .Z(PRODUCT[243]) );
  AND U246 ( .A(A[244]), .B(B[0]), .Z(PRODUCT[244]) );
  AND U247 ( .A(A[245]), .B(B[0]), .Z(PRODUCT[245]) );
  AND U248 ( .A(A[246]), .B(B[0]), .Z(PRODUCT[246]) );
  AND U249 ( .A(A[247]), .B(B[0]), .Z(PRODUCT[247]) );
  AND U250 ( .A(A[248]), .B(B[0]), .Z(PRODUCT[248]) );
  AND U251 ( .A(A[249]), .B(B[0]), .Z(PRODUCT[249]) );
  AND U252 ( .A(A[250]), .B(B[0]), .Z(PRODUCT[250]) );
  AND U253 ( .A(A[251]), .B(B[0]), .Z(PRODUCT[251]) );
  AND U254 ( .A(A[252]), .B(B[0]), .Z(PRODUCT[252]) );
  AND U255 ( .A(A[253]), .B(B[0]), .Z(PRODUCT[253]) );
  AND U256 ( .A(A[254]), .B(B[0]), .Z(PRODUCT[254]) );
  AND U257 ( .A(A[255]), .B(B[0]), .Z(PRODUCT[255]) );
  AND U258 ( .A(A[256]), .B(B[0]), .Z(PRODUCT[256]) );
  AND U259 ( .A(A[257]), .B(B[0]), .Z(PRODUCT[257]) );
  AND U260 ( .A(A[258]), .B(B[0]), .Z(PRODUCT[258]) );
  AND U261 ( .A(A[259]), .B(B[0]), .Z(PRODUCT[259]) );
  AND U262 ( .A(A[260]), .B(B[0]), .Z(PRODUCT[260]) );
  AND U263 ( .A(A[261]), .B(B[0]), .Z(PRODUCT[261]) );
  AND U264 ( .A(A[262]), .B(B[0]), .Z(PRODUCT[262]) );
  AND U265 ( .A(A[263]), .B(B[0]), .Z(PRODUCT[263]) );
  AND U266 ( .A(A[264]), .B(B[0]), .Z(PRODUCT[264]) );
  AND U267 ( .A(A[265]), .B(B[0]), .Z(PRODUCT[265]) );
  AND U268 ( .A(A[266]), .B(B[0]), .Z(PRODUCT[266]) );
  AND U269 ( .A(A[267]), .B(B[0]), .Z(PRODUCT[267]) );
  AND U270 ( .A(A[268]), .B(B[0]), .Z(PRODUCT[268]) );
  AND U271 ( .A(A[269]), .B(B[0]), .Z(PRODUCT[269]) );
  AND U272 ( .A(A[270]), .B(B[0]), .Z(PRODUCT[270]) );
  AND U273 ( .A(A[271]), .B(B[0]), .Z(PRODUCT[271]) );
  AND U274 ( .A(A[272]), .B(B[0]), .Z(PRODUCT[272]) );
  AND U275 ( .A(A[273]), .B(B[0]), .Z(PRODUCT[273]) );
  AND U276 ( .A(A[274]), .B(B[0]), .Z(PRODUCT[274]) );
  AND U277 ( .A(A[275]), .B(B[0]), .Z(PRODUCT[275]) );
  AND U278 ( .A(A[276]), .B(B[0]), .Z(PRODUCT[276]) );
  AND U279 ( .A(A[277]), .B(B[0]), .Z(PRODUCT[277]) );
  AND U280 ( .A(A[278]), .B(B[0]), .Z(PRODUCT[278]) );
  AND U281 ( .A(A[279]), .B(B[0]), .Z(PRODUCT[279]) );
  AND U282 ( .A(A[280]), .B(B[0]), .Z(PRODUCT[280]) );
  AND U283 ( .A(A[281]), .B(B[0]), .Z(PRODUCT[281]) );
  AND U284 ( .A(A[282]), .B(B[0]), .Z(PRODUCT[282]) );
  AND U285 ( .A(A[283]), .B(B[0]), .Z(PRODUCT[283]) );
  AND U286 ( .A(A[284]), .B(B[0]), .Z(PRODUCT[284]) );
  AND U287 ( .A(A[285]), .B(B[0]), .Z(PRODUCT[285]) );
  AND U288 ( .A(A[286]), .B(B[0]), .Z(PRODUCT[286]) );
  AND U289 ( .A(A[287]), .B(B[0]), .Z(PRODUCT[287]) );
  AND U290 ( .A(A[288]), .B(B[0]), .Z(PRODUCT[288]) );
  AND U291 ( .A(A[289]), .B(B[0]), .Z(PRODUCT[289]) );
  AND U292 ( .A(A[290]), .B(B[0]), .Z(PRODUCT[290]) );
  AND U293 ( .A(A[291]), .B(B[0]), .Z(PRODUCT[291]) );
  AND U294 ( .A(A[292]), .B(B[0]), .Z(PRODUCT[292]) );
  AND U295 ( .A(A[293]), .B(B[0]), .Z(PRODUCT[293]) );
  AND U296 ( .A(A[294]), .B(B[0]), .Z(PRODUCT[294]) );
  AND U297 ( .A(A[295]), .B(B[0]), .Z(PRODUCT[295]) );
  AND U298 ( .A(A[296]), .B(B[0]), .Z(PRODUCT[296]) );
  AND U299 ( .A(A[297]), .B(B[0]), .Z(PRODUCT[297]) );
  AND U300 ( .A(A[298]), .B(B[0]), .Z(PRODUCT[298]) );
  AND U301 ( .A(A[299]), .B(B[0]), .Z(PRODUCT[299]) );
  AND U302 ( .A(A[300]), .B(B[0]), .Z(PRODUCT[300]) );
  AND U303 ( .A(A[301]), .B(B[0]), .Z(PRODUCT[301]) );
  AND U304 ( .A(A[302]), .B(B[0]), .Z(PRODUCT[302]) );
  AND U305 ( .A(A[303]), .B(B[0]), .Z(PRODUCT[303]) );
  AND U306 ( .A(A[304]), .B(B[0]), .Z(PRODUCT[304]) );
  AND U307 ( .A(A[305]), .B(B[0]), .Z(PRODUCT[305]) );
  AND U308 ( .A(A[306]), .B(B[0]), .Z(PRODUCT[306]) );
  AND U309 ( .A(A[307]), .B(B[0]), .Z(PRODUCT[307]) );
  AND U310 ( .A(A[308]), .B(B[0]), .Z(PRODUCT[308]) );
  AND U311 ( .A(A[309]), .B(B[0]), .Z(PRODUCT[309]) );
  AND U312 ( .A(A[310]), .B(B[0]), .Z(PRODUCT[310]) );
  AND U313 ( .A(A[311]), .B(B[0]), .Z(PRODUCT[311]) );
  AND U314 ( .A(A[312]), .B(B[0]), .Z(PRODUCT[312]) );
  AND U315 ( .A(A[313]), .B(B[0]), .Z(PRODUCT[313]) );
  AND U316 ( .A(A[314]), .B(B[0]), .Z(PRODUCT[314]) );
  AND U317 ( .A(A[315]), .B(B[0]), .Z(PRODUCT[315]) );
  AND U318 ( .A(A[316]), .B(B[0]), .Z(PRODUCT[316]) );
  AND U319 ( .A(A[317]), .B(B[0]), .Z(PRODUCT[317]) );
  AND U320 ( .A(A[318]), .B(B[0]), .Z(PRODUCT[318]) );
  AND U321 ( .A(A[319]), .B(B[0]), .Z(PRODUCT[319]) );
  AND U322 ( .A(A[320]), .B(B[0]), .Z(PRODUCT[320]) );
  AND U323 ( .A(A[321]), .B(B[0]), .Z(PRODUCT[321]) );
  AND U324 ( .A(A[322]), .B(B[0]), .Z(PRODUCT[322]) );
  AND U325 ( .A(A[323]), .B(B[0]), .Z(PRODUCT[323]) );
  AND U326 ( .A(A[324]), .B(B[0]), .Z(PRODUCT[324]) );
  AND U327 ( .A(A[325]), .B(B[0]), .Z(PRODUCT[325]) );
  AND U328 ( .A(A[326]), .B(B[0]), .Z(PRODUCT[326]) );
  AND U329 ( .A(A[327]), .B(B[0]), .Z(PRODUCT[327]) );
  AND U330 ( .A(A[328]), .B(B[0]), .Z(PRODUCT[328]) );
  AND U331 ( .A(A[329]), .B(B[0]), .Z(PRODUCT[329]) );
  AND U332 ( .A(A[330]), .B(B[0]), .Z(PRODUCT[330]) );
  AND U333 ( .A(A[331]), .B(B[0]), .Z(PRODUCT[331]) );
  AND U334 ( .A(A[332]), .B(B[0]), .Z(PRODUCT[332]) );
  AND U335 ( .A(A[333]), .B(B[0]), .Z(PRODUCT[333]) );
  AND U336 ( .A(A[334]), .B(B[0]), .Z(PRODUCT[334]) );
  AND U337 ( .A(A[335]), .B(B[0]), .Z(PRODUCT[335]) );
  AND U338 ( .A(A[336]), .B(B[0]), .Z(PRODUCT[336]) );
  AND U339 ( .A(A[337]), .B(B[0]), .Z(PRODUCT[337]) );
  AND U340 ( .A(A[338]), .B(B[0]), .Z(PRODUCT[338]) );
  AND U341 ( .A(A[339]), .B(B[0]), .Z(PRODUCT[339]) );
  AND U342 ( .A(A[340]), .B(B[0]), .Z(PRODUCT[340]) );
  AND U343 ( .A(A[341]), .B(B[0]), .Z(PRODUCT[341]) );
  AND U344 ( .A(A[342]), .B(B[0]), .Z(PRODUCT[342]) );
  AND U345 ( .A(A[343]), .B(B[0]), .Z(PRODUCT[343]) );
  AND U346 ( .A(A[344]), .B(B[0]), .Z(PRODUCT[344]) );
  AND U347 ( .A(A[345]), .B(B[0]), .Z(PRODUCT[345]) );
  AND U348 ( .A(A[346]), .B(B[0]), .Z(PRODUCT[346]) );
  AND U349 ( .A(A[347]), .B(B[0]), .Z(PRODUCT[347]) );
  AND U350 ( .A(A[348]), .B(B[0]), .Z(PRODUCT[348]) );
  AND U351 ( .A(A[349]), .B(B[0]), .Z(PRODUCT[349]) );
  AND U352 ( .A(A[350]), .B(B[0]), .Z(PRODUCT[350]) );
  AND U353 ( .A(A[351]), .B(B[0]), .Z(PRODUCT[351]) );
  AND U354 ( .A(A[352]), .B(B[0]), .Z(PRODUCT[352]) );
  AND U355 ( .A(A[353]), .B(B[0]), .Z(PRODUCT[353]) );
  AND U356 ( .A(A[354]), .B(B[0]), .Z(PRODUCT[354]) );
  AND U357 ( .A(A[355]), .B(B[0]), .Z(PRODUCT[355]) );
  AND U358 ( .A(A[356]), .B(B[0]), .Z(PRODUCT[356]) );
  AND U359 ( .A(A[357]), .B(B[0]), .Z(PRODUCT[357]) );
  AND U360 ( .A(A[358]), .B(B[0]), .Z(PRODUCT[358]) );
  AND U361 ( .A(A[359]), .B(B[0]), .Z(PRODUCT[359]) );
  AND U362 ( .A(A[360]), .B(B[0]), .Z(PRODUCT[360]) );
  AND U363 ( .A(A[361]), .B(B[0]), .Z(PRODUCT[361]) );
  AND U364 ( .A(A[362]), .B(B[0]), .Z(PRODUCT[362]) );
  AND U365 ( .A(A[363]), .B(B[0]), .Z(PRODUCT[363]) );
  AND U366 ( .A(A[364]), .B(B[0]), .Z(PRODUCT[364]) );
  AND U367 ( .A(A[365]), .B(B[0]), .Z(PRODUCT[365]) );
  AND U368 ( .A(A[366]), .B(B[0]), .Z(PRODUCT[366]) );
  AND U369 ( .A(A[367]), .B(B[0]), .Z(PRODUCT[367]) );
  AND U370 ( .A(A[368]), .B(B[0]), .Z(PRODUCT[368]) );
  AND U371 ( .A(A[369]), .B(B[0]), .Z(PRODUCT[369]) );
  AND U372 ( .A(A[370]), .B(B[0]), .Z(PRODUCT[370]) );
  AND U373 ( .A(A[371]), .B(B[0]), .Z(PRODUCT[371]) );
  AND U374 ( .A(A[372]), .B(B[0]), .Z(PRODUCT[372]) );
  AND U375 ( .A(A[373]), .B(B[0]), .Z(PRODUCT[373]) );
  AND U376 ( .A(A[374]), .B(B[0]), .Z(PRODUCT[374]) );
  AND U377 ( .A(A[375]), .B(B[0]), .Z(PRODUCT[375]) );
  AND U378 ( .A(A[376]), .B(B[0]), .Z(PRODUCT[376]) );
  AND U379 ( .A(A[377]), .B(B[0]), .Z(PRODUCT[377]) );
  AND U380 ( .A(A[378]), .B(B[0]), .Z(PRODUCT[378]) );
  AND U381 ( .A(A[379]), .B(B[0]), .Z(PRODUCT[379]) );
  AND U382 ( .A(A[380]), .B(B[0]), .Z(PRODUCT[380]) );
  AND U383 ( .A(A[381]), .B(B[0]), .Z(PRODUCT[381]) );
  AND U384 ( .A(A[382]), .B(B[0]), .Z(PRODUCT[382]) );
  AND U385 ( .A(A[383]), .B(B[0]), .Z(PRODUCT[383]) );
  AND U386 ( .A(A[384]), .B(B[0]), .Z(PRODUCT[384]) );
  AND U387 ( .A(A[385]), .B(B[0]), .Z(PRODUCT[385]) );
  AND U388 ( .A(A[386]), .B(B[0]), .Z(PRODUCT[386]) );
  AND U389 ( .A(A[387]), .B(B[0]), .Z(PRODUCT[387]) );
  AND U390 ( .A(A[388]), .B(B[0]), .Z(PRODUCT[388]) );
  AND U391 ( .A(A[389]), .B(B[0]), .Z(PRODUCT[389]) );
  AND U392 ( .A(A[390]), .B(B[0]), .Z(PRODUCT[390]) );
  AND U393 ( .A(A[391]), .B(B[0]), .Z(PRODUCT[391]) );
  AND U394 ( .A(A[392]), .B(B[0]), .Z(PRODUCT[392]) );
  AND U395 ( .A(A[393]), .B(B[0]), .Z(PRODUCT[393]) );
  AND U396 ( .A(A[394]), .B(B[0]), .Z(PRODUCT[394]) );
  AND U397 ( .A(A[395]), .B(B[0]), .Z(PRODUCT[395]) );
  AND U398 ( .A(A[396]), .B(B[0]), .Z(PRODUCT[396]) );
  AND U399 ( .A(A[397]), .B(B[0]), .Z(PRODUCT[397]) );
  AND U400 ( .A(A[398]), .B(B[0]), .Z(PRODUCT[398]) );
  AND U401 ( .A(A[399]), .B(B[0]), .Z(PRODUCT[399]) );
  AND U402 ( .A(A[400]), .B(B[0]), .Z(PRODUCT[400]) );
  AND U403 ( .A(A[401]), .B(B[0]), .Z(PRODUCT[401]) );
  AND U404 ( .A(A[402]), .B(B[0]), .Z(PRODUCT[402]) );
  AND U405 ( .A(A[403]), .B(B[0]), .Z(PRODUCT[403]) );
  AND U406 ( .A(A[404]), .B(B[0]), .Z(PRODUCT[404]) );
  AND U407 ( .A(A[405]), .B(B[0]), .Z(PRODUCT[405]) );
  AND U408 ( .A(A[406]), .B(B[0]), .Z(PRODUCT[406]) );
  AND U409 ( .A(A[407]), .B(B[0]), .Z(PRODUCT[407]) );
  AND U410 ( .A(A[408]), .B(B[0]), .Z(PRODUCT[408]) );
  AND U411 ( .A(A[409]), .B(B[0]), .Z(PRODUCT[409]) );
  AND U412 ( .A(A[410]), .B(B[0]), .Z(PRODUCT[410]) );
  AND U413 ( .A(A[411]), .B(B[0]), .Z(PRODUCT[411]) );
  AND U414 ( .A(A[412]), .B(B[0]), .Z(PRODUCT[412]) );
  AND U415 ( .A(A[413]), .B(B[0]), .Z(PRODUCT[413]) );
  AND U416 ( .A(A[414]), .B(B[0]), .Z(PRODUCT[414]) );
  AND U417 ( .A(A[415]), .B(B[0]), .Z(PRODUCT[415]) );
  AND U418 ( .A(A[416]), .B(B[0]), .Z(PRODUCT[416]) );
  AND U419 ( .A(A[417]), .B(B[0]), .Z(PRODUCT[417]) );
  AND U420 ( .A(A[418]), .B(B[0]), .Z(PRODUCT[418]) );
  AND U421 ( .A(A[419]), .B(B[0]), .Z(PRODUCT[419]) );
  AND U422 ( .A(A[420]), .B(B[0]), .Z(PRODUCT[420]) );
  AND U423 ( .A(A[421]), .B(B[0]), .Z(PRODUCT[421]) );
  AND U424 ( .A(A[422]), .B(B[0]), .Z(PRODUCT[422]) );
  AND U425 ( .A(A[423]), .B(B[0]), .Z(PRODUCT[423]) );
  AND U426 ( .A(A[424]), .B(B[0]), .Z(PRODUCT[424]) );
  AND U427 ( .A(A[425]), .B(B[0]), .Z(PRODUCT[425]) );
  AND U428 ( .A(A[426]), .B(B[0]), .Z(PRODUCT[426]) );
  AND U429 ( .A(A[427]), .B(B[0]), .Z(PRODUCT[427]) );
  AND U430 ( .A(A[428]), .B(B[0]), .Z(PRODUCT[428]) );
  AND U431 ( .A(A[429]), .B(B[0]), .Z(PRODUCT[429]) );
  AND U432 ( .A(A[430]), .B(B[0]), .Z(PRODUCT[430]) );
  AND U433 ( .A(A[431]), .B(B[0]), .Z(PRODUCT[431]) );
  AND U434 ( .A(A[432]), .B(B[0]), .Z(PRODUCT[432]) );
  AND U435 ( .A(A[433]), .B(B[0]), .Z(PRODUCT[433]) );
  AND U436 ( .A(A[434]), .B(B[0]), .Z(PRODUCT[434]) );
  AND U437 ( .A(A[435]), .B(B[0]), .Z(PRODUCT[435]) );
  AND U438 ( .A(A[436]), .B(B[0]), .Z(PRODUCT[436]) );
  AND U439 ( .A(A[437]), .B(B[0]), .Z(PRODUCT[437]) );
  AND U440 ( .A(A[438]), .B(B[0]), .Z(PRODUCT[438]) );
  AND U441 ( .A(A[439]), .B(B[0]), .Z(PRODUCT[439]) );
  AND U442 ( .A(A[440]), .B(B[0]), .Z(PRODUCT[440]) );
  AND U443 ( .A(A[441]), .B(B[0]), .Z(PRODUCT[441]) );
  AND U444 ( .A(A[442]), .B(B[0]), .Z(PRODUCT[442]) );
  AND U445 ( .A(A[443]), .B(B[0]), .Z(PRODUCT[443]) );
  AND U446 ( .A(A[444]), .B(B[0]), .Z(PRODUCT[444]) );
  AND U447 ( .A(A[445]), .B(B[0]), .Z(PRODUCT[445]) );
  AND U448 ( .A(A[446]), .B(B[0]), .Z(PRODUCT[446]) );
  AND U449 ( .A(A[447]), .B(B[0]), .Z(PRODUCT[447]) );
  AND U450 ( .A(A[448]), .B(B[0]), .Z(PRODUCT[448]) );
  AND U451 ( .A(A[449]), .B(B[0]), .Z(PRODUCT[449]) );
  AND U452 ( .A(A[450]), .B(B[0]), .Z(PRODUCT[450]) );
  AND U453 ( .A(A[451]), .B(B[0]), .Z(PRODUCT[451]) );
  AND U454 ( .A(A[452]), .B(B[0]), .Z(PRODUCT[452]) );
  AND U455 ( .A(A[453]), .B(B[0]), .Z(PRODUCT[453]) );
  AND U456 ( .A(A[454]), .B(B[0]), .Z(PRODUCT[454]) );
  AND U457 ( .A(A[455]), .B(B[0]), .Z(PRODUCT[455]) );
  AND U458 ( .A(A[456]), .B(B[0]), .Z(PRODUCT[456]) );
  AND U459 ( .A(A[457]), .B(B[0]), .Z(PRODUCT[457]) );
  AND U460 ( .A(A[458]), .B(B[0]), .Z(PRODUCT[458]) );
  AND U461 ( .A(A[459]), .B(B[0]), .Z(PRODUCT[459]) );
  AND U462 ( .A(A[460]), .B(B[0]), .Z(PRODUCT[460]) );
  AND U463 ( .A(A[461]), .B(B[0]), .Z(PRODUCT[461]) );
  AND U464 ( .A(A[462]), .B(B[0]), .Z(PRODUCT[462]) );
  AND U465 ( .A(A[463]), .B(B[0]), .Z(PRODUCT[463]) );
  AND U466 ( .A(A[464]), .B(B[0]), .Z(PRODUCT[464]) );
  AND U467 ( .A(A[465]), .B(B[0]), .Z(PRODUCT[465]) );
  AND U468 ( .A(A[466]), .B(B[0]), .Z(PRODUCT[466]) );
  AND U469 ( .A(A[467]), .B(B[0]), .Z(PRODUCT[467]) );
  AND U470 ( .A(A[468]), .B(B[0]), .Z(PRODUCT[468]) );
  AND U471 ( .A(A[469]), .B(B[0]), .Z(PRODUCT[469]) );
  AND U472 ( .A(A[470]), .B(B[0]), .Z(PRODUCT[470]) );
  AND U473 ( .A(A[471]), .B(B[0]), .Z(PRODUCT[471]) );
  AND U474 ( .A(A[472]), .B(B[0]), .Z(PRODUCT[472]) );
  AND U475 ( .A(A[473]), .B(B[0]), .Z(PRODUCT[473]) );
  AND U476 ( .A(A[474]), .B(B[0]), .Z(PRODUCT[474]) );
  AND U477 ( .A(A[475]), .B(B[0]), .Z(PRODUCT[475]) );
  AND U478 ( .A(A[476]), .B(B[0]), .Z(PRODUCT[476]) );
  AND U479 ( .A(A[477]), .B(B[0]), .Z(PRODUCT[477]) );
  AND U480 ( .A(A[478]), .B(B[0]), .Z(PRODUCT[478]) );
  AND U481 ( .A(A[479]), .B(B[0]), .Z(PRODUCT[479]) );
  AND U482 ( .A(A[480]), .B(B[0]), .Z(PRODUCT[480]) );
  AND U483 ( .A(A[481]), .B(B[0]), .Z(PRODUCT[481]) );
  AND U484 ( .A(A[482]), .B(B[0]), .Z(PRODUCT[482]) );
  AND U485 ( .A(A[483]), .B(B[0]), .Z(PRODUCT[483]) );
  AND U486 ( .A(A[484]), .B(B[0]), .Z(PRODUCT[484]) );
  AND U487 ( .A(A[485]), .B(B[0]), .Z(PRODUCT[485]) );
  AND U488 ( .A(A[486]), .B(B[0]), .Z(PRODUCT[486]) );
  AND U489 ( .A(A[487]), .B(B[0]), .Z(PRODUCT[487]) );
  AND U490 ( .A(A[488]), .B(B[0]), .Z(PRODUCT[488]) );
  AND U491 ( .A(A[489]), .B(B[0]), .Z(PRODUCT[489]) );
  AND U492 ( .A(A[490]), .B(B[0]), .Z(PRODUCT[490]) );
  AND U493 ( .A(A[491]), .B(B[0]), .Z(PRODUCT[491]) );
  AND U494 ( .A(A[492]), .B(B[0]), .Z(PRODUCT[492]) );
  AND U495 ( .A(A[493]), .B(B[0]), .Z(PRODUCT[493]) );
  AND U496 ( .A(A[494]), .B(B[0]), .Z(PRODUCT[494]) );
  AND U497 ( .A(A[495]), .B(B[0]), .Z(PRODUCT[495]) );
  AND U498 ( .A(A[496]), .B(B[0]), .Z(PRODUCT[496]) );
  AND U499 ( .A(A[497]), .B(B[0]), .Z(PRODUCT[497]) );
  AND U500 ( .A(A[498]), .B(B[0]), .Z(PRODUCT[498]) );
  AND U501 ( .A(A[499]), .B(B[0]), .Z(PRODUCT[499]) );
  AND U502 ( .A(A[500]), .B(B[0]), .Z(PRODUCT[500]) );
  AND U503 ( .A(A[501]), .B(B[0]), .Z(PRODUCT[501]) );
  AND U504 ( .A(A[502]), .B(B[0]), .Z(PRODUCT[502]) );
  AND U505 ( .A(A[503]), .B(B[0]), .Z(PRODUCT[503]) );
  AND U506 ( .A(A[504]), .B(B[0]), .Z(PRODUCT[504]) );
  AND U507 ( .A(A[505]), .B(B[0]), .Z(PRODUCT[505]) );
  AND U508 ( .A(A[506]), .B(B[0]), .Z(PRODUCT[506]) );
  AND U509 ( .A(A[507]), .B(B[0]), .Z(PRODUCT[507]) );
  AND U510 ( .A(A[508]), .B(B[0]), .Z(PRODUCT[508]) );
  AND U511 ( .A(A[509]), .B(B[0]), .Z(PRODUCT[509]) );
  AND U512 ( .A(A[510]), .B(B[0]), .Z(PRODUCT[510]) );
  AND U513 ( .A(A[511]), .B(B[0]), .Z(PRODUCT[511]) );
  AND U514 ( .A(A[512]), .B(B[0]), .Z(PRODUCT[512]) );
  AND U515 ( .A(A[513]), .B(B[0]), .Z(PRODUCT[513]) );
  AND U516 ( .A(A[514]), .B(B[0]), .Z(PRODUCT[514]) );
  AND U517 ( .A(A[515]), .B(B[0]), .Z(PRODUCT[515]) );
  AND U518 ( .A(A[516]), .B(B[0]), .Z(PRODUCT[516]) );
  AND U519 ( .A(A[517]), .B(B[0]), .Z(PRODUCT[517]) );
  AND U520 ( .A(A[518]), .B(B[0]), .Z(PRODUCT[518]) );
  AND U521 ( .A(A[519]), .B(B[0]), .Z(PRODUCT[519]) );
  AND U522 ( .A(A[520]), .B(B[0]), .Z(PRODUCT[520]) );
  AND U523 ( .A(A[521]), .B(B[0]), .Z(PRODUCT[521]) );
  AND U524 ( .A(A[522]), .B(B[0]), .Z(PRODUCT[522]) );
  AND U525 ( .A(A[523]), .B(B[0]), .Z(PRODUCT[523]) );
  AND U526 ( .A(A[524]), .B(B[0]), .Z(PRODUCT[524]) );
  AND U527 ( .A(A[525]), .B(B[0]), .Z(PRODUCT[525]) );
  AND U528 ( .A(A[526]), .B(B[0]), .Z(PRODUCT[526]) );
  AND U529 ( .A(A[527]), .B(B[0]), .Z(PRODUCT[527]) );
  AND U530 ( .A(A[528]), .B(B[0]), .Z(PRODUCT[528]) );
  AND U531 ( .A(A[529]), .B(B[0]), .Z(PRODUCT[529]) );
  AND U532 ( .A(A[530]), .B(B[0]), .Z(PRODUCT[530]) );
  AND U533 ( .A(A[531]), .B(B[0]), .Z(PRODUCT[531]) );
  AND U534 ( .A(A[532]), .B(B[0]), .Z(PRODUCT[532]) );
  AND U535 ( .A(A[533]), .B(B[0]), .Z(PRODUCT[533]) );
  AND U536 ( .A(A[534]), .B(B[0]), .Z(PRODUCT[534]) );
  AND U537 ( .A(A[535]), .B(B[0]), .Z(PRODUCT[535]) );
  AND U538 ( .A(A[536]), .B(B[0]), .Z(PRODUCT[536]) );
  AND U539 ( .A(A[537]), .B(B[0]), .Z(PRODUCT[537]) );
  AND U540 ( .A(A[538]), .B(B[0]), .Z(PRODUCT[538]) );
  AND U541 ( .A(A[539]), .B(B[0]), .Z(PRODUCT[539]) );
  AND U542 ( .A(A[540]), .B(B[0]), .Z(PRODUCT[540]) );
  AND U543 ( .A(A[541]), .B(B[0]), .Z(PRODUCT[541]) );
  AND U544 ( .A(A[542]), .B(B[0]), .Z(PRODUCT[542]) );
  AND U545 ( .A(A[543]), .B(B[0]), .Z(PRODUCT[543]) );
  AND U546 ( .A(A[544]), .B(B[0]), .Z(PRODUCT[544]) );
  AND U547 ( .A(A[545]), .B(B[0]), .Z(PRODUCT[545]) );
  AND U548 ( .A(A[546]), .B(B[0]), .Z(PRODUCT[546]) );
  AND U549 ( .A(A[547]), .B(B[0]), .Z(PRODUCT[547]) );
  AND U550 ( .A(A[548]), .B(B[0]), .Z(PRODUCT[548]) );
  AND U551 ( .A(A[549]), .B(B[0]), .Z(PRODUCT[549]) );
  AND U552 ( .A(A[550]), .B(B[0]), .Z(PRODUCT[550]) );
  AND U553 ( .A(A[551]), .B(B[0]), .Z(PRODUCT[551]) );
  AND U554 ( .A(A[552]), .B(B[0]), .Z(PRODUCT[552]) );
  AND U555 ( .A(A[553]), .B(B[0]), .Z(PRODUCT[553]) );
  AND U556 ( .A(A[554]), .B(B[0]), .Z(PRODUCT[554]) );
  AND U557 ( .A(A[555]), .B(B[0]), .Z(PRODUCT[555]) );
  AND U558 ( .A(A[556]), .B(B[0]), .Z(PRODUCT[556]) );
  AND U559 ( .A(A[557]), .B(B[0]), .Z(PRODUCT[557]) );
  AND U560 ( .A(A[558]), .B(B[0]), .Z(PRODUCT[558]) );
  AND U561 ( .A(A[559]), .B(B[0]), .Z(PRODUCT[559]) );
  AND U562 ( .A(A[560]), .B(B[0]), .Z(PRODUCT[560]) );
  AND U563 ( .A(A[561]), .B(B[0]), .Z(PRODUCT[561]) );
  AND U564 ( .A(A[562]), .B(B[0]), .Z(PRODUCT[562]) );
  AND U565 ( .A(A[563]), .B(B[0]), .Z(PRODUCT[563]) );
  AND U566 ( .A(A[564]), .B(B[0]), .Z(PRODUCT[564]) );
  AND U567 ( .A(A[565]), .B(B[0]), .Z(PRODUCT[565]) );
  AND U568 ( .A(A[566]), .B(B[0]), .Z(PRODUCT[566]) );
  AND U569 ( .A(A[567]), .B(B[0]), .Z(PRODUCT[567]) );
  AND U570 ( .A(A[568]), .B(B[0]), .Z(PRODUCT[568]) );
  AND U571 ( .A(A[569]), .B(B[0]), .Z(PRODUCT[569]) );
  AND U572 ( .A(A[570]), .B(B[0]), .Z(PRODUCT[570]) );
  AND U573 ( .A(A[571]), .B(B[0]), .Z(PRODUCT[571]) );
  AND U574 ( .A(A[572]), .B(B[0]), .Z(PRODUCT[572]) );
  AND U575 ( .A(A[573]), .B(B[0]), .Z(PRODUCT[573]) );
  AND U576 ( .A(A[574]), .B(B[0]), .Z(PRODUCT[574]) );
  AND U577 ( .A(A[575]), .B(B[0]), .Z(PRODUCT[575]) );
  AND U578 ( .A(A[576]), .B(B[0]), .Z(PRODUCT[576]) );
  AND U579 ( .A(A[577]), .B(B[0]), .Z(PRODUCT[577]) );
  AND U580 ( .A(A[578]), .B(B[0]), .Z(PRODUCT[578]) );
  AND U581 ( .A(A[579]), .B(B[0]), .Z(PRODUCT[579]) );
  AND U582 ( .A(A[580]), .B(B[0]), .Z(PRODUCT[580]) );
  AND U583 ( .A(A[581]), .B(B[0]), .Z(PRODUCT[581]) );
  AND U584 ( .A(A[582]), .B(B[0]), .Z(PRODUCT[582]) );
  AND U585 ( .A(A[583]), .B(B[0]), .Z(PRODUCT[583]) );
  AND U586 ( .A(A[584]), .B(B[0]), .Z(PRODUCT[584]) );
  AND U587 ( .A(A[585]), .B(B[0]), .Z(PRODUCT[585]) );
  AND U588 ( .A(A[586]), .B(B[0]), .Z(PRODUCT[586]) );
  AND U589 ( .A(A[587]), .B(B[0]), .Z(PRODUCT[587]) );
  AND U590 ( .A(A[588]), .B(B[0]), .Z(PRODUCT[588]) );
  AND U591 ( .A(A[589]), .B(B[0]), .Z(PRODUCT[589]) );
  AND U592 ( .A(A[590]), .B(B[0]), .Z(PRODUCT[590]) );
  AND U593 ( .A(A[591]), .B(B[0]), .Z(PRODUCT[591]) );
  AND U594 ( .A(A[592]), .B(B[0]), .Z(PRODUCT[592]) );
  AND U595 ( .A(A[593]), .B(B[0]), .Z(PRODUCT[593]) );
  AND U596 ( .A(A[594]), .B(B[0]), .Z(PRODUCT[594]) );
  AND U597 ( .A(A[595]), .B(B[0]), .Z(PRODUCT[595]) );
  AND U598 ( .A(A[596]), .B(B[0]), .Z(PRODUCT[596]) );
  AND U599 ( .A(A[597]), .B(B[0]), .Z(PRODUCT[597]) );
  AND U600 ( .A(A[598]), .B(B[0]), .Z(PRODUCT[598]) );
  AND U601 ( .A(A[599]), .B(B[0]), .Z(PRODUCT[599]) );
  AND U602 ( .A(A[600]), .B(B[0]), .Z(PRODUCT[600]) );
  AND U603 ( .A(A[601]), .B(B[0]), .Z(PRODUCT[601]) );
  AND U604 ( .A(A[602]), .B(B[0]), .Z(PRODUCT[602]) );
  AND U605 ( .A(A[603]), .B(B[0]), .Z(PRODUCT[603]) );
  AND U606 ( .A(A[604]), .B(B[0]), .Z(PRODUCT[604]) );
  AND U607 ( .A(A[605]), .B(B[0]), .Z(PRODUCT[605]) );
  AND U608 ( .A(A[606]), .B(B[0]), .Z(PRODUCT[606]) );
  AND U609 ( .A(A[607]), .B(B[0]), .Z(PRODUCT[607]) );
  AND U610 ( .A(A[608]), .B(B[0]), .Z(PRODUCT[608]) );
  AND U611 ( .A(A[609]), .B(B[0]), .Z(PRODUCT[609]) );
  AND U612 ( .A(A[610]), .B(B[0]), .Z(PRODUCT[610]) );
  AND U613 ( .A(A[611]), .B(B[0]), .Z(PRODUCT[611]) );
  AND U614 ( .A(A[612]), .B(B[0]), .Z(PRODUCT[612]) );
  AND U615 ( .A(A[613]), .B(B[0]), .Z(PRODUCT[613]) );
  AND U616 ( .A(A[614]), .B(B[0]), .Z(PRODUCT[614]) );
  AND U617 ( .A(A[615]), .B(B[0]), .Z(PRODUCT[615]) );
  AND U618 ( .A(A[616]), .B(B[0]), .Z(PRODUCT[616]) );
  AND U619 ( .A(A[617]), .B(B[0]), .Z(PRODUCT[617]) );
  AND U620 ( .A(A[618]), .B(B[0]), .Z(PRODUCT[618]) );
  AND U621 ( .A(A[619]), .B(B[0]), .Z(PRODUCT[619]) );
  AND U622 ( .A(A[620]), .B(B[0]), .Z(PRODUCT[620]) );
  AND U623 ( .A(A[621]), .B(B[0]), .Z(PRODUCT[621]) );
  AND U624 ( .A(A[622]), .B(B[0]), .Z(PRODUCT[622]) );
  AND U625 ( .A(A[623]), .B(B[0]), .Z(PRODUCT[623]) );
  AND U626 ( .A(A[624]), .B(B[0]), .Z(PRODUCT[624]) );
  AND U627 ( .A(A[625]), .B(B[0]), .Z(PRODUCT[625]) );
  AND U628 ( .A(A[626]), .B(B[0]), .Z(PRODUCT[626]) );
  AND U629 ( .A(A[627]), .B(B[0]), .Z(PRODUCT[627]) );
  AND U630 ( .A(A[628]), .B(B[0]), .Z(PRODUCT[628]) );
  AND U631 ( .A(A[629]), .B(B[0]), .Z(PRODUCT[629]) );
  AND U632 ( .A(A[630]), .B(B[0]), .Z(PRODUCT[630]) );
  AND U633 ( .A(A[631]), .B(B[0]), .Z(PRODUCT[631]) );
  AND U634 ( .A(A[632]), .B(B[0]), .Z(PRODUCT[632]) );
  AND U635 ( .A(A[633]), .B(B[0]), .Z(PRODUCT[633]) );
  AND U636 ( .A(A[634]), .B(B[0]), .Z(PRODUCT[634]) );
  AND U637 ( .A(A[635]), .B(B[0]), .Z(PRODUCT[635]) );
  AND U638 ( .A(A[636]), .B(B[0]), .Z(PRODUCT[636]) );
  AND U639 ( .A(A[637]), .B(B[0]), .Z(PRODUCT[637]) );
  AND U640 ( .A(A[638]), .B(B[0]), .Z(PRODUCT[638]) );
  AND U641 ( .A(A[639]), .B(B[0]), .Z(PRODUCT[639]) );
  AND U642 ( .A(A[640]), .B(B[0]), .Z(PRODUCT[640]) );
  AND U643 ( .A(A[641]), .B(B[0]), .Z(PRODUCT[641]) );
  AND U644 ( .A(A[642]), .B(B[0]), .Z(PRODUCT[642]) );
  AND U645 ( .A(A[643]), .B(B[0]), .Z(PRODUCT[643]) );
  AND U646 ( .A(A[644]), .B(B[0]), .Z(PRODUCT[644]) );
  AND U647 ( .A(A[645]), .B(B[0]), .Z(PRODUCT[645]) );
  AND U648 ( .A(A[646]), .B(B[0]), .Z(PRODUCT[646]) );
  AND U649 ( .A(A[647]), .B(B[0]), .Z(PRODUCT[647]) );
  AND U650 ( .A(A[648]), .B(B[0]), .Z(PRODUCT[648]) );
  AND U651 ( .A(A[649]), .B(B[0]), .Z(PRODUCT[649]) );
  AND U652 ( .A(A[650]), .B(B[0]), .Z(PRODUCT[650]) );
  AND U653 ( .A(A[651]), .B(B[0]), .Z(PRODUCT[651]) );
  AND U654 ( .A(A[652]), .B(B[0]), .Z(PRODUCT[652]) );
  AND U655 ( .A(A[653]), .B(B[0]), .Z(PRODUCT[653]) );
  AND U656 ( .A(A[654]), .B(B[0]), .Z(PRODUCT[654]) );
  AND U657 ( .A(A[655]), .B(B[0]), .Z(PRODUCT[655]) );
  AND U658 ( .A(A[656]), .B(B[0]), .Z(PRODUCT[656]) );
  AND U659 ( .A(A[657]), .B(B[0]), .Z(PRODUCT[657]) );
  AND U660 ( .A(A[658]), .B(B[0]), .Z(PRODUCT[658]) );
  AND U661 ( .A(A[659]), .B(B[0]), .Z(PRODUCT[659]) );
  AND U662 ( .A(A[660]), .B(B[0]), .Z(PRODUCT[660]) );
  AND U663 ( .A(A[661]), .B(B[0]), .Z(PRODUCT[661]) );
  AND U664 ( .A(A[662]), .B(B[0]), .Z(PRODUCT[662]) );
  AND U665 ( .A(A[663]), .B(B[0]), .Z(PRODUCT[663]) );
  AND U666 ( .A(A[664]), .B(B[0]), .Z(PRODUCT[664]) );
  AND U667 ( .A(A[665]), .B(B[0]), .Z(PRODUCT[665]) );
  AND U668 ( .A(A[666]), .B(B[0]), .Z(PRODUCT[666]) );
  AND U669 ( .A(A[667]), .B(B[0]), .Z(PRODUCT[667]) );
  AND U670 ( .A(A[668]), .B(B[0]), .Z(PRODUCT[668]) );
  AND U671 ( .A(A[669]), .B(B[0]), .Z(PRODUCT[669]) );
  AND U672 ( .A(A[670]), .B(B[0]), .Z(PRODUCT[670]) );
  AND U673 ( .A(A[671]), .B(B[0]), .Z(PRODUCT[671]) );
  AND U674 ( .A(A[672]), .B(B[0]), .Z(PRODUCT[672]) );
  AND U675 ( .A(A[673]), .B(B[0]), .Z(PRODUCT[673]) );
  AND U676 ( .A(A[674]), .B(B[0]), .Z(PRODUCT[674]) );
  AND U677 ( .A(A[675]), .B(B[0]), .Z(PRODUCT[675]) );
  AND U678 ( .A(A[676]), .B(B[0]), .Z(PRODUCT[676]) );
  AND U679 ( .A(A[677]), .B(B[0]), .Z(PRODUCT[677]) );
  AND U680 ( .A(A[678]), .B(B[0]), .Z(PRODUCT[678]) );
  AND U681 ( .A(A[679]), .B(B[0]), .Z(PRODUCT[679]) );
  AND U682 ( .A(A[680]), .B(B[0]), .Z(PRODUCT[680]) );
  AND U683 ( .A(A[681]), .B(B[0]), .Z(PRODUCT[681]) );
  AND U684 ( .A(A[682]), .B(B[0]), .Z(PRODUCT[682]) );
  AND U685 ( .A(A[683]), .B(B[0]), .Z(PRODUCT[683]) );
  AND U686 ( .A(A[684]), .B(B[0]), .Z(PRODUCT[684]) );
  AND U687 ( .A(A[685]), .B(B[0]), .Z(PRODUCT[685]) );
  AND U688 ( .A(A[686]), .B(B[0]), .Z(PRODUCT[686]) );
  AND U689 ( .A(A[687]), .B(B[0]), .Z(PRODUCT[687]) );
  AND U690 ( .A(A[688]), .B(B[0]), .Z(PRODUCT[688]) );
  AND U691 ( .A(A[689]), .B(B[0]), .Z(PRODUCT[689]) );
  AND U692 ( .A(A[690]), .B(B[0]), .Z(PRODUCT[690]) );
  AND U693 ( .A(A[691]), .B(B[0]), .Z(PRODUCT[691]) );
  AND U694 ( .A(A[692]), .B(B[0]), .Z(PRODUCT[692]) );
  AND U695 ( .A(A[693]), .B(B[0]), .Z(PRODUCT[693]) );
  AND U696 ( .A(A[694]), .B(B[0]), .Z(PRODUCT[694]) );
  AND U697 ( .A(A[695]), .B(B[0]), .Z(PRODUCT[695]) );
  AND U698 ( .A(A[696]), .B(B[0]), .Z(PRODUCT[696]) );
  AND U699 ( .A(A[697]), .B(B[0]), .Z(PRODUCT[697]) );
  AND U700 ( .A(A[698]), .B(B[0]), .Z(PRODUCT[698]) );
  AND U701 ( .A(A[699]), .B(B[0]), .Z(PRODUCT[699]) );
  AND U702 ( .A(A[700]), .B(B[0]), .Z(PRODUCT[700]) );
  AND U703 ( .A(A[701]), .B(B[0]), .Z(PRODUCT[701]) );
  AND U704 ( .A(A[702]), .B(B[0]), .Z(PRODUCT[702]) );
  AND U705 ( .A(A[703]), .B(B[0]), .Z(PRODUCT[703]) );
  AND U706 ( .A(A[704]), .B(B[0]), .Z(PRODUCT[704]) );
  AND U707 ( .A(A[705]), .B(B[0]), .Z(PRODUCT[705]) );
  AND U708 ( .A(A[706]), .B(B[0]), .Z(PRODUCT[706]) );
  AND U709 ( .A(A[707]), .B(B[0]), .Z(PRODUCT[707]) );
  AND U710 ( .A(A[708]), .B(B[0]), .Z(PRODUCT[708]) );
  AND U711 ( .A(A[709]), .B(B[0]), .Z(PRODUCT[709]) );
  AND U712 ( .A(A[710]), .B(B[0]), .Z(PRODUCT[710]) );
  AND U713 ( .A(A[711]), .B(B[0]), .Z(PRODUCT[711]) );
  AND U714 ( .A(A[712]), .B(B[0]), .Z(PRODUCT[712]) );
  AND U715 ( .A(A[713]), .B(B[0]), .Z(PRODUCT[713]) );
  AND U716 ( .A(A[714]), .B(B[0]), .Z(PRODUCT[714]) );
  AND U717 ( .A(A[715]), .B(B[0]), .Z(PRODUCT[715]) );
  AND U718 ( .A(A[716]), .B(B[0]), .Z(PRODUCT[716]) );
  AND U719 ( .A(A[717]), .B(B[0]), .Z(PRODUCT[717]) );
  AND U720 ( .A(A[718]), .B(B[0]), .Z(PRODUCT[718]) );
  AND U721 ( .A(A[719]), .B(B[0]), .Z(PRODUCT[719]) );
  AND U722 ( .A(A[720]), .B(B[0]), .Z(PRODUCT[720]) );
  AND U723 ( .A(A[721]), .B(B[0]), .Z(PRODUCT[721]) );
  AND U724 ( .A(A[722]), .B(B[0]), .Z(PRODUCT[722]) );
  AND U725 ( .A(A[723]), .B(B[0]), .Z(PRODUCT[723]) );
  AND U726 ( .A(A[724]), .B(B[0]), .Z(PRODUCT[724]) );
  AND U727 ( .A(A[725]), .B(B[0]), .Z(PRODUCT[725]) );
  AND U728 ( .A(A[726]), .B(B[0]), .Z(PRODUCT[726]) );
  AND U729 ( .A(A[727]), .B(B[0]), .Z(PRODUCT[727]) );
  AND U730 ( .A(A[728]), .B(B[0]), .Z(PRODUCT[728]) );
  AND U731 ( .A(A[729]), .B(B[0]), .Z(PRODUCT[729]) );
  AND U732 ( .A(A[730]), .B(B[0]), .Z(PRODUCT[730]) );
  AND U733 ( .A(A[731]), .B(B[0]), .Z(PRODUCT[731]) );
  AND U734 ( .A(A[732]), .B(B[0]), .Z(PRODUCT[732]) );
  AND U735 ( .A(A[733]), .B(B[0]), .Z(PRODUCT[733]) );
  AND U736 ( .A(A[734]), .B(B[0]), .Z(PRODUCT[734]) );
  AND U737 ( .A(A[735]), .B(B[0]), .Z(PRODUCT[735]) );
  AND U738 ( .A(A[736]), .B(B[0]), .Z(PRODUCT[736]) );
  AND U739 ( .A(A[737]), .B(B[0]), .Z(PRODUCT[737]) );
  AND U740 ( .A(A[738]), .B(B[0]), .Z(PRODUCT[738]) );
  AND U741 ( .A(A[739]), .B(B[0]), .Z(PRODUCT[739]) );
  AND U742 ( .A(A[740]), .B(B[0]), .Z(PRODUCT[740]) );
  AND U743 ( .A(A[741]), .B(B[0]), .Z(PRODUCT[741]) );
  AND U744 ( .A(A[742]), .B(B[0]), .Z(PRODUCT[742]) );
  AND U745 ( .A(A[743]), .B(B[0]), .Z(PRODUCT[743]) );
  AND U746 ( .A(A[744]), .B(B[0]), .Z(PRODUCT[744]) );
  AND U747 ( .A(A[745]), .B(B[0]), .Z(PRODUCT[745]) );
  AND U748 ( .A(A[746]), .B(B[0]), .Z(PRODUCT[746]) );
  AND U749 ( .A(A[747]), .B(B[0]), .Z(PRODUCT[747]) );
  AND U750 ( .A(A[748]), .B(B[0]), .Z(PRODUCT[748]) );
  AND U751 ( .A(A[749]), .B(B[0]), .Z(PRODUCT[749]) );
  AND U752 ( .A(A[750]), .B(B[0]), .Z(PRODUCT[750]) );
  AND U753 ( .A(A[751]), .B(B[0]), .Z(PRODUCT[751]) );
  AND U754 ( .A(A[752]), .B(B[0]), .Z(PRODUCT[752]) );
  AND U755 ( .A(A[753]), .B(B[0]), .Z(PRODUCT[753]) );
  AND U756 ( .A(A[754]), .B(B[0]), .Z(PRODUCT[754]) );
  AND U757 ( .A(A[755]), .B(B[0]), .Z(PRODUCT[755]) );
  AND U758 ( .A(A[756]), .B(B[0]), .Z(PRODUCT[756]) );
  AND U759 ( .A(A[757]), .B(B[0]), .Z(PRODUCT[757]) );
  AND U760 ( .A(A[758]), .B(B[0]), .Z(PRODUCT[758]) );
  AND U761 ( .A(A[759]), .B(B[0]), .Z(PRODUCT[759]) );
  AND U762 ( .A(A[760]), .B(B[0]), .Z(PRODUCT[760]) );
  AND U763 ( .A(A[761]), .B(B[0]), .Z(PRODUCT[761]) );
  AND U764 ( .A(A[762]), .B(B[0]), .Z(PRODUCT[762]) );
  AND U765 ( .A(A[763]), .B(B[0]), .Z(PRODUCT[763]) );
  AND U766 ( .A(A[764]), .B(B[0]), .Z(PRODUCT[764]) );
  AND U767 ( .A(A[765]), .B(B[0]), .Z(PRODUCT[765]) );
  AND U768 ( .A(A[766]), .B(B[0]), .Z(PRODUCT[766]) );
  AND U769 ( .A(A[767]), .B(B[0]), .Z(PRODUCT[767]) );
  AND U770 ( .A(A[768]), .B(B[0]), .Z(PRODUCT[768]) );
  AND U771 ( .A(A[769]), .B(B[0]), .Z(PRODUCT[769]) );
  AND U772 ( .A(A[770]), .B(B[0]), .Z(PRODUCT[770]) );
  AND U773 ( .A(A[771]), .B(B[0]), .Z(PRODUCT[771]) );
  AND U774 ( .A(A[772]), .B(B[0]), .Z(PRODUCT[772]) );
  AND U775 ( .A(A[773]), .B(B[0]), .Z(PRODUCT[773]) );
  AND U776 ( .A(A[774]), .B(B[0]), .Z(PRODUCT[774]) );
  AND U777 ( .A(A[775]), .B(B[0]), .Z(PRODUCT[775]) );
  AND U778 ( .A(A[776]), .B(B[0]), .Z(PRODUCT[776]) );
  AND U779 ( .A(A[777]), .B(B[0]), .Z(PRODUCT[777]) );
  AND U780 ( .A(A[778]), .B(B[0]), .Z(PRODUCT[778]) );
  AND U781 ( .A(A[779]), .B(B[0]), .Z(PRODUCT[779]) );
  AND U782 ( .A(A[780]), .B(B[0]), .Z(PRODUCT[780]) );
  AND U783 ( .A(A[781]), .B(B[0]), .Z(PRODUCT[781]) );
  AND U784 ( .A(A[782]), .B(B[0]), .Z(PRODUCT[782]) );
  AND U785 ( .A(A[783]), .B(B[0]), .Z(PRODUCT[783]) );
  AND U786 ( .A(A[784]), .B(B[0]), .Z(PRODUCT[784]) );
  AND U787 ( .A(A[785]), .B(B[0]), .Z(PRODUCT[785]) );
  AND U788 ( .A(A[786]), .B(B[0]), .Z(PRODUCT[786]) );
  AND U789 ( .A(A[787]), .B(B[0]), .Z(PRODUCT[787]) );
  AND U790 ( .A(A[788]), .B(B[0]), .Z(PRODUCT[788]) );
  AND U791 ( .A(A[789]), .B(B[0]), .Z(PRODUCT[789]) );
  AND U792 ( .A(A[790]), .B(B[0]), .Z(PRODUCT[790]) );
  AND U793 ( .A(A[791]), .B(B[0]), .Z(PRODUCT[791]) );
  AND U794 ( .A(A[792]), .B(B[0]), .Z(PRODUCT[792]) );
  AND U795 ( .A(A[793]), .B(B[0]), .Z(PRODUCT[793]) );
  AND U796 ( .A(A[794]), .B(B[0]), .Z(PRODUCT[794]) );
  AND U797 ( .A(A[795]), .B(B[0]), .Z(PRODUCT[795]) );
  AND U798 ( .A(A[796]), .B(B[0]), .Z(PRODUCT[796]) );
  AND U799 ( .A(A[797]), .B(B[0]), .Z(PRODUCT[797]) );
  AND U800 ( .A(A[798]), .B(B[0]), .Z(PRODUCT[798]) );
  AND U801 ( .A(A[799]), .B(B[0]), .Z(PRODUCT[799]) );
  AND U802 ( .A(A[800]), .B(B[0]), .Z(PRODUCT[800]) );
  AND U803 ( .A(A[801]), .B(B[0]), .Z(PRODUCT[801]) );
  AND U804 ( .A(A[802]), .B(B[0]), .Z(PRODUCT[802]) );
  AND U805 ( .A(A[803]), .B(B[0]), .Z(PRODUCT[803]) );
  AND U806 ( .A(A[804]), .B(B[0]), .Z(PRODUCT[804]) );
  AND U807 ( .A(A[805]), .B(B[0]), .Z(PRODUCT[805]) );
  AND U808 ( .A(A[806]), .B(B[0]), .Z(PRODUCT[806]) );
  AND U809 ( .A(A[807]), .B(B[0]), .Z(PRODUCT[807]) );
  AND U810 ( .A(A[808]), .B(B[0]), .Z(PRODUCT[808]) );
  AND U811 ( .A(A[809]), .B(B[0]), .Z(PRODUCT[809]) );
  AND U812 ( .A(A[810]), .B(B[0]), .Z(PRODUCT[810]) );
  AND U813 ( .A(A[811]), .B(B[0]), .Z(PRODUCT[811]) );
  AND U814 ( .A(A[812]), .B(B[0]), .Z(PRODUCT[812]) );
  AND U815 ( .A(A[813]), .B(B[0]), .Z(PRODUCT[813]) );
  AND U816 ( .A(A[814]), .B(B[0]), .Z(PRODUCT[814]) );
  AND U817 ( .A(A[815]), .B(B[0]), .Z(PRODUCT[815]) );
  AND U818 ( .A(A[816]), .B(B[0]), .Z(PRODUCT[816]) );
  AND U819 ( .A(A[817]), .B(B[0]), .Z(PRODUCT[817]) );
  AND U820 ( .A(A[818]), .B(B[0]), .Z(PRODUCT[818]) );
  AND U821 ( .A(A[819]), .B(B[0]), .Z(PRODUCT[819]) );
  AND U822 ( .A(A[820]), .B(B[0]), .Z(PRODUCT[820]) );
  AND U823 ( .A(A[821]), .B(B[0]), .Z(PRODUCT[821]) );
  AND U824 ( .A(A[822]), .B(B[0]), .Z(PRODUCT[822]) );
  AND U825 ( .A(A[823]), .B(B[0]), .Z(PRODUCT[823]) );
  AND U826 ( .A(A[824]), .B(B[0]), .Z(PRODUCT[824]) );
  AND U827 ( .A(A[825]), .B(B[0]), .Z(PRODUCT[825]) );
  AND U828 ( .A(A[826]), .B(B[0]), .Z(PRODUCT[826]) );
  AND U829 ( .A(A[827]), .B(B[0]), .Z(PRODUCT[827]) );
  AND U830 ( .A(A[828]), .B(B[0]), .Z(PRODUCT[828]) );
  AND U831 ( .A(A[829]), .B(B[0]), .Z(PRODUCT[829]) );
  AND U832 ( .A(A[830]), .B(B[0]), .Z(PRODUCT[830]) );
  AND U833 ( .A(A[831]), .B(B[0]), .Z(PRODUCT[831]) );
  AND U834 ( .A(A[832]), .B(B[0]), .Z(PRODUCT[832]) );
  AND U835 ( .A(A[833]), .B(B[0]), .Z(PRODUCT[833]) );
  AND U836 ( .A(A[834]), .B(B[0]), .Z(PRODUCT[834]) );
  AND U837 ( .A(A[835]), .B(B[0]), .Z(PRODUCT[835]) );
  AND U838 ( .A(A[836]), .B(B[0]), .Z(PRODUCT[836]) );
  AND U839 ( .A(A[837]), .B(B[0]), .Z(PRODUCT[837]) );
  AND U840 ( .A(A[838]), .B(B[0]), .Z(PRODUCT[838]) );
  AND U841 ( .A(A[839]), .B(B[0]), .Z(PRODUCT[839]) );
  AND U842 ( .A(A[840]), .B(B[0]), .Z(PRODUCT[840]) );
  AND U843 ( .A(A[841]), .B(B[0]), .Z(PRODUCT[841]) );
  AND U844 ( .A(A[842]), .B(B[0]), .Z(PRODUCT[842]) );
  AND U845 ( .A(A[843]), .B(B[0]), .Z(PRODUCT[843]) );
  AND U846 ( .A(A[844]), .B(B[0]), .Z(PRODUCT[844]) );
  AND U847 ( .A(A[845]), .B(B[0]), .Z(PRODUCT[845]) );
  AND U848 ( .A(A[846]), .B(B[0]), .Z(PRODUCT[846]) );
  AND U849 ( .A(A[847]), .B(B[0]), .Z(PRODUCT[847]) );
  AND U850 ( .A(A[848]), .B(B[0]), .Z(PRODUCT[848]) );
  AND U851 ( .A(A[849]), .B(B[0]), .Z(PRODUCT[849]) );
  AND U852 ( .A(A[850]), .B(B[0]), .Z(PRODUCT[850]) );
  AND U853 ( .A(A[851]), .B(B[0]), .Z(PRODUCT[851]) );
  AND U854 ( .A(A[852]), .B(B[0]), .Z(PRODUCT[852]) );
  AND U855 ( .A(A[853]), .B(B[0]), .Z(PRODUCT[853]) );
  AND U856 ( .A(A[854]), .B(B[0]), .Z(PRODUCT[854]) );
  AND U857 ( .A(A[855]), .B(B[0]), .Z(PRODUCT[855]) );
  AND U858 ( .A(A[856]), .B(B[0]), .Z(PRODUCT[856]) );
  AND U859 ( .A(A[857]), .B(B[0]), .Z(PRODUCT[857]) );
  AND U860 ( .A(A[858]), .B(B[0]), .Z(PRODUCT[858]) );
  AND U861 ( .A(A[859]), .B(B[0]), .Z(PRODUCT[859]) );
  AND U862 ( .A(A[860]), .B(B[0]), .Z(PRODUCT[860]) );
  AND U863 ( .A(A[861]), .B(B[0]), .Z(PRODUCT[861]) );
  AND U864 ( .A(A[862]), .B(B[0]), .Z(PRODUCT[862]) );
  AND U865 ( .A(A[863]), .B(B[0]), .Z(PRODUCT[863]) );
  AND U866 ( .A(A[864]), .B(B[0]), .Z(PRODUCT[864]) );
  AND U867 ( .A(A[865]), .B(B[0]), .Z(PRODUCT[865]) );
  AND U868 ( .A(A[866]), .B(B[0]), .Z(PRODUCT[866]) );
  AND U869 ( .A(A[867]), .B(B[0]), .Z(PRODUCT[867]) );
  AND U870 ( .A(A[868]), .B(B[0]), .Z(PRODUCT[868]) );
  AND U871 ( .A(A[869]), .B(B[0]), .Z(PRODUCT[869]) );
  AND U872 ( .A(A[870]), .B(B[0]), .Z(PRODUCT[870]) );
  AND U873 ( .A(A[871]), .B(B[0]), .Z(PRODUCT[871]) );
  AND U874 ( .A(A[872]), .B(B[0]), .Z(PRODUCT[872]) );
  AND U875 ( .A(A[873]), .B(B[0]), .Z(PRODUCT[873]) );
  AND U876 ( .A(A[874]), .B(B[0]), .Z(PRODUCT[874]) );
  AND U877 ( .A(A[875]), .B(B[0]), .Z(PRODUCT[875]) );
  AND U878 ( .A(A[876]), .B(B[0]), .Z(PRODUCT[876]) );
  AND U879 ( .A(A[877]), .B(B[0]), .Z(PRODUCT[877]) );
  AND U880 ( .A(A[878]), .B(B[0]), .Z(PRODUCT[878]) );
  AND U881 ( .A(A[879]), .B(B[0]), .Z(PRODUCT[879]) );
  AND U882 ( .A(A[880]), .B(B[0]), .Z(PRODUCT[880]) );
  AND U883 ( .A(A[881]), .B(B[0]), .Z(PRODUCT[881]) );
  AND U884 ( .A(A[882]), .B(B[0]), .Z(PRODUCT[882]) );
  AND U885 ( .A(A[883]), .B(B[0]), .Z(PRODUCT[883]) );
  AND U886 ( .A(A[884]), .B(B[0]), .Z(PRODUCT[884]) );
  AND U887 ( .A(A[885]), .B(B[0]), .Z(PRODUCT[885]) );
  AND U888 ( .A(A[886]), .B(B[0]), .Z(PRODUCT[886]) );
  AND U889 ( .A(A[887]), .B(B[0]), .Z(PRODUCT[887]) );
  AND U890 ( .A(A[888]), .B(B[0]), .Z(PRODUCT[888]) );
  AND U891 ( .A(A[889]), .B(B[0]), .Z(PRODUCT[889]) );
  AND U892 ( .A(A[890]), .B(B[0]), .Z(PRODUCT[890]) );
  AND U893 ( .A(A[891]), .B(B[0]), .Z(PRODUCT[891]) );
  AND U894 ( .A(A[892]), .B(B[0]), .Z(PRODUCT[892]) );
  AND U895 ( .A(A[893]), .B(B[0]), .Z(PRODUCT[893]) );
  AND U896 ( .A(A[894]), .B(B[0]), .Z(PRODUCT[894]) );
  AND U897 ( .A(A[895]), .B(B[0]), .Z(PRODUCT[895]) );
  AND U898 ( .A(A[896]), .B(B[0]), .Z(PRODUCT[896]) );
  AND U899 ( .A(A[897]), .B(B[0]), .Z(PRODUCT[897]) );
  AND U900 ( .A(A[898]), .B(B[0]), .Z(PRODUCT[898]) );
  AND U901 ( .A(A[899]), .B(B[0]), .Z(PRODUCT[899]) );
  AND U902 ( .A(A[900]), .B(B[0]), .Z(PRODUCT[900]) );
  AND U903 ( .A(A[901]), .B(B[0]), .Z(PRODUCT[901]) );
  AND U904 ( .A(A[902]), .B(B[0]), .Z(PRODUCT[902]) );
  AND U905 ( .A(A[903]), .B(B[0]), .Z(PRODUCT[903]) );
  AND U906 ( .A(A[904]), .B(B[0]), .Z(PRODUCT[904]) );
  AND U907 ( .A(A[905]), .B(B[0]), .Z(PRODUCT[905]) );
  AND U908 ( .A(A[906]), .B(B[0]), .Z(PRODUCT[906]) );
  AND U909 ( .A(A[907]), .B(B[0]), .Z(PRODUCT[907]) );
  AND U910 ( .A(A[908]), .B(B[0]), .Z(PRODUCT[908]) );
  AND U911 ( .A(A[909]), .B(B[0]), .Z(PRODUCT[909]) );
  AND U912 ( .A(A[910]), .B(B[0]), .Z(PRODUCT[910]) );
  AND U913 ( .A(A[911]), .B(B[0]), .Z(PRODUCT[911]) );
  AND U914 ( .A(A[912]), .B(B[0]), .Z(PRODUCT[912]) );
  AND U915 ( .A(A[913]), .B(B[0]), .Z(PRODUCT[913]) );
  AND U916 ( .A(A[914]), .B(B[0]), .Z(PRODUCT[914]) );
  AND U917 ( .A(A[915]), .B(B[0]), .Z(PRODUCT[915]) );
  AND U918 ( .A(A[916]), .B(B[0]), .Z(PRODUCT[916]) );
  AND U919 ( .A(A[917]), .B(B[0]), .Z(PRODUCT[917]) );
  AND U920 ( .A(A[918]), .B(B[0]), .Z(PRODUCT[918]) );
  AND U921 ( .A(A[919]), .B(B[0]), .Z(PRODUCT[919]) );
  AND U922 ( .A(A[920]), .B(B[0]), .Z(PRODUCT[920]) );
  AND U923 ( .A(A[921]), .B(B[0]), .Z(PRODUCT[921]) );
  AND U924 ( .A(A[922]), .B(B[0]), .Z(PRODUCT[922]) );
  AND U925 ( .A(A[923]), .B(B[0]), .Z(PRODUCT[923]) );
  AND U926 ( .A(A[924]), .B(B[0]), .Z(PRODUCT[924]) );
  AND U927 ( .A(A[925]), .B(B[0]), .Z(PRODUCT[925]) );
  AND U928 ( .A(A[926]), .B(B[0]), .Z(PRODUCT[926]) );
  AND U929 ( .A(A[927]), .B(B[0]), .Z(PRODUCT[927]) );
  AND U930 ( .A(A[928]), .B(B[0]), .Z(PRODUCT[928]) );
  AND U931 ( .A(A[929]), .B(B[0]), .Z(PRODUCT[929]) );
  AND U932 ( .A(A[930]), .B(B[0]), .Z(PRODUCT[930]) );
  AND U933 ( .A(A[931]), .B(B[0]), .Z(PRODUCT[931]) );
  AND U934 ( .A(A[932]), .B(B[0]), .Z(PRODUCT[932]) );
  AND U935 ( .A(A[933]), .B(B[0]), .Z(PRODUCT[933]) );
  AND U936 ( .A(A[934]), .B(B[0]), .Z(PRODUCT[934]) );
  AND U937 ( .A(A[935]), .B(B[0]), .Z(PRODUCT[935]) );
  AND U938 ( .A(A[936]), .B(B[0]), .Z(PRODUCT[936]) );
  AND U939 ( .A(A[937]), .B(B[0]), .Z(PRODUCT[937]) );
  AND U940 ( .A(A[938]), .B(B[0]), .Z(PRODUCT[938]) );
  AND U941 ( .A(A[939]), .B(B[0]), .Z(PRODUCT[939]) );
  AND U942 ( .A(A[940]), .B(B[0]), .Z(PRODUCT[940]) );
  AND U943 ( .A(A[941]), .B(B[0]), .Z(PRODUCT[941]) );
  AND U944 ( .A(A[942]), .B(B[0]), .Z(PRODUCT[942]) );
  AND U945 ( .A(A[943]), .B(B[0]), .Z(PRODUCT[943]) );
  AND U946 ( .A(A[944]), .B(B[0]), .Z(PRODUCT[944]) );
  AND U947 ( .A(A[945]), .B(B[0]), .Z(PRODUCT[945]) );
  AND U948 ( .A(A[946]), .B(B[0]), .Z(PRODUCT[946]) );
  AND U949 ( .A(A[947]), .B(B[0]), .Z(PRODUCT[947]) );
  AND U950 ( .A(A[948]), .B(B[0]), .Z(PRODUCT[948]) );
  AND U951 ( .A(A[949]), .B(B[0]), .Z(PRODUCT[949]) );
  AND U952 ( .A(A[950]), .B(B[0]), .Z(PRODUCT[950]) );
  AND U953 ( .A(A[951]), .B(B[0]), .Z(PRODUCT[951]) );
  AND U954 ( .A(A[952]), .B(B[0]), .Z(PRODUCT[952]) );
  AND U955 ( .A(A[953]), .B(B[0]), .Z(PRODUCT[953]) );
  AND U956 ( .A(A[954]), .B(B[0]), .Z(PRODUCT[954]) );
  AND U957 ( .A(A[955]), .B(B[0]), .Z(PRODUCT[955]) );
  AND U958 ( .A(A[956]), .B(B[0]), .Z(PRODUCT[956]) );
  AND U959 ( .A(A[957]), .B(B[0]), .Z(PRODUCT[957]) );
  AND U960 ( .A(A[958]), .B(B[0]), .Z(PRODUCT[958]) );
  AND U961 ( .A(A[959]), .B(B[0]), .Z(PRODUCT[959]) );
  AND U962 ( .A(A[960]), .B(B[0]), .Z(PRODUCT[960]) );
  AND U963 ( .A(A[961]), .B(B[0]), .Z(PRODUCT[961]) );
  AND U964 ( .A(A[962]), .B(B[0]), .Z(PRODUCT[962]) );
  AND U965 ( .A(A[963]), .B(B[0]), .Z(PRODUCT[963]) );
  AND U966 ( .A(A[964]), .B(B[0]), .Z(PRODUCT[964]) );
  AND U967 ( .A(A[965]), .B(B[0]), .Z(PRODUCT[965]) );
  AND U968 ( .A(A[966]), .B(B[0]), .Z(PRODUCT[966]) );
  AND U969 ( .A(A[967]), .B(B[0]), .Z(PRODUCT[967]) );
  AND U970 ( .A(A[968]), .B(B[0]), .Z(PRODUCT[968]) );
  AND U971 ( .A(A[969]), .B(B[0]), .Z(PRODUCT[969]) );
  AND U972 ( .A(A[970]), .B(B[0]), .Z(PRODUCT[970]) );
  AND U973 ( .A(A[971]), .B(B[0]), .Z(PRODUCT[971]) );
  AND U974 ( .A(A[972]), .B(B[0]), .Z(PRODUCT[972]) );
  AND U975 ( .A(A[973]), .B(B[0]), .Z(PRODUCT[973]) );
  AND U976 ( .A(A[974]), .B(B[0]), .Z(PRODUCT[974]) );
  AND U977 ( .A(A[975]), .B(B[0]), .Z(PRODUCT[975]) );
  AND U978 ( .A(A[976]), .B(B[0]), .Z(PRODUCT[976]) );
  AND U979 ( .A(A[977]), .B(B[0]), .Z(PRODUCT[977]) );
  AND U980 ( .A(A[978]), .B(B[0]), .Z(PRODUCT[978]) );
  AND U981 ( .A(A[979]), .B(B[0]), .Z(PRODUCT[979]) );
  AND U982 ( .A(A[980]), .B(B[0]), .Z(PRODUCT[980]) );
  AND U983 ( .A(A[981]), .B(B[0]), .Z(PRODUCT[981]) );
  AND U984 ( .A(A[982]), .B(B[0]), .Z(PRODUCT[982]) );
  AND U985 ( .A(A[983]), .B(B[0]), .Z(PRODUCT[983]) );
  AND U986 ( .A(A[984]), .B(B[0]), .Z(PRODUCT[984]) );
  AND U987 ( .A(A[985]), .B(B[0]), .Z(PRODUCT[985]) );
  AND U988 ( .A(A[986]), .B(B[0]), .Z(PRODUCT[986]) );
  AND U989 ( .A(A[987]), .B(B[0]), .Z(PRODUCT[987]) );
  AND U990 ( .A(A[988]), .B(B[0]), .Z(PRODUCT[988]) );
  AND U991 ( .A(A[989]), .B(B[0]), .Z(PRODUCT[989]) );
  AND U992 ( .A(A[990]), .B(B[0]), .Z(PRODUCT[990]) );
  AND U993 ( .A(A[991]), .B(B[0]), .Z(PRODUCT[991]) );
  AND U994 ( .A(A[992]), .B(B[0]), .Z(PRODUCT[992]) );
  AND U995 ( .A(A[993]), .B(B[0]), .Z(PRODUCT[993]) );
  AND U996 ( .A(A[994]), .B(B[0]), .Z(PRODUCT[994]) );
  AND U997 ( .A(A[995]), .B(B[0]), .Z(PRODUCT[995]) );
  AND U998 ( .A(A[996]), .B(B[0]), .Z(PRODUCT[996]) );
  AND U999 ( .A(A[997]), .B(B[0]), .Z(PRODUCT[997]) );
  AND U1000 ( .A(A[998]), .B(B[0]), .Z(PRODUCT[998]) );
  AND U1001 ( .A(A[999]), .B(B[0]), .Z(PRODUCT[999]) );
  AND U1002 ( .A(A[1000]), .B(B[0]), .Z(PRODUCT[1000]) );
  AND U1003 ( .A(A[1001]), .B(B[0]), .Z(PRODUCT[1001]) );
  AND U1004 ( .A(A[1002]), .B(B[0]), .Z(PRODUCT[1002]) );
  AND U1005 ( .A(A[1003]), .B(B[0]), .Z(PRODUCT[1003]) );
  AND U1006 ( .A(A[1004]), .B(B[0]), .Z(PRODUCT[1004]) );
  AND U1007 ( .A(A[1005]), .B(B[0]), .Z(PRODUCT[1005]) );
  AND U1008 ( .A(A[1006]), .B(B[0]), .Z(PRODUCT[1006]) );
  AND U1009 ( .A(A[1007]), .B(B[0]), .Z(PRODUCT[1007]) );
  AND U1010 ( .A(A[1008]), .B(B[0]), .Z(PRODUCT[1008]) );
  AND U1011 ( .A(A[1009]), .B(B[0]), .Z(PRODUCT[1009]) );
  AND U1012 ( .A(A[1010]), .B(B[0]), .Z(PRODUCT[1010]) );
  AND U1013 ( .A(A[1011]), .B(B[0]), .Z(PRODUCT[1011]) );
  AND U1014 ( .A(A[1012]), .B(B[0]), .Z(PRODUCT[1012]) );
  AND U1015 ( .A(A[1013]), .B(B[0]), .Z(PRODUCT[1013]) );
  AND U1016 ( .A(A[1014]), .B(B[0]), .Z(PRODUCT[1014]) );
  AND U1017 ( .A(A[1015]), .B(B[0]), .Z(PRODUCT[1015]) );
  AND U1018 ( .A(A[1016]), .B(B[0]), .Z(PRODUCT[1016]) );
  AND U1019 ( .A(A[1017]), .B(B[0]), .Z(PRODUCT[1017]) );
  AND U1020 ( .A(A[1018]), .B(B[0]), .Z(PRODUCT[1018]) );
  AND U1021 ( .A(A[1019]), .B(B[0]), .Z(PRODUCT[1019]) );
  AND U1022 ( .A(A[1020]), .B(B[0]), .Z(PRODUCT[1020]) );
  AND U1023 ( .A(A[1021]), .B(B[0]), .Z(PRODUCT[1021]) );
  AND U1024 ( .A(A[1022]), .B(B[0]), .Z(PRODUCT[1022]) );
  AND U1025 ( .A(A[1023]), .B(B[0]), .Z(PRODUCT[1023]) );
endmodule


module mult_N1024_CC1024 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [0:0] b;
  output [1023:0] c;
  input clk, rst;

  wire   [1023:1] swire;
  wire   [1023:0] clocal;
  wire   [2047:1024] sreg;
  wire   SYNOPSYS_UNCONNECTED__0;

  DFF \sreg_reg[1024]  ( .D(swire[1]), .CLK(clk), .RST(rst), .Q(sreg[1024]) );
  DFF \sreg_reg[1025]  ( .D(swire[2]), .CLK(clk), .RST(rst), .Q(sreg[1025]) );
  DFF \sreg_reg[1026]  ( .D(swire[3]), .CLK(clk), .RST(rst), .Q(sreg[1026]) );
  DFF \sreg_reg[1027]  ( .D(swire[4]), .CLK(clk), .RST(rst), .Q(sreg[1027]) );
  DFF \sreg_reg[1028]  ( .D(swire[5]), .CLK(clk), .RST(rst), .Q(sreg[1028]) );
  DFF \sreg_reg[1029]  ( .D(swire[6]), .CLK(clk), .RST(rst), .Q(sreg[1029]) );
  DFF \sreg_reg[1030]  ( .D(swire[7]), .CLK(clk), .RST(rst), .Q(sreg[1030]) );
  DFF \sreg_reg[1031]  ( .D(swire[8]), .CLK(clk), .RST(rst), .Q(sreg[1031]) );
  DFF \sreg_reg[1032]  ( .D(swire[9]), .CLK(clk), .RST(rst), .Q(sreg[1032]) );
  DFF \sreg_reg[1033]  ( .D(swire[10]), .CLK(clk), .RST(rst), .Q(sreg[1033])
         );
  DFF \sreg_reg[1034]  ( .D(swire[11]), .CLK(clk), .RST(rst), .Q(sreg[1034])
         );
  DFF \sreg_reg[1035]  ( .D(swire[12]), .CLK(clk), .RST(rst), .Q(sreg[1035])
         );
  DFF \sreg_reg[1036]  ( .D(swire[13]), .CLK(clk), .RST(rst), .Q(sreg[1036])
         );
  DFF \sreg_reg[1037]  ( .D(swire[14]), .CLK(clk), .RST(rst), .Q(sreg[1037])
         );
  DFF \sreg_reg[1038]  ( .D(swire[15]), .CLK(clk), .RST(rst), .Q(sreg[1038])
         );
  DFF \sreg_reg[1039]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[1039])
         );
  DFF \sreg_reg[1040]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[1040])
         );
  DFF \sreg_reg[1041]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[1041])
         );
  DFF \sreg_reg[1042]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[1042])
         );
  DFF \sreg_reg[1043]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[1043])
         );
  DFF \sreg_reg[1044]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[1044])
         );
  DFF \sreg_reg[1045]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[1045])
         );
  DFF \sreg_reg[1046]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[1046])
         );
  DFF \sreg_reg[1047]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[1047])
         );
  DFF \sreg_reg[1048]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[1048])
         );
  DFF \sreg_reg[1049]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[1049])
         );
  DFF \sreg_reg[1050]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[1050])
         );
  DFF \sreg_reg[1051]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[1051])
         );
  DFF \sreg_reg[1052]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[1052])
         );
  DFF \sreg_reg[1053]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[1053])
         );
  DFF \sreg_reg[1054]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[1054])
         );
  DFF \sreg_reg[1055]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[1055])
         );
  DFF \sreg_reg[1056]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[1056])
         );
  DFF \sreg_reg[1057]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[1057])
         );
  DFF \sreg_reg[1058]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[1058])
         );
  DFF \sreg_reg[1059]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[1059])
         );
  DFF \sreg_reg[1060]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[1060])
         );
  DFF \sreg_reg[1061]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[1061])
         );
  DFF \sreg_reg[1062]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[1062])
         );
  DFF \sreg_reg[1063]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[1063])
         );
  DFF \sreg_reg[1064]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[1064])
         );
  DFF \sreg_reg[1065]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[1065])
         );
  DFF \sreg_reg[1066]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[1066])
         );
  DFF \sreg_reg[1067]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[1067])
         );
  DFF \sreg_reg[1068]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[1068])
         );
  DFF \sreg_reg[1069]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[1069])
         );
  DFF \sreg_reg[1070]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[1070])
         );
  DFF \sreg_reg[1071]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[1071])
         );
  DFF \sreg_reg[1072]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[1072])
         );
  DFF \sreg_reg[1073]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[1073])
         );
  DFF \sreg_reg[1074]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[1074])
         );
  DFF \sreg_reg[1075]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[1075])
         );
  DFF \sreg_reg[1076]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[1076])
         );
  DFF \sreg_reg[1077]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[1077])
         );
  DFF \sreg_reg[1078]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[1078])
         );
  DFF \sreg_reg[1079]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[1079])
         );
  DFF \sreg_reg[1080]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[1080])
         );
  DFF \sreg_reg[1081]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[1081])
         );
  DFF \sreg_reg[1082]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[1082])
         );
  DFF \sreg_reg[1083]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[1083])
         );
  DFF \sreg_reg[1084]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[1084])
         );
  DFF \sreg_reg[1085]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[1085])
         );
  DFF \sreg_reg[1086]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[1086])
         );
  DFF \sreg_reg[1087]  ( .D(swire[64]), .CLK(clk), .RST(rst), .Q(sreg[1087])
         );
  DFF \sreg_reg[1088]  ( .D(swire[65]), .CLK(clk), .RST(rst), .Q(sreg[1088])
         );
  DFF \sreg_reg[1089]  ( .D(swire[66]), .CLK(clk), .RST(rst), .Q(sreg[1089])
         );
  DFF \sreg_reg[1090]  ( .D(swire[67]), .CLK(clk), .RST(rst), .Q(sreg[1090])
         );
  DFF \sreg_reg[1091]  ( .D(swire[68]), .CLK(clk), .RST(rst), .Q(sreg[1091])
         );
  DFF \sreg_reg[1092]  ( .D(swire[69]), .CLK(clk), .RST(rst), .Q(sreg[1092])
         );
  DFF \sreg_reg[1093]  ( .D(swire[70]), .CLK(clk), .RST(rst), .Q(sreg[1093])
         );
  DFF \sreg_reg[1094]  ( .D(swire[71]), .CLK(clk), .RST(rst), .Q(sreg[1094])
         );
  DFF \sreg_reg[1095]  ( .D(swire[72]), .CLK(clk), .RST(rst), .Q(sreg[1095])
         );
  DFF \sreg_reg[1096]  ( .D(swire[73]), .CLK(clk), .RST(rst), .Q(sreg[1096])
         );
  DFF \sreg_reg[1097]  ( .D(swire[74]), .CLK(clk), .RST(rst), .Q(sreg[1097])
         );
  DFF \sreg_reg[1098]  ( .D(swire[75]), .CLK(clk), .RST(rst), .Q(sreg[1098])
         );
  DFF \sreg_reg[1099]  ( .D(swire[76]), .CLK(clk), .RST(rst), .Q(sreg[1099])
         );
  DFF \sreg_reg[1100]  ( .D(swire[77]), .CLK(clk), .RST(rst), .Q(sreg[1100])
         );
  DFF \sreg_reg[1101]  ( .D(swire[78]), .CLK(clk), .RST(rst), .Q(sreg[1101])
         );
  DFF \sreg_reg[1102]  ( .D(swire[79]), .CLK(clk), .RST(rst), .Q(sreg[1102])
         );
  DFF \sreg_reg[1103]  ( .D(swire[80]), .CLK(clk), .RST(rst), .Q(sreg[1103])
         );
  DFF \sreg_reg[1104]  ( .D(swire[81]), .CLK(clk), .RST(rst), .Q(sreg[1104])
         );
  DFF \sreg_reg[1105]  ( .D(swire[82]), .CLK(clk), .RST(rst), .Q(sreg[1105])
         );
  DFF \sreg_reg[1106]  ( .D(swire[83]), .CLK(clk), .RST(rst), .Q(sreg[1106])
         );
  DFF \sreg_reg[1107]  ( .D(swire[84]), .CLK(clk), .RST(rst), .Q(sreg[1107])
         );
  DFF \sreg_reg[1108]  ( .D(swire[85]), .CLK(clk), .RST(rst), .Q(sreg[1108])
         );
  DFF \sreg_reg[1109]  ( .D(swire[86]), .CLK(clk), .RST(rst), .Q(sreg[1109])
         );
  DFF \sreg_reg[1110]  ( .D(swire[87]), .CLK(clk), .RST(rst), .Q(sreg[1110])
         );
  DFF \sreg_reg[1111]  ( .D(swire[88]), .CLK(clk), .RST(rst), .Q(sreg[1111])
         );
  DFF \sreg_reg[1112]  ( .D(swire[89]), .CLK(clk), .RST(rst), .Q(sreg[1112])
         );
  DFF \sreg_reg[1113]  ( .D(swire[90]), .CLK(clk), .RST(rst), .Q(sreg[1113])
         );
  DFF \sreg_reg[1114]  ( .D(swire[91]), .CLK(clk), .RST(rst), .Q(sreg[1114])
         );
  DFF \sreg_reg[1115]  ( .D(swire[92]), .CLK(clk), .RST(rst), .Q(sreg[1115])
         );
  DFF \sreg_reg[1116]  ( .D(swire[93]), .CLK(clk), .RST(rst), .Q(sreg[1116])
         );
  DFF \sreg_reg[1117]  ( .D(swire[94]), .CLK(clk), .RST(rst), .Q(sreg[1117])
         );
  DFF \sreg_reg[1118]  ( .D(swire[95]), .CLK(clk), .RST(rst), .Q(sreg[1118])
         );
  DFF \sreg_reg[1119]  ( .D(swire[96]), .CLK(clk), .RST(rst), .Q(sreg[1119])
         );
  DFF \sreg_reg[1120]  ( .D(swire[97]), .CLK(clk), .RST(rst), .Q(sreg[1120])
         );
  DFF \sreg_reg[1121]  ( .D(swire[98]), .CLK(clk), .RST(rst), .Q(sreg[1121])
         );
  DFF \sreg_reg[1122]  ( .D(swire[99]), .CLK(clk), .RST(rst), .Q(sreg[1122])
         );
  DFF \sreg_reg[1123]  ( .D(swire[100]), .CLK(clk), .RST(rst), .Q(sreg[1123])
         );
  DFF \sreg_reg[1124]  ( .D(swire[101]), .CLK(clk), .RST(rst), .Q(sreg[1124])
         );
  DFF \sreg_reg[1125]  ( .D(swire[102]), .CLK(clk), .RST(rst), .Q(sreg[1125])
         );
  DFF \sreg_reg[1126]  ( .D(swire[103]), .CLK(clk), .RST(rst), .Q(sreg[1126])
         );
  DFF \sreg_reg[1127]  ( .D(swire[104]), .CLK(clk), .RST(rst), .Q(sreg[1127])
         );
  DFF \sreg_reg[1128]  ( .D(swire[105]), .CLK(clk), .RST(rst), .Q(sreg[1128])
         );
  DFF \sreg_reg[1129]  ( .D(swire[106]), .CLK(clk), .RST(rst), .Q(sreg[1129])
         );
  DFF \sreg_reg[1130]  ( .D(swire[107]), .CLK(clk), .RST(rst), .Q(sreg[1130])
         );
  DFF \sreg_reg[1131]  ( .D(swire[108]), .CLK(clk), .RST(rst), .Q(sreg[1131])
         );
  DFF \sreg_reg[1132]  ( .D(swire[109]), .CLK(clk), .RST(rst), .Q(sreg[1132])
         );
  DFF \sreg_reg[1133]  ( .D(swire[110]), .CLK(clk), .RST(rst), .Q(sreg[1133])
         );
  DFF \sreg_reg[1134]  ( .D(swire[111]), .CLK(clk), .RST(rst), .Q(sreg[1134])
         );
  DFF \sreg_reg[1135]  ( .D(swire[112]), .CLK(clk), .RST(rst), .Q(sreg[1135])
         );
  DFF \sreg_reg[1136]  ( .D(swire[113]), .CLK(clk), .RST(rst), .Q(sreg[1136])
         );
  DFF \sreg_reg[1137]  ( .D(swire[114]), .CLK(clk), .RST(rst), .Q(sreg[1137])
         );
  DFF \sreg_reg[1138]  ( .D(swire[115]), .CLK(clk), .RST(rst), .Q(sreg[1138])
         );
  DFF \sreg_reg[1139]  ( .D(swire[116]), .CLK(clk), .RST(rst), .Q(sreg[1139])
         );
  DFF \sreg_reg[1140]  ( .D(swire[117]), .CLK(clk), .RST(rst), .Q(sreg[1140])
         );
  DFF \sreg_reg[1141]  ( .D(swire[118]), .CLK(clk), .RST(rst), .Q(sreg[1141])
         );
  DFF \sreg_reg[1142]  ( .D(swire[119]), .CLK(clk), .RST(rst), .Q(sreg[1142])
         );
  DFF \sreg_reg[1143]  ( .D(swire[120]), .CLK(clk), .RST(rst), .Q(sreg[1143])
         );
  DFF \sreg_reg[1144]  ( .D(swire[121]), .CLK(clk), .RST(rst), .Q(sreg[1144])
         );
  DFF \sreg_reg[1145]  ( .D(swire[122]), .CLK(clk), .RST(rst), .Q(sreg[1145])
         );
  DFF \sreg_reg[1146]  ( .D(swire[123]), .CLK(clk), .RST(rst), .Q(sreg[1146])
         );
  DFF \sreg_reg[1147]  ( .D(swire[124]), .CLK(clk), .RST(rst), .Q(sreg[1147])
         );
  DFF \sreg_reg[1148]  ( .D(swire[125]), .CLK(clk), .RST(rst), .Q(sreg[1148])
         );
  DFF \sreg_reg[1149]  ( .D(swire[126]), .CLK(clk), .RST(rst), .Q(sreg[1149])
         );
  DFF \sreg_reg[1150]  ( .D(swire[127]), .CLK(clk), .RST(rst), .Q(sreg[1150])
         );
  DFF \sreg_reg[1151]  ( .D(swire[128]), .CLK(clk), .RST(rst), .Q(sreg[1151])
         );
  DFF \sreg_reg[1152]  ( .D(swire[129]), .CLK(clk), .RST(rst), .Q(sreg[1152])
         );
  DFF \sreg_reg[1153]  ( .D(swire[130]), .CLK(clk), .RST(rst), .Q(sreg[1153])
         );
  DFF \sreg_reg[1154]  ( .D(swire[131]), .CLK(clk), .RST(rst), .Q(sreg[1154])
         );
  DFF \sreg_reg[1155]  ( .D(swire[132]), .CLK(clk), .RST(rst), .Q(sreg[1155])
         );
  DFF \sreg_reg[1156]  ( .D(swire[133]), .CLK(clk), .RST(rst), .Q(sreg[1156])
         );
  DFF \sreg_reg[1157]  ( .D(swire[134]), .CLK(clk), .RST(rst), .Q(sreg[1157])
         );
  DFF \sreg_reg[1158]  ( .D(swire[135]), .CLK(clk), .RST(rst), .Q(sreg[1158])
         );
  DFF \sreg_reg[1159]  ( .D(swire[136]), .CLK(clk), .RST(rst), .Q(sreg[1159])
         );
  DFF \sreg_reg[1160]  ( .D(swire[137]), .CLK(clk), .RST(rst), .Q(sreg[1160])
         );
  DFF \sreg_reg[1161]  ( .D(swire[138]), .CLK(clk), .RST(rst), .Q(sreg[1161])
         );
  DFF \sreg_reg[1162]  ( .D(swire[139]), .CLK(clk), .RST(rst), .Q(sreg[1162])
         );
  DFF \sreg_reg[1163]  ( .D(swire[140]), .CLK(clk), .RST(rst), .Q(sreg[1163])
         );
  DFF \sreg_reg[1164]  ( .D(swire[141]), .CLK(clk), .RST(rst), .Q(sreg[1164])
         );
  DFF \sreg_reg[1165]  ( .D(swire[142]), .CLK(clk), .RST(rst), .Q(sreg[1165])
         );
  DFF \sreg_reg[1166]  ( .D(swire[143]), .CLK(clk), .RST(rst), .Q(sreg[1166])
         );
  DFF \sreg_reg[1167]  ( .D(swire[144]), .CLK(clk), .RST(rst), .Q(sreg[1167])
         );
  DFF \sreg_reg[1168]  ( .D(swire[145]), .CLK(clk), .RST(rst), .Q(sreg[1168])
         );
  DFF \sreg_reg[1169]  ( .D(swire[146]), .CLK(clk), .RST(rst), .Q(sreg[1169])
         );
  DFF \sreg_reg[1170]  ( .D(swire[147]), .CLK(clk), .RST(rst), .Q(sreg[1170])
         );
  DFF \sreg_reg[1171]  ( .D(swire[148]), .CLK(clk), .RST(rst), .Q(sreg[1171])
         );
  DFF \sreg_reg[1172]  ( .D(swire[149]), .CLK(clk), .RST(rst), .Q(sreg[1172])
         );
  DFF \sreg_reg[1173]  ( .D(swire[150]), .CLK(clk), .RST(rst), .Q(sreg[1173])
         );
  DFF \sreg_reg[1174]  ( .D(swire[151]), .CLK(clk), .RST(rst), .Q(sreg[1174])
         );
  DFF \sreg_reg[1175]  ( .D(swire[152]), .CLK(clk), .RST(rst), .Q(sreg[1175])
         );
  DFF \sreg_reg[1176]  ( .D(swire[153]), .CLK(clk), .RST(rst), .Q(sreg[1176])
         );
  DFF \sreg_reg[1177]  ( .D(swire[154]), .CLK(clk), .RST(rst), .Q(sreg[1177])
         );
  DFF \sreg_reg[1178]  ( .D(swire[155]), .CLK(clk), .RST(rst), .Q(sreg[1178])
         );
  DFF \sreg_reg[1179]  ( .D(swire[156]), .CLK(clk), .RST(rst), .Q(sreg[1179])
         );
  DFF \sreg_reg[1180]  ( .D(swire[157]), .CLK(clk), .RST(rst), .Q(sreg[1180])
         );
  DFF \sreg_reg[1181]  ( .D(swire[158]), .CLK(clk), .RST(rst), .Q(sreg[1181])
         );
  DFF \sreg_reg[1182]  ( .D(swire[159]), .CLK(clk), .RST(rst), .Q(sreg[1182])
         );
  DFF \sreg_reg[1183]  ( .D(swire[160]), .CLK(clk), .RST(rst), .Q(sreg[1183])
         );
  DFF \sreg_reg[1184]  ( .D(swire[161]), .CLK(clk), .RST(rst), .Q(sreg[1184])
         );
  DFF \sreg_reg[1185]  ( .D(swire[162]), .CLK(clk), .RST(rst), .Q(sreg[1185])
         );
  DFF \sreg_reg[1186]  ( .D(swire[163]), .CLK(clk), .RST(rst), .Q(sreg[1186])
         );
  DFF \sreg_reg[1187]  ( .D(swire[164]), .CLK(clk), .RST(rst), .Q(sreg[1187])
         );
  DFF \sreg_reg[1188]  ( .D(swire[165]), .CLK(clk), .RST(rst), .Q(sreg[1188])
         );
  DFF \sreg_reg[1189]  ( .D(swire[166]), .CLK(clk), .RST(rst), .Q(sreg[1189])
         );
  DFF \sreg_reg[1190]  ( .D(swire[167]), .CLK(clk), .RST(rst), .Q(sreg[1190])
         );
  DFF \sreg_reg[1191]  ( .D(swire[168]), .CLK(clk), .RST(rst), .Q(sreg[1191])
         );
  DFF \sreg_reg[1192]  ( .D(swire[169]), .CLK(clk), .RST(rst), .Q(sreg[1192])
         );
  DFF \sreg_reg[1193]  ( .D(swire[170]), .CLK(clk), .RST(rst), .Q(sreg[1193])
         );
  DFF \sreg_reg[1194]  ( .D(swire[171]), .CLK(clk), .RST(rst), .Q(sreg[1194])
         );
  DFF \sreg_reg[1195]  ( .D(swire[172]), .CLK(clk), .RST(rst), .Q(sreg[1195])
         );
  DFF \sreg_reg[1196]  ( .D(swire[173]), .CLK(clk), .RST(rst), .Q(sreg[1196])
         );
  DFF \sreg_reg[1197]  ( .D(swire[174]), .CLK(clk), .RST(rst), .Q(sreg[1197])
         );
  DFF \sreg_reg[1198]  ( .D(swire[175]), .CLK(clk), .RST(rst), .Q(sreg[1198])
         );
  DFF \sreg_reg[1199]  ( .D(swire[176]), .CLK(clk), .RST(rst), .Q(sreg[1199])
         );
  DFF \sreg_reg[1200]  ( .D(swire[177]), .CLK(clk), .RST(rst), .Q(sreg[1200])
         );
  DFF \sreg_reg[1201]  ( .D(swire[178]), .CLK(clk), .RST(rst), .Q(sreg[1201])
         );
  DFF \sreg_reg[1202]  ( .D(swire[179]), .CLK(clk), .RST(rst), .Q(sreg[1202])
         );
  DFF \sreg_reg[1203]  ( .D(swire[180]), .CLK(clk), .RST(rst), .Q(sreg[1203])
         );
  DFF \sreg_reg[1204]  ( .D(swire[181]), .CLK(clk), .RST(rst), .Q(sreg[1204])
         );
  DFF \sreg_reg[1205]  ( .D(swire[182]), .CLK(clk), .RST(rst), .Q(sreg[1205])
         );
  DFF \sreg_reg[1206]  ( .D(swire[183]), .CLK(clk), .RST(rst), .Q(sreg[1206])
         );
  DFF \sreg_reg[1207]  ( .D(swire[184]), .CLK(clk), .RST(rst), .Q(sreg[1207])
         );
  DFF \sreg_reg[1208]  ( .D(swire[185]), .CLK(clk), .RST(rst), .Q(sreg[1208])
         );
  DFF \sreg_reg[1209]  ( .D(swire[186]), .CLK(clk), .RST(rst), .Q(sreg[1209])
         );
  DFF \sreg_reg[1210]  ( .D(swire[187]), .CLK(clk), .RST(rst), .Q(sreg[1210])
         );
  DFF \sreg_reg[1211]  ( .D(swire[188]), .CLK(clk), .RST(rst), .Q(sreg[1211])
         );
  DFF \sreg_reg[1212]  ( .D(swire[189]), .CLK(clk), .RST(rst), .Q(sreg[1212])
         );
  DFF \sreg_reg[1213]  ( .D(swire[190]), .CLK(clk), .RST(rst), .Q(sreg[1213])
         );
  DFF \sreg_reg[1214]  ( .D(swire[191]), .CLK(clk), .RST(rst), .Q(sreg[1214])
         );
  DFF \sreg_reg[1215]  ( .D(swire[192]), .CLK(clk), .RST(rst), .Q(sreg[1215])
         );
  DFF \sreg_reg[1216]  ( .D(swire[193]), .CLK(clk), .RST(rst), .Q(sreg[1216])
         );
  DFF \sreg_reg[1217]  ( .D(swire[194]), .CLK(clk), .RST(rst), .Q(sreg[1217])
         );
  DFF \sreg_reg[1218]  ( .D(swire[195]), .CLK(clk), .RST(rst), .Q(sreg[1218])
         );
  DFF \sreg_reg[1219]  ( .D(swire[196]), .CLK(clk), .RST(rst), .Q(sreg[1219])
         );
  DFF \sreg_reg[1220]  ( .D(swire[197]), .CLK(clk), .RST(rst), .Q(sreg[1220])
         );
  DFF \sreg_reg[1221]  ( .D(swire[198]), .CLK(clk), .RST(rst), .Q(sreg[1221])
         );
  DFF \sreg_reg[1222]  ( .D(swire[199]), .CLK(clk), .RST(rst), .Q(sreg[1222])
         );
  DFF \sreg_reg[1223]  ( .D(swire[200]), .CLK(clk), .RST(rst), .Q(sreg[1223])
         );
  DFF \sreg_reg[1224]  ( .D(swire[201]), .CLK(clk), .RST(rst), .Q(sreg[1224])
         );
  DFF \sreg_reg[1225]  ( .D(swire[202]), .CLK(clk), .RST(rst), .Q(sreg[1225])
         );
  DFF \sreg_reg[1226]  ( .D(swire[203]), .CLK(clk), .RST(rst), .Q(sreg[1226])
         );
  DFF \sreg_reg[1227]  ( .D(swire[204]), .CLK(clk), .RST(rst), .Q(sreg[1227])
         );
  DFF \sreg_reg[1228]  ( .D(swire[205]), .CLK(clk), .RST(rst), .Q(sreg[1228])
         );
  DFF \sreg_reg[1229]  ( .D(swire[206]), .CLK(clk), .RST(rst), .Q(sreg[1229])
         );
  DFF \sreg_reg[1230]  ( .D(swire[207]), .CLK(clk), .RST(rst), .Q(sreg[1230])
         );
  DFF \sreg_reg[1231]  ( .D(swire[208]), .CLK(clk), .RST(rst), .Q(sreg[1231])
         );
  DFF \sreg_reg[1232]  ( .D(swire[209]), .CLK(clk), .RST(rst), .Q(sreg[1232])
         );
  DFF \sreg_reg[1233]  ( .D(swire[210]), .CLK(clk), .RST(rst), .Q(sreg[1233])
         );
  DFF \sreg_reg[1234]  ( .D(swire[211]), .CLK(clk), .RST(rst), .Q(sreg[1234])
         );
  DFF \sreg_reg[1235]  ( .D(swire[212]), .CLK(clk), .RST(rst), .Q(sreg[1235])
         );
  DFF \sreg_reg[1236]  ( .D(swire[213]), .CLK(clk), .RST(rst), .Q(sreg[1236])
         );
  DFF \sreg_reg[1237]  ( .D(swire[214]), .CLK(clk), .RST(rst), .Q(sreg[1237])
         );
  DFF \sreg_reg[1238]  ( .D(swire[215]), .CLK(clk), .RST(rst), .Q(sreg[1238])
         );
  DFF \sreg_reg[1239]  ( .D(swire[216]), .CLK(clk), .RST(rst), .Q(sreg[1239])
         );
  DFF \sreg_reg[1240]  ( .D(swire[217]), .CLK(clk), .RST(rst), .Q(sreg[1240])
         );
  DFF \sreg_reg[1241]  ( .D(swire[218]), .CLK(clk), .RST(rst), .Q(sreg[1241])
         );
  DFF \sreg_reg[1242]  ( .D(swire[219]), .CLK(clk), .RST(rst), .Q(sreg[1242])
         );
  DFF \sreg_reg[1243]  ( .D(swire[220]), .CLK(clk), .RST(rst), .Q(sreg[1243])
         );
  DFF \sreg_reg[1244]  ( .D(swire[221]), .CLK(clk), .RST(rst), .Q(sreg[1244])
         );
  DFF \sreg_reg[1245]  ( .D(swire[222]), .CLK(clk), .RST(rst), .Q(sreg[1245])
         );
  DFF \sreg_reg[1246]  ( .D(swire[223]), .CLK(clk), .RST(rst), .Q(sreg[1246])
         );
  DFF \sreg_reg[1247]  ( .D(swire[224]), .CLK(clk), .RST(rst), .Q(sreg[1247])
         );
  DFF \sreg_reg[1248]  ( .D(swire[225]), .CLK(clk), .RST(rst), .Q(sreg[1248])
         );
  DFF \sreg_reg[1249]  ( .D(swire[226]), .CLK(clk), .RST(rst), .Q(sreg[1249])
         );
  DFF \sreg_reg[1250]  ( .D(swire[227]), .CLK(clk), .RST(rst), .Q(sreg[1250])
         );
  DFF \sreg_reg[1251]  ( .D(swire[228]), .CLK(clk), .RST(rst), .Q(sreg[1251])
         );
  DFF \sreg_reg[1252]  ( .D(swire[229]), .CLK(clk), .RST(rst), .Q(sreg[1252])
         );
  DFF \sreg_reg[1253]  ( .D(swire[230]), .CLK(clk), .RST(rst), .Q(sreg[1253])
         );
  DFF \sreg_reg[1254]  ( .D(swire[231]), .CLK(clk), .RST(rst), .Q(sreg[1254])
         );
  DFF \sreg_reg[1255]  ( .D(swire[232]), .CLK(clk), .RST(rst), .Q(sreg[1255])
         );
  DFF \sreg_reg[1256]  ( .D(swire[233]), .CLK(clk), .RST(rst), .Q(sreg[1256])
         );
  DFF \sreg_reg[1257]  ( .D(swire[234]), .CLK(clk), .RST(rst), .Q(sreg[1257])
         );
  DFF \sreg_reg[1258]  ( .D(swire[235]), .CLK(clk), .RST(rst), .Q(sreg[1258])
         );
  DFF \sreg_reg[1259]  ( .D(swire[236]), .CLK(clk), .RST(rst), .Q(sreg[1259])
         );
  DFF \sreg_reg[1260]  ( .D(swire[237]), .CLK(clk), .RST(rst), .Q(sreg[1260])
         );
  DFF \sreg_reg[1261]  ( .D(swire[238]), .CLK(clk), .RST(rst), .Q(sreg[1261])
         );
  DFF \sreg_reg[1262]  ( .D(swire[239]), .CLK(clk), .RST(rst), .Q(sreg[1262])
         );
  DFF \sreg_reg[1263]  ( .D(swire[240]), .CLK(clk), .RST(rst), .Q(sreg[1263])
         );
  DFF \sreg_reg[1264]  ( .D(swire[241]), .CLK(clk), .RST(rst), .Q(sreg[1264])
         );
  DFF \sreg_reg[1265]  ( .D(swire[242]), .CLK(clk), .RST(rst), .Q(sreg[1265])
         );
  DFF \sreg_reg[1266]  ( .D(swire[243]), .CLK(clk), .RST(rst), .Q(sreg[1266])
         );
  DFF \sreg_reg[1267]  ( .D(swire[244]), .CLK(clk), .RST(rst), .Q(sreg[1267])
         );
  DFF \sreg_reg[1268]  ( .D(swire[245]), .CLK(clk), .RST(rst), .Q(sreg[1268])
         );
  DFF \sreg_reg[1269]  ( .D(swire[246]), .CLK(clk), .RST(rst), .Q(sreg[1269])
         );
  DFF \sreg_reg[1270]  ( .D(swire[247]), .CLK(clk), .RST(rst), .Q(sreg[1270])
         );
  DFF \sreg_reg[1271]  ( .D(swire[248]), .CLK(clk), .RST(rst), .Q(sreg[1271])
         );
  DFF \sreg_reg[1272]  ( .D(swire[249]), .CLK(clk), .RST(rst), .Q(sreg[1272])
         );
  DFF \sreg_reg[1273]  ( .D(swire[250]), .CLK(clk), .RST(rst), .Q(sreg[1273])
         );
  DFF \sreg_reg[1274]  ( .D(swire[251]), .CLK(clk), .RST(rst), .Q(sreg[1274])
         );
  DFF \sreg_reg[1275]  ( .D(swire[252]), .CLK(clk), .RST(rst), .Q(sreg[1275])
         );
  DFF \sreg_reg[1276]  ( .D(swire[253]), .CLK(clk), .RST(rst), .Q(sreg[1276])
         );
  DFF \sreg_reg[1277]  ( .D(swire[254]), .CLK(clk), .RST(rst), .Q(sreg[1277])
         );
  DFF \sreg_reg[1278]  ( .D(swire[255]), .CLK(clk), .RST(rst), .Q(sreg[1278])
         );
  DFF \sreg_reg[1279]  ( .D(swire[256]), .CLK(clk), .RST(rst), .Q(sreg[1279])
         );
  DFF \sreg_reg[1280]  ( .D(swire[257]), .CLK(clk), .RST(rst), .Q(sreg[1280])
         );
  DFF \sreg_reg[1281]  ( .D(swire[258]), .CLK(clk), .RST(rst), .Q(sreg[1281])
         );
  DFF \sreg_reg[1282]  ( .D(swire[259]), .CLK(clk), .RST(rst), .Q(sreg[1282])
         );
  DFF \sreg_reg[1283]  ( .D(swire[260]), .CLK(clk), .RST(rst), .Q(sreg[1283])
         );
  DFF \sreg_reg[1284]  ( .D(swire[261]), .CLK(clk), .RST(rst), .Q(sreg[1284])
         );
  DFF \sreg_reg[1285]  ( .D(swire[262]), .CLK(clk), .RST(rst), .Q(sreg[1285])
         );
  DFF \sreg_reg[1286]  ( .D(swire[263]), .CLK(clk), .RST(rst), .Q(sreg[1286])
         );
  DFF \sreg_reg[1287]  ( .D(swire[264]), .CLK(clk), .RST(rst), .Q(sreg[1287])
         );
  DFF \sreg_reg[1288]  ( .D(swire[265]), .CLK(clk), .RST(rst), .Q(sreg[1288])
         );
  DFF \sreg_reg[1289]  ( .D(swire[266]), .CLK(clk), .RST(rst), .Q(sreg[1289])
         );
  DFF \sreg_reg[1290]  ( .D(swire[267]), .CLK(clk), .RST(rst), .Q(sreg[1290])
         );
  DFF \sreg_reg[1291]  ( .D(swire[268]), .CLK(clk), .RST(rst), .Q(sreg[1291])
         );
  DFF \sreg_reg[1292]  ( .D(swire[269]), .CLK(clk), .RST(rst), .Q(sreg[1292])
         );
  DFF \sreg_reg[1293]  ( .D(swire[270]), .CLK(clk), .RST(rst), .Q(sreg[1293])
         );
  DFF \sreg_reg[1294]  ( .D(swire[271]), .CLK(clk), .RST(rst), .Q(sreg[1294])
         );
  DFF \sreg_reg[1295]  ( .D(swire[272]), .CLK(clk), .RST(rst), .Q(sreg[1295])
         );
  DFF \sreg_reg[1296]  ( .D(swire[273]), .CLK(clk), .RST(rst), .Q(sreg[1296])
         );
  DFF \sreg_reg[1297]  ( .D(swire[274]), .CLK(clk), .RST(rst), .Q(sreg[1297])
         );
  DFF \sreg_reg[1298]  ( .D(swire[275]), .CLK(clk), .RST(rst), .Q(sreg[1298])
         );
  DFF \sreg_reg[1299]  ( .D(swire[276]), .CLK(clk), .RST(rst), .Q(sreg[1299])
         );
  DFF \sreg_reg[1300]  ( .D(swire[277]), .CLK(clk), .RST(rst), .Q(sreg[1300])
         );
  DFF \sreg_reg[1301]  ( .D(swire[278]), .CLK(clk), .RST(rst), .Q(sreg[1301])
         );
  DFF \sreg_reg[1302]  ( .D(swire[279]), .CLK(clk), .RST(rst), .Q(sreg[1302])
         );
  DFF \sreg_reg[1303]  ( .D(swire[280]), .CLK(clk), .RST(rst), .Q(sreg[1303])
         );
  DFF \sreg_reg[1304]  ( .D(swire[281]), .CLK(clk), .RST(rst), .Q(sreg[1304])
         );
  DFF \sreg_reg[1305]  ( .D(swire[282]), .CLK(clk), .RST(rst), .Q(sreg[1305])
         );
  DFF \sreg_reg[1306]  ( .D(swire[283]), .CLK(clk), .RST(rst), .Q(sreg[1306])
         );
  DFF \sreg_reg[1307]  ( .D(swire[284]), .CLK(clk), .RST(rst), .Q(sreg[1307])
         );
  DFF \sreg_reg[1308]  ( .D(swire[285]), .CLK(clk), .RST(rst), .Q(sreg[1308])
         );
  DFF \sreg_reg[1309]  ( .D(swire[286]), .CLK(clk), .RST(rst), .Q(sreg[1309])
         );
  DFF \sreg_reg[1310]  ( .D(swire[287]), .CLK(clk), .RST(rst), .Q(sreg[1310])
         );
  DFF \sreg_reg[1311]  ( .D(swire[288]), .CLK(clk), .RST(rst), .Q(sreg[1311])
         );
  DFF \sreg_reg[1312]  ( .D(swire[289]), .CLK(clk), .RST(rst), .Q(sreg[1312])
         );
  DFF \sreg_reg[1313]  ( .D(swire[290]), .CLK(clk), .RST(rst), .Q(sreg[1313])
         );
  DFF \sreg_reg[1314]  ( .D(swire[291]), .CLK(clk), .RST(rst), .Q(sreg[1314])
         );
  DFF \sreg_reg[1315]  ( .D(swire[292]), .CLK(clk), .RST(rst), .Q(sreg[1315])
         );
  DFF \sreg_reg[1316]  ( .D(swire[293]), .CLK(clk), .RST(rst), .Q(sreg[1316])
         );
  DFF \sreg_reg[1317]  ( .D(swire[294]), .CLK(clk), .RST(rst), .Q(sreg[1317])
         );
  DFF \sreg_reg[1318]  ( .D(swire[295]), .CLK(clk), .RST(rst), .Q(sreg[1318])
         );
  DFF \sreg_reg[1319]  ( .D(swire[296]), .CLK(clk), .RST(rst), .Q(sreg[1319])
         );
  DFF \sreg_reg[1320]  ( .D(swire[297]), .CLK(clk), .RST(rst), .Q(sreg[1320])
         );
  DFF \sreg_reg[1321]  ( .D(swire[298]), .CLK(clk), .RST(rst), .Q(sreg[1321])
         );
  DFF \sreg_reg[1322]  ( .D(swire[299]), .CLK(clk), .RST(rst), .Q(sreg[1322])
         );
  DFF \sreg_reg[1323]  ( .D(swire[300]), .CLK(clk), .RST(rst), .Q(sreg[1323])
         );
  DFF \sreg_reg[1324]  ( .D(swire[301]), .CLK(clk), .RST(rst), .Q(sreg[1324])
         );
  DFF \sreg_reg[1325]  ( .D(swire[302]), .CLK(clk), .RST(rst), .Q(sreg[1325])
         );
  DFF \sreg_reg[1326]  ( .D(swire[303]), .CLK(clk), .RST(rst), .Q(sreg[1326])
         );
  DFF \sreg_reg[1327]  ( .D(swire[304]), .CLK(clk), .RST(rst), .Q(sreg[1327])
         );
  DFF \sreg_reg[1328]  ( .D(swire[305]), .CLK(clk), .RST(rst), .Q(sreg[1328])
         );
  DFF \sreg_reg[1329]  ( .D(swire[306]), .CLK(clk), .RST(rst), .Q(sreg[1329])
         );
  DFF \sreg_reg[1330]  ( .D(swire[307]), .CLK(clk), .RST(rst), .Q(sreg[1330])
         );
  DFF \sreg_reg[1331]  ( .D(swire[308]), .CLK(clk), .RST(rst), .Q(sreg[1331])
         );
  DFF \sreg_reg[1332]  ( .D(swire[309]), .CLK(clk), .RST(rst), .Q(sreg[1332])
         );
  DFF \sreg_reg[1333]  ( .D(swire[310]), .CLK(clk), .RST(rst), .Q(sreg[1333])
         );
  DFF \sreg_reg[1334]  ( .D(swire[311]), .CLK(clk), .RST(rst), .Q(sreg[1334])
         );
  DFF \sreg_reg[1335]  ( .D(swire[312]), .CLK(clk), .RST(rst), .Q(sreg[1335])
         );
  DFF \sreg_reg[1336]  ( .D(swire[313]), .CLK(clk), .RST(rst), .Q(sreg[1336])
         );
  DFF \sreg_reg[1337]  ( .D(swire[314]), .CLK(clk), .RST(rst), .Q(sreg[1337])
         );
  DFF \sreg_reg[1338]  ( .D(swire[315]), .CLK(clk), .RST(rst), .Q(sreg[1338])
         );
  DFF \sreg_reg[1339]  ( .D(swire[316]), .CLK(clk), .RST(rst), .Q(sreg[1339])
         );
  DFF \sreg_reg[1340]  ( .D(swire[317]), .CLK(clk), .RST(rst), .Q(sreg[1340])
         );
  DFF \sreg_reg[1341]  ( .D(swire[318]), .CLK(clk), .RST(rst), .Q(sreg[1341])
         );
  DFF \sreg_reg[1342]  ( .D(swire[319]), .CLK(clk), .RST(rst), .Q(sreg[1342])
         );
  DFF \sreg_reg[1343]  ( .D(swire[320]), .CLK(clk), .RST(rst), .Q(sreg[1343])
         );
  DFF \sreg_reg[1344]  ( .D(swire[321]), .CLK(clk), .RST(rst), .Q(sreg[1344])
         );
  DFF \sreg_reg[1345]  ( .D(swire[322]), .CLK(clk), .RST(rst), .Q(sreg[1345])
         );
  DFF \sreg_reg[1346]  ( .D(swire[323]), .CLK(clk), .RST(rst), .Q(sreg[1346])
         );
  DFF \sreg_reg[1347]  ( .D(swire[324]), .CLK(clk), .RST(rst), .Q(sreg[1347])
         );
  DFF \sreg_reg[1348]  ( .D(swire[325]), .CLK(clk), .RST(rst), .Q(sreg[1348])
         );
  DFF \sreg_reg[1349]  ( .D(swire[326]), .CLK(clk), .RST(rst), .Q(sreg[1349])
         );
  DFF \sreg_reg[1350]  ( .D(swire[327]), .CLK(clk), .RST(rst), .Q(sreg[1350])
         );
  DFF \sreg_reg[1351]  ( .D(swire[328]), .CLK(clk), .RST(rst), .Q(sreg[1351])
         );
  DFF \sreg_reg[1352]  ( .D(swire[329]), .CLK(clk), .RST(rst), .Q(sreg[1352])
         );
  DFF \sreg_reg[1353]  ( .D(swire[330]), .CLK(clk), .RST(rst), .Q(sreg[1353])
         );
  DFF \sreg_reg[1354]  ( .D(swire[331]), .CLK(clk), .RST(rst), .Q(sreg[1354])
         );
  DFF \sreg_reg[1355]  ( .D(swire[332]), .CLK(clk), .RST(rst), .Q(sreg[1355])
         );
  DFF \sreg_reg[1356]  ( .D(swire[333]), .CLK(clk), .RST(rst), .Q(sreg[1356])
         );
  DFF \sreg_reg[1357]  ( .D(swire[334]), .CLK(clk), .RST(rst), .Q(sreg[1357])
         );
  DFF \sreg_reg[1358]  ( .D(swire[335]), .CLK(clk), .RST(rst), .Q(sreg[1358])
         );
  DFF \sreg_reg[1359]  ( .D(swire[336]), .CLK(clk), .RST(rst), .Q(sreg[1359])
         );
  DFF \sreg_reg[1360]  ( .D(swire[337]), .CLK(clk), .RST(rst), .Q(sreg[1360])
         );
  DFF \sreg_reg[1361]  ( .D(swire[338]), .CLK(clk), .RST(rst), .Q(sreg[1361])
         );
  DFF \sreg_reg[1362]  ( .D(swire[339]), .CLK(clk), .RST(rst), .Q(sreg[1362])
         );
  DFF \sreg_reg[1363]  ( .D(swire[340]), .CLK(clk), .RST(rst), .Q(sreg[1363])
         );
  DFF \sreg_reg[1364]  ( .D(swire[341]), .CLK(clk), .RST(rst), .Q(sreg[1364])
         );
  DFF \sreg_reg[1365]  ( .D(swire[342]), .CLK(clk), .RST(rst), .Q(sreg[1365])
         );
  DFF \sreg_reg[1366]  ( .D(swire[343]), .CLK(clk), .RST(rst), .Q(sreg[1366])
         );
  DFF \sreg_reg[1367]  ( .D(swire[344]), .CLK(clk), .RST(rst), .Q(sreg[1367])
         );
  DFF \sreg_reg[1368]  ( .D(swire[345]), .CLK(clk), .RST(rst), .Q(sreg[1368])
         );
  DFF \sreg_reg[1369]  ( .D(swire[346]), .CLK(clk), .RST(rst), .Q(sreg[1369])
         );
  DFF \sreg_reg[1370]  ( .D(swire[347]), .CLK(clk), .RST(rst), .Q(sreg[1370])
         );
  DFF \sreg_reg[1371]  ( .D(swire[348]), .CLK(clk), .RST(rst), .Q(sreg[1371])
         );
  DFF \sreg_reg[1372]  ( .D(swire[349]), .CLK(clk), .RST(rst), .Q(sreg[1372])
         );
  DFF \sreg_reg[1373]  ( .D(swire[350]), .CLK(clk), .RST(rst), .Q(sreg[1373])
         );
  DFF \sreg_reg[1374]  ( .D(swire[351]), .CLK(clk), .RST(rst), .Q(sreg[1374])
         );
  DFF \sreg_reg[1375]  ( .D(swire[352]), .CLK(clk), .RST(rst), .Q(sreg[1375])
         );
  DFF \sreg_reg[1376]  ( .D(swire[353]), .CLK(clk), .RST(rst), .Q(sreg[1376])
         );
  DFF \sreg_reg[1377]  ( .D(swire[354]), .CLK(clk), .RST(rst), .Q(sreg[1377])
         );
  DFF \sreg_reg[1378]  ( .D(swire[355]), .CLK(clk), .RST(rst), .Q(sreg[1378])
         );
  DFF \sreg_reg[1379]  ( .D(swire[356]), .CLK(clk), .RST(rst), .Q(sreg[1379])
         );
  DFF \sreg_reg[1380]  ( .D(swire[357]), .CLK(clk), .RST(rst), .Q(sreg[1380])
         );
  DFF \sreg_reg[1381]  ( .D(swire[358]), .CLK(clk), .RST(rst), .Q(sreg[1381])
         );
  DFF \sreg_reg[1382]  ( .D(swire[359]), .CLK(clk), .RST(rst), .Q(sreg[1382])
         );
  DFF \sreg_reg[1383]  ( .D(swire[360]), .CLK(clk), .RST(rst), .Q(sreg[1383])
         );
  DFF \sreg_reg[1384]  ( .D(swire[361]), .CLK(clk), .RST(rst), .Q(sreg[1384])
         );
  DFF \sreg_reg[1385]  ( .D(swire[362]), .CLK(clk), .RST(rst), .Q(sreg[1385])
         );
  DFF \sreg_reg[1386]  ( .D(swire[363]), .CLK(clk), .RST(rst), .Q(sreg[1386])
         );
  DFF \sreg_reg[1387]  ( .D(swire[364]), .CLK(clk), .RST(rst), .Q(sreg[1387])
         );
  DFF \sreg_reg[1388]  ( .D(swire[365]), .CLK(clk), .RST(rst), .Q(sreg[1388])
         );
  DFF \sreg_reg[1389]  ( .D(swire[366]), .CLK(clk), .RST(rst), .Q(sreg[1389])
         );
  DFF \sreg_reg[1390]  ( .D(swire[367]), .CLK(clk), .RST(rst), .Q(sreg[1390])
         );
  DFF \sreg_reg[1391]  ( .D(swire[368]), .CLK(clk), .RST(rst), .Q(sreg[1391])
         );
  DFF \sreg_reg[1392]  ( .D(swire[369]), .CLK(clk), .RST(rst), .Q(sreg[1392])
         );
  DFF \sreg_reg[1393]  ( .D(swire[370]), .CLK(clk), .RST(rst), .Q(sreg[1393])
         );
  DFF \sreg_reg[1394]  ( .D(swire[371]), .CLK(clk), .RST(rst), .Q(sreg[1394])
         );
  DFF \sreg_reg[1395]  ( .D(swire[372]), .CLK(clk), .RST(rst), .Q(sreg[1395])
         );
  DFF \sreg_reg[1396]  ( .D(swire[373]), .CLK(clk), .RST(rst), .Q(sreg[1396])
         );
  DFF \sreg_reg[1397]  ( .D(swire[374]), .CLK(clk), .RST(rst), .Q(sreg[1397])
         );
  DFF \sreg_reg[1398]  ( .D(swire[375]), .CLK(clk), .RST(rst), .Q(sreg[1398])
         );
  DFF \sreg_reg[1399]  ( .D(swire[376]), .CLK(clk), .RST(rst), .Q(sreg[1399])
         );
  DFF \sreg_reg[1400]  ( .D(swire[377]), .CLK(clk), .RST(rst), .Q(sreg[1400])
         );
  DFF \sreg_reg[1401]  ( .D(swire[378]), .CLK(clk), .RST(rst), .Q(sreg[1401])
         );
  DFF \sreg_reg[1402]  ( .D(swire[379]), .CLK(clk), .RST(rst), .Q(sreg[1402])
         );
  DFF \sreg_reg[1403]  ( .D(swire[380]), .CLK(clk), .RST(rst), .Q(sreg[1403])
         );
  DFF \sreg_reg[1404]  ( .D(swire[381]), .CLK(clk), .RST(rst), .Q(sreg[1404])
         );
  DFF \sreg_reg[1405]  ( .D(swire[382]), .CLK(clk), .RST(rst), .Q(sreg[1405])
         );
  DFF \sreg_reg[1406]  ( .D(swire[383]), .CLK(clk), .RST(rst), .Q(sreg[1406])
         );
  DFF \sreg_reg[1407]  ( .D(swire[384]), .CLK(clk), .RST(rst), .Q(sreg[1407])
         );
  DFF \sreg_reg[1408]  ( .D(swire[385]), .CLK(clk), .RST(rst), .Q(sreg[1408])
         );
  DFF \sreg_reg[1409]  ( .D(swire[386]), .CLK(clk), .RST(rst), .Q(sreg[1409])
         );
  DFF \sreg_reg[1410]  ( .D(swire[387]), .CLK(clk), .RST(rst), .Q(sreg[1410])
         );
  DFF \sreg_reg[1411]  ( .D(swire[388]), .CLK(clk), .RST(rst), .Q(sreg[1411])
         );
  DFF \sreg_reg[1412]  ( .D(swire[389]), .CLK(clk), .RST(rst), .Q(sreg[1412])
         );
  DFF \sreg_reg[1413]  ( .D(swire[390]), .CLK(clk), .RST(rst), .Q(sreg[1413])
         );
  DFF \sreg_reg[1414]  ( .D(swire[391]), .CLK(clk), .RST(rst), .Q(sreg[1414])
         );
  DFF \sreg_reg[1415]  ( .D(swire[392]), .CLK(clk), .RST(rst), .Q(sreg[1415])
         );
  DFF \sreg_reg[1416]  ( .D(swire[393]), .CLK(clk), .RST(rst), .Q(sreg[1416])
         );
  DFF \sreg_reg[1417]  ( .D(swire[394]), .CLK(clk), .RST(rst), .Q(sreg[1417])
         );
  DFF \sreg_reg[1418]  ( .D(swire[395]), .CLK(clk), .RST(rst), .Q(sreg[1418])
         );
  DFF \sreg_reg[1419]  ( .D(swire[396]), .CLK(clk), .RST(rst), .Q(sreg[1419])
         );
  DFF \sreg_reg[1420]  ( .D(swire[397]), .CLK(clk), .RST(rst), .Q(sreg[1420])
         );
  DFF \sreg_reg[1421]  ( .D(swire[398]), .CLK(clk), .RST(rst), .Q(sreg[1421])
         );
  DFF \sreg_reg[1422]  ( .D(swire[399]), .CLK(clk), .RST(rst), .Q(sreg[1422])
         );
  DFF \sreg_reg[1423]  ( .D(swire[400]), .CLK(clk), .RST(rst), .Q(sreg[1423])
         );
  DFF \sreg_reg[1424]  ( .D(swire[401]), .CLK(clk), .RST(rst), .Q(sreg[1424])
         );
  DFF \sreg_reg[1425]  ( .D(swire[402]), .CLK(clk), .RST(rst), .Q(sreg[1425])
         );
  DFF \sreg_reg[1426]  ( .D(swire[403]), .CLK(clk), .RST(rst), .Q(sreg[1426])
         );
  DFF \sreg_reg[1427]  ( .D(swire[404]), .CLK(clk), .RST(rst), .Q(sreg[1427])
         );
  DFF \sreg_reg[1428]  ( .D(swire[405]), .CLK(clk), .RST(rst), .Q(sreg[1428])
         );
  DFF \sreg_reg[1429]  ( .D(swire[406]), .CLK(clk), .RST(rst), .Q(sreg[1429])
         );
  DFF \sreg_reg[1430]  ( .D(swire[407]), .CLK(clk), .RST(rst), .Q(sreg[1430])
         );
  DFF \sreg_reg[1431]  ( .D(swire[408]), .CLK(clk), .RST(rst), .Q(sreg[1431])
         );
  DFF \sreg_reg[1432]  ( .D(swire[409]), .CLK(clk), .RST(rst), .Q(sreg[1432])
         );
  DFF \sreg_reg[1433]  ( .D(swire[410]), .CLK(clk), .RST(rst), .Q(sreg[1433])
         );
  DFF \sreg_reg[1434]  ( .D(swire[411]), .CLK(clk), .RST(rst), .Q(sreg[1434])
         );
  DFF \sreg_reg[1435]  ( .D(swire[412]), .CLK(clk), .RST(rst), .Q(sreg[1435])
         );
  DFF \sreg_reg[1436]  ( .D(swire[413]), .CLK(clk), .RST(rst), .Q(sreg[1436])
         );
  DFF \sreg_reg[1437]  ( .D(swire[414]), .CLK(clk), .RST(rst), .Q(sreg[1437])
         );
  DFF \sreg_reg[1438]  ( .D(swire[415]), .CLK(clk), .RST(rst), .Q(sreg[1438])
         );
  DFF \sreg_reg[1439]  ( .D(swire[416]), .CLK(clk), .RST(rst), .Q(sreg[1439])
         );
  DFF \sreg_reg[1440]  ( .D(swire[417]), .CLK(clk), .RST(rst), .Q(sreg[1440])
         );
  DFF \sreg_reg[1441]  ( .D(swire[418]), .CLK(clk), .RST(rst), .Q(sreg[1441])
         );
  DFF \sreg_reg[1442]  ( .D(swire[419]), .CLK(clk), .RST(rst), .Q(sreg[1442])
         );
  DFF \sreg_reg[1443]  ( .D(swire[420]), .CLK(clk), .RST(rst), .Q(sreg[1443])
         );
  DFF \sreg_reg[1444]  ( .D(swire[421]), .CLK(clk), .RST(rst), .Q(sreg[1444])
         );
  DFF \sreg_reg[1445]  ( .D(swire[422]), .CLK(clk), .RST(rst), .Q(sreg[1445])
         );
  DFF \sreg_reg[1446]  ( .D(swire[423]), .CLK(clk), .RST(rst), .Q(sreg[1446])
         );
  DFF \sreg_reg[1447]  ( .D(swire[424]), .CLK(clk), .RST(rst), .Q(sreg[1447])
         );
  DFF \sreg_reg[1448]  ( .D(swire[425]), .CLK(clk), .RST(rst), .Q(sreg[1448])
         );
  DFF \sreg_reg[1449]  ( .D(swire[426]), .CLK(clk), .RST(rst), .Q(sreg[1449])
         );
  DFF \sreg_reg[1450]  ( .D(swire[427]), .CLK(clk), .RST(rst), .Q(sreg[1450])
         );
  DFF \sreg_reg[1451]  ( .D(swire[428]), .CLK(clk), .RST(rst), .Q(sreg[1451])
         );
  DFF \sreg_reg[1452]  ( .D(swire[429]), .CLK(clk), .RST(rst), .Q(sreg[1452])
         );
  DFF \sreg_reg[1453]  ( .D(swire[430]), .CLK(clk), .RST(rst), .Q(sreg[1453])
         );
  DFF \sreg_reg[1454]  ( .D(swire[431]), .CLK(clk), .RST(rst), .Q(sreg[1454])
         );
  DFF \sreg_reg[1455]  ( .D(swire[432]), .CLK(clk), .RST(rst), .Q(sreg[1455])
         );
  DFF \sreg_reg[1456]  ( .D(swire[433]), .CLK(clk), .RST(rst), .Q(sreg[1456])
         );
  DFF \sreg_reg[1457]  ( .D(swire[434]), .CLK(clk), .RST(rst), .Q(sreg[1457])
         );
  DFF \sreg_reg[1458]  ( .D(swire[435]), .CLK(clk), .RST(rst), .Q(sreg[1458])
         );
  DFF \sreg_reg[1459]  ( .D(swire[436]), .CLK(clk), .RST(rst), .Q(sreg[1459])
         );
  DFF \sreg_reg[1460]  ( .D(swire[437]), .CLK(clk), .RST(rst), .Q(sreg[1460])
         );
  DFF \sreg_reg[1461]  ( .D(swire[438]), .CLK(clk), .RST(rst), .Q(sreg[1461])
         );
  DFF \sreg_reg[1462]  ( .D(swire[439]), .CLK(clk), .RST(rst), .Q(sreg[1462])
         );
  DFF \sreg_reg[1463]  ( .D(swire[440]), .CLK(clk), .RST(rst), .Q(sreg[1463])
         );
  DFF \sreg_reg[1464]  ( .D(swire[441]), .CLK(clk), .RST(rst), .Q(sreg[1464])
         );
  DFF \sreg_reg[1465]  ( .D(swire[442]), .CLK(clk), .RST(rst), .Q(sreg[1465])
         );
  DFF \sreg_reg[1466]  ( .D(swire[443]), .CLK(clk), .RST(rst), .Q(sreg[1466])
         );
  DFF \sreg_reg[1467]  ( .D(swire[444]), .CLK(clk), .RST(rst), .Q(sreg[1467])
         );
  DFF \sreg_reg[1468]  ( .D(swire[445]), .CLK(clk), .RST(rst), .Q(sreg[1468])
         );
  DFF \sreg_reg[1469]  ( .D(swire[446]), .CLK(clk), .RST(rst), .Q(sreg[1469])
         );
  DFF \sreg_reg[1470]  ( .D(swire[447]), .CLK(clk), .RST(rst), .Q(sreg[1470])
         );
  DFF \sreg_reg[1471]  ( .D(swire[448]), .CLK(clk), .RST(rst), .Q(sreg[1471])
         );
  DFF \sreg_reg[1472]  ( .D(swire[449]), .CLK(clk), .RST(rst), .Q(sreg[1472])
         );
  DFF \sreg_reg[1473]  ( .D(swire[450]), .CLK(clk), .RST(rst), .Q(sreg[1473])
         );
  DFF \sreg_reg[1474]  ( .D(swire[451]), .CLK(clk), .RST(rst), .Q(sreg[1474])
         );
  DFF \sreg_reg[1475]  ( .D(swire[452]), .CLK(clk), .RST(rst), .Q(sreg[1475])
         );
  DFF \sreg_reg[1476]  ( .D(swire[453]), .CLK(clk), .RST(rst), .Q(sreg[1476])
         );
  DFF \sreg_reg[1477]  ( .D(swire[454]), .CLK(clk), .RST(rst), .Q(sreg[1477])
         );
  DFF \sreg_reg[1478]  ( .D(swire[455]), .CLK(clk), .RST(rst), .Q(sreg[1478])
         );
  DFF \sreg_reg[1479]  ( .D(swire[456]), .CLK(clk), .RST(rst), .Q(sreg[1479])
         );
  DFF \sreg_reg[1480]  ( .D(swire[457]), .CLK(clk), .RST(rst), .Q(sreg[1480])
         );
  DFF \sreg_reg[1481]  ( .D(swire[458]), .CLK(clk), .RST(rst), .Q(sreg[1481])
         );
  DFF \sreg_reg[1482]  ( .D(swire[459]), .CLK(clk), .RST(rst), .Q(sreg[1482])
         );
  DFF \sreg_reg[1483]  ( .D(swire[460]), .CLK(clk), .RST(rst), .Q(sreg[1483])
         );
  DFF \sreg_reg[1484]  ( .D(swire[461]), .CLK(clk), .RST(rst), .Q(sreg[1484])
         );
  DFF \sreg_reg[1485]  ( .D(swire[462]), .CLK(clk), .RST(rst), .Q(sreg[1485])
         );
  DFF \sreg_reg[1486]  ( .D(swire[463]), .CLK(clk), .RST(rst), .Q(sreg[1486])
         );
  DFF \sreg_reg[1487]  ( .D(swire[464]), .CLK(clk), .RST(rst), .Q(sreg[1487])
         );
  DFF \sreg_reg[1488]  ( .D(swire[465]), .CLK(clk), .RST(rst), .Q(sreg[1488])
         );
  DFF \sreg_reg[1489]  ( .D(swire[466]), .CLK(clk), .RST(rst), .Q(sreg[1489])
         );
  DFF \sreg_reg[1490]  ( .D(swire[467]), .CLK(clk), .RST(rst), .Q(sreg[1490])
         );
  DFF \sreg_reg[1491]  ( .D(swire[468]), .CLK(clk), .RST(rst), .Q(sreg[1491])
         );
  DFF \sreg_reg[1492]  ( .D(swire[469]), .CLK(clk), .RST(rst), .Q(sreg[1492])
         );
  DFF \sreg_reg[1493]  ( .D(swire[470]), .CLK(clk), .RST(rst), .Q(sreg[1493])
         );
  DFF \sreg_reg[1494]  ( .D(swire[471]), .CLK(clk), .RST(rst), .Q(sreg[1494])
         );
  DFF \sreg_reg[1495]  ( .D(swire[472]), .CLK(clk), .RST(rst), .Q(sreg[1495])
         );
  DFF \sreg_reg[1496]  ( .D(swire[473]), .CLK(clk), .RST(rst), .Q(sreg[1496])
         );
  DFF \sreg_reg[1497]  ( .D(swire[474]), .CLK(clk), .RST(rst), .Q(sreg[1497])
         );
  DFF \sreg_reg[1498]  ( .D(swire[475]), .CLK(clk), .RST(rst), .Q(sreg[1498])
         );
  DFF \sreg_reg[1499]  ( .D(swire[476]), .CLK(clk), .RST(rst), .Q(sreg[1499])
         );
  DFF \sreg_reg[1500]  ( .D(swire[477]), .CLK(clk), .RST(rst), .Q(sreg[1500])
         );
  DFF \sreg_reg[1501]  ( .D(swire[478]), .CLK(clk), .RST(rst), .Q(sreg[1501])
         );
  DFF \sreg_reg[1502]  ( .D(swire[479]), .CLK(clk), .RST(rst), .Q(sreg[1502])
         );
  DFF \sreg_reg[1503]  ( .D(swire[480]), .CLK(clk), .RST(rst), .Q(sreg[1503])
         );
  DFF \sreg_reg[1504]  ( .D(swire[481]), .CLK(clk), .RST(rst), .Q(sreg[1504])
         );
  DFF \sreg_reg[1505]  ( .D(swire[482]), .CLK(clk), .RST(rst), .Q(sreg[1505])
         );
  DFF \sreg_reg[1506]  ( .D(swire[483]), .CLK(clk), .RST(rst), .Q(sreg[1506])
         );
  DFF \sreg_reg[1507]  ( .D(swire[484]), .CLK(clk), .RST(rst), .Q(sreg[1507])
         );
  DFF \sreg_reg[1508]  ( .D(swire[485]), .CLK(clk), .RST(rst), .Q(sreg[1508])
         );
  DFF \sreg_reg[1509]  ( .D(swire[486]), .CLK(clk), .RST(rst), .Q(sreg[1509])
         );
  DFF \sreg_reg[1510]  ( .D(swire[487]), .CLK(clk), .RST(rst), .Q(sreg[1510])
         );
  DFF \sreg_reg[1511]  ( .D(swire[488]), .CLK(clk), .RST(rst), .Q(sreg[1511])
         );
  DFF \sreg_reg[1512]  ( .D(swire[489]), .CLK(clk), .RST(rst), .Q(sreg[1512])
         );
  DFF \sreg_reg[1513]  ( .D(swire[490]), .CLK(clk), .RST(rst), .Q(sreg[1513])
         );
  DFF \sreg_reg[1514]  ( .D(swire[491]), .CLK(clk), .RST(rst), .Q(sreg[1514])
         );
  DFF \sreg_reg[1515]  ( .D(swire[492]), .CLK(clk), .RST(rst), .Q(sreg[1515])
         );
  DFF \sreg_reg[1516]  ( .D(swire[493]), .CLK(clk), .RST(rst), .Q(sreg[1516])
         );
  DFF \sreg_reg[1517]  ( .D(swire[494]), .CLK(clk), .RST(rst), .Q(sreg[1517])
         );
  DFF \sreg_reg[1518]  ( .D(swire[495]), .CLK(clk), .RST(rst), .Q(sreg[1518])
         );
  DFF \sreg_reg[1519]  ( .D(swire[496]), .CLK(clk), .RST(rst), .Q(sreg[1519])
         );
  DFF \sreg_reg[1520]  ( .D(swire[497]), .CLK(clk), .RST(rst), .Q(sreg[1520])
         );
  DFF \sreg_reg[1521]  ( .D(swire[498]), .CLK(clk), .RST(rst), .Q(sreg[1521])
         );
  DFF \sreg_reg[1522]  ( .D(swire[499]), .CLK(clk), .RST(rst), .Q(sreg[1522])
         );
  DFF \sreg_reg[1523]  ( .D(swire[500]), .CLK(clk), .RST(rst), .Q(sreg[1523])
         );
  DFF \sreg_reg[1524]  ( .D(swire[501]), .CLK(clk), .RST(rst), .Q(sreg[1524])
         );
  DFF \sreg_reg[1525]  ( .D(swire[502]), .CLK(clk), .RST(rst), .Q(sreg[1525])
         );
  DFF \sreg_reg[1526]  ( .D(swire[503]), .CLK(clk), .RST(rst), .Q(sreg[1526])
         );
  DFF \sreg_reg[1527]  ( .D(swire[504]), .CLK(clk), .RST(rst), .Q(sreg[1527])
         );
  DFF \sreg_reg[1528]  ( .D(swire[505]), .CLK(clk), .RST(rst), .Q(sreg[1528])
         );
  DFF \sreg_reg[1529]  ( .D(swire[506]), .CLK(clk), .RST(rst), .Q(sreg[1529])
         );
  DFF \sreg_reg[1530]  ( .D(swire[507]), .CLK(clk), .RST(rst), .Q(sreg[1530])
         );
  DFF \sreg_reg[1531]  ( .D(swire[508]), .CLK(clk), .RST(rst), .Q(sreg[1531])
         );
  DFF \sreg_reg[1532]  ( .D(swire[509]), .CLK(clk), .RST(rst), .Q(sreg[1532])
         );
  DFF \sreg_reg[1533]  ( .D(swire[510]), .CLK(clk), .RST(rst), .Q(sreg[1533])
         );
  DFF \sreg_reg[1534]  ( .D(swire[511]), .CLK(clk), .RST(rst), .Q(sreg[1534])
         );
  DFF \sreg_reg[1535]  ( .D(swire[512]), .CLK(clk), .RST(rst), .Q(sreg[1535])
         );
  DFF \sreg_reg[1536]  ( .D(swire[513]), .CLK(clk), .RST(rst), .Q(sreg[1536])
         );
  DFF \sreg_reg[1537]  ( .D(swire[514]), .CLK(clk), .RST(rst), .Q(sreg[1537])
         );
  DFF \sreg_reg[1538]  ( .D(swire[515]), .CLK(clk), .RST(rst), .Q(sreg[1538])
         );
  DFF \sreg_reg[1539]  ( .D(swire[516]), .CLK(clk), .RST(rst), .Q(sreg[1539])
         );
  DFF \sreg_reg[1540]  ( .D(swire[517]), .CLK(clk), .RST(rst), .Q(sreg[1540])
         );
  DFF \sreg_reg[1541]  ( .D(swire[518]), .CLK(clk), .RST(rst), .Q(sreg[1541])
         );
  DFF \sreg_reg[1542]  ( .D(swire[519]), .CLK(clk), .RST(rst), .Q(sreg[1542])
         );
  DFF \sreg_reg[1543]  ( .D(swire[520]), .CLK(clk), .RST(rst), .Q(sreg[1543])
         );
  DFF \sreg_reg[1544]  ( .D(swire[521]), .CLK(clk), .RST(rst), .Q(sreg[1544])
         );
  DFF \sreg_reg[1545]  ( .D(swire[522]), .CLK(clk), .RST(rst), .Q(sreg[1545])
         );
  DFF \sreg_reg[1546]  ( .D(swire[523]), .CLK(clk), .RST(rst), .Q(sreg[1546])
         );
  DFF \sreg_reg[1547]  ( .D(swire[524]), .CLK(clk), .RST(rst), .Q(sreg[1547])
         );
  DFF \sreg_reg[1548]  ( .D(swire[525]), .CLK(clk), .RST(rst), .Q(sreg[1548])
         );
  DFF \sreg_reg[1549]  ( .D(swire[526]), .CLK(clk), .RST(rst), .Q(sreg[1549])
         );
  DFF \sreg_reg[1550]  ( .D(swire[527]), .CLK(clk), .RST(rst), .Q(sreg[1550])
         );
  DFF \sreg_reg[1551]  ( .D(swire[528]), .CLK(clk), .RST(rst), .Q(sreg[1551])
         );
  DFF \sreg_reg[1552]  ( .D(swire[529]), .CLK(clk), .RST(rst), .Q(sreg[1552])
         );
  DFF \sreg_reg[1553]  ( .D(swire[530]), .CLK(clk), .RST(rst), .Q(sreg[1553])
         );
  DFF \sreg_reg[1554]  ( .D(swire[531]), .CLK(clk), .RST(rst), .Q(sreg[1554])
         );
  DFF \sreg_reg[1555]  ( .D(swire[532]), .CLK(clk), .RST(rst), .Q(sreg[1555])
         );
  DFF \sreg_reg[1556]  ( .D(swire[533]), .CLK(clk), .RST(rst), .Q(sreg[1556])
         );
  DFF \sreg_reg[1557]  ( .D(swire[534]), .CLK(clk), .RST(rst), .Q(sreg[1557])
         );
  DFF \sreg_reg[1558]  ( .D(swire[535]), .CLK(clk), .RST(rst), .Q(sreg[1558])
         );
  DFF \sreg_reg[1559]  ( .D(swire[536]), .CLK(clk), .RST(rst), .Q(sreg[1559])
         );
  DFF \sreg_reg[1560]  ( .D(swire[537]), .CLK(clk), .RST(rst), .Q(sreg[1560])
         );
  DFF \sreg_reg[1561]  ( .D(swire[538]), .CLK(clk), .RST(rst), .Q(sreg[1561])
         );
  DFF \sreg_reg[1562]  ( .D(swire[539]), .CLK(clk), .RST(rst), .Q(sreg[1562])
         );
  DFF \sreg_reg[1563]  ( .D(swire[540]), .CLK(clk), .RST(rst), .Q(sreg[1563])
         );
  DFF \sreg_reg[1564]  ( .D(swire[541]), .CLK(clk), .RST(rst), .Q(sreg[1564])
         );
  DFF \sreg_reg[1565]  ( .D(swire[542]), .CLK(clk), .RST(rst), .Q(sreg[1565])
         );
  DFF \sreg_reg[1566]  ( .D(swire[543]), .CLK(clk), .RST(rst), .Q(sreg[1566])
         );
  DFF \sreg_reg[1567]  ( .D(swire[544]), .CLK(clk), .RST(rst), .Q(sreg[1567])
         );
  DFF \sreg_reg[1568]  ( .D(swire[545]), .CLK(clk), .RST(rst), .Q(sreg[1568])
         );
  DFF \sreg_reg[1569]  ( .D(swire[546]), .CLK(clk), .RST(rst), .Q(sreg[1569])
         );
  DFF \sreg_reg[1570]  ( .D(swire[547]), .CLK(clk), .RST(rst), .Q(sreg[1570])
         );
  DFF \sreg_reg[1571]  ( .D(swire[548]), .CLK(clk), .RST(rst), .Q(sreg[1571])
         );
  DFF \sreg_reg[1572]  ( .D(swire[549]), .CLK(clk), .RST(rst), .Q(sreg[1572])
         );
  DFF \sreg_reg[1573]  ( .D(swire[550]), .CLK(clk), .RST(rst), .Q(sreg[1573])
         );
  DFF \sreg_reg[1574]  ( .D(swire[551]), .CLK(clk), .RST(rst), .Q(sreg[1574])
         );
  DFF \sreg_reg[1575]  ( .D(swire[552]), .CLK(clk), .RST(rst), .Q(sreg[1575])
         );
  DFF \sreg_reg[1576]  ( .D(swire[553]), .CLK(clk), .RST(rst), .Q(sreg[1576])
         );
  DFF \sreg_reg[1577]  ( .D(swire[554]), .CLK(clk), .RST(rst), .Q(sreg[1577])
         );
  DFF \sreg_reg[1578]  ( .D(swire[555]), .CLK(clk), .RST(rst), .Q(sreg[1578])
         );
  DFF \sreg_reg[1579]  ( .D(swire[556]), .CLK(clk), .RST(rst), .Q(sreg[1579])
         );
  DFF \sreg_reg[1580]  ( .D(swire[557]), .CLK(clk), .RST(rst), .Q(sreg[1580])
         );
  DFF \sreg_reg[1581]  ( .D(swire[558]), .CLK(clk), .RST(rst), .Q(sreg[1581])
         );
  DFF \sreg_reg[1582]  ( .D(swire[559]), .CLK(clk), .RST(rst), .Q(sreg[1582])
         );
  DFF \sreg_reg[1583]  ( .D(swire[560]), .CLK(clk), .RST(rst), .Q(sreg[1583])
         );
  DFF \sreg_reg[1584]  ( .D(swire[561]), .CLK(clk), .RST(rst), .Q(sreg[1584])
         );
  DFF \sreg_reg[1585]  ( .D(swire[562]), .CLK(clk), .RST(rst), .Q(sreg[1585])
         );
  DFF \sreg_reg[1586]  ( .D(swire[563]), .CLK(clk), .RST(rst), .Q(sreg[1586])
         );
  DFF \sreg_reg[1587]  ( .D(swire[564]), .CLK(clk), .RST(rst), .Q(sreg[1587])
         );
  DFF \sreg_reg[1588]  ( .D(swire[565]), .CLK(clk), .RST(rst), .Q(sreg[1588])
         );
  DFF \sreg_reg[1589]  ( .D(swire[566]), .CLK(clk), .RST(rst), .Q(sreg[1589])
         );
  DFF \sreg_reg[1590]  ( .D(swire[567]), .CLK(clk), .RST(rst), .Q(sreg[1590])
         );
  DFF \sreg_reg[1591]  ( .D(swire[568]), .CLK(clk), .RST(rst), .Q(sreg[1591])
         );
  DFF \sreg_reg[1592]  ( .D(swire[569]), .CLK(clk), .RST(rst), .Q(sreg[1592])
         );
  DFF \sreg_reg[1593]  ( .D(swire[570]), .CLK(clk), .RST(rst), .Q(sreg[1593])
         );
  DFF \sreg_reg[1594]  ( .D(swire[571]), .CLK(clk), .RST(rst), .Q(sreg[1594])
         );
  DFF \sreg_reg[1595]  ( .D(swire[572]), .CLK(clk), .RST(rst), .Q(sreg[1595])
         );
  DFF \sreg_reg[1596]  ( .D(swire[573]), .CLK(clk), .RST(rst), .Q(sreg[1596])
         );
  DFF \sreg_reg[1597]  ( .D(swire[574]), .CLK(clk), .RST(rst), .Q(sreg[1597])
         );
  DFF \sreg_reg[1598]  ( .D(swire[575]), .CLK(clk), .RST(rst), .Q(sreg[1598])
         );
  DFF \sreg_reg[1599]  ( .D(swire[576]), .CLK(clk), .RST(rst), .Q(sreg[1599])
         );
  DFF \sreg_reg[1600]  ( .D(swire[577]), .CLK(clk), .RST(rst), .Q(sreg[1600])
         );
  DFF \sreg_reg[1601]  ( .D(swire[578]), .CLK(clk), .RST(rst), .Q(sreg[1601])
         );
  DFF \sreg_reg[1602]  ( .D(swire[579]), .CLK(clk), .RST(rst), .Q(sreg[1602])
         );
  DFF \sreg_reg[1603]  ( .D(swire[580]), .CLK(clk), .RST(rst), .Q(sreg[1603])
         );
  DFF \sreg_reg[1604]  ( .D(swire[581]), .CLK(clk), .RST(rst), .Q(sreg[1604])
         );
  DFF \sreg_reg[1605]  ( .D(swire[582]), .CLK(clk), .RST(rst), .Q(sreg[1605])
         );
  DFF \sreg_reg[1606]  ( .D(swire[583]), .CLK(clk), .RST(rst), .Q(sreg[1606])
         );
  DFF \sreg_reg[1607]  ( .D(swire[584]), .CLK(clk), .RST(rst), .Q(sreg[1607])
         );
  DFF \sreg_reg[1608]  ( .D(swire[585]), .CLK(clk), .RST(rst), .Q(sreg[1608])
         );
  DFF \sreg_reg[1609]  ( .D(swire[586]), .CLK(clk), .RST(rst), .Q(sreg[1609])
         );
  DFF \sreg_reg[1610]  ( .D(swire[587]), .CLK(clk), .RST(rst), .Q(sreg[1610])
         );
  DFF \sreg_reg[1611]  ( .D(swire[588]), .CLK(clk), .RST(rst), .Q(sreg[1611])
         );
  DFF \sreg_reg[1612]  ( .D(swire[589]), .CLK(clk), .RST(rst), .Q(sreg[1612])
         );
  DFF \sreg_reg[1613]  ( .D(swire[590]), .CLK(clk), .RST(rst), .Q(sreg[1613])
         );
  DFF \sreg_reg[1614]  ( .D(swire[591]), .CLK(clk), .RST(rst), .Q(sreg[1614])
         );
  DFF \sreg_reg[1615]  ( .D(swire[592]), .CLK(clk), .RST(rst), .Q(sreg[1615])
         );
  DFF \sreg_reg[1616]  ( .D(swire[593]), .CLK(clk), .RST(rst), .Q(sreg[1616])
         );
  DFF \sreg_reg[1617]  ( .D(swire[594]), .CLK(clk), .RST(rst), .Q(sreg[1617])
         );
  DFF \sreg_reg[1618]  ( .D(swire[595]), .CLK(clk), .RST(rst), .Q(sreg[1618])
         );
  DFF \sreg_reg[1619]  ( .D(swire[596]), .CLK(clk), .RST(rst), .Q(sreg[1619])
         );
  DFF \sreg_reg[1620]  ( .D(swire[597]), .CLK(clk), .RST(rst), .Q(sreg[1620])
         );
  DFF \sreg_reg[1621]  ( .D(swire[598]), .CLK(clk), .RST(rst), .Q(sreg[1621])
         );
  DFF \sreg_reg[1622]  ( .D(swire[599]), .CLK(clk), .RST(rst), .Q(sreg[1622])
         );
  DFF \sreg_reg[1623]  ( .D(swire[600]), .CLK(clk), .RST(rst), .Q(sreg[1623])
         );
  DFF \sreg_reg[1624]  ( .D(swire[601]), .CLK(clk), .RST(rst), .Q(sreg[1624])
         );
  DFF \sreg_reg[1625]  ( .D(swire[602]), .CLK(clk), .RST(rst), .Q(sreg[1625])
         );
  DFF \sreg_reg[1626]  ( .D(swire[603]), .CLK(clk), .RST(rst), .Q(sreg[1626])
         );
  DFF \sreg_reg[1627]  ( .D(swire[604]), .CLK(clk), .RST(rst), .Q(sreg[1627])
         );
  DFF \sreg_reg[1628]  ( .D(swire[605]), .CLK(clk), .RST(rst), .Q(sreg[1628])
         );
  DFF \sreg_reg[1629]  ( .D(swire[606]), .CLK(clk), .RST(rst), .Q(sreg[1629])
         );
  DFF \sreg_reg[1630]  ( .D(swire[607]), .CLK(clk), .RST(rst), .Q(sreg[1630])
         );
  DFF \sreg_reg[1631]  ( .D(swire[608]), .CLK(clk), .RST(rst), .Q(sreg[1631])
         );
  DFF \sreg_reg[1632]  ( .D(swire[609]), .CLK(clk), .RST(rst), .Q(sreg[1632])
         );
  DFF \sreg_reg[1633]  ( .D(swire[610]), .CLK(clk), .RST(rst), .Q(sreg[1633])
         );
  DFF \sreg_reg[1634]  ( .D(swire[611]), .CLK(clk), .RST(rst), .Q(sreg[1634])
         );
  DFF \sreg_reg[1635]  ( .D(swire[612]), .CLK(clk), .RST(rst), .Q(sreg[1635])
         );
  DFF \sreg_reg[1636]  ( .D(swire[613]), .CLK(clk), .RST(rst), .Q(sreg[1636])
         );
  DFF \sreg_reg[1637]  ( .D(swire[614]), .CLK(clk), .RST(rst), .Q(sreg[1637])
         );
  DFF \sreg_reg[1638]  ( .D(swire[615]), .CLK(clk), .RST(rst), .Q(sreg[1638])
         );
  DFF \sreg_reg[1639]  ( .D(swire[616]), .CLK(clk), .RST(rst), .Q(sreg[1639])
         );
  DFF \sreg_reg[1640]  ( .D(swire[617]), .CLK(clk), .RST(rst), .Q(sreg[1640])
         );
  DFF \sreg_reg[1641]  ( .D(swire[618]), .CLK(clk), .RST(rst), .Q(sreg[1641])
         );
  DFF \sreg_reg[1642]  ( .D(swire[619]), .CLK(clk), .RST(rst), .Q(sreg[1642])
         );
  DFF \sreg_reg[1643]  ( .D(swire[620]), .CLK(clk), .RST(rst), .Q(sreg[1643])
         );
  DFF \sreg_reg[1644]  ( .D(swire[621]), .CLK(clk), .RST(rst), .Q(sreg[1644])
         );
  DFF \sreg_reg[1645]  ( .D(swire[622]), .CLK(clk), .RST(rst), .Q(sreg[1645])
         );
  DFF \sreg_reg[1646]  ( .D(swire[623]), .CLK(clk), .RST(rst), .Q(sreg[1646])
         );
  DFF \sreg_reg[1647]  ( .D(swire[624]), .CLK(clk), .RST(rst), .Q(sreg[1647])
         );
  DFF \sreg_reg[1648]  ( .D(swire[625]), .CLK(clk), .RST(rst), .Q(sreg[1648])
         );
  DFF \sreg_reg[1649]  ( .D(swire[626]), .CLK(clk), .RST(rst), .Q(sreg[1649])
         );
  DFF \sreg_reg[1650]  ( .D(swire[627]), .CLK(clk), .RST(rst), .Q(sreg[1650])
         );
  DFF \sreg_reg[1651]  ( .D(swire[628]), .CLK(clk), .RST(rst), .Q(sreg[1651])
         );
  DFF \sreg_reg[1652]  ( .D(swire[629]), .CLK(clk), .RST(rst), .Q(sreg[1652])
         );
  DFF \sreg_reg[1653]  ( .D(swire[630]), .CLK(clk), .RST(rst), .Q(sreg[1653])
         );
  DFF \sreg_reg[1654]  ( .D(swire[631]), .CLK(clk), .RST(rst), .Q(sreg[1654])
         );
  DFF \sreg_reg[1655]  ( .D(swire[632]), .CLK(clk), .RST(rst), .Q(sreg[1655])
         );
  DFF \sreg_reg[1656]  ( .D(swire[633]), .CLK(clk), .RST(rst), .Q(sreg[1656])
         );
  DFF \sreg_reg[1657]  ( .D(swire[634]), .CLK(clk), .RST(rst), .Q(sreg[1657])
         );
  DFF \sreg_reg[1658]  ( .D(swire[635]), .CLK(clk), .RST(rst), .Q(sreg[1658])
         );
  DFF \sreg_reg[1659]  ( .D(swire[636]), .CLK(clk), .RST(rst), .Q(sreg[1659])
         );
  DFF \sreg_reg[1660]  ( .D(swire[637]), .CLK(clk), .RST(rst), .Q(sreg[1660])
         );
  DFF \sreg_reg[1661]  ( .D(swire[638]), .CLK(clk), .RST(rst), .Q(sreg[1661])
         );
  DFF \sreg_reg[1662]  ( .D(swire[639]), .CLK(clk), .RST(rst), .Q(sreg[1662])
         );
  DFF \sreg_reg[1663]  ( .D(swire[640]), .CLK(clk), .RST(rst), .Q(sreg[1663])
         );
  DFF \sreg_reg[1664]  ( .D(swire[641]), .CLK(clk), .RST(rst), .Q(sreg[1664])
         );
  DFF \sreg_reg[1665]  ( .D(swire[642]), .CLK(clk), .RST(rst), .Q(sreg[1665])
         );
  DFF \sreg_reg[1666]  ( .D(swire[643]), .CLK(clk), .RST(rst), .Q(sreg[1666])
         );
  DFF \sreg_reg[1667]  ( .D(swire[644]), .CLK(clk), .RST(rst), .Q(sreg[1667])
         );
  DFF \sreg_reg[1668]  ( .D(swire[645]), .CLK(clk), .RST(rst), .Q(sreg[1668])
         );
  DFF \sreg_reg[1669]  ( .D(swire[646]), .CLK(clk), .RST(rst), .Q(sreg[1669])
         );
  DFF \sreg_reg[1670]  ( .D(swire[647]), .CLK(clk), .RST(rst), .Q(sreg[1670])
         );
  DFF \sreg_reg[1671]  ( .D(swire[648]), .CLK(clk), .RST(rst), .Q(sreg[1671])
         );
  DFF \sreg_reg[1672]  ( .D(swire[649]), .CLK(clk), .RST(rst), .Q(sreg[1672])
         );
  DFF \sreg_reg[1673]  ( .D(swire[650]), .CLK(clk), .RST(rst), .Q(sreg[1673])
         );
  DFF \sreg_reg[1674]  ( .D(swire[651]), .CLK(clk), .RST(rst), .Q(sreg[1674])
         );
  DFF \sreg_reg[1675]  ( .D(swire[652]), .CLK(clk), .RST(rst), .Q(sreg[1675])
         );
  DFF \sreg_reg[1676]  ( .D(swire[653]), .CLK(clk), .RST(rst), .Q(sreg[1676])
         );
  DFF \sreg_reg[1677]  ( .D(swire[654]), .CLK(clk), .RST(rst), .Q(sreg[1677])
         );
  DFF \sreg_reg[1678]  ( .D(swire[655]), .CLK(clk), .RST(rst), .Q(sreg[1678])
         );
  DFF \sreg_reg[1679]  ( .D(swire[656]), .CLK(clk), .RST(rst), .Q(sreg[1679])
         );
  DFF \sreg_reg[1680]  ( .D(swire[657]), .CLK(clk), .RST(rst), .Q(sreg[1680])
         );
  DFF \sreg_reg[1681]  ( .D(swire[658]), .CLK(clk), .RST(rst), .Q(sreg[1681])
         );
  DFF \sreg_reg[1682]  ( .D(swire[659]), .CLK(clk), .RST(rst), .Q(sreg[1682])
         );
  DFF \sreg_reg[1683]  ( .D(swire[660]), .CLK(clk), .RST(rst), .Q(sreg[1683])
         );
  DFF \sreg_reg[1684]  ( .D(swire[661]), .CLK(clk), .RST(rst), .Q(sreg[1684])
         );
  DFF \sreg_reg[1685]  ( .D(swire[662]), .CLK(clk), .RST(rst), .Q(sreg[1685])
         );
  DFF \sreg_reg[1686]  ( .D(swire[663]), .CLK(clk), .RST(rst), .Q(sreg[1686])
         );
  DFF \sreg_reg[1687]  ( .D(swire[664]), .CLK(clk), .RST(rst), .Q(sreg[1687])
         );
  DFF \sreg_reg[1688]  ( .D(swire[665]), .CLK(clk), .RST(rst), .Q(sreg[1688])
         );
  DFF \sreg_reg[1689]  ( .D(swire[666]), .CLK(clk), .RST(rst), .Q(sreg[1689])
         );
  DFF \sreg_reg[1690]  ( .D(swire[667]), .CLK(clk), .RST(rst), .Q(sreg[1690])
         );
  DFF \sreg_reg[1691]  ( .D(swire[668]), .CLK(clk), .RST(rst), .Q(sreg[1691])
         );
  DFF \sreg_reg[1692]  ( .D(swire[669]), .CLK(clk), .RST(rst), .Q(sreg[1692])
         );
  DFF \sreg_reg[1693]  ( .D(swire[670]), .CLK(clk), .RST(rst), .Q(sreg[1693])
         );
  DFF \sreg_reg[1694]  ( .D(swire[671]), .CLK(clk), .RST(rst), .Q(sreg[1694])
         );
  DFF \sreg_reg[1695]  ( .D(swire[672]), .CLK(clk), .RST(rst), .Q(sreg[1695])
         );
  DFF \sreg_reg[1696]  ( .D(swire[673]), .CLK(clk), .RST(rst), .Q(sreg[1696])
         );
  DFF \sreg_reg[1697]  ( .D(swire[674]), .CLK(clk), .RST(rst), .Q(sreg[1697])
         );
  DFF \sreg_reg[1698]  ( .D(swire[675]), .CLK(clk), .RST(rst), .Q(sreg[1698])
         );
  DFF \sreg_reg[1699]  ( .D(swire[676]), .CLK(clk), .RST(rst), .Q(sreg[1699])
         );
  DFF \sreg_reg[1700]  ( .D(swire[677]), .CLK(clk), .RST(rst), .Q(sreg[1700])
         );
  DFF \sreg_reg[1701]  ( .D(swire[678]), .CLK(clk), .RST(rst), .Q(sreg[1701])
         );
  DFF \sreg_reg[1702]  ( .D(swire[679]), .CLK(clk), .RST(rst), .Q(sreg[1702])
         );
  DFF \sreg_reg[1703]  ( .D(swire[680]), .CLK(clk), .RST(rst), .Q(sreg[1703])
         );
  DFF \sreg_reg[1704]  ( .D(swire[681]), .CLK(clk), .RST(rst), .Q(sreg[1704])
         );
  DFF \sreg_reg[1705]  ( .D(swire[682]), .CLK(clk), .RST(rst), .Q(sreg[1705])
         );
  DFF \sreg_reg[1706]  ( .D(swire[683]), .CLK(clk), .RST(rst), .Q(sreg[1706])
         );
  DFF \sreg_reg[1707]  ( .D(swire[684]), .CLK(clk), .RST(rst), .Q(sreg[1707])
         );
  DFF \sreg_reg[1708]  ( .D(swire[685]), .CLK(clk), .RST(rst), .Q(sreg[1708])
         );
  DFF \sreg_reg[1709]  ( .D(swire[686]), .CLK(clk), .RST(rst), .Q(sreg[1709])
         );
  DFF \sreg_reg[1710]  ( .D(swire[687]), .CLK(clk), .RST(rst), .Q(sreg[1710])
         );
  DFF \sreg_reg[1711]  ( .D(swire[688]), .CLK(clk), .RST(rst), .Q(sreg[1711])
         );
  DFF \sreg_reg[1712]  ( .D(swire[689]), .CLK(clk), .RST(rst), .Q(sreg[1712])
         );
  DFF \sreg_reg[1713]  ( .D(swire[690]), .CLK(clk), .RST(rst), .Q(sreg[1713])
         );
  DFF \sreg_reg[1714]  ( .D(swire[691]), .CLK(clk), .RST(rst), .Q(sreg[1714])
         );
  DFF \sreg_reg[1715]  ( .D(swire[692]), .CLK(clk), .RST(rst), .Q(sreg[1715])
         );
  DFF \sreg_reg[1716]  ( .D(swire[693]), .CLK(clk), .RST(rst), .Q(sreg[1716])
         );
  DFF \sreg_reg[1717]  ( .D(swire[694]), .CLK(clk), .RST(rst), .Q(sreg[1717])
         );
  DFF \sreg_reg[1718]  ( .D(swire[695]), .CLK(clk), .RST(rst), .Q(sreg[1718])
         );
  DFF \sreg_reg[1719]  ( .D(swire[696]), .CLK(clk), .RST(rst), .Q(sreg[1719])
         );
  DFF \sreg_reg[1720]  ( .D(swire[697]), .CLK(clk), .RST(rst), .Q(sreg[1720])
         );
  DFF \sreg_reg[1721]  ( .D(swire[698]), .CLK(clk), .RST(rst), .Q(sreg[1721])
         );
  DFF \sreg_reg[1722]  ( .D(swire[699]), .CLK(clk), .RST(rst), .Q(sreg[1722])
         );
  DFF \sreg_reg[1723]  ( .D(swire[700]), .CLK(clk), .RST(rst), .Q(sreg[1723])
         );
  DFF \sreg_reg[1724]  ( .D(swire[701]), .CLK(clk), .RST(rst), .Q(sreg[1724])
         );
  DFF \sreg_reg[1725]  ( .D(swire[702]), .CLK(clk), .RST(rst), .Q(sreg[1725])
         );
  DFF \sreg_reg[1726]  ( .D(swire[703]), .CLK(clk), .RST(rst), .Q(sreg[1726])
         );
  DFF \sreg_reg[1727]  ( .D(swire[704]), .CLK(clk), .RST(rst), .Q(sreg[1727])
         );
  DFF \sreg_reg[1728]  ( .D(swire[705]), .CLK(clk), .RST(rst), .Q(sreg[1728])
         );
  DFF \sreg_reg[1729]  ( .D(swire[706]), .CLK(clk), .RST(rst), .Q(sreg[1729])
         );
  DFF \sreg_reg[1730]  ( .D(swire[707]), .CLK(clk), .RST(rst), .Q(sreg[1730])
         );
  DFF \sreg_reg[1731]  ( .D(swire[708]), .CLK(clk), .RST(rst), .Q(sreg[1731])
         );
  DFF \sreg_reg[1732]  ( .D(swire[709]), .CLK(clk), .RST(rst), .Q(sreg[1732])
         );
  DFF \sreg_reg[1733]  ( .D(swire[710]), .CLK(clk), .RST(rst), .Q(sreg[1733])
         );
  DFF \sreg_reg[1734]  ( .D(swire[711]), .CLK(clk), .RST(rst), .Q(sreg[1734])
         );
  DFF \sreg_reg[1735]  ( .D(swire[712]), .CLK(clk), .RST(rst), .Q(sreg[1735])
         );
  DFF \sreg_reg[1736]  ( .D(swire[713]), .CLK(clk), .RST(rst), .Q(sreg[1736])
         );
  DFF \sreg_reg[1737]  ( .D(swire[714]), .CLK(clk), .RST(rst), .Q(sreg[1737])
         );
  DFF \sreg_reg[1738]  ( .D(swire[715]), .CLK(clk), .RST(rst), .Q(sreg[1738])
         );
  DFF \sreg_reg[1739]  ( .D(swire[716]), .CLK(clk), .RST(rst), .Q(sreg[1739])
         );
  DFF \sreg_reg[1740]  ( .D(swire[717]), .CLK(clk), .RST(rst), .Q(sreg[1740])
         );
  DFF \sreg_reg[1741]  ( .D(swire[718]), .CLK(clk), .RST(rst), .Q(sreg[1741])
         );
  DFF \sreg_reg[1742]  ( .D(swire[719]), .CLK(clk), .RST(rst), .Q(sreg[1742])
         );
  DFF \sreg_reg[1743]  ( .D(swire[720]), .CLK(clk), .RST(rst), .Q(sreg[1743])
         );
  DFF \sreg_reg[1744]  ( .D(swire[721]), .CLK(clk), .RST(rst), .Q(sreg[1744])
         );
  DFF \sreg_reg[1745]  ( .D(swire[722]), .CLK(clk), .RST(rst), .Q(sreg[1745])
         );
  DFF \sreg_reg[1746]  ( .D(swire[723]), .CLK(clk), .RST(rst), .Q(sreg[1746])
         );
  DFF \sreg_reg[1747]  ( .D(swire[724]), .CLK(clk), .RST(rst), .Q(sreg[1747])
         );
  DFF \sreg_reg[1748]  ( .D(swire[725]), .CLK(clk), .RST(rst), .Q(sreg[1748])
         );
  DFF \sreg_reg[1749]  ( .D(swire[726]), .CLK(clk), .RST(rst), .Q(sreg[1749])
         );
  DFF \sreg_reg[1750]  ( .D(swire[727]), .CLK(clk), .RST(rst), .Q(sreg[1750])
         );
  DFF \sreg_reg[1751]  ( .D(swire[728]), .CLK(clk), .RST(rst), .Q(sreg[1751])
         );
  DFF \sreg_reg[1752]  ( .D(swire[729]), .CLK(clk), .RST(rst), .Q(sreg[1752])
         );
  DFF \sreg_reg[1753]  ( .D(swire[730]), .CLK(clk), .RST(rst), .Q(sreg[1753])
         );
  DFF \sreg_reg[1754]  ( .D(swire[731]), .CLK(clk), .RST(rst), .Q(sreg[1754])
         );
  DFF \sreg_reg[1755]  ( .D(swire[732]), .CLK(clk), .RST(rst), .Q(sreg[1755])
         );
  DFF \sreg_reg[1756]  ( .D(swire[733]), .CLK(clk), .RST(rst), .Q(sreg[1756])
         );
  DFF \sreg_reg[1757]  ( .D(swire[734]), .CLK(clk), .RST(rst), .Q(sreg[1757])
         );
  DFF \sreg_reg[1758]  ( .D(swire[735]), .CLK(clk), .RST(rst), .Q(sreg[1758])
         );
  DFF \sreg_reg[1759]  ( .D(swire[736]), .CLK(clk), .RST(rst), .Q(sreg[1759])
         );
  DFF \sreg_reg[1760]  ( .D(swire[737]), .CLK(clk), .RST(rst), .Q(sreg[1760])
         );
  DFF \sreg_reg[1761]  ( .D(swire[738]), .CLK(clk), .RST(rst), .Q(sreg[1761])
         );
  DFF \sreg_reg[1762]  ( .D(swire[739]), .CLK(clk), .RST(rst), .Q(sreg[1762])
         );
  DFF \sreg_reg[1763]  ( .D(swire[740]), .CLK(clk), .RST(rst), .Q(sreg[1763])
         );
  DFF \sreg_reg[1764]  ( .D(swire[741]), .CLK(clk), .RST(rst), .Q(sreg[1764])
         );
  DFF \sreg_reg[1765]  ( .D(swire[742]), .CLK(clk), .RST(rst), .Q(sreg[1765])
         );
  DFF \sreg_reg[1766]  ( .D(swire[743]), .CLK(clk), .RST(rst), .Q(sreg[1766])
         );
  DFF \sreg_reg[1767]  ( .D(swire[744]), .CLK(clk), .RST(rst), .Q(sreg[1767])
         );
  DFF \sreg_reg[1768]  ( .D(swire[745]), .CLK(clk), .RST(rst), .Q(sreg[1768])
         );
  DFF \sreg_reg[1769]  ( .D(swire[746]), .CLK(clk), .RST(rst), .Q(sreg[1769])
         );
  DFF \sreg_reg[1770]  ( .D(swire[747]), .CLK(clk), .RST(rst), .Q(sreg[1770])
         );
  DFF \sreg_reg[1771]  ( .D(swire[748]), .CLK(clk), .RST(rst), .Q(sreg[1771])
         );
  DFF \sreg_reg[1772]  ( .D(swire[749]), .CLK(clk), .RST(rst), .Q(sreg[1772])
         );
  DFF \sreg_reg[1773]  ( .D(swire[750]), .CLK(clk), .RST(rst), .Q(sreg[1773])
         );
  DFF \sreg_reg[1774]  ( .D(swire[751]), .CLK(clk), .RST(rst), .Q(sreg[1774])
         );
  DFF \sreg_reg[1775]  ( .D(swire[752]), .CLK(clk), .RST(rst), .Q(sreg[1775])
         );
  DFF \sreg_reg[1776]  ( .D(swire[753]), .CLK(clk), .RST(rst), .Q(sreg[1776])
         );
  DFF \sreg_reg[1777]  ( .D(swire[754]), .CLK(clk), .RST(rst), .Q(sreg[1777])
         );
  DFF \sreg_reg[1778]  ( .D(swire[755]), .CLK(clk), .RST(rst), .Q(sreg[1778])
         );
  DFF \sreg_reg[1779]  ( .D(swire[756]), .CLK(clk), .RST(rst), .Q(sreg[1779])
         );
  DFF \sreg_reg[1780]  ( .D(swire[757]), .CLK(clk), .RST(rst), .Q(sreg[1780])
         );
  DFF \sreg_reg[1781]  ( .D(swire[758]), .CLK(clk), .RST(rst), .Q(sreg[1781])
         );
  DFF \sreg_reg[1782]  ( .D(swire[759]), .CLK(clk), .RST(rst), .Q(sreg[1782])
         );
  DFF \sreg_reg[1783]  ( .D(swire[760]), .CLK(clk), .RST(rst), .Q(sreg[1783])
         );
  DFF \sreg_reg[1784]  ( .D(swire[761]), .CLK(clk), .RST(rst), .Q(sreg[1784])
         );
  DFF \sreg_reg[1785]  ( .D(swire[762]), .CLK(clk), .RST(rst), .Q(sreg[1785])
         );
  DFF \sreg_reg[1786]  ( .D(swire[763]), .CLK(clk), .RST(rst), .Q(sreg[1786])
         );
  DFF \sreg_reg[1787]  ( .D(swire[764]), .CLK(clk), .RST(rst), .Q(sreg[1787])
         );
  DFF \sreg_reg[1788]  ( .D(swire[765]), .CLK(clk), .RST(rst), .Q(sreg[1788])
         );
  DFF \sreg_reg[1789]  ( .D(swire[766]), .CLK(clk), .RST(rst), .Q(sreg[1789])
         );
  DFF \sreg_reg[1790]  ( .D(swire[767]), .CLK(clk), .RST(rst), .Q(sreg[1790])
         );
  DFF \sreg_reg[1791]  ( .D(swire[768]), .CLK(clk), .RST(rst), .Q(sreg[1791])
         );
  DFF \sreg_reg[1792]  ( .D(swire[769]), .CLK(clk), .RST(rst), .Q(sreg[1792])
         );
  DFF \sreg_reg[1793]  ( .D(swire[770]), .CLK(clk), .RST(rst), .Q(sreg[1793])
         );
  DFF \sreg_reg[1794]  ( .D(swire[771]), .CLK(clk), .RST(rst), .Q(sreg[1794])
         );
  DFF \sreg_reg[1795]  ( .D(swire[772]), .CLK(clk), .RST(rst), .Q(sreg[1795])
         );
  DFF \sreg_reg[1796]  ( .D(swire[773]), .CLK(clk), .RST(rst), .Q(sreg[1796])
         );
  DFF \sreg_reg[1797]  ( .D(swire[774]), .CLK(clk), .RST(rst), .Q(sreg[1797])
         );
  DFF \sreg_reg[1798]  ( .D(swire[775]), .CLK(clk), .RST(rst), .Q(sreg[1798])
         );
  DFF \sreg_reg[1799]  ( .D(swire[776]), .CLK(clk), .RST(rst), .Q(sreg[1799])
         );
  DFF \sreg_reg[1800]  ( .D(swire[777]), .CLK(clk), .RST(rst), .Q(sreg[1800])
         );
  DFF \sreg_reg[1801]  ( .D(swire[778]), .CLK(clk), .RST(rst), .Q(sreg[1801])
         );
  DFF \sreg_reg[1802]  ( .D(swire[779]), .CLK(clk), .RST(rst), .Q(sreg[1802])
         );
  DFF \sreg_reg[1803]  ( .D(swire[780]), .CLK(clk), .RST(rst), .Q(sreg[1803])
         );
  DFF \sreg_reg[1804]  ( .D(swire[781]), .CLK(clk), .RST(rst), .Q(sreg[1804])
         );
  DFF \sreg_reg[1805]  ( .D(swire[782]), .CLK(clk), .RST(rst), .Q(sreg[1805])
         );
  DFF \sreg_reg[1806]  ( .D(swire[783]), .CLK(clk), .RST(rst), .Q(sreg[1806])
         );
  DFF \sreg_reg[1807]  ( .D(swire[784]), .CLK(clk), .RST(rst), .Q(sreg[1807])
         );
  DFF \sreg_reg[1808]  ( .D(swire[785]), .CLK(clk), .RST(rst), .Q(sreg[1808])
         );
  DFF \sreg_reg[1809]  ( .D(swire[786]), .CLK(clk), .RST(rst), .Q(sreg[1809])
         );
  DFF \sreg_reg[1810]  ( .D(swire[787]), .CLK(clk), .RST(rst), .Q(sreg[1810])
         );
  DFF \sreg_reg[1811]  ( .D(swire[788]), .CLK(clk), .RST(rst), .Q(sreg[1811])
         );
  DFF \sreg_reg[1812]  ( .D(swire[789]), .CLK(clk), .RST(rst), .Q(sreg[1812])
         );
  DFF \sreg_reg[1813]  ( .D(swire[790]), .CLK(clk), .RST(rst), .Q(sreg[1813])
         );
  DFF \sreg_reg[1814]  ( .D(swire[791]), .CLK(clk), .RST(rst), .Q(sreg[1814])
         );
  DFF \sreg_reg[1815]  ( .D(swire[792]), .CLK(clk), .RST(rst), .Q(sreg[1815])
         );
  DFF \sreg_reg[1816]  ( .D(swire[793]), .CLK(clk), .RST(rst), .Q(sreg[1816])
         );
  DFF \sreg_reg[1817]  ( .D(swire[794]), .CLK(clk), .RST(rst), .Q(sreg[1817])
         );
  DFF \sreg_reg[1818]  ( .D(swire[795]), .CLK(clk), .RST(rst), .Q(sreg[1818])
         );
  DFF \sreg_reg[1819]  ( .D(swire[796]), .CLK(clk), .RST(rst), .Q(sreg[1819])
         );
  DFF \sreg_reg[1820]  ( .D(swire[797]), .CLK(clk), .RST(rst), .Q(sreg[1820])
         );
  DFF \sreg_reg[1821]  ( .D(swire[798]), .CLK(clk), .RST(rst), .Q(sreg[1821])
         );
  DFF \sreg_reg[1822]  ( .D(swire[799]), .CLK(clk), .RST(rst), .Q(sreg[1822])
         );
  DFF \sreg_reg[1823]  ( .D(swire[800]), .CLK(clk), .RST(rst), .Q(sreg[1823])
         );
  DFF \sreg_reg[1824]  ( .D(swire[801]), .CLK(clk), .RST(rst), .Q(sreg[1824])
         );
  DFF \sreg_reg[1825]  ( .D(swire[802]), .CLK(clk), .RST(rst), .Q(sreg[1825])
         );
  DFF \sreg_reg[1826]  ( .D(swire[803]), .CLK(clk), .RST(rst), .Q(sreg[1826])
         );
  DFF \sreg_reg[1827]  ( .D(swire[804]), .CLK(clk), .RST(rst), .Q(sreg[1827])
         );
  DFF \sreg_reg[1828]  ( .D(swire[805]), .CLK(clk), .RST(rst), .Q(sreg[1828])
         );
  DFF \sreg_reg[1829]  ( .D(swire[806]), .CLK(clk), .RST(rst), .Q(sreg[1829])
         );
  DFF \sreg_reg[1830]  ( .D(swire[807]), .CLK(clk), .RST(rst), .Q(sreg[1830])
         );
  DFF \sreg_reg[1831]  ( .D(swire[808]), .CLK(clk), .RST(rst), .Q(sreg[1831])
         );
  DFF \sreg_reg[1832]  ( .D(swire[809]), .CLK(clk), .RST(rst), .Q(sreg[1832])
         );
  DFF \sreg_reg[1833]  ( .D(swire[810]), .CLK(clk), .RST(rst), .Q(sreg[1833])
         );
  DFF \sreg_reg[1834]  ( .D(swire[811]), .CLK(clk), .RST(rst), .Q(sreg[1834])
         );
  DFF \sreg_reg[1835]  ( .D(swire[812]), .CLK(clk), .RST(rst), .Q(sreg[1835])
         );
  DFF \sreg_reg[1836]  ( .D(swire[813]), .CLK(clk), .RST(rst), .Q(sreg[1836])
         );
  DFF \sreg_reg[1837]  ( .D(swire[814]), .CLK(clk), .RST(rst), .Q(sreg[1837])
         );
  DFF \sreg_reg[1838]  ( .D(swire[815]), .CLK(clk), .RST(rst), .Q(sreg[1838])
         );
  DFF \sreg_reg[1839]  ( .D(swire[816]), .CLK(clk), .RST(rst), .Q(sreg[1839])
         );
  DFF \sreg_reg[1840]  ( .D(swire[817]), .CLK(clk), .RST(rst), .Q(sreg[1840])
         );
  DFF \sreg_reg[1841]  ( .D(swire[818]), .CLK(clk), .RST(rst), .Q(sreg[1841])
         );
  DFF \sreg_reg[1842]  ( .D(swire[819]), .CLK(clk), .RST(rst), .Q(sreg[1842])
         );
  DFF \sreg_reg[1843]  ( .D(swire[820]), .CLK(clk), .RST(rst), .Q(sreg[1843])
         );
  DFF \sreg_reg[1844]  ( .D(swire[821]), .CLK(clk), .RST(rst), .Q(sreg[1844])
         );
  DFF \sreg_reg[1845]  ( .D(swire[822]), .CLK(clk), .RST(rst), .Q(sreg[1845])
         );
  DFF \sreg_reg[1846]  ( .D(swire[823]), .CLK(clk), .RST(rst), .Q(sreg[1846])
         );
  DFF \sreg_reg[1847]  ( .D(swire[824]), .CLK(clk), .RST(rst), .Q(sreg[1847])
         );
  DFF \sreg_reg[1848]  ( .D(swire[825]), .CLK(clk), .RST(rst), .Q(sreg[1848])
         );
  DFF \sreg_reg[1849]  ( .D(swire[826]), .CLK(clk), .RST(rst), .Q(sreg[1849])
         );
  DFF \sreg_reg[1850]  ( .D(swire[827]), .CLK(clk), .RST(rst), .Q(sreg[1850])
         );
  DFF \sreg_reg[1851]  ( .D(swire[828]), .CLK(clk), .RST(rst), .Q(sreg[1851])
         );
  DFF \sreg_reg[1852]  ( .D(swire[829]), .CLK(clk), .RST(rst), .Q(sreg[1852])
         );
  DFF \sreg_reg[1853]  ( .D(swire[830]), .CLK(clk), .RST(rst), .Q(sreg[1853])
         );
  DFF \sreg_reg[1854]  ( .D(swire[831]), .CLK(clk), .RST(rst), .Q(sreg[1854])
         );
  DFF \sreg_reg[1855]  ( .D(swire[832]), .CLK(clk), .RST(rst), .Q(sreg[1855])
         );
  DFF \sreg_reg[1856]  ( .D(swire[833]), .CLK(clk), .RST(rst), .Q(sreg[1856])
         );
  DFF \sreg_reg[1857]  ( .D(swire[834]), .CLK(clk), .RST(rst), .Q(sreg[1857])
         );
  DFF \sreg_reg[1858]  ( .D(swire[835]), .CLK(clk), .RST(rst), .Q(sreg[1858])
         );
  DFF \sreg_reg[1859]  ( .D(swire[836]), .CLK(clk), .RST(rst), .Q(sreg[1859])
         );
  DFF \sreg_reg[1860]  ( .D(swire[837]), .CLK(clk), .RST(rst), .Q(sreg[1860])
         );
  DFF \sreg_reg[1861]  ( .D(swire[838]), .CLK(clk), .RST(rst), .Q(sreg[1861])
         );
  DFF \sreg_reg[1862]  ( .D(swire[839]), .CLK(clk), .RST(rst), .Q(sreg[1862])
         );
  DFF \sreg_reg[1863]  ( .D(swire[840]), .CLK(clk), .RST(rst), .Q(sreg[1863])
         );
  DFF \sreg_reg[1864]  ( .D(swire[841]), .CLK(clk), .RST(rst), .Q(sreg[1864])
         );
  DFF \sreg_reg[1865]  ( .D(swire[842]), .CLK(clk), .RST(rst), .Q(sreg[1865])
         );
  DFF \sreg_reg[1866]  ( .D(swire[843]), .CLK(clk), .RST(rst), .Q(sreg[1866])
         );
  DFF \sreg_reg[1867]  ( .D(swire[844]), .CLK(clk), .RST(rst), .Q(sreg[1867])
         );
  DFF \sreg_reg[1868]  ( .D(swire[845]), .CLK(clk), .RST(rst), .Q(sreg[1868])
         );
  DFF \sreg_reg[1869]  ( .D(swire[846]), .CLK(clk), .RST(rst), .Q(sreg[1869])
         );
  DFF \sreg_reg[1870]  ( .D(swire[847]), .CLK(clk), .RST(rst), .Q(sreg[1870])
         );
  DFF \sreg_reg[1871]  ( .D(swire[848]), .CLK(clk), .RST(rst), .Q(sreg[1871])
         );
  DFF \sreg_reg[1872]  ( .D(swire[849]), .CLK(clk), .RST(rst), .Q(sreg[1872])
         );
  DFF \sreg_reg[1873]  ( .D(swire[850]), .CLK(clk), .RST(rst), .Q(sreg[1873])
         );
  DFF \sreg_reg[1874]  ( .D(swire[851]), .CLK(clk), .RST(rst), .Q(sreg[1874])
         );
  DFF \sreg_reg[1875]  ( .D(swire[852]), .CLK(clk), .RST(rst), .Q(sreg[1875])
         );
  DFF \sreg_reg[1876]  ( .D(swire[853]), .CLK(clk), .RST(rst), .Q(sreg[1876])
         );
  DFF \sreg_reg[1877]  ( .D(swire[854]), .CLK(clk), .RST(rst), .Q(sreg[1877])
         );
  DFF \sreg_reg[1878]  ( .D(swire[855]), .CLK(clk), .RST(rst), .Q(sreg[1878])
         );
  DFF \sreg_reg[1879]  ( .D(swire[856]), .CLK(clk), .RST(rst), .Q(sreg[1879])
         );
  DFF \sreg_reg[1880]  ( .D(swire[857]), .CLK(clk), .RST(rst), .Q(sreg[1880])
         );
  DFF \sreg_reg[1881]  ( .D(swire[858]), .CLK(clk), .RST(rst), .Q(sreg[1881])
         );
  DFF \sreg_reg[1882]  ( .D(swire[859]), .CLK(clk), .RST(rst), .Q(sreg[1882])
         );
  DFF \sreg_reg[1883]  ( .D(swire[860]), .CLK(clk), .RST(rst), .Q(sreg[1883])
         );
  DFF \sreg_reg[1884]  ( .D(swire[861]), .CLK(clk), .RST(rst), .Q(sreg[1884])
         );
  DFF \sreg_reg[1885]  ( .D(swire[862]), .CLK(clk), .RST(rst), .Q(sreg[1885])
         );
  DFF \sreg_reg[1886]  ( .D(swire[863]), .CLK(clk), .RST(rst), .Q(sreg[1886])
         );
  DFF \sreg_reg[1887]  ( .D(swire[864]), .CLK(clk), .RST(rst), .Q(sreg[1887])
         );
  DFF \sreg_reg[1888]  ( .D(swire[865]), .CLK(clk), .RST(rst), .Q(sreg[1888])
         );
  DFF \sreg_reg[1889]  ( .D(swire[866]), .CLK(clk), .RST(rst), .Q(sreg[1889])
         );
  DFF \sreg_reg[1890]  ( .D(swire[867]), .CLK(clk), .RST(rst), .Q(sreg[1890])
         );
  DFF \sreg_reg[1891]  ( .D(swire[868]), .CLK(clk), .RST(rst), .Q(sreg[1891])
         );
  DFF \sreg_reg[1892]  ( .D(swire[869]), .CLK(clk), .RST(rst), .Q(sreg[1892])
         );
  DFF \sreg_reg[1893]  ( .D(swire[870]), .CLK(clk), .RST(rst), .Q(sreg[1893])
         );
  DFF \sreg_reg[1894]  ( .D(swire[871]), .CLK(clk), .RST(rst), .Q(sreg[1894])
         );
  DFF \sreg_reg[1895]  ( .D(swire[872]), .CLK(clk), .RST(rst), .Q(sreg[1895])
         );
  DFF \sreg_reg[1896]  ( .D(swire[873]), .CLK(clk), .RST(rst), .Q(sreg[1896])
         );
  DFF \sreg_reg[1897]  ( .D(swire[874]), .CLK(clk), .RST(rst), .Q(sreg[1897])
         );
  DFF \sreg_reg[1898]  ( .D(swire[875]), .CLK(clk), .RST(rst), .Q(sreg[1898])
         );
  DFF \sreg_reg[1899]  ( .D(swire[876]), .CLK(clk), .RST(rst), .Q(sreg[1899])
         );
  DFF \sreg_reg[1900]  ( .D(swire[877]), .CLK(clk), .RST(rst), .Q(sreg[1900])
         );
  DFF \sreg_reg[1901]  ( .D(swire[878]), .CLK(clk), .RST(rst), .Q(sreg[1901])
         );
  DFF \sreg_reg[1902]  ( .D(swire[879]), .CLK(clk), .RST(rst), .Q(sreg[1902])
         );
  DFF \sreg_reg[1903]  ( .D(swire[880]), .CLK(clk), .RST(rst), .Q(sreg[1903])
         );
  DFF \sreg_reg[1904]  ( .D(swire[881]), .CLK(clk), .RST(rst), .Q(sreg[1904])
         );
  DFF \sreg_reg[1905]  ( .D(swire[882]), .CLK(clk), .RST(rst), .Q(sreg[1905])
         );
  DFF \sreg_reg[1906]  ( .D(swire[883]), .CLK(clk), .RST(rst), .Q(sreg[1906])
         );
  DFF \sreg_reg[1907]  ( .D(swire[884]), .CLK(clk), .RST(rst), .Q(sreg[1907])
         );
  DFF \sreg_reg[1908]  ( .D(swire[885]), .CLK(clk), .RST(rst), .Q(sreg[1908])
         );
  DFF \sreg_reg[1909]  ( .D(swire[886]), .CLK(clk), .RST(rst), .Q(sreg[1909])
         );
  DFF \sreg_reg[1910]  ( .D(swire[887]), .CLK(clk), .RST(rst), .Q(sreg[1910])
         );
  DFF \sreg_reg[1911]  ( .D(swire[888]), .CLK(clk), .RST(rst), .Q(sreg[1911])
         );
  DFF \sreg_reg[1912]  ( .D(swire[889]), .CLK(clk), .RST(rst), .Q(sreg[1912])
         );
  DFF \sreg_reg[1913]  ( .D(swire[890]), .CLK(clk), .RST(rst), .Q(sreg[1913])
         );
  DFF \sreg_reg[1914]  ( .D(swire[891]), .CLK(clk), .RST(rst), .Q(sreg[1914])
         );
  DFF \sreg_reg[1915]  ( .D(swire[892]), .CLK(clk), .RST(rst), .Q(sreg[1915])
         );
  DFF \sreg_reg[1916]  ( .D(swire[893]), .CLK(clk), .RST(rst), .Q(sreg[1916])
         );
  DFF \sreg_reg[1917]  ( .D(swire[894]), .CLK(clk), .RST(rst), .Q(sreg[1917])
         );
  DFF \sreg_reg[1918]  ( .D(swire[895]), .CLK(clk), .RST(rst), .Q(sreg[1918])
         );
  DFF \sreg_reg[1919]  ( .D(swire[896]), .CLK(clk), .RST(rst), .Q(sreg[1919])
         );
  DFF \sreg_reg[1920]  ( .D(swire[897]), .CLK(clk), .RST(rst), .Q(sreg[1920])
         );
  DFF \sreg_reg[1921]  ( .D(swire[898]), .CLK(clk), .RST(rst), .Q(sreg[1921])
         );
  DFF \sreg_reg[1922]  ( .D(swire[899]), .CLK(clk), .RST(rst), .Q(sreg[1922])
         );
  DFF \sreg_reg[1923]  ( .D(swire[900]), .CLK(clk), .RST(rst), .Q(sreg[1923])
         );
  DFF \sreg_reg[1924]  ( .D(swire[901]), .CLK(clk), .RST(rst), .Q(sreg[1924])
         );
  DFF \sreg_reg[1925]  ( .D(swire[902]), .CLK(clk), .RST(rst), .Q(sreg[1925])
         );
  DFF \sreg_reg[1926]  ( .D(swire[903]), .CLK(clk), .RST(rst), .Q(sreg[1926])
         );
  DFF \sreg_reg[1927]  ( .D(swire[904]), .CLK(clk), .RST(rst), .Q(sreg[1927])
         );
  DFF \sreg_reg[1928]  ( .D(swire[905]), .CLK(clk), .RST(rst), .Q(sreg[1928])
         );
  DFF \sreg_reg[1929]  ( .D(swire[906]), .CLK(clk), .RST(rst), .Q(sreg[1929])
         );
  DFF \sreg_reg[1930]  ( .D(swire[907]), .CLK(clk), .RST(rst), .Q(sreg[1930])
         );
  DFF \sreg_reg[1931]  ( .D(swire[908]), .CLK(clk), .RST(rst), .Q(sreg[1931])
         );
  DFF \sreg_reg[1932]  ( .D(swire[909]), .CLK(clk), .RST(rst), .Q(sreg[1932])
         );
  DFF \sreg_reg[1933]  ( .D(swire[910]), .CLK(clk), .RST(rst), .Q(sreg[1933])
         );
  DFF \sreg_reg[1934]  ( .D(swire[911]), .CLK(clk), .RST(rst), .Q(sreg[1934])
         );
  DFF \sreg_reg[1935]  ( .D(swire[912]), .CLK(clk), .RST(rst), .Q(sreg[1935])
         );
  DFF \sreg_reg[1936]  ( .D(swire[913]), .CLK(clk), .RST(rst), .Q(sreg[1936])
         );
  DFF \sreg_reg[1937]  ( .D(swire[914]), .CLK(clk), .RST(rst), .Q(sreg[1937])
         );
  DFF \sreg_reg[1938]  ( .D(swire[915]), .CLK(clk), .RST(rst), .Q(sreg[1938])
         );
  DFF \sreg_reg[1939]  ( .D(swire[916]), .CLK(clk), .RST(rst), .Q(sreg[1939])
         );
  DFF \sreg_reg[1940]  ( .D(swire[917]), .CLK(clk), .RST(rst), .Q(sreg[1940])
         );
  DFF \sreg_reg[1941]  ( .D(swire[918]), .CLK(clk), .RST(rst), .Q(sreg[1941])
         );
  DFF \sreg_reg[1942]  ( .D(swire[919]), .CLK(clk), .RST(rst), .Q(sreg[1942])
         );
  DFF \sreg_reg[1943]  ( .D(swire[920]), .CLK(clk), .RST(rst), .Q(sreg[1943])
         );
  DFF \sreg_reg[1944]  ( .D(swire[921]), .CLK(clk), .RST(rst), .Q(sreg[1944])
         );
  DFF \sreg_reg[1945]  ( .D(swire[922]), .CLK(clk), .RST(rst), .Q(sreg[1945])
         );
  DFF \sreg_reg[1946]  ( .D(swire[923]), .CLK(clk), .RST(rst), .Q(sreg[1946])
         );
  DFF \sreg_reg[1947]  ( .D(swire[924]), .CLK(clk), .RST(rst), .Q(sreg[1947])
         );
  DFF \sreg_reg[1948]  ( .D(swire[925]), .CLK(clk), .RST(rst), .Q(sreg[1948])
         );
  DFF \sreg_reg[1949]  ( .D(swire[926]), .CLK(clk), .RST(rst), .Q(sreg[1949])
         );
  DFF \sreg_reg[1950]  ( .D(swire[927]), .CLK(clk), .RST(rst), .Q(sreg[1950])
         );
  DFF \sreg_reg[1951]  ( .D(swire[928]), .CLK(clk), .RST(rst), .Q(sreg[1951])
         );
  DFF \sreg_reg[1952]  ( .D(swire[929]), .CLK(clk), .RST(rst), .Q(sreg[1952])
         );
  DFF \sreg_reg[1953]  ( .D(swire[930]), .CLK(clk), .RST(rst), .Q(sreg[1953])
         );
  DFF \sreg_reg[1954]  ( .D(swire[931]), .CLK(clk), .RST(rst), .Q(sreg[1954])
         );
  DFF \sreg_reg[1955]  ( .D(swire[932]), .CLK(clk), .RST(rst), .Q(sreg[1955])
         );
  DFF \sreg_reg[1956]  ( .D(swire[933]), .CLK(clk), .RST(rst), .Q(sreg[1956])
         );
  DFF \sreg_reg[1957]  ( .D(swire[934]), .CLK(clk), .RST(rst), .Q(sreg[1957])
         );
  DFF \sreg_reg[1958]  ( .D(swire[935]), .CLK(clk), .RST(rst), .Q(sreg[1958])
         );
  DFF \sreg_reg[1959]  ( .D(swire[936]), .CLK(clk), .RST(rst), .Q(sreg[1959])
         );
  DFF \sreg_reg[1960]  ( .D(swire[937]), .CLK(clk), .RST(rst), .Q(sreg[1960])
         );
  DFF \sreg_reg[1961]  ( .D(swire[938]), .CLK(clk), .RST(rst), .Q(sreg[1961])
         );
  DFF \sreg_reg[1962]  ( .D(swire[939]), .CLK(clk), .RST(rst), .Q(sreg[1962])
         );
  DFF \sreg_reg[1963]  ( .D(swire[940]), .CLK(clk), .RST(rst), .Q(sreg[1963])
         );
  DFF \sreg_reg[1964]  ( .D(swire[941]), .CLK(clk), .RST(rst), .Q(sreg[1964])
         );
  DFF \sreg_reg[1965]  ( .D(swire[942]), .CLK(clk), .RST(rst), .Q(sreg[1965])
         );
  DFF \sreg_reg[1966]  ( .D(swire[943]), .CLK(clk), .RST(rst), .Q(sreg[1966])
         );
  DFF \sreg_reg[1967]  ( .D(swire[944]), .CLK(clk), .RST(rst), .Q(sreg[1967])
         );
  DFF \sreg_reg[1968]  ( .D(swire[945]), .CLK(clk), .RST(rst), .Q(sreg[1968])
         );
  DFF \sreg_reg[1969]  ( .D(swire[946]), .CLK(clk), .RST(rst), .Q(sreg[1969])
         );
  DFF \sreg_reg[1970]  ( .D(swire[947]), .CLK(clk), .RST(rst), .Q(sreg[1970])
         );
  DFF \sreg_reg[1971]  ( .D(swire[948]), .CLK(clk), .RST(rst), .Q(sreg[1971])
         );
  DFF \sreg_reg[1972]  ( .D(swire[949]), .CLK(clk), .RST(rst), .Q(sreg[1972])
         );
  DFF \sreg_reg[1973]  ( .D(swire[950]), .CLK(clk), .RST(rst), .Q(sreg[1973])
         );
  DFF \sreg_reg[1974]  ( .D(swire[951]), .CLK(clk), .RST(rst), .Q(sreg[1974])
         );
  DFF \sreg_reg[1975]  ( .D(swire[952]), .CLK(clk), .RST(rst), .Q(sreg[1975])
         );
  DFF \sreg_reg[1976]  ( .D(swire[953]), .CLK(clk), .RST(rst), .Q(sreg[1976])
         );
  DFF \sreg_reg[1977]  ( .D(swire[954]), .CLK(clk), .RST(rst), .Q(sreg[1977])
         );
  DFF \sreg_reg[1978]  ( .D(swire[955]), .CLK(clk), .RST(rst), .Q(sreg[1978])
         );
  DFF \sreg_reg[1979]  ( .D(swire[956]), .CLK(clk), .RST(rst), .Q(sreg[1979])
         );
  DFF \sreg_reg[1980]  ( .D(swire[957]), .CLK(clk), .RST(rst), .Q(sreg[1980])
         );
  DFF \sreg_reg[1981]  ( .D(swire[958]), .CLK(clk), .RST(rst), .Q(sreg[1981])
         );
  DFF \sreg_reg[1982]  ( .D(swire[959]), .CLK(clk), .RST(rst), .Q(sreg[1982])
         );
  DFF \sreg_reg[1983]  ( .D(swire[960]), .CLK(clk), .RST(rst), .Q(sreg[1983])
         );
  DFF \sreg_reg[1984]  ( .D(swire[961]), .CLK(clk), .RST(rst), .Q(sreg[1984])
         );
  DFF \sreg_reg[1985]  ( .D(swire[962]), .CLK(clk), .RST(rst), .Q(sreg[1985])
         );
  DFF \sreg_reg[1986]  ( .D(swire[963]), .CLK(clk), .RST(rst), .Q(sreg[1986])
         );
  DFF \sreg_reg[1987]  ( .D(swire[964]), .CLK(clk), .RST(rst), .Q(sreg[1987])
         );
  DFF \sreg_reg[1988]  ( .D(swire[965]), .CLK(clk), .RST(rst), .Q(sreg[1988])
         );
  DFF \sreg_reg[1989]  ( .D(swire[966]), .CLK(clk), .RST(rst), .Q(sreg[1989])
         );
  DFF \sreg_reg[1990]  ( .D(swire[967]), .CLK(clk), .RST(rst), .Q(sreg[1990])
         );
  DFF \sreg_reg[1991]  ( .D(swire[968]), .CLK(clk), .RST(rst), .Q(sreg[1991])
         );
  DFF \sreg_reg[1992]  ( .D(swire[969]), .CLK(clk), .RST(rst), .Q(sreg[1992])
         );
  DFF \sreg_reg[1993]  ( .D(swire[970]), .CLK(clk), .RST(rst), .Q(sreg[1993])
         );
  DFF \sreg_reg[1994]  ( .D(swire[971]), .CLK(clk), .RST(rst), .Q(sreg[1994])
         );
  DFF \sreg_reg[1995]  ( .D(swire[972]), .CLK(clk), .RST(rst), .Q(sreg[1995])
         );
  DFF \sreg_reg[1996]  ( .D(swire[973]), .CLK(clk), .RST(rst), .Q(sreg[1996])
         );
  DFF \sreg_reg[1997]  ( .D(swire[974]), .CLK(clk), .RST(rst), .Q(sreg[1997])
         );
  DFF \sreg_reg[1998]  ( .D(swire[975]), .CLK(clk), .RST(rst), .Q(sreg[1998])
         );
  DFF \sreg_reg[1999]  ( .D(swire[976]), .CLK(clk), .RST(rst), .Q(sreg[1999])
         );
  DFF \sreg_reg[2000]  ( .D(swire[977]), .CLK(clk), .RST(rst), .Q(sreg[2000])
         );
  DFF \sreg_reg[2001]  ( .D(swire[978]), .CLK(clk), .RST(rst), .Q(sreg[2001])
         );
  DFF \sreg_reg[2002]  ( .D(swire[979]), .CLK(clk), .RST(rst), .Q(sreg[2002])
         );
  DFF \sreg_reg[2003]  ( .D(swire[980]), .CLK(clk), .RST(rst), .Q(sreg[2003])
         );
  DFF \sreg_reg[2004]  ( .D(swire[981]), .CLK(clk), .RST(rst), .Q(sreg[2004])
         );
  DFF \sreg_reg[2005]  ( .D(swire[982]), .CLK(clk), .RST(rst), .Q(sreg[2005])
         );
  DFF \sreg_reg[2006]  ( .D(swire[983]), .CLK(clk), .RST(rst), .Q(sreg[2006])
         );
  DFF \sreg_reg[2007]  ( .D(swire[984]), .CLK(clk), .RST(rst), .Q(sreg[2007])
         );
  DFF \sreg_reg[2008]  ( .D(swire[985]), .CLK(clk), .RST(rst), .Q(sreg[2008])
         );
  DFF \sreg_reg[2009]  ( .D(swire[986]), .CLK(clk), .RST(rst), .Q(sreg[2009])
         );
  DFF \sreg_reg[2010]  ( .D(swire[987]), .CLK(clk), .RST(rst), .Q(sreg[2010])
         );
  DFF \sreg_reg[2011]  ( .D(swire[988]), .CLK(clk), .RST(rst), .Q(sreg[2011])
         );
  DFF \sreg_reg[2012]  ( .D(swire[989]), .CLK(clk), .RST(rst), .Q(sreg[2012])
         );
  DFF \sreg_reg[2013]  ( .D(swire[990]), .CLK(clk), .RST(rst), .Q(sreg[2013])
         );
  DFF \sreg_reg[2014]  ( .D(swire[991]), .CLK(clk), .RST(rst), .Q(sreg[2014])
         );
  DFF \sreg_reg[2015]  ( .D(swire[992]), .CLK(clk), .RST(rst), .Q(sreg[2015])
         );
  DFF \sreg_reg[2016]  ( .D(swire[993]), .CLK(clk), .RST(rst), .Q(sreg[2016])
         );
  DFF \sreg_reg[2017]  ( .D(swire[994]), .CLK(clk), .RST(rst), .Q(sreg[2017])
         );
  DFF \sreg_reg[2018]  ( .D(swire[995]), .CLK(clk), .RST(rst), .Q(sreg[2018])
         );
  DFF \sreg_reg[2019]  ( .D(swire[996]), .CLK(clk), .RST(rst), .Q(sreg[2019])
         );
  DFF \sreg_reg[2020]  ( .D(swire[997]), .CLK(clk), .RST(rst), .Q(sreg[2020])
         );
  DFF \sreg_reg[2021]  ( .D(swire[998]), .CLK(clk), .RST(rst), .Q(sreg[2021])
         );
  DFF \sreg_reg[2022]  ( .D(swire[999]), .CLK(clk), .RST(rst), .Q(sreg[2022])
         );
  DFF \sreg_reg[2023]  ( .D(swire[1000]), .CLK(clk), .RST(rst), .Q(sreg[2023])
         );
  DFF \sreg_reg[2024]  ( .D(swire[1001]), .CLK(clk), .RST(rst), .Q(sreg[2024])
         );
  DFF \sreg_reg[2025]  ( .D(swire[1002]), .CLK(clk), .RST(rst), .Q(sreg[2025])
         );
  DFF \sreg_reg[2026]  ( .D(swire[1003]), .CLK(clk), .RST(rst), .Q(sreg[2026])
         );
  DFF \sreg_reg[2027]  ( .D(swire[1004]), .CLK(clk), .RST(rst), .Q(sreg[2027])
         );
  DFF \sreg_reg[2028]  ( .D(swire[1005]), .CLK(clk), .RST(rst), .Q(sreg[2028])
         );
  DFF \sreg_reg[2029]  ( .D(swire[1006]), .CLK(clk), .RST(rst), .Q(sreg[2029])
         );
  DFF \sreg_reg[2030]  ( .D(swire[1007]), .CLK(clk), .RST(rst), .Q(sreg[2030])
         );
  DFF \sreg_reg[2031]  ( .D(swire[1008]), .CLK(clk), .RST(rst), .Q(sreg[2031])
         );
  DFF \sreg_reg[2032]  ( .D(swire[1009]), .CLK(clk), .RST(rst), .Q(sreg[2032])
         );
  DFF \sreg_reg[2033]  ( .D(swire[1010]), .CLK(clk), .RST(rst), .Q(sreg[2033])
         );
  DFF \sreg_reg[2034]  ( .D(swire[1011]), .CLK(clk), .RST(rst), .Q(sreg[2034])
         );
  DFF \sreg_reg[2035]  ( .D(swire[1012]), .CLK(clk), .RST(rst), .Q(sreg[2035])
         );
  DFF \sreg_reg[2036]  ( .D(swire[1013]), .CLK(clk), .RST(rst), .Q(sreg[2036])
         );
  DFF \sreg_reg[2037]  ( .D(swire[1014]), .CLK(clk), .RST(rst), .Q(sreg[2037])
         );
  DFF \sreg_reg[2038]  ( .D(swire[1015]), .CLK(clk), .RST(rst), .Q(sreg[2038])
         );
  DFF \sreg_reg[2039]  ( .D(swire[1016]), .CLK(clk), .RST(rst), .Q(sreg[2039])
         );
  DFF \sreg_reg[2040]  ( .D(swire[1017]), .CLK(clk), .RST(rst), .Q(sreg[2040])
         );
  DFF \sreg_reg[2041]  ( .D(swire[1018]), .CLK(clk), .RST(rst), .Q(sreg[2041])
         );
  DFF \sreg_reg[2042]  ( .D(swire[1019]), .CLK(clk), .RST(rst), .Q(sreg[2042])
         );
  DFF \sreg_reg[2043]  ( .D(swire[1020]), .CLK(clk), .RST(rst), .Q(sreg[2043])
         );
  DFF \sreg_reg[2044]  ( .D(swire[1021]), .CLK(clk), .RST(rst), .Q(sreg[2044])
         );
  DFF \sreg_reg[2045]  ( .D(swire[1022]), .CLK(clk), .RST(rst), .Q(sreg[2045])
         );
  DFF \sreg_reg[2046]  ( .D(swire[1023]), .CLK(clk), .RST(rst), .Q(sreg[2046])
         );
  DFF \sreg_reg[1023]  ( .D(c[1023]), .CLK(clk), .RST(rst), .Q(c[1022]) );
  DFF \sreg_reg[1022]  ( .D(c[1022]), .CLK(clk), .RST(rst), .Q(c[1021]) );
  DFF \sreg_reg[1021]  ( .D(c[1021]), .CLK(clk), .RST(rst), .Q(c[1020]) );
  DFF \sreg_reg[1020]  ( .D(c[1020]), .CLK(clk), .RST(rst), .Q(c[1019]) );
  DFF \sreg_reg[1019]  ( .D(c[1019]), .CLK(clk), .RST(rst), .Q(c[1018]) );
  DFF \sreg_reg[1018]  ( .D(c[1018]), .CLK(clk), .RST(rst), .Q(c[1017]) );
  DFF \sreg_reg[1017]  ( .D(c[1017]), .CLK(clk), .RST(rst), .Q(c[1016]) );
  DFF \sreg_reg[1016]  ( .D(c[1016]), .CLK(clk), .RST(rst), .Q(c[1015]) );
  DFF \sreg_reg[1015]  ( .D(c[1015]), .CLK(clk), .RST(rst), .Q(c[1014]) );
  DFF \sreg_reg[1014]  ( .D(c[1014]), .CLK(clk), .RST(rst), .Q(c[1013]) );
  DFF \sreg_reg[1013]  ( .D(c[1013]), .CLK(clk), .RST(rst), .Q(c[1012]) );
  DFF \sreg_reg[1012]  ( .D(c[1012]), .CLK(clk), .RST(rst), .Q(c[1011]) );
  DFF \sreg_reg[1011]  ( .D(c[1011]), .CLK(clk), .RST(rst), .Q(c[1010]) );
  DFF \sreg_reg[1010]  ( .D(c[1010]), .CLK(clk), .RST(rst), .Q(c[1009]) );
  DFF \sreg_reg[1009]  ( .D(c[1009]), .CLK(clk), .RST(rst), .Q(c[1008]) );
  DFF \sreg_reg[1008]  ( .D(c[1008]), .CLK(clk), .RST(rst), .Q(c[1007]) );
  DFF \sreg_reg[1007]  ( .D(c[1007]), .CLK(clk), .RST(rst), .Q(c[1006]) );
  DFF \sreg_reg[1006]  ( .D(c[1006]), .CLK(clk), .RST(rst), .Q(c[1005]) );
  DFF \sreg_reg[1005]  ( .D(c[1005]), .CLK(clk), .RST(rst), .Q(c[1004]) );
  DFF \sreg_reg[1004]  ( .D(c[1004]), .CLK(clk), .RST(rst), .Q(c[1003]) );
  DFF \sreg_reg[1003]  ( .D(c[1003]), .CLK(clk), .RST(rst), .Q(c[1002]) );
  DFF \sreg_reg[1002]  ( .D(c[1002]), .CLK(clk), .RST(rst), .Q(c[1001]) );
  DFF \sreg_reg[1001]  ( .D(c[1001]), .CLK(clk), .RST(rst), .Q(c[1000]) );
  DFF \sreg_reg[1000]  ( .D(c[1000]), .CLK(clk), .RST(rst), .Q(c[999]) );
  DFF \sreg_reg[999]  ( .D(c[999]), .CLK(clk), .RST(rst), .Q(c[998]) );
  DFF \sreg_reg[998]  ( .D(c[998]), .CLK(clk), .RST(rst), .Q(c[997]) );
  DFF \sreg_reg[997]  ( .D(c[997]), .CLK(clk), .RST(rst), .Q(c[996]) );
  DFF \sreg_reg[996]  ( .D(c[996]), .CLK(clk), .RST(rst), .Q(c[995]) );
  DFF \sreg_reg[995]  ( .D(c[995]), .CLK(clk), .RST(rst), .Q(c[994]) );
  DFF \sreg_reg[994]  ( .D(c[994]), .CLK(clk), .RST(rst), .Q(c[993]) );
  DFF \sreg_reg[993]  ( .D(c[993]), .CLK(clk), .RST(rst), .Q(c[992]) );
  DFF \sreg_reg[992]  ( .D(c[992]), .CLK(clk), .RST(rst), .Q(c[991]) );
  DFF \sreg_reg[991]  ( .D(c[991]), .CLK(clk), .RST(rst), .Q(c[990]) );
  DFF \sreg_reg[990]  ( .D(c[990]), .CLK(clk), .RST(rst), .Q(c[989]) );
  DFF \sreg_reg[989]  ( .D(c[989]), .CLK(clk), .RST(rst), .Q(c[988]) );
  DFF \sreg_reg[988]  ( .D(c[988]), .CLK(clk), .RST(rst), .Q(c[987]) );
  DFF \sreg_reg[987]  ( .D(c[987]), .CLK(clk), .RST(rst), .Q(c[986]) );
  DFF \sreg_reg[986]  ( .D(c[986]), .CLK(clk), .RST(rst), .Q(c[985]) );
  DFF \sreg_reg[985]  ( .D(c[985]), .CLK(clk), .RST(rst), .Q(c[984]) );
  DFF \sreg_reg[984]  ( .D(c[984]), .CLK(clk), .RST(rst), .Q(c[983]) );
  DFF \sreg_reg[983]  ( .D(c[983]), .CLK(clk), .RST(rst), .Q(c[982]) );
  DFF \sreg_reg[982]  ( .D(c[982]), .CLK(clk), .RST(rst), .Q(c[981]) );
  DFF \sreg_reg[981]  ( .D(c[981]), .CLK(clk), .RST(rst), .Q(c[980]) );
  DFF \sreg_reg[980]  ( .D(c[980]), .CLK(clk), .RST(rst), .Q(c[979]) );
  DFF \sreg_reg[979]  ( .D(c[979]), .CLK(clk), .RST(rst), .Q(c[978]) );
  DFF \sreg_reg[978]  ( .D(c[978]), .CLK(clk), .RST(rst), .Q(c[977]) );
  DFF \sreg_reg[977]  ( .D(c[977]), .CLK(clk), .RST(rst), .Q(c[976]) );
  DFF \sreg_reg[976]  ( .D(c[976]), .CLK(clk), .RST(rst), .Q(c[975]) );
  DFF \sreg_reg[975]  ( .D(c[975]), .CLK(clk), .RST(rst), .Q(c[974]) );
  DFF \sreg_reg[974]  ( .D(c[974]), .CLK(clk), .RST(rst), .Q(c[973]) );
  DFF \sreg_reg[973]  ( .D(c[973]), .CLK(clk), .RST(rst), .Q(c[972]) );
  DFF \sreg_reg[972]  ( .D(c[972]), .CLK(clk), .RST(rst), .Q(c[971]) );
  DFF \sreg_reg[971]  ( .D(c[971]), .CLK(clk), .RST(rst), .Q(c[970]) );
  DFF \sreg_reg[970]  ( .D(c[970]), .CLK(clk), .RST(rst), .Q(c[969]) );
  DFF \sreg_reg[969]  ( .D(c[969]), .CLK(clk), .RST(rst), .Q(c[968]) );
  DFF \sreg_reg[968]  ( .D(c[968]), .CLK(clk), .RST(rst), .Q(c[967]) );
  DFF \sreg_reg[967]  ( .D(c[967]), .CLK(clk), .RST(rst), .Q(c[966]) );
  DFF \sreg_reg[966]  ( .D(c[966]), .CLK(clk), .RST(rst), .Q(c[965]) );
  DFF \sreg_reg[965]  ( .D(c[965]), .CLK(clk), .RST(rst), .Q(c[964]) );
  DFF \sreg_reg[964]  ( .D(c[964]), .CLK(clk), .RST(rst), .Q(c[963]) );
  DFF \sreg_reg[963]  ( .D(c[963]), .CLK(clk), .RST(rst), .Q(c[962]) );
  DFF \sreg_reg[962]  ( .D(c[962]), .CLK(clk), .RST(rst), .Q(c[961]) );
  DFF \sreg_reg[961]  ( .D(c[961]), .CLK(clk), .RST(rst), .Q(c[960]) );
  DFF \sreg_reg[960]  ( .D(c[960]), .CLK(clk), .RST(rst), .Q(c[959]) );
  DFF \sreg_reg[959]  ( .D(c[959]), .CLK(clk), .RST(rst), .Q(c[958]) );
  DFF \sreg_reg[958]  ( .D(c[958]), .CLK(clk), .RST(rst), .Q(c[957]) );
  DFF \sreg_reg[957]  ( .D(c[957]), .CLK(clk), .RST(rst), .Q(c[956]) );
  DFF \sreg_reg[956]  ( .D(c[956]), .CLK(clk), .RST(rst), .Q(c[955]) );
  DFF \sreg_reg[955]  ( .D(c[955]), .CLK(clk), .RST(rst), .Q(c[954]) );
  DFF \sreg_reg[954]  ( .D(c[954]), .CLK(clk), .RST(rst), .Q(c[953]) );
  DFF \sreg_reg[953]  ( .D(c[953]), .CLK(clk), .RST(rst), .Q(c[952]) );
  DFF \sreg_reg[952]  ( .D(c[952]), .CLK(clk), .RST(rst), .Q(c[951]) );
  DFF \sreg_reg[951]  ( .D(c[951]), .CLK(clk), .RST(rst), .Q(c[950]) );
  DFF \sreg_reg[950]  ( .D(c[950]), .CLK(clk), .RST(rst), .Q(c[949]) );
  DFF \sreg_reg[949]  ( .D(c[949]), .CLK(clk), .RST(rst), .Q(c[948]) );
  DFF \sreg_reg[948]  ( .D(c[948]), .CLK(clk), .RST(rst), .Q(c[947]) );
  DFF \sreg_reg[947]  ( .D(c[947]), .CLK(clk), .RST(rst), .Q(c[946]) );
  DFF \sreg_reg[946]  ( .D(c[946]), .CLK(clk), .RST(rst), .Q(c[945]) );
  DFF \sreg_reg[945]  ( .D(c[945]), .CLK(clk), .RST(rst), .Q(c[944]) );
  DFF \sreg_reg[944]  ( .D(c[944]), .CLK(clk), .RST(rst), .Q(c[943]) );
  DFF \sreg_reg[943]  ( .D(c[943]), .CLK(clk), .RST(rst), .Q(c[942]) );
  DFF \sreg_reg[942]  ( .D(c[942]), .CLK(clk), .RST(rst), .Q(c[941]) );
  DFF \sreg_reg[941]  ( .D(c[941]), .CLK(clk), .RST(rst), .Q(c[940]) );
  DFF \sreg_reg[940]  ( .D(c[940]), .CLK(clk), .RST(rst), .Q(c[939]) );
  DFF \sreg_reg[939]  ( .D(c[939]), .CLK(clk), .RST(rst), .Q(c[938]) );
  DFF \sreg_reg[938]  ( .D(c[938]), .CLK(clk), .RST(rst), .Q(c[937]) );
  DFF \sreg_reg[937]  ( .D(c[937]), .CLK(clk), .RST(rst), .Q(c[936]) );
  DFF \sreg_reg[936]  ( .D(c[936]), .CLK(clk), .RST(rst), .Q(c[935]) );
  DFF \sreg_reg[935]  ( .D(c[935]), .CLK(clk), .RST(rst), .Q(c[934]) );
  DFF \sreg_reg[934]  ( .D(c[934]), .CLK(clk), .RST(rst), .Q(c[933]) );
  DFF \sreg_reg[933]  ( .D(c[933]), .CLK(clk), .RST(rst), .Q(c[932]) );
  DFF \sreg_reg[932]  ( .D(c[932]), .CLK(clk), .RST(rst), .Q(c[931]) );
  DFF \sreg_reg[931]  ( .D(c[931]), .CLK(clk), .RST(rst), .Q(c[930]) );
  DFF \sreg_reg[930]  ( .D(c[930]), .CLK(clk), .RST(rst), .Q(c[929]) );
  DFF \sreg_reg[929]  ( .D(c[929]), .CLK(clk), .RST(rst), .Q(c[928]) );
  DFF \sreg_reg[928]  ( .D(c[928]), .CLK(clk), .RST(rst), .Q(c[927]) );
  DFF \sreg_reg[927]  ( .D(c[927]), .CLK(clk), .RST(rst), .Q(c[926]) );
  DFF \sreg_reg[926]  ( .D(c[926]), .CLK(clk), .RST(rst), .Q(c[925]) );
  DFF \sreg_reg[925]  ( .D(c[925]), .CLK(clk), .RST(rst), .Q(c[924]) );
  DFF \sreg_reg[924]  ( .D(c[924]), .CLK(clk), .RST(rst), .Q(c[923]) );
  DFF \sreg_reg[923]  ( .D(c[923]), .CLK(clk), .RST(rst), .Q(c[922]) );
  DFF \sreg_reg[922]  ( .D(c[922]), .CLK(clk), .RST(rst), .Q(c[921]) );
  DFF \sreg_reg[921]  ( .D(c[921]), .CLK(clk), .RST(rst), .Q(c[920]) );
  DFF \sreg_reg[920]  ( .D(c[920]), .CLK(clk), .RST(rst), .Q(c[919]) );
  DFF \sreg_reg[919]  ( .D(c[919]), .CLK(clk), .RST(rst), .Q(c[918]) );
  DFF \sreg_reg[918]  ( .D(c[918]), .CLK(clk), .RST(rst), .Q(c[917]) );
  DFF \sreg_reg[917]  ( .D(c[917]), .CLK(clk), .RST(rst), .Q(c[916]) );
  DFF \sreg_reg[916]  ( .D(c[916]), .CLK(clk), .RST(rst), .Q(c[915]) );
  DFF \sreg_reg[915]  ( .D(c[915]), .CLK(clk), .RST(rst), .Q(c[914]) );
  DFF \sreg_reg[914]  ( .D(c[914]), .CLK(clk), .RST(rst), .Q(c[913]) );
  DFF \sreg_reg[913]  ( .D(c[913]), .CLK(clk), .RST(rst), .Q(c[912]) );
  DFF \sreg_reg[912]  ( .D(c[912]), .CLK(clk), .RST(rst), .Q(c[911]) );
  DFF \sreg_reg[911]  ( .D(c[911]), .CLK(clk), .RST(rst), .Q(c[910]) );
  DFF \sreg_reg[910]  ( .D(c[910]), .CLK(clk), .RST(rst), .Q(c[909]) );
  DFF \sreg_reg[909]  ( .D(c[909]), .CLK(clk), .RST(rst), .Q(c[908]) );
  DFF \sreg_reg[908]  ( .D(c[908]), .CLK(clk), .RST(rst), .Q(c[907]) );
  DFF \sreg_reg[907]  ( .D(c[907]), .CLK(clk), .RST(rst), .Q(c[906]) );
  DFF \sreg_reg[906]  ( .D(c[906]), .CLK(clk), .RST(rst), .Q(c[905]) );
  DFF \sreg_reg[905]  ( .D(c[905]), .CLK(clk), .RST(rst), .Q(c[904]) );
  DFF \sreg_reg[904]  ( .D(c[904]), .CLK(clk), .RST(rst), .Q(c[903]) );
  DFF \sreg_reg[903]  ( .D(c[903]), .CLK(clk), .RST(rst), .Q(c[902]) );
  DFF \sreg_reg[902]  ( .D(c[902]), .CLK(clk), .RST(rst), .Q(c[901]) );
  DFF \sreg_reg[901]  ( .D(c[901]), .CLK(clk), .RST(rst), .Q(c[900]) );
  DFF \sreg_reg[900]  ( .D(c[900]), .CLK(clk), .RST(rst), .Q(c[899]) );
  DFF \sreg_reg[899]  ( .D(c[899]), .CLK(clk), .RST(rst), .Q(c[898]) );
  DFF \sreg_reg[898]  ( .D(c[898]), .CLK(clk), .RST(rst), .Q(c[897]) );
  DFF \sreg_reg[897]  ( .D(c[897]), .CLK(clk), .RST(rst), .Q(c[896]) );
  DFF \sreg_reg[896]  ( .D(c[896]), .CLK(clk), .RST(rst), .Q(c[895]) );
  DFF \sreg_reg[895]  ( .D(c[895]), .CLK(clk), .RST(rst), .Q(c[894]) );
  DFF \sreg_reg[894]  ( .D(c[894]), .CLK(clk), .RST(rst), .Q(c[893]) );
  DFF \sreg_reg[893]  ( .D(c[893]), .CLK(clk), .RST(rst), .Q(c[892]) );
  DFF \sreg_reg[892]  ( .D(c[892]), .CLK(clk), .RST(rst), .Q(c[891]) );
  DFF \sreg_reg[891]  ( .D(c[891]), .CLK(clk), .RST(rst), .Q(c[890]) );
  DFF \sreg_reg[890]  ( .D(c[890]), .CLK(clk), .RST(rst), .Q(c[889]) );
  DFF \sreg_reg[889]  ( .D(c[889]), .CLK(clk), .RST(rst), .Q(c[888]) );
  DFF \sreg_reg[888]  ( .D(c[888]), .CLK(clk), .RST(rst), .Q(c[887]) );
  DFF \sreg_reg[887]  ( .D(c[887]), .CLK(clk), .RST(rst), .Q(c[886]) );
  DFF \sreg_reg[886]  ( .D(c[886]), .CLK(clk), .RST(rst), .Q(c[885]) );
  DFF \sreg_reg[885]  ( .D(c[885]), .CLK(clk), .RST(rst), .Q(c[884]) );
  DFF \sreg_reg[884]  ( .D(c[884]), .CLK(clk), .RST(rst), .Q(c[883]) );
  DFF \sreg_reg[883]  ( .D(c[883]), .CLK(clk), .RST(rst), .Q(c[882]) );
  DFF \sreg_reg[882]  ( .D(c[882]), .CLK(clk), .RST(rst), .Q(c[881]) );
  DFF \sreg_reg[881]  ( .D(c[881]), .CLK(clk), .RST(rst), .Q(c[880]) );
  DFF \sreg_reg[880]  ( .D(c[880]), .CLK(clk), .RST(rst), .Q(c[879]) );
  DFF \sreg_reg[879]  ( .D(c[879]), .CLK(clk), .RST(rst), .Q(c[878]) );
  DFF \sreg_reg[878]  ( .D(c[878]), .CLK(clk), .RST(rst), .Q(c[877]) );
  DFF \sreg_reg[877]  ( .D(c[877]), .CLK(clk), .RST(rst), .Q(c[876]) );
  DFF \sreg_reg[876]  ( .D(c[876]), .CLK(clk), .RST(rst), .Q(c[875]) );
  DFF \sreg_reg[875]  ( .D(c[875]), .CLK(clk), .RST(rst), .Q(c[874]) );
  DFF \sreg_reg[874]  ( .D(c[874]), .CLK(clk), .RST(rst), .Q(c[873]) );
  DFF \sreg_reg[873]  ( .D(c[873]), .CLK(clk), .RST(rst), .Q(c[872]) );
  DFF \sreg_reg[872]  ( .D(c[872]), .CLK(clk), .RST(rst), .Q(c[871]) );
  DFF \sreg_reg[871]  ( .D(c[871]), .CLK(clk), .RST(rst), .Q(c[870]) );
  DFF \sreg_reg[870]  ( .D(c[870]), .CLK(clk), .RST(rst), .Q(c[869]) );
  DFF \sreg_reg[869]  ( .D(c[869]), .CLK(clk), .RST(rst), .Q(c[868]) );
  DFF \sreg_reg[868]  ( .D(c[868]), .CLK(clk), .RST(rst), .Q(c[867]) );
  DFF \sreg_reg[867]  ( .D(c[867]), .CLK(clk), .RST(rst), .Q(c[866]) );
  DFF \sreg_reg[866]  ( .D(c[866]), .CLK(clk), .RST(rst), .Q(c[865]) );
  DFF \sreg_reg[865]  ( .D(c[865]), .CLK(clk), .RST(rst), .Q(c[864]) );
  DFF \sreg_reg[864]  ( .D(c[864]), .CLK(clk), .RST(rst), .Q(c[863]) );
  DFF \sreg_reg[863]  ( .D(c[863]), .CLK(clk), .RST(rst), .Q(c[862]) );
  DFF \sreg_reg[862]  ( .D(c[862]), .CLK(clk), .RST(rst), .Q(c[861]) );
  DFF \sreg_reg[861]  ( .D(c[861]), .CLK(clk), .RST(rst), .Q(c[860]) );
  DFF \sreg_reg[860]  ( .D(c[860]), .CLK(clk), .RST(rst), .Q(c[859]) );
  DFF \sreg_reg[859]  ( .D(c[859]), .CLK(clk), .RST(rst), .Q(c[858]) );
  DFF \sreg_reg[858]  ( .D(c[858]), .CLK(clk), .RST(rst), .Q(c[857]) );
  DFF \sreg_reg[857]  ( .D(c[857]), .CLK(clk), .RST(rst), .Q(c[856]) );
  DFF \sreg_reg[856]  ( .D(c[856]), .CLK(clk), .RST(rst), .Q(c[855]) );
  DFF \sreg_reg[855]  ( .D(c[855]), .CLK(clk), .RST(rst), .Q(c[854]) );
  DFF \sreg_reg[854]  ( .D(c[854]), .CLK(clk), .RST(rst), .Q(c[853]) );
  DFF \sreg_reg[853]  ( .D(c[853]), .CLK(clk), .RST(rst), .Q(c[852]) );
  DFF \sreg_reg[852]  ( .D(c[852]), .CLK(clk), .RST(rst), .Q(c[851]) );
  DFF \sreg_reg[851]  ( .D(c[851]), .CLK(clk), .RST(rst), .Q(c[850]) );
  DFF \sreg_reg[850]  ( .D(c[850]), .CLK(clk), .RST(rst), .Q(c[849]) );
  DFF \sreg_reg[849]  ( .D(c[849]), .CLK(clk), .RST(rst), .Q(c[848]) );
  DFF \sreg_reg[848]  ( .D(c[848]), .CLK(clk), .RST(rst), .Q(c[847]) );
  DFF \sreg_reg[847]  ( .D(c[847]), .CLK(clk), .RST(rst), .Q(c[846]) );
  DFF \sreg_reg[846]  ( .D(c[846]), .CLK(clk), .RST(rst), .Q(c[845]) );
  DFF \sreg_reg[845]  ( .D(c[845]), .CLK(clk), .RST(rst), .Q(c[844]) );
  DFF \sreg_reg[844]  ( .D(c[844]), .CLK(clk), .RST(rst), .Q(c[843]) );
  DFF \sreg_reg[843]  ( .D(c[843]), .CLK(clk), .RST(rst), .Q(c[842]) );
  DFF \sreg_reg[842]  ( .D(c[842]), .CLK(clk), .RST(rst), .Q(c[841]) );
  DFF \sreg_reg[841]  ( .D(c[841]), .CLK(clk), .RST(rst), .Q(c[840]) );
  DFF \sreg_reg[840]  ( .D(c[840]), .CLK(clk), .RST(rst), .Q(c[839]) );
  DFF \sreg_reg[839]  ( .D(c[839]), .CLK(clk), .RST(rst), .Q(c[838]) );
  DFF \sreg_reg[838]  ( .D(c[838]), .CLK(clk), .RST(rst), .Q(c[837]) );
  DFF \sreg_reg[837]  ( .D(c[837]), .CLK(clk), .RST(rst), .Q(c[836]) );
  DFF \sreg_reg[836]  ( .D(c[836]), .CLK(clk), .RST(rst), .Q(c[835]) );
  DFF \sreg_reg[835]  ( .D(c[835]), .CLK(clk), .RST(rst), .Q(c[834]) );
  DFF \sreg_reg[834]  ( .D(c[834]), .CLK(clk), .RST(rst), .Q(c[833]) );
  DFF \sreg_reg[833]  ( .D(c[833]), .CLK(clk), .RST(rst), .Q(c[832]) );
  DFF \sreg_reg[832]  ( .D(c[832]), .CLK(clk), .RST(rst), .Q(c[831]) );
  DFF \sreg_reg[831]  ( .D(c[831]), .CLK(clk), .RST(rst), .Q(c[830]) );
  DFF \sreg_reg[830]  ( .D(c[830]), .CLK(clk), .RST(rst), .Q(c[829]) );
  DFF \sreg_reg[829]  ( .D(c[829]), .CLK(clk), .RST(rst), .Q(c[828]) );
  DFF \sreg_reg[828]  ( .D(c[828]), .CLK(clk), .RST(rst), .Q(c[827]) );
  DFF \sreg_reg[827]  ( .D(c[827]), .CLK(clk), .RST(rst), .Q(c[826]) );
  DFF \sreg_reg[826]  ( .D(c[826]), .CLK(clk), .RST(rst), .Q(c[825]) );
  DFF \sreg_reg[825]  ( .D(c[825]), .CLK(clk), .RST(rst), .Q(c[824]) );
  DFF \sreg_reg[824]  ( .D(c[824]), .CLK(clk), .RST(rst), .Q(c[823]) );
  DFF \sreg_reg[823]  ( .D(c[823]), .CLK(clk), .RST(rst), .Q(c[822]) );
  DFF \sreg_reg[822]  ( .D(c[822]), .CLK(clk), .RST(rst), .Q(c[821]) );
  DFF \sreg_reg[821]  ( .D(c[821]), .CLK(clk), .RST(rst), .Q(c[820]) );
  DFF \sreg_reg[820]  ( .D(c[820]), .CLK(clk), .RST(rst), .Q(c[819]) );
  DFF \sreg_reg[819]  ( .D(c[819]), .CLK(clk), .RST(rst), .Q(c[818]) );
  DFF \sreg_reg[818]  ( .D(c[818]), .CLK(clk), .RST(rst), .Q(c[817]) );
  DFF \sreg_reg[817]  ( .D(c[817]), .CLK(clk), .RST(rst), .Q(c[816]) );
  DFF \sreg_reg[816]  ( .D(c[816]), .CLK(clk), .RST(rst), .Q(c[815]) );
  DFF \sreg_reg[815]  ( .D(c[815]), .CLK(clk), .RST(rst), .Q(c[814]) );
  DFF \sreg_reg[814]  ( .D(c[814]), .CLK(clk), .RST(rst), .Q(c[813]) );
  DFF \sreg_reg[813]  ( .D(c[813]), .CLK(clk), .RST(rst), .Q(c[812]) );
  DFF \sreg_reg[812]  ( .D(c[812]), .CLK(clk), .RST(rst), .Q(c[811]) );
  DFF \sreg_reg[811]  ( .D(c[811]), .CLK(clk), .RST(rst), .Q(c[810]) );
  DFF \sreg_reg[810]  ( .D(c[810]), .CLK(clk), .RST(rst), .Q(c[809]) );
  DFF \sreg_reg[809]  ( .D(c[809]), .CLK(clk), .RST(rst), .Q(c[808]) );
  DFF \sreg_reg[808]  ( .D(c[808]), .CLK(clk), .RST(rst), .Q(c[807]) );
  DFF \sreg_reg[807]  ( .D(c[807]), .CLK(clk), .RST(rst), .Q(c[806]) );
  DFF \sreg_reg[806]  ( .D(c[806]), .CLK(clk), .RST(rst), .Q(c[805]) );
  DFF \sreg_reg[805]  ( .D(c[805]), .CLK(clk), .RST(rst), .Q(c[804]) );
  DFF \sreg_reg[804]  ( .D(c[804]), .CLK(clk), .RST(rst), .Q(c[803]) );
  DFF \sreg_reg[803]  ( .D(c[803]), .CLK(clk), .RST(rst), .Q(c[802]) );
  DFF \sreg_reg[802]  ( .D(c[802]), .CLK(clk), .RST(rst), .Q(c[801]) );
  DFF \sreg_reg[801]  ( .D(c[801]), .CLK(clk), .RST(rst), .Q(c[800]) );
  DFF \sreg_reg[800]  ( .D(c[800]), .CLK(clk), .RST(rst), .Q(c[799]) );
  DFF \sreg_reg[799]  ( .D(c[799]), .CLK(clk), .RST(rst), .Q(c[798]) );
  DFF \sreg_reg[798]  ( .D(c[798]), .CLK(clk), .RST(rst), .Q(c[797]) );
  DFF \sreg_reg[797]  ( .D(c[797]), .CLK(clk), .RST(rst), .Q(c[796]) );
  DFF \sreg_reg[796]  ( .D(c[796]), .CLK(clk), .RST(rst), .Q(c[795]) );
  DFF \sreg_reg[795]  ( .D(c[795]), .CLK(clk), .RST(rst), .Q(c[794]) );
  DFF \sreg_reg[794]  ( .D(c[794]), .CLK(clk), .RST(rst), .Q(c[793]) );
  DFF \sreg_reg[793]  ( .D(c[793]), .CLK(clk), .RST(rst), .Q(c[792]) );
  DFF \sreg_reg[792]  ( .D(c[792]), .CLK(clk), .RST(rst), .Q(c[791]) );
  DFF \sreg_reg[791]  ( .D(c[791]), .CLK(clk), .RST(rst), .Q(c[790]) );
  DFF \sreg_reg[790]  ( .D(c[790]), .CLK(clk), .RST(rst), .Q(c[789]) );
  DFF \sreg_reg[789]  ( .D(c[789]), .CLK(clk), .RST(rst), .Q(c[788]) );
  DFF \sreg_reg[788]  ( .D(c[788]), .CLK(clk), .RST(rst), .Q(c[787]) );
  DFF \sreg_reg[787]  ( .D(c[787]), .CLK(clk), .RST(rst), .Q(c[786]) );
  DFF \sreg_reg[786]  ( .D(c[786]), .CLK(clk), .RST(rst), .Q(c[785]) );
  DFF \sreg_reg[785]  ( .D(c[785]), .CLK(clk), .RST(rst), .Q(c[784]) );
  DFF \sreg_reg[784]  ( .D(c[784]), .CLK(clk), .RST(rst), .Q(c[783]) );
  DFF \sreg_reg[783]  ( .D(c[783]), .CLK(clk), .RST(rst), .Q(c[782]) );
  DFF \sreg_reg[782]  ( .D(c[782]), .CLK(clk), .RST(rst), .Q(c[781]) );
  DFF \sreg_reg[781]  ( .D(c[781]), .CLK(clk), .RST(rst), .Q(c[780]) );
  DFF \sreg_reg[780]  ( .D(c[780]), .CLK(clk), .RST(rst), .Q(c[779]) );
  DFF \sreg_reg[779]  ( .D(c[779]), .CLK(clk), .RST(rst), .Q(c[778]) );
  DFF \sreg_reg[778]  ( .D(c[778]), .CLK(clk), .RST(rst), .Q(c[777]) );
  DFF \sreg_reg[777]  ( .D(c[777]), .CLK(clk), .RST(rst), .Q(c[776]) );
  DFF \sreg_reg[776]  ( .D(c[776]), .CLK(clk), .RST(rst), .Q(c[775]) );
  DFF \sreg_reg[775]  ( .D(c[775]), .CLK(clk), .RST(rst), .Q(c[774]) );
  DFF \sreg_reg[774]  ( .D(c[774]), .CLK(clk), .RST(rst), .Q(c[773]) );
  DFF \sreg_reg[773]  ( .D(c[773]), .CLK(clk), .RST(rst), .Q(c[772]) );
  DFF \sreg_reg[772]  ( .D(c[772]), .CLK(clk), .RST(rst), .Q(c[771]) );
  DFF \sreg_reg[771]  ( .D(c[771]), .CLK(clk), .RST(rst), .Q(c[770]) );
  DFF \sreg_reg[770]  ( .D(c[770]), .CLK(clk), .RST(rst), .Q(c[769]) );
  DFF \sreg_reg[769]  ( .D(c[769]), .CLK(clk), .RST(rst), .Q(c[768]) );
  DFF \sreg_reg[768]  ( .D(c[768]), .CLK(clk), .RST(rst), .Q(c[767]) );
  DFF \sreg_reg[767]  ( .D(c[767]), .CLK(clk), .RST(rst), .Q(c[766]) );
  DFF \sreg_reg[766]  ( .D(c[766]), .CLK(clk), .RST(rst), .Q(c[765]) );
  DFF \sreg_reg[765]  ( .D(c[765]), .CLK(clk), .RST(rst), .Q(c[764]) );
  DFF \sreg_reg[764]  ( .D(c[764]), .CLK(clk), .RST(rst), .Q(c[763]) );
  DFF \sreg_reg[763]  ( .D(c[763]), .CLK(clk), .RST(rst), .Q(c[762]) );
  DFF \sreg_reg[762]  ( .D(c[762]), .CLK(clk), .RST(rst), .Q(c[761]) );
  DFF \sreg_reg[761]  ( .D(c[761]), .CLK(clk), .RST(rst), .Q(c[760]) );
  DFF \sreg_reg[760]  ( .D(c[760]), .CLK(clk), .RST(rst), .Q(c[759]) );
  DFF \sreg_reg[759]  ( .D(c[759]), .CLK(clk), .RST(rst), .Q(c[758]) );
  DFF \sreg_reg[758]  ( .D(c[758]), .CLK(clk), .RST(rst), .Q(c[757]) );
  DFF \sreg_reg[757]  ( .D(c[757]), .CLK(clk), .RST(rst), .Q(c[756]) );
  DFF \sreg_reg[756]  ( .D(c[756]), .CLK(clk), .RST(rst), .Q(c[755]) );
  DFF \sreg_reg[755]  ( .D(c[755]), .CLK(clk), .RST(rst), .Q(c[754]) );
  DFF \sreg_reg[754]  ( .D(c[754]), .CLK(clk), .RST(rst), .Q(c[753]) );
  DFF \sreg_reg[753]  ( .D(c[753]), .CLK(clk), .RST(rst), .Q(c[752]) );
  DFF \sreg_reg[752]  ( .D(c[752]), .CLK(clk), .RST(rst), .Q(c[751]) );
  DFF \sreg_reg[751]  ( .D(c[751]), .CLK(clk), .RST(rst), .Q(c[750]) );
  DFF \sreg_reg[750]  ( .D(c[750]), .CLK(clk), .RST(rst), .Q(c[749]) );
  DFF \sreg_reg[749]  ( .D(c[749]), .CLK(clk), .RST(rst), .Q(c[748]) );
  DFF \sreg_reg[748]  ( .D(c[748]), .CLK(clk), .RST(rst), .Q(c[747]) );
  DFF \sreg_reg[747]  ( .D(c[747]), .CLK(clk), .RST(rst), .Q(c[746]) );
  DFF \sreg_reg[746]  ( .D(c[746]), .CLK(clk), .RST(rst), .Q(c[745]) );
  DFF \sreg_reg[745]  ( .D(c[745]), .CLK(clk), .RST(rst), .Q(c[744]) );
  DFF \sreg_reg[744]  ( .D(c[744]), .CLK(clk), .RST(rst), .Q(c[743]) );
  DFF \sreg_reg[743]  ( .D(c[743]), .CLK(clk), .RST(rst), .Q(c[742]) );
  DFF \sreg_reg[742]  ( .D(c[742]), .CLK(clk), .RST(rst), .Q(c[741]) );
  DFF \sreg_reg[741]  ( .D(c[741]), .CLK(clk), .RST(rst), .Q(c[740]) );
  DFF \sreg_reg[740]  ( .D(c[740]), .CLK(clk), .RST(rst), .Q(c[739]) );
  DFF \sreg_reg[739]  ( .D(c[739]), .CLK(clk), .RST(rst), .Q(c[738]) );
  DFF \sreg_reg[738]  ( .D(c[738]), .CLK(clk), .RST(rst), .Q(c[737]) );
  DFF \sreg_reg[737]  ( .D(c[737]), .CLK(clk), .RST(rst), .Q(c[736]) );
  DFF \sreg_reg[736]  ( .D(c[736]), .CLK(clk), .RST(rst), .Q(c[735]) );
  DFF \sreg_reg[735]  ( .D(c[735]), .CLK(clk), .RST(rst), .Q(c[734]) );
  DFF \sreg_reg[734]  ( .D(c[734]), .CLK(clk), .RST(rst), .Q(c[733]) );
  DFF \sreg_reg[733]  ( .D(c[733]), .CLK(clk), .RST(rst), .Q(c[732]) );
  DFF \sreg_reg[732]  ( .D(c[732]), .CLK(clk), .RST(rst), .Q(c[731]) );
  DFF \sreg_reg[731]  ( .D(c[731]), .CLK(clk), .RST(rst), .Q(c[730]) );
  DFF \sreg_reg[730]  ( .D(c[730]), .CLK(clk), .RST(rst), .Q(c[729]) );
  DFF \sreg_reg[729]  ( .D(c[729]), .CLK(clk), .RST(rst), .Q(c[728]) );
  DFF \sreg_reg[728]  ( .D(c[728]), .CLK(clk), .RST(rst), .Q(c[727]) );
  DFF \sreg_reg[727]  ( .D(c[727]), .CLK(clk), .RST(rst), .Q(c[726]) );
  DFF \sreg_reg[726]  ( .D(c[726]), .CLK(clk), .RST(rst), .Q(c[725]) );
  DFF \sreg_reg[725]  ( .D(c[725]), .CLK(clk), .RST(rst), .Q(c[724]) );
  DFF \sreg_reg[724]  ( .D(c[724]), .CLK(clk), .RST(rst), .Q(c[723]) );
  DFF \sreg_reg[723]  ( .D(c[723]), .CLK(clk), .RST(rst), .Q(c[722]) );
  DFF \sreg_reg[722]  ( .D(c[722]), .CLK(clk), .RST(rst), .Q(c[721]) );
  DFF \sreg_reg[721]  ( .D(c[721]), .CLK(clk), .RST(rst), .Q(c[720]) );
  DFF \sreg_reg[720]  ( .D(c[720]), .CLK(clk), .RST(rst), .Q(c[719]) );
  DFF \sreg_reg[719]  ( .D(c[719]), .CLK(clk), .RST(rst), .Q(c[718]) );
  DFF \sreg_reg[718]  ( .D(c[718]), .CLK(clk), .RST(rst), .Q(c[717]) );
  DFF \sreg_reg[717]  ( .D(c[717]), .CLK(clk), .RST(rst), .Q(c[716]) );
  DFF \sreg_reg[716]  ( .D(c[716]), .CLK(clk), .RST(rst), .Q(c[715]) );
  DFF \sreg_reg[715]  ( .D(c[715]), .CLK(clk), .RST(rst), .Q(c[714]) );
  DFF \sreg_reg[714]  ( .D(c[714]), .CLK(clk), .RST(rst), .Q(c[713]) );
  DFF \sreg_reg[713]  ( .D(c[713]), .CLK(clk), .RST(rst), .Q(c[712]) );
  DFF \sreg_reg[712]  ( .D(c[712]), .CLK(clk), .RST(rst), .Q(c[711]) );
  DFF \sreg_reg[711]  ( .D(c[711]), .CLK(clk), .RST(rst), .Q(c[710]) );
  DFF \sreg_reg[710]  ( .D(c[710]), .CLK(clk), .RST(rst), .Q(c[709]) );
  DFF \sreg_reg[709]  ( .D(c[709]), .CLK(clk), .RST(rst), .Q(c[708]) );
  DFF \sreg_reg[708]  ( .D(c[708]), .CLK(clk), .RST(rst), .Q(c[707]) );
  DFF \sreg_reg[707]  ( .D(c[707]), .CLK(clk), .RST(rst), .Q(c[706]) );
  DFF \sreg_reg[706]  ( .D(c[706]), .CLK(clk), .RST(rst), .Q(c[705]) );
  DFF \sreg_reg[705]  ( .D(c[705]), .CLK(clk), .RST(rst), .Q(c[704]) );
  DFF \sreg_reg[704]  ( .D(c[704]), .CLK(clk), .RST(rst), .Q(c[703]) );
  DFF \sreg_reg[703]  ( .D(c[703]), .CLK(clk), .RST(rst), .Q(c[702]) );
  DFF \sreg_reg[702]  ( .D(c[702]), .CLK(clk), .RST(rst), .Q(c[701]) );
  DFF \sreg_reg[701]  ( .D(c[701]), .CLK(clk), .RST(rst), .Q(c[700]) );
  DFF \sreg_reg[700]  ( .D(c[700]), .CLK(clk), .RST(rst), .Q(c[699]) );
  DFF \sreg_reg[699]  ( .D(c[699]), .CLK(clk), .RST(rst), .Q(c[698]) );
  DFF \sreg_reg[698]  ( .D(c[698]), .CLK(clk), .RST(rst), .Q(c[697]) );
  DFF \sreg_reg[697]  ( .D(c[697]), .CLK(clk), .RST(rst), .Q(c[696]) );
  DFF \sreg_reg[696]  ( .D(c[696]), .CLK(clk), .RST(rst), .Q(c[695]) );
  DFF \sreg_reg[695]  ( .D(c[695]), .CLK(clk), .RST(rst), .Q(c[694]) );
  DFF \sreg_reg[694]  ( .D(c[694]), .CLK(clk), .RST(rst), .Q(c[693]) );
  DFF \sreg_reg[693]  ( .D(c[693]), .CLK(clk), .RST(rst), .Q(c[692]) );
  DFF \sreg_reg[692]  ( .D(c[692]), .CLK(clk), .RST(rst), .Q(c[691]) );
  DFF \sreg_reg[691]  ( .D(c[691]), .CLK(clk), .RST(rst), .Q(c[690]) );
  DFF \sreg_reg[690]  ( .D(c[690]), .CLK(clk), .RST(rst), .Q(c[689]) );
  DFF \sreg_reg[689]  ( .D(c[689]), .CLK(clk), .RST(rst), .Q(c[688]) );
  DFF \sreg_reg[688]  ( .D(c[688]), .CLK(clk), .RST(rst), .Q(c[687]) );
  DFF \sreg_reg[687]  ( .D(c[687]), .CLK(clk), .RST(rst), .Q(c[686]) );
  DFF \sreg_reg[686]  ( .D(c[686]), .CLK(clk), .RST(rst), .Q(c[685]) );
  DFF \sreg_reg[685]  ( .D(c[685]), .CLK(clk), .RST(rst), .Q(c[684]) );
  DFF \sreg_reg[684]  ( .D(c[684]), .CLK(clk), .RST(rst), .Q(c[683]) );
  DFF \sreg_reg[683]  ( .D(c[683]), .CLK(clk), .RST(rst), .Q(c[682]) );
  DFF \sreg_reg[682]  ( .D(c[682]), .CLK(clk), .RST(rst), .Q(c[681]) );
  DFF \sreg_reg[681]  ( .D(c[681]), .CLK(clk), .RST(rst), .Q(c[680]) );
  DFF \sreg_reg[680]  ( .D(c[680]), .CLK(clk), .RST(rst), .Q(c[679]) );
  DFF \sreg_reg[679]  ( .D(c[679]), .CLK(clk), .RST(rst), .Q(c[678]) );
  DFF \sreg_reg[678]  ( .D(c[678]), .CLK(clk), .RST(rst), .Q(c[677]) );
  DFF \sreg_reg[677]  ( .D(c[677]), .CLK(clk), .RST(rst), .Q(c[676]) );
  DFF \sreg_reg[676]  ( .D(c[676]), .CLK(clk), .RST(rst), .Q(c[675]) );
  DFF \sreg_reg[675]  ( .D(c[675]), .CLK(clk), .RST(rst), .Q(c[674]) );
  DFF \sreg_reg[674]  ( .D(c[674]), .CLK(clk), .RST(rst), .Q(c[673]) );
  DFF \sreg_reg[673]  ( .D(c[673]), .CLK(clk), .RST(rst), .Q(c[672]) );
  DFF \sreg_reg[672]  ( .D(c[672]), .CLK(clk), .RST(rst), .Q(c[671]) );
  DFF \sreg_reg[671]  ( .D(c[671]), .CLK(clk), .RST(rst), .Q(c[670]) );
  DFF \sreg_reg[670]  ( .D(c[670]), .CLK(clk), .RST(rst), .Q(c[669]) );
  DFF \sreg_reg[669]  ( .D(c[669]), .CLK(clk), .RST(rst), .Q(c[668]) );
  DFF \sreg_reg[668]  ( .D(c[668]), .CLK(clk), .RST(rst), .Q(c[667]) );
  DFF \sreg_reg[667]  ( .D(c[667]), .CLK(clk), .RST(rst), .Q(c[666]) );
  DFF \sreg_reg[666]  ( .D(c[666]), .CLK(clk), .RST(rst), .Q(c[665]) );
  DFF \sreg_reg[665]  ( .D(c[665]), .CLK(clk), .RST(rst), .Q(c[664]) );
  DFF \sreg_reg[664]  ( .D(c[664]), .CLK(clk), .RST(rst), .Q(c[663]) );
  DFF \sreg_reg[663]  ( .D(c[663]), .CLK(clk), .RST(rst), .Q(c[662]) );
  DFF \sreg_reg[662]  ( .D(c[662]), .CLK(clk), .RST(rst), .Q(c[661]) );
  DFF \sreg_reg[661]  ( .D(c[661]), .CLK(clk), .RST(rst), .Q(c[660]) );
  DFF \sreg_reg[660]  ( .D(c[660]), .CLK(clk), .RST(rst), .Q(c[659]) );
  DFF \sreg_reg[659]  ( .D(c[659]), .CLK(clk), .RST(rst), .Q(c[658]) );
  DFF \sreg_reg[658]  ( .D(c[658]), .CLK(clk), .RST(rst), .Q(c[657]) );
  DFF \sreg_reg[657]  ( .D(c[657]), .CLK(clk), .RST(rst), .Q(c[656]) );
  DFF \sreg_reg[656]  ( .D(c[656]), .CLK(clk), .RST(rst), .Q(c[655]) );
  DFF \sreg_reg[655]  ( .D(c[655]), .CLK(clk), .RST(rst), .Q(c[654]) );
  DFF \sreg_reg[654]  ( .D(c[654]), .CLK(clk), .RST(rst), .Q(c[653]) );
  DFF \sreg_reg[653]  ( .D(c[653]), .CLK(clk), .RST(rst), .Q(c[652]) );
  DFF \sreg_reg[652]  ( .D(c[652]), .CLK(clk), .RST(rst), .Q(c[651]) );
  DFF \sreg_reg[651]  ( .D(c[651]), .CLK(clk), .RST(rst), .Q(c[650]) );
  DFF \sreg_reg[650]  ( .D(c[650]), .CLK(clk), .RST(rst), .Q(c[649]) );
  DFF \sreg_reg[649]  ( .D(c[649]), .CLK(clk), .RST(rst), .Q(c[648]) );
  DFF \sreg_reg[648]  ( .D(c[648]), .CLK(clk), .RST(rst), .Q(c[647]) );
  DFF \sreg_reg[647]  ( .D(c[647]), .CLK(clk), .RST(rst), .Q(c[646]) );
  DFF \sreg_reg[646]  ( .D(c[646]), .CLK(clk), .RST(rst), .Q(c[645]) );
  DFF \sreg_reg[645]  ( .D(c[645]), .CLK(clk), .RST(rst), .Q(c[644]) );
  DFF \sreg_reg[644]  ( .D(c[644]), .CLK(clk), .RST(rst), .Q(c[643]) );
  DFF \sreg_reg[643]  ( .D(c[643]), .CLK(clk), .RST(rst), .Q(c[642]) );
  DFF \sreg_reg[642]  ( .D(c[642]), .CLK(clk), .RST(rst), .Q(c[641]) );
  DFF \sreg_reg[641]  ( .D(c[641]), .CLK(clk), .RST(rst), .Q(c[640]) );
  DFF \sreg_reg[640]  ( .D(c[640]), .CLK(clk), .RST(rst), .Q(c[639]) );
  DFF \sreg_reg[639]  ( .D(c[639]), .CLK(clk), .RST(rst), .Q(c[638]) );
  DFF \sreg_reg[638]  ( .D(c[638]), .CLK(clk), .RST(rst), .Q(c[637]) );
  DFF \sreg_reg[637]  ( .D(c[637]), .CLK(clk), .RST(rst), .Q(c[636]) );
  DFF \sreg_reg[636]  ( .D(c[636]), .CLK(clk), .RST(rst), .Q(c[635]) );
  DFF \sreg_reg[635]  ( .D(c[635]), .CLK(clk), .RST(rst), .Q(c[634]) );
  DFF \sreg_reg[634]  ( .D(c[634]), .CLK(clk), .RST(rst), .Q(c[633]) );
  DFF \sreg_reg[633]  ( .D(c[633]), .CLK(clk), .RST(rst), .Q(c[632]) );
  DFF \sreg_reg[632]  ( .D(c[632]), .CLK(clk), .RST(rst), .Q(c[631]) );
  DFF \sreg_reg[631]  ( .D(c[631]), .CLK(clk), .RST(rst), .Q(c[630]) );
  DFF \sreg_reg[630]  ( .D(c[630]), .CLK(clk), .RST(rst), .Q(c[629]) );
  DFF \sreg_reg[629]  ( .D(c[629]), .CLK(clk), .RST(rst), .Q(c[628]) );
  DFF \sreg_reg[628]  ( .D(c[628]), .CLK(clk), .RST(rst), .Q(c[627]) );
  DFF \sreg_reg[627]  ( .D(c[627]), .CLK(clk), .RST(rst), .Q(c[626]) );
  DFF \sreg_reg[626]  ( .D(c[626]), .CLK(clk), .RST(rst), .Q(c[625]) );
  DFF \sreg_reg[625]  ( .D(c[625]), .CLK(clk), .RST(rst), .Q(c[624]) );
  DFF \sreg_reg[624]  ( .D(c[624]), .CLK(clk), .RST(rst), .Q(c[623]) );
  DFF \sreg_reg[623]  ( .D(c[623]), .CLK(clk), .RST(rst), .Q(c[622]) );
  DFF \sreg_reg[622]  ( .D(c[622]), .CLK(clk), .RST(rst), .Q(c[621]) );
  DFF \sreg_reg[621]  ( .D(c[621]), .CLK(clk), .RST(rst), .Q(c[620]) );
  DFF \sreg_reg[620]  ( .D(c[620]), .CLK(clk), .RST(rst), .Q(c[619]) );
  DFF \sreg_reg[619]  ( .D(c[619]), .CLK(clk), .RST(rst), .Q(c[618]) );
  DFF \sreg_reg[618]  ( .D(c[618]), .CLK(clk), .RST(rst), .Q(c[617]) );
  DFF \sreg_reg[617]  ( .D(c[617]), .CLK(clk), .RST(rst), .Q(c[616]) );
  DFF \sreg_reg[616]  ( .D(c[616]), .CLK(clk), .RST(rst), .Q(c[615]) );
  DFF \sreg_reg[615]  ( .D(c[615]), .CLK(clk), .RST(rst), .Q(c[614]) );
  DFF \sreg_reg[614]  ( .D(c[614]), .CLK(clk), .RST(rst), .Q(c[613]) );
  DFF \sreg_reg[613]  ( .D(c[613]), .CLK(clk), .RST(rst), .Q(c[612]) );
  DFF \sreg_reg[612]  ( .D(c[612]), .CLK(clk), .RST(rst), .Q(c[611]) );
  DFF \sreg_reg[611]  ( .D(c[611]), .CLK(clk), .RST(rst), .Q(c[610]) );
  DFF \sreg_reg[610]  ( .D(c[610]), .CLK(clk), .RST(rst), .Q(c[609]) );
  DFF \sreg_reg[609]  ( .D(c[609]), .CLK(clk), .RST(rst), .Q(c[608]) );
  DFF \sreg_reg[608]  ( .D(c[608]), .CLK(clk), .RST(rst), .Q(c[607]) );
  DFF \sreg_reg[607]  ( .D(c[607]), .CLK(clk), .RST(rst), .Q(c[606]) );
  DFF \sreg_reg[606]  ( .D(c[606]), .CLK(clk), .RST(rst), .Q(c[605]) );
  DFF \sreg_reg[605]  ( .D(c[605]), .CLK(clk), .RST(rst), .Q(c[604]) );
  DFF \sreg_reg[604]  ( .D(c[604]), .CLK(clk), .RST(rst), .Q(c[603]) );
  DFF \sreg_reg[603]  ( .D(c[603]), .CLK(clk), .RST(rst), .Q(c[602]) );
  DFF \sreg_reg[602]  ( .D(c[602]), .CLK(clk), .RST(rst), .Q(c[601]) );
  DFF \sreg_reg[601]  ( .D(c[601]), .CLK(clk), .RST(rst), .Q(c[600]) );
  DFF \sreg_reg[600]  ( .D(c[600]), .CLK(clk), .RST(rst), .Q(c[599]) );
  DFF \sreg_reg[599]  ( .D(c[599]), .CLK(clk), .RST(rst), .Q(c[598]) );
  DFF \sreg_reg[598]  ( .D(c[598]), .CLK(clk), .RST(rst), .Q(c[597]) );
  DFF \sreg_reg[597]  ( .D(c[597]), .CLK(clk), .RST(rst), .Q(c[596]) );
  DFF \sreg_reg[596]  ( .D(c[596]), .CLK(clk), .RST(rst), .Q(c[595]) );
  DFF \sreg_reg[595]  ( .D(c[595]), .CLK(clk), .RST(rst), .Q(c[594]) );
  DFF \sreg_reg[594]  ( .D(c[594]), .CLK(clk), .RST(rst), .Q(c[593]) );
  DFF \sreg_reg[593]  ( .D(c[593]), .CLK(clk), .RST(rst), .Q(c[592]) );
  DFF \sreg_reg[592]  ( .D(c[592]), .CLK(clk), .RST(rst), .Q(c[591]) );
  DFF \sreg_reg[591]  ( .D(c[591]), .CLK(clk), .RST(rst), .Q(c[590]) );
  DFF \sreg_reg[590]  ( .D(c[590]), .CLK(clk), .RST(rst), .Q(c[589]) );
  DFF \sreg_reg[589]  ( .D(c[589]), .CLK(clk), .RST(rst), .Q(c[588]) );
  DFF \sreg_reg[588]  ( .D(c[588]), .CLK(clk), .RST(rst), .Q(c[587]) );
  DFF \sreg_reg[587]  ( .D(c[587]), .CLK(clk), .RST(rst), .Q(c[586]) );
  DFF \sreg_reg[586]  ( .D(c[586]), .CLK(clk), .RST(rst), .Q(c[585]) );
  DFF \sreg_reg[585]  ( .D(c[585]), .CLK(clk), .RST(rst), .Q(c[584]) );
  DFF \sreg_reg[584]  ( .D(c[584]), .CLK(clk), .RST(rst), .Q(c[583]) );
  DFF \sreg_reg[583]  ( .D(c[583]), .CLK(clk), .RST(rst), .Q(c[582]) );
  DFF \sreg_reg[582]  ( .D(c[582]), .CLK(clk), .RST(rst), .Q(c[581]) );
  DFF \sreg_reg[581]  ( .D(c[581]), .CLK(clk), .RST(rst), .Q(c[580]) );
  DFF \sreg_reg[580]  ( .D(c[580]), .CLK(clk), .RST(rst), .Q(c[579]) );
  DFF \sreg_reg[579]  ( .D(c[579]), .CLK(clk), .RST(rst), .Q(c[578]) );
  DFF \sreg_reg[578]  ( .D(c[578]), .CLK(clk), .RST(rst), .Q(c[577]) );
  DFF \sreg_reg[577]  ( .D(c[577]), .CLK(clk), .RST(rst), .Q(c[576]) );
  DFF \sreg_reg[576]  ( .D(c[576]), .CLK(clk), .RST(rst), .Q(c[575]) );
  DFF \sreg_reg[575]  ( .D(c[575]), .CLK(clk), .RST(rst), .Q(c[574]) );
  DFF \sreg_reg[574]  ( .D(c[574]), .CLK(clk), .RST(rst), .Q(c[573]) );
  DFF \sreg_reg[573]  ( .D(c[573]), .CLK(clk), .RST(rst), .Q(c[572]) );
  DFF \sreg_reg[572]  ( .D(c[572]), .CLK(clk), .RST(rst), .Q(c[571]) );
  DFF \sreg_reg[571]  ( .D(c[571]), .CLK(clk), .RST(rst), .Q(c[570]) );
  DFF \sreg_reg[570]  ( .D(c[570]), .CLK(clk), .RST(rst), .Q(c[569]) );
  DFF \sreg_reg[569]  ( .D(c[569]), .CLK(clk), .RST(rst), .Q(c[568]) );
  DFF \sreg_reg[568]  ( .D(c[568]), .CLK(clk), .RST(rst), .Q(c[567]) );
  DFF \sreg_reg[567]  ( .D(c[567]), .CLK(clk), .RST(rst), .Q(c[566]) );
  DFF \sreg_reg[566]  ( .D(c[566]), .CLK(clk), .RST(rst), .Q(c[565]) );
  DFF \sreg_reg[565]  ( .D(c[565]), .CLK(clk), .RST(rst), .Q(c[564]) );
  DFF \sreg_reg[564]  ( .D(c[564]), .CLK(clk), .RST(rst), .Q(c[563]) );
  DFF \sreg_reg[563]  ( .D(c[563]), .CLK(clk), .RST(rst), .Q(c[562]) );
  DFF \sreg_reg[562]  ( .D(c[562]), .CLK(clk), .RST(rst), .Q(c[561]) );
  DFF \sreg_reg[561]  ( .D(c[561]), .CLK(clk), .RST(rst), .Q(c[560]) );
  DFF \sreg_reg[560]  ( .D(c[560]), .CLK(clk), .RST(rst), .Q(c[559]) );
  DFF \sreg_reg[559]  ( .D(c[559]), .CLK(clk), .RST(rst), .Q(c[558]) );
  DFF \sreg_reg[558]  ( .D(c[558]), .CLK(clk), .RST(rst), .Q(c[557]) );
  DFF \sreg_reg[557]  ( .D(c[557]), .CLK(clk), .RST(rst), .Q(c[556]) );
  DFF \sreg_reg[556]  ( .D(c[556]), .CLK(clk), .RST(rst), .Q(c[555]) );
  DFF \sreg_reg[555]  ( .D(c[555]), .CLK(clk), .RST(rst), .Q(c[554]) );
  DFF \sreg_reg[554]  ( .D(c[554]), .CLK(clk), .RST(rst), .Q(c[553]) );
  DFF \sreg_reg[553]  ( .D(c[553]), .CLK(clk), .RST(rst), .Q(c[552]) );
  DFF \sreg_reg[552]  ( .D(c[552]), .CLK(clk), .RST(rst), .Q(c[551]) );
  DFF \sreg_reg[551]  ( .D(c[551]), .CLK(clk), .RST(rst), .Q(c[550]) );
  DFF \sreg_reg[550]  ( .D(c[550]), .CLK(clk), .RST(rst), .Q(c[549]) );
  DFF \sreg_reg[549]  ( .D(c[549]), .CLK(clk), .RST(rst), .Q(c[548]) );
  DFF \sreg_reg[548]  ( .D(c[548]), .CLK(clk), .RST(rst), .Q(c[547]) );
  DFF \sreg_reg[547]  ( .D(c[547]), .CLK(clk), .RST(rst), .Q(c[546]) );
  DFF \sreg_reg[546]  ( .D(c[546]), .CLK(clk), .RST(rst), .Q(c[545]) );
  DFF \sreg_reg[545]  ( .D(c[545]), .CLK(clk), .RST(rst), .Q(c[544]) );
  DFF \sreg_reg[544]  ( .D(c[544]), .CLK(clk), .RST(rst), .Q(c[543]) );
  DFF \sreg_reg[543]  ( .D(c[543]), .CLK(clk), .RST(rst), .Q(c[542]) );
  DFF \sreg_reg[542]  ( .D(c[542]), .CLK(clk), .RST(rst), .Q(c[541]) );
  DFF \sreg_reg[541]  ( .D(c[541]), .CLK(clk), .RST(rst), .Q(c[540]) );
  DFF \sreg_reg[540]  ( .D(c[540]), .CLK(clk), .RST(rst), .Q(c[539]) );
  DFF \sreg_reg[539]  ( .D(c[539]), .CLK(clk), .RST(rst), .Q(c[538]) );
  DFF \sreg_reg[538]  ( .D(c[538]), .CLK(clk), .RST(rst), .Q(c[537]) );
  DFF \sreg_reg[537]  ( .D(c[537]), .CLK(clk), .RST(rst), .Q(c[536]) );
  DFF \sreg_reg[536]  ( .D(c[536]), .CLK(clk), .RST(rst), .Q(c[535]) );
  DFF \sreg_reg[535]  ( .D(c[535]), .CLK(clk), .RST(rst), .Q(c[534]) );
  DFF \sreg_reg[534]  ( .D(c[534]), .CLK(clk), .RST(rst), .Q(c[533]) );
  DFF \sreg_reg[533]  ( .D(c[533]), .CLK(clk), .RST(rst), .Q(c[532]) );
  DFF \sreg_reg[532]  ( .D(c[532]), .CLK(clk), .RST(rst), .Q(c[531]) );
  DFF \sreg_reg[531]  ( .D(c[531]), .CLK(clk), .RST(rst), .Q(c[530]) );
  DFF \sreg_reg[530]  ( .D(c[530]), .CLK(clk), .RST(rst), .Q(c[529]) );
  DFF \sreg_reg[529]  ( .D(c[529]), .CLK(clk), .RST(rst), .Q(c[528]) );
  DFF \sreg_reg[528]  ( .D(c[528]), .CLK(clk), .RST(rst), .Q(c[527]) );
  DFF \sreg_reg[527]  ( .D(c[527]), .CLK(clk), .RST(rst), .Q(c[526]) );
  DFF \sreg_reg[526]  ( .D(c[526]), .CLK(clk), .RST(rst), .Q(c[525]) );
  DFF \sreg_reg[525]  ( .D(c[525]), .CLK(clk), .RST(rst), .Q(c[524]) );
  DFF \sreg_reg[524]  ( .D(c[524]), .CLK(clk), .RST(rst), .Q(c[523]) );
  DFF \sreg_reg[523]  ( .D(c[523]), .CLK(clk), .RST(rst), .Q(c[522]) );
  DFF \sreg_reg[522]  ( .D(c[522]), .CLK(clk), .RST(rst), .Q(c[521]) );
  DFF \sreg_reg[521]  ( .D(c[521]), .CLK(clk), .RST(rst), .Q(c[520]) );
  DFF \sreg_reg[520]  ( .D(c[520]), .CLK(clk), .RST(rst), .Q(c[519]) );
  DFF \sreg_reg[519]  ( .D(c[519]), .CLK(clk), .RST(rst), .Q(c[518]) );
  DFF \sreg_reg[518]  ( .D(c[518]), .CLK(clk), .RST(rst), .Q(c[517]) );
  DFF \sreg_reg[517]  ( .D(c[517]), .CLK(clk), .RST(rst), .Q(c[516]) );
  DFF \sreg_reg[516]  ( .D(c[516]), .CLK(clk), .RST(rst), .Q(c[515]) );
  DFF \sreg_reg[515]  ( .D(c[515]), .CLK(clk), .RST(rst), .Q(c[514]) );
  DFF \sreg_reg[514]  ( .D(c[514]), .CLK(clk), .RST(rst), .Q(c[513]) );
  DFF \sreg_reg[513]  ( .D(c[513]), .CLK(clk), .RST(rst), .Q(c[512]) );
  DFF \sreg_reg[512]  ( .D(c[512]), .CLK(clk), .RST(rst), .Q(c[511]) );
  DFF \sreg_reg[511]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(c[510]) );
  DFF \sreg_reg[510]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(c[509]) );
  DFF \sreg_reg[509]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(c[508]) );
  DFF \sreg_reg[508]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(c[507]) );
  DFF \sreg_reg[507]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(c[506]) );
  DFF \sreg_reg[506]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(c[505]) );
  DFF \sreg_reg[505]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(c[504]) );
  DFF \sreg_reg[504]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(c[503]) );
  DFF \sreg_reg[503]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(c[502]) );
  DFF \sreg_reg[502]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(c[501]) );
  DFF \sreg_reg[501]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(c[500]) );
  DFF \sreg_reg[500]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(c[499]) );
  DFF \sreg_reg[499]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(c[498]) );
  DFF \sreg_reg[498]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(c[497]) );
  DFF \sreg_reg[497]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(c[496]) );
  DFF \sreg_reg[496]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(c[495]) );
  DFF \sreg_reg[495]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(c[494]) );
  DFF \sreg_reg[494]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(c[493]) );
  DFF \sreg_reg[493]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(c[492]) );
  DFF \sreg_reg[492]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(c[491]) );
  DFF \sreg_reg[491]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(c[490]) );
  DFF \sreg_reg[490]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(c[489]) );
  DFF \sreg_reg[489]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(c[488]) );
  DFF \sreg_reg[488]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(c[487]) );
  DFF \sreg_reg[487]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(c[486]) );
  DFF \sreg_reg[486]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(c[485]) );
  DFF \sreg_reg[485]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(c[484]) );
  DFF \sreg_reg[484]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(c[483]) );
  DFF \sreg_reg[483]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(c[482]) );
  DFF \sreg_reg[482]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(c[481]) );
  DFF \sreg_reg[481]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(c[480]) );
  DFF \sreg_reg[480]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(c[479]) );
  DFF \sreg_reg[479]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(c[478]) );
  DFF \sreg_reg[478]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(c[477]) );
  DFF \sreg_reg[477]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(c[476]) );
  DFF \sreg_reg[476]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(c[475]) );
  DFF \sreg_reg[475]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(c[474]) );
  DFF \sreg_reg[474]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(c[473]) );
  DFF \sreg_reg[473]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(c[472]) );
  DFF \sreg_reg[472]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(c[471]) );
  DFF \sreg_reg[471]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(c[470]) );
  DFF \sreg_reg[470]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(c[469]) );
  DFF \sreg_reg[469]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(c[468]) );
  DFF \sreg_reg[468]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(c[467]) );
  DFF \sreg_reg[467]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(c[466]) );
  DFF \sreg_reg[466]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(c[465]) );
  DFF \sreg_reg[465]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(c[464]) );
  DFF \sreg_reg[464]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(c[463]) );
  DFF \sreg_reg[463]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(c[462]) );
  DFF \sreg_reg[462]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(c[461]) );
  DFF \sreg_reg[461]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(c[460]) );
  DFF \sreg_reg[460]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(c[459]) );
  DFF \sreg_reg[459]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(c[458]) );
  DFF \sreg_reg[458]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(c[457]) );
  DFF \sreg_reg[457]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(c[456]) );
  DFF \sreg_reg[456]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(c[455]) );
  DFF \sreg_reg[455]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(c[454]) );
  DFF \sreg_reg[454]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(c[453]) );
  DFF \sreg_reg[453]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(c[452]) );
  DFF \sreg_reg[452]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(c[451]) );
  DFF \sreg_reg[451]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(c[450]) );
  DFF \sreg_reg[450]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(c[449]) );
  DFF \sreg_reg[449]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(c[448]) );
  DFF \sreg_reg[448]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(c[447]) );
  DFF \sreg_reg[447]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(c[446]) );
  DFF \sreg_reg[446]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(c[445]) );
  DFF \sreg_reg[445]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(c[444]) );
  DFF \sreg_reg[444]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(c[443]) );
  DFF \sreg_reg[443]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(c[442]) );
  DFF \sreg_reg[442]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(c[441]) );
  DFF \sreg_reg[441]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(c[440]) );
  DFF \sreg_reg[440]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(c[439]) );
  DFF \sreg_reg[439]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(c[438]) );
  DFF \sreg_reg[438]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(c[437]) );
  DFF \sreg_reg[437]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(c[436]) );
  DFF \sreg_reg[436]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(c[435]) );
  DFF \sreg_reg[435]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(c[434]) );
  DFF \sreg_reg[434]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(c[433]) );
  DFF \sreg_reg[433]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(c[432]) );
  DFF \sreg_reg[432]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(c[431]) );
  DFF \sreg_reg[431]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(c[430]) );
  DFF \sreg_reg[430]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(c[429]) );
  DFF \sreg_reg[429]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(c[428]) );
  DFF \sreg_reg[428]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(c[427]) );
  DFF \sreg_reg[427]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(c[426]) );
  DFF \sreg_reg[426]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(c[425]) );
  DFF \sreg_reg[425]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(c[424]) );
  DFF \sreg_reg[424]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(c[423]) );
  DFF \sreg_reg[423]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(c[422]) );
  DFF \sreg_reg[422]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(c[421]) );
  DFF \sreg_reg[421]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(c[420]) );
  DFF \sreg_reg[420]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(c[419]) );
  DFF \sreg_reg[419]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(c[418]) );
  DFF \sreg_reg[418]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(c[417]) );
  DFF \sreg_reg[417]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(c[416]) );
  DFF \sreg_reg[416]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(c[415]) );
  DFF \sreg_reg[415]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(c[414]) );
  DFF \sreg_reg[414]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(c[413]) );
  DFF \sreg_reg[413]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(c[412]) );
  DFF \sreg_reg[412]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(c[411]) );
  DFF \sreg_reg[411]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(c[410]) );
  DFF \sreg_reg[410]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(c[409]) );
  DFF \sreg_reg[409]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(c[408]) );
  DFF \sreg_reg[408]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(c[407]) );
  DFF \sreg_reg[407]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(c[406]) );
  DFF \sreg_reg[406]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(c[405]) );
  DFF \sreg_reg[405]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(c[404]) );
  DFF \sreg_reg[404]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(c[403]) );
  DFF \sreg_reg[403]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(c[402]) );
  DFF \sreg_reg[402]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(c[401]) );
  DFF \sreg_reg[401]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(c[400]) );
  DFF \sreg_reg[400]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(c[399]) );
  DFF \sreg_reg[399]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(c[398]) );
  DFF \sreg_reg[398]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(c[397]) );
  DFF \sreg_reg[397]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(c[396]) );
  DFF \sreg_reg[396]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(c[395]) );
  DFF \sreg_reg[395]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(c[394]) );
  DFF \sreg_reg[394]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(c[393]) );
  DFF \sreg_reg[393]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(c[392]) );
  DFF \sreg_reg[392]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(c[391]) );
  DFF \sreg_reg[391]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(c[390]) );
  DFF \sreg_reg[390]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(c[389]) );
  DFF \sreg_reg[389]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(c[388]) );
  DFF \sreg_reg[388]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(c[387]) );
  DFF \sreg_reg[387]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(c[386]) );
  DFF \sreg_reg[386]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(c[385]) );
  DFF \sreg_reg[385]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(c[384]) );
  DFF \sreg_reg[384]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(c[383]) );
  DFF \sreg_reg[383]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(c[382]) );
  DFF \sreg_reg[382]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(c[381]) );
  DFF \sreg_reg[381]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(c[380]) );
  DFF \sreg_reg[380]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(c[379]) );
  DFF \sreg_reg[379]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(c[378]) );
  DFF \sreg_reg[378]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(c[377]) );
  DFF \sreg_reg[377]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(c[376]) );
  DFF \sreg_reg[376]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(c[375]) );
  DFF \sreg_reg[375]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(c[374]) );
  DFF \sreg_reg[374]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(c[373]) );
  DFF \sreg_reg[373]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(c[372]) );
  DFF \sreg_reg[372]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(c[371]) );
  DFF \sreg_reg[371]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(c[370]) );
  DFF \sreg_reg[370]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(c[369]) );
  DFF \sreg_reg[369]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(c[368]) );
  DFF \sreg_reg[368]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(c[367]) );
  DFF \sreg_reg[367]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(c[366]) );
  DFF \sreg_reg[366]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(c[365]) );
  DFF \sreg_reg[365]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(c[364]) );
  DFF \sreg_reg[364]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(c[363]) );
  DFF \sreg_reg[363]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(c[362]) );
  DFF \sreg_reg[362]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(c[361]) );
  DFF \sreg_reg[361]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(c[360]) );
  DFF \sreg_reg[360]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(c[359]) );
  DFF \sreg_reg[359]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(c[358]) );
  DFF \sreg_reg[358]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(c[357]) );
  DFF \sreg_reg[357]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(c[356]) );
  DFF \sreg_reg[356]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(c[355]) );
  DFF \sreg_reg[355]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(c[354]) );
  DFF \sreg_reg[354]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(c[353]) );
  DFF \sreg_reg[353]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(c[352]) );
  DFF \sreg_reg[352]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(c[351]) );
  DFF \sreg_reg[351]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(c[350]) );
  DFF \sreg_reg[350]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(c[349]) );
  DFF \sreg_reg[349]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(c[348]) );
  DFF \sreg_reg[348]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(c[347]) );
  DFF \sreg_reg[347]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(c[346]) );
  DFF \sreg_reg[346]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(c[345]) );
  DFF \sreg_reg[345]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(c[344]) );
  DFF \sreg_reg[344]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(c[343]) );
  DFF \sreg_reg[343]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(c[342]) );
  DFF \sreg_reg[342]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(c[341]) );
  DFF \sreg_reg[341]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(c[340]) );
  DFF \sreg_reg[340]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(c[339]) );
  DFF \sreg_reg[339]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(c[338]) );
  DFF \sreg_reg[338]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(c[337]) );
  DFF \sreg_reg[337]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(c[336]) );
  DFF \sreg_reg[336]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(c[335]) );
  DFF \sreg_reg[335]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(c[334]) );
  DFF \sreg_reg[334]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(c[333]) );
  DFF \sreg_reg[333]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(c[332]) );
  DFF \sreg_reg[332]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(c[331]) );
  DFF \sreg_reg[331]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(c[330]) );
  DFF \sreg_reg[330]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(c[329]) );
  DFF \sreg_reg[329]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(c[328]) );
  DFF \sreg_reg[328]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(c[327]) );
  DFF \sreg_reg[327]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(c[326]) );
  DFF \sreg_reg[326]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(c[325]) );
  DFF \sreg_reg[325]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(c[324]) );
  DFF \sreg_reg[324]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(c[323]) );
  DFF \sreg_reg[323]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(c[322]) );
  DFF \sreg_reg[322]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(c[321]) );
  DFF \sreg_reg[321]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(c[320]) );
  DFF \sreg_reg[320]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(c[319]) );
  DFF \sreg_reg[319]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(c[318]) );
  DFF \sreg_reg[318]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(c[317]) );
  DFF \sreg_reg[317]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(c[316]) );
  DFF \sreg_reg[316]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(c[315]) );
  DFF \sreg_reg[315]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(c[314]) );
  DFF \sreg_reg[314]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(c[313]) );
  DFF \sreg_reg[313]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(c[312]) );
  DFF \sreg_reg[312]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(c[311]) );
  DFF \sreg_reg[311]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(c[310]) );
  DFF \sreg_reg[310]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(c[309]) );
  DFF \sreg_reg[309]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(c[308]) );
  DFF \sreg_reg[308]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(c[307]) );
  DFF \sreg_reg[307]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(c[306]) );
  DFF \sreg_reg[306]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(c[305]) );
  DFF \sreg_reg[305]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(c[304]) );
  DFF \sreg_reg[304]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(c[303]) );
  DFF \sreg_reg[303]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(c[302]) );
  DFF \sreg_reg[302]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(c[301]) );
  DFF \sreg_reg[301]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(c[300]) );
  DFF \sreg_reg[300]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(c[299]) );
  DFF \sreg_reg[299]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(c[298]) );
  DFF \sreg_reg[298]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(c[297]) );
  DFF \sreg_reg[297]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(c[296]) );
  DFF \sreg_reg[296]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(c[295]) );
  DFF \sreg_reg[295]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(c[294]) );
  DFF \sreg_reg[294]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(c[293]) );
  DFF \sreg_reg[293]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(c[292]) );
  DFF \sreg_reg[292]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(c[291]) );
  DFF \sreg_reg[291]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(c[290]) );
  DFF \sreg_reg[290]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(c[289]) );
  DFF \sreg_reg[289]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(c[288]) );
  DFF \sreg_reg[288]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(c[287]) );
  DFF \sreg_reg[287]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(c[286]) );
  DFF \sreg_reg[286]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(c[285]) );
  DFF \sreg_reg[285]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(c[284]) );
  DFF \sreg_reg[284]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(c[283]) );
  DFF \sreg_reg[283]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(c[282]) );
  DFF \sreg_reg[282]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(c[281]) );
  DFF \sreg_reg[281]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(c[280]) );
  DFF \sreg_reg[280]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(c[279]) );
  DFF \sreg_reg[279]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(c[278]) );
  DFF \sreg_reg[278]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(c[277]) );
  DFF \sreg_reg[277]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(c[276]) );
  DFF \sreg_reg[276]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(c[275]) );
  DFF \sreg_reg[275]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(c[274]) );
  DFF \sreg_reg[274]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(c[273]) );
  DFF \sreg_reg[273]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(c[272]) );
  DFF \sreg_reg[272]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(c[271]) );
  DFF \sreg_reg[271]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(c[270]) );
  DFF \sreg_reg[270]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(c[269]) );
  DFF \sreg_reg[269]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(c[268]) );
  DFF \sreg_reg[268]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(c[267]) );
  DFF \sreg_reg[267]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(c[266]) );
  DFF \sreg_reg[266]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(c[265]) );
  DFF \sreg_reg[265]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(c[264]) );
  DFF \sreg_reg[264]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(c[263]) );
  DFF \sreg_reg[263]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(c[262]) );
  DFF \sreg_reg[262]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(c[261]) );
  DFF \sreg_reg[261]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(c[260]) );
  DFF \sreg_reg[260]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(c[259]) );
  DFF \sreg_reg[259]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(c[258]) );
  DFF \sreg_reg[258]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(c[257]) );
  DFF \sreg_reg[257]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(c[256]) );
  DFF \sreg_reg[256]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(c[255]) );
  DFF \sreg_reg[255]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[254]) );
  DFF \sreg_reg[254]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[253]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[252]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[251]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[250]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[249]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[248]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[247]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[246]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[245]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[244]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[243]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[242]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[241]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[240]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[239]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[238]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[237]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[236]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[235]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[234]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[233]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[232]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[231]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[230]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[229]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[228]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[227]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[226]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[225]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[224]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[223]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[222]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[221]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[220]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[219]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[218]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[217]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[216]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[215]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[214]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[213]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[212]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[211]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[210]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[209]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[208]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[207]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[206]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[205]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[204]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[203]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[202]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[201]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[200]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[199]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[198]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[197]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[196]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[195]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[194]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[193]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[192]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[191]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[190]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[189]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[188]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[187]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[186]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[185]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[184]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[183]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[182]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[181]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[180]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[179]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[178]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[177]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[176]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[175]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[174]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[173]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[172]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[171]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[170]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[169]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[168]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[167]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[166]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[165]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[164]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[163]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[162]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[161]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[160]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[159]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[158]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[157]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[156]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[155]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[154]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[153]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[152]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[151]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[150]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[149]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[148]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[147]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[146]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[145]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[144]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[143]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[142]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[141]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[140]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[139]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[138]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[137]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[136]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[135]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[134]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[133]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[132]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[131]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[130]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[129]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[128]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[7]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[6]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[5]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[4]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[3]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[2]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[1]  ( .D(c[1]), .CLK(clk), .RST(rst), .Q(c[0]) );
  ADD_N1024 ADD_ ( .A({1'b0, sreg[2046:1024]}), .B(clocal), .CI(1'b0), .S({
        swire, c[1023]}) );
  mult_N1024_CC1024_DW02_mult_0 mult_44 ( .A(a), .B(b[0]), .TC(1'b0), 
        .PRODUCT({SYNOPSYS_UNCONNECTED__0, clocal}) );
endmodule

