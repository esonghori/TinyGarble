
module FA_1985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_63 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_2015 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2014 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2013 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2012 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2011 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2010 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2009 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2008 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2007 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2006 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2005 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2004 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2003 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2002 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2001 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2000 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1999 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1998 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1997 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1996 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1995 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1994 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1993 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1992 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1991 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_1990 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_1989 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_1988 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_1987 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_1986 \FAINST[30].FA_  ( .A(1'b0), .B(B[30]), .CI(1'b0), .S(S[30]) );
  FA_1985 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(1'b0), .S(S[31]) );
endmodule


module FA_2017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_64 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;
  wire   \C[31] ;

  FA_2047 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2046 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2045 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2044 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2043 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2042 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2041 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2040 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2039 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2038 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2037 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2036 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2035 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2034 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2033 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2032 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2031 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2030 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2029 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2028 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_2027 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_2026 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_2025 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_2024 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_2023 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_2022 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_2021 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_2020 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_2019 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_2018 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(1'b0), .S(S[30]), .CO(
        \C[31] ) );
  FA_2017 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(\C[31] ), .S(S[31]) );
endmodule


module FA_2049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_65 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2079 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2078 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2077 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2076 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2075 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2074 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2073 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2072 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2071 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2070 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2069 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2068 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2067 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2066 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2065 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2064 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2063 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2062 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2061 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2060 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_2059 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_2058 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_2057 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_2056 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_2055 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_2054 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_2053 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_2052 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_2051 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(1'b0), .S(S[29]), .CO(
        C[30]) );
  FA_2050 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2049 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_66 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2111 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2110 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2109 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2108 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2107 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2106 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2105 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2104 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2103 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2102 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2101 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2100 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2099 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2098 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2097 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2096 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2095 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2094 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2093 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2092 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_2091 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_2090 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_2089 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_2088 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_2087 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_2086 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_2085 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_2084 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(1'b0), .S(S[28]), .CO(
        C[29]) );
  FA_2083 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2082 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2081 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_67 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2143 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2142 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2141 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2140 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2139 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2138 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2137 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2136 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2135 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2134 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2133 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2132 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2131 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2130 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2129 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2128 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2127 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2126 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2125 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2124 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_2123 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_2122 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_2121 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_2120 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_2119 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_2118 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_2117 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(1'b0), .S(S[27]), .CO(
        C[28]) );
  FA_2116 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2115 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2114 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2113 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_68 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2175 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2174 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2173 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2172 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2171 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2170 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2169 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2168 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2167 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2166 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2165 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2164 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2163 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2162 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2161 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2160 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2159 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2158 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2157 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2156 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_2155 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_2154 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_2153 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_2152 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_2151 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_2150 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(1'b0), .S(S[26]), .CO(
        C[27]) );
  FA_2149 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2148 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2147 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2146 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2145 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_69 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2207 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2206 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2205 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2204 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2203 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2202 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2201 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2200 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2199 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2198 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2197 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2196 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2195 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2194 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2193 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2192 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2191 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2190 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2189 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2188 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_2187 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_2186 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_2185 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_2184 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_2183 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(1'b0), .S(S[25]), .CO(
        C[26]) );
  FA_2182 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2181 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2180 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2179 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2178 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2177 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_70 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2239 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2238 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2237 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2236 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2235 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2234 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2233 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2232 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2231 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2230 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2229 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2228 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2227 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2226 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2225 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2224 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2223 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2222 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2221 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2220 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_2219 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_2218 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_2217 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_2216 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(1'b0), .S(S[24]), .CO(
        C[25]) );
  FA_2215 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2214 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2213 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2212 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2211 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2210 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2209 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_71 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2271 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2270 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2269 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2268 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2267 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2266 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2265 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2264 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2263 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2262 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2261 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2260 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2259 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2258 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2257 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2256 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2255 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2254 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2253 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2252 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_2251 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_2250 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_2249 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(1'b0), .S(S[23]), .CO(
        C[24]) );
  FA_2248 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2247 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2246 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2245 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2244 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2243 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2242 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2241 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_72 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2303 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2302 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2301 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2300 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2299 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2298 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2297 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2296 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2295 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2294 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2293 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2292 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2291 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2290 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2289 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2288 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2287 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2286 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2285 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2284 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_2283 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_2282 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(1'b0), .S(S[22]), .CO(
        C[23]) );
  FA_2281 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2280 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2279 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2278 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2277 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2276 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2275 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2274 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2273 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_73 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2335 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2334 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2333 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2332 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2331 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2330 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2329 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2328 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2327 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2326 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2325 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2324 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2323 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2322 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2321 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2320 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2319 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2318 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2317 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2316 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_2315 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(1'b0), .S(S[21]), .CO(
        C[22]) );
  FA_2314 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2313 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2312 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2311 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2310 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2309 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2308 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2307 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2306 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2305 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_74 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2367 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2366 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2365 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2364 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2363 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2362 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2361 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2360 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2359 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2358 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2357 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2356 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2355 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2354 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2353 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2352 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2351 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2350 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2349 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2348 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(1'b0), .S(S[20]), .CO(
        C[21]) );
  FA_2347 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2346 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2345 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2344 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2343 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2342 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2341 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2340 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2339 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2338 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2337 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_75 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2399 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2398 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2397 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2396 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2395 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2394 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2393 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2392 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2391 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2390 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2389 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2388 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2387 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2386 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2385 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2384 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2383 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2382 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2381 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(1'b0), .S(S[19]), .CO(
        C[20]) );
  FA_2380 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2379 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2378 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2377 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2376 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2375 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2374 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2373 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2372 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2371 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2370 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2369 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_76 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2431 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2430 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2429 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2428 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2427 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2426 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2425 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2424 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2423 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2422 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2421 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2420 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2419 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2418 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2417 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2416 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2415 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2414 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(1'b0), .S(S[18]), .CO(
        C[19]) );
  FA_2413 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2412 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2411 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2410 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2409 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2408 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2407 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2406 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2405 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2404 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2403 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2402 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2401 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_77 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2463 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2462 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2461 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2460 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2459 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2458 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2457 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2456 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2455 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2454 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2453 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2452 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2451 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2450 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2449 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2448 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2447 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(1'b0), .S(S[17]), .CO(
        C[18]) );
  FA_2446 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2445 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2444 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2443 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2442 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2441 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2440 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2439 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2438 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2437 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2436 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2435 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2434 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2433 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_78 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2495 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2494 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2493 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2492 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2491 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2490 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2489 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2488 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2487 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2486 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2485 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2484 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2483 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2482 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2481 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2480 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(1'b0), .S(S[16]), .CO(
        C[17]) );
  FA_2479 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2478 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2477 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2476 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2475 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2474 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2473 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2472 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2471 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2470 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2469 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2468 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2467 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2466 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2465 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_79 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2527 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2526 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2525 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2524 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2523 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2522 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2521 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2520 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2519 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2518 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2517 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2516 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2515 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2514 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2513 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(1'b0), .S(S[15]), .CO(
        C[16]) );
  FA_2512 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2511 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2510 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2509 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2508 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2507 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2506 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2505 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2504 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2503 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2502 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2501 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2500 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2499 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2498 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2497 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_80 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2559 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2558 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2557 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2556 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2555 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2554 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2553 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2552 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2551 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2550 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2549 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2548 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2547 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2546 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(1'b0), .S(S[14]), .CO(
        C[15]) );
  FA_2545 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2544 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2543 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2542 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2541 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2540 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2539 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2538 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2537 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2536 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2535 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2534 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2533 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2532 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2531 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2530 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2529 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_81 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2591 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2590 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2589 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2588 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2587 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2586 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2585 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2584 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2583 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2582 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2581 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2580 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2579 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(1'b0), .S(S[13]), .CO(
        C[14]) );
  FA_2578 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2577 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2576 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2575 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2574 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2573 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2572 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2571 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2570 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2569 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2568 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2567 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2566 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2565 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2564 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2563 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2562 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2561 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_82 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2623 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2622 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2621 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2620 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2619 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2618 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2617 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2616 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2615 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2614 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2613 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2612 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(1'b0), .S(S[12]), .CO(
        C[13]) );
  FA_2611 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2610 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2609 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2608 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2607 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2606 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2605 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2604 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2603 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2602 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2601 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2600 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2599 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2598 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2597 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2596 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2595 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2594 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2593 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_83 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2655 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2654 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2653 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2652 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2651 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2650 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2649 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2648 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2647 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2646 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2645 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(1'b0), .S(S[11]), .CO(
        C[12]) );
  FA_2644 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2643 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2642 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2641 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2640 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2639 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2638 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2637 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2636 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2635 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2634 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2633 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2632 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2631 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2630 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2629 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2628 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2627 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2626 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2625 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_84 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2687 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2686 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2685 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2684 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2683 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2682 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2681 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2680 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2679 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2678 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(1'b0), .S(S[10]), .CO(
        C[11]) );
  FA_2677 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2676 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2675 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2674 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2673 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2672 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2671 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2670 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2669 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2668 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2667 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2666 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2665 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2664 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2663 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2662 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2661 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2660 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2659 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2658 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2657 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_85 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2719 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2718 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2717 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2716 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2715 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2714 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2713 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2712 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2711 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(1'b0), .S(S[9]), .CO(C[10]) );
  FA_2710 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2709 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2708 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2707 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2706 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2705 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2704 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2703 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2702 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2701 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2700 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2699 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2698 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2697 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2696 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2695 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2694 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2693 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2692 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2691 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2690 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2689 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_86 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2751 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2750 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2749 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2748 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2747 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2746 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2745 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2744 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(1'b0), .S(S[8]), .CO(C[9])
         );
  FA_2743 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_2742 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2741 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2740 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2739 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2738 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2737 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2736 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2735 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2734 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2733 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2732 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2731 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2730 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2729 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2728 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2727 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2726 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2725 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2724 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2723 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2722 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2721 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_87 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2783 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2782 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2781 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2780 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2779 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2778 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2777 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(1'b0), .S(S[7]), .CO(C[8])
         );
  FA_2776 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_2775 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_2774 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2773 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2772 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2771 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2770 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2769 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2768 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2767 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2766 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2765 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2764 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2763 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2762 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2761 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2760 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2759 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2758 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2757 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2756 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2755 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2754 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2753 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_88 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2815 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2814 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2813 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2812 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2811 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2810 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(1'b0), .S(S[6]), .CO(C[7])
         );
  FA_2809 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_2808 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_2807 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_2806 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2805 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2804 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2803 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2802 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2801 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2800 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2799 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2798 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2797 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2796 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2795 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2794 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2793 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2792 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2791 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2790 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2789 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2788 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2787 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2786 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2785 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_89 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2847 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2846 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2845 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2844 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2843 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(1'b0), .S(S[5]), .CO(C[6])
         );
  FA_2842 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_2841 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_2840 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_2839 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_2838 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2837 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2836 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2835 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2834 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2833 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2832 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2831 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2830 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2829 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2828 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2827 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2826 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2825 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2824 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2823 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2822 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2821 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2820 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2819 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2818 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2817 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_90 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2879 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2878 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2877 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2876 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(1'b0), .S(S[4]), .CO(C[5])
         );
  FA_2875 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_2874 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_2873 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_2872 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_2871 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_2870 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2869 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2868 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2867 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2866 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2865 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2864 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2863 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2862 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2861 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2860 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2859 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2858 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2857 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2856 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2855 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2854 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2853 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2852 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2851 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2850 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2849 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_91 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2911 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2910 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2909 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(1'b0), .S(S[3]), .CO(C[4])
         );
  FA_2908 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_2907 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_2906 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_2905 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_2904 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_2903 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_2902 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2901 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2900 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2899 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2898 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2897 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2896 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2895 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2894 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2893 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2892 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2891 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2890 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2889 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2888 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2887 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2886 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2885 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2884 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2883 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2882 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2881 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_92 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2943 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2942 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(1'b0), .S(S[2]), .CO(C[3])
         );
  FA_2941 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_2940 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_2939 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_2938 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_2937 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_2936 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_2935 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_2934 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2933 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2932 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2931 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2930 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2929 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2928 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2927 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2926 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2925 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2924 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2923 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2922 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2921 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2920 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2919 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2918 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2917 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2916 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2915 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2914 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2913 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_2945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_2975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module ADD_N32_93 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_2975 \FAINST[1].FA_  ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(S[1]) );
  FA_2974 \FAINST[2].FA_  ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(S[2]) );
  FA_2973 \FAINST[3].FA_  ( .A(A[3]), .B(1'b0), .CI(1'b0), .S(S[3]) );
  FA_2972 \FAINST[4].FA_  ( .A(A[4]), .B(1'b0), .CI(1'b0), .S(S[4]) );
  FA_2971 \FAINST[5].FA_  ( .A(A[5]), .B(1'b0), .CI(1'b0), .S(S[5]) );
  FA_2970 \FAINST[6].FA_  ( .A(A[6]), .B(1'b0), .CI(1'b0), .S(S[6]) );
  FA_2969 \FAINST[7].FA_  ( .A(A[7]), .B(1'b0), .CI(1'b0), .S(S[7]) );
  FA_2968 \FAINST[8].FA_  ( .A(A[8]), .B(1'b0), .CI(1'b0), .S(S[8]) );
  FA_2967 \FAINST[9].FA_  ( .A(A[9]), .B(1'b0), .CI(1'b0), .S(S[9]) );
  FA_2966 \FAINST[10].FA_  ( .A(A[10]), .B(1'b0), .CI(1'b0), .S(S[10]) );
  FA_2965 \FAINST[11].FA_  ( .A(A[11]), .B(1'b0), .CI(1'b0), .S(S[11]) );
  FA_2964 \FAINST[12].FA_  ( .A(A[12]), .B(1'b0), .CI(1'b0), .S(S[12]) );
  FA_2963 \FAINST[13].FA_  ( .A(A[13]), .B(1'b0), .CI(1'b0), .S(S[13]) );
  FA_2962 \FAINST[14].FA_  ( .A(A[14]), .B(1'b0), .CI(1'b0), .S(S[14]) );
  FA_2961 \FAINST[15].FA_  ( .A(A[15]), .B(1'b0), .CI(1'b0), .S(S[15]) );
  FA_2960 \FAINST[16].FA_  ( .A(A[16]), .B(1'b0), .CI(1'b0), .S(S[16]) );
  FA_2959 \FAINST[17].FA_  ( .A(A[17]), .B(1'b0), .CI(1'b0), .S(S[17]) );
  FA_2958 \FAINST[18].FA_  ( .A(A[18]), .B(1'b0), .CI(1'b0), .S(S[18]) );
  FA_2957 \FAINST[19].FA_  ( .A(A[19]), .B(1'b0), .CI(1'b0), .S(S[19]) );
  FA_2956 \FAINST[20].FA_  ( .A(A[20]), .B(1'b0), .CI(1'b0), .S(S[20]) );
  FA_2955 \FAINST[21].FA_  ( .A(A[21]), .B(1'b0), .CI(1'b0), .S(S[21]) );
  FA_2954 \FAINST[22].FA_  ( .A(A[22]), .B(1'b0), .CI(1'b0), .S(S[22]) );
  FA_2953 \FAINST[23].FA_  ( .A(A[23]), .B(1'b0), .CI(1'b0), .S(S[23]) );
  FA_2952 \FAINST[24].FA_  ( .A(A[24]), .B(1'b0), .CI(1'b0), .S(S[24]) );
  FA_2951 \FAINST[25].FA_  ( .A(A[25]), .B(1'b0), .CI(1'b0), .S(S[25]) );
  FA_2950 \FAINST[26].FA_  ( .A(A[26]), .B(1'b0), .CI(1'b0), .S(S[26]) );
  FA_2949 \FAINST[27].FA_  ( .A(A[27]), .B(1'b0), .CI(1'b0), .S(S[27]) );
  FA_2948 \FAINST[28].FA_  ( .A(A[28]), .B(1'b0), .CI(1'b0), .S(S[28]) );
  FA_2947 \FAINST[29].FA_  ( .A(A[29]), .B(1'b0), .CI(1'b0), .S(S[29]) );
  FA_2946 \FAINST[30].FA_  ( .A(A[30]), .B(1'b0), .CI(1'b0), .S(S[30]) );
  FA_2945 \FAINST[31].FA_  ( .A(A[31]), .B(1'b0), .CI(1'b0), .S(S[31]) );
endmodule


module MULT_N32_0 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   \w[31][31] , \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] ,
         \w[31][26] , \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] ,
         \w[31][21] , \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] ,
         \w[31][16] , \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] ,
         \w[31][11] , \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] ,
         \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] ,
         \w[31][1] , \w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] ,
         \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] ,
         \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] ,
         \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] ,
         \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] ,
         \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] ,
         \w[30][2] , \w[30][1] , \w[29][31] , \w[29][30] , \w[29][29] ,
         \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] ,
         \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] ,
         \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] ,
         \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] ,
         \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] ,
         \w[29][3] , \w[29][2] , \w[29][1] , \w[28][31] , \w[28][30] ,
         \w[28][29] , \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] ,
         \w[28][24] , \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] ,
         \w[28][19] , \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] ,
         \w[28][14] , \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] ,
         \w[28][9] , \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] ,
         \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , \w[27][31] ,
         \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] ,
         \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] ,
         \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] ,
         \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] ,
         \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] ,
         \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] ,
         \w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] ,
         \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] ,
         \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] ,
         \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] ,
         \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] ,
         \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] ,
         \w[26][1] , \w[25][31] , \w[25][30] , \w[25][29] , \w[25][28] ,
         \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , \w[25][23] ,
         \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , \w[25][18] ,
         \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , \w[25][13] ,
         \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , \w[25][8] ,
         \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] ,
         \w[25][2] , \w[25][1] , \w[24][31] , \w[24][30] , \w[24][29] ,
         \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] ,
         \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] ,
         \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] ,
         \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] ,
         \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] ,
         \w[24][3] , \w[24][2] , \w[24][1] , \w[23][31] , \w[23][30] ,
         \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] ,
         \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] ,
         \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] ,
         \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] ,
         \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] ,
         \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , \w[22][31] ,
         \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , \w[22][26] ,
         \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , \w[22][21] ,
         \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , \w[22][16] ,
         \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , \w[22][11] ,
         \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , \w[22][6] ,
         \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] ,
         \w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] ,
         \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] ,
         \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] ,
         \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] ,
         \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] ,
         \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] ,
         \w[21][1] , \w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] ,
         \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] ,
         \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] ,
         \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] ,
         \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] ,
         \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] ,
         \w[20][2] , \w[20][1] , \w[19][31] , \w[19][30] , \w[19][29] ,
         \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] ,
         \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] ,
         \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] ,
         \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] ,
         \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] ,
         \w[19][3] , \w[19][2] , \w[19][1] , \w[18][31] , \w[18][30] ,
         \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] ,
         \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] ,
         \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] ,
         \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] ,
         \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] ,
         \w[18][4] , \w[18][3] , \w[18][2] , \w[18][1] , \w[17][31] ,
         \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] ,
         \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] ,
         \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] ,
         \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] ,
         \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] ,
         \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] ,
         \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] ,
         \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] ,
         \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] ,
         \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] ,
         \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] ,
         \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] ,
         \w[16][1] , \w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] ,
         \w[15][27] , \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] ,
         \w[15][22] , \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] ,
         \w[15][17] , \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] ,
         \w[15][12] , \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] ,
         \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] ,
         \w[15][2] , \w[15][1] , \w[14][31] , \w[14][30] , \w[14][29] ,
         \w[14][28] , \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] ,
         \w[14][23] , \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] ,
         \w[14][18] , \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] ,
         \w[14][13] , \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] ,
         \w[14][8] , \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] ,
         \w[14][3] , \w[14][2] , \w[14][1] , \w[13][31] , \w[13][30] ,
         \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] ,
         \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] ,
         \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] ,
         \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] ,
         \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] ,
         \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , \w[12][31] ,
         \w[12][30] , \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] ,
         \w[12][25] , \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] ,
         \w[12][20] , \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] ,
         \w[12][15] , \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] ,
         \w[12][10] , \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] ,
         \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , \w[12][1] ,
         \w[11][31] , \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] ,
         \w[11][26] , \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] ,
         \w[11][21] , \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] ,
         \w[11][16] , \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] ,
         \w[11][11] , \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] ,
         \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] ,
         \w[11][1] , \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] ,
         \w[10][27] , \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] ,
         \w[10][22] , \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] ,
         \w[10][17] , \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] ,
         \w[10][12] , \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] ,
         \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] ,
         \w[10][2] , \w[10][1] , \w[9][31] , \w[9][30] , \w[9][29] ,
         \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] ,
         \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] ,
         \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] ,
         \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] ,
         \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] ,
         \w[9][1] , \w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] ,
         \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] ,
         \w[8][21] , \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] ,
         \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , \w[8][12] ,
         \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , \w[8][6] ,
         \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , \w[7][31] ,
         \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] ,
         \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] ,
         \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] ,
         \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] ,
         \w[7][10] , \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] ,
         \w[7][4] , \w[7][3] , \w[7][2] , \w[7][1] , \w[6][31] , \w[6][30] ,
         \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] ,
         \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] ,
         \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] ,
         \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] ,
         \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] ,
         \w[6][2] , \w[6][1] , \w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] ,
         \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] ,
         \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] ,
         \w[5][17] , \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] ,
         \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] ,
         \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] ,
         \w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] ,
         \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] ,
         \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] ,
         \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] ,
         \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] ,
         \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , \w[3][31] ,
         \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] ,
         \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] ,
         \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] ,
         \w[3][15] , \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] ,
         \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] ,
         \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , \w[2][31] , \w[2][30] ,
         \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] ,
         \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] ,
         \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] ,
         \w[2][14] , \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] ,
         \w[2][8] , \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] ,
         \w[2][2] , \w[2][1] , \_0_net_[31] , \_0_net_[30] , \_0_net_[29] ,
         \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , \_0_net_[25] ,
         \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , \_0_net_[21] ,
         \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , \_0_net_[17] ,
         \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , \_0_net_[13] ,
         \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , \_0_net_[9] ,
         \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] ,
         \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_2_net_[31] ,
         \_2_net_[30] , \_2_net_[29] , \_2_net_[28] , \_2_net_[27] ,
         \_2_net_[26] , \_2_net_[25] , \_2_net_[24] , \_2_net_[23] ,
         \_2_net_[22] , \_2_net_[21] , \_2_net_[20] , \_2_net_[19] ,
         \_2_net_[18] , \_2_net_[17] , \_2_net_[16] , \_2_net_[15] ,
         \_2_net_[14] , \_2_net_[13] , \_2_net_[12] , \_2_net_[11] ,
         \_2_net_[10] , \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] ,
         \_2_net_[5] , \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , \_4_net_[31] ,
         \_4_net_[30] , \_4_net_[29] , \_4_net_[28] , \_4_net_[27] ,
         \_4_net_[26] , \_4_net_[25] , \_4_net_[24] , \_4_net_[23] ,
         \_4_net_[22] , \_4_net_[21] , \_4_net_[20] , \_4_net_[19] ,
         \_4_net_[18] , \_4_net_[17] , \_4_net_[16] , \_4_net_[15] ,
         \_4_net_[14] , \_4_net_[13] , \_4_net_[12] , \_4_net_[11] ,
         \_4_net_[10] , \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] ,
         \_4_net_[5] , \_4_net_[4] , \_4_net_[3] , \_6_net_[31] ,
         \_6_net_[30] , \_6_net_[29] , \_6_net_[28] , \_6_net_[27] ,
         \_6_net_[26] , \_6_net_[25] , \_6_net_[24] , \_6_net_[23] ,
         \_6_net_[22] , \_6_net_[21] , \_6_net_[20] , \_6_net_[19] ,
         \_6_net_[18] , \_6_net_[17] , \_6_net_[16] , \_6_net_[15] ,
         \_6_net_[14] , \_6_net_[13] , \_6_net_[12] , \_6_net_[11] ,
         \_6_net_[10] , \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] ,
         \_6_net_[5] , \_6_net_[4] , \_8_net_[31] , \_8_net_[30] ,
         \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] ,
         \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] ,
         \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] ,
         \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] ,
         \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] ,
         \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] ,
         \_10_net_[31] , \_10_net_[30] , \_10_net_[29] , \_10_net_[28] ,
         \_10_net_[27] , \_10_net_[26] , \_10_net_[25] , \_10_net_[24] ,
         \_10_net_[23] , \_10_net_[22] , \_10_net_[21] , \_10_net_[20] ,
         \_10_net_[19] , \_10_net_[18] , \_10_net_[17] , \_10_net_[16] ,
         \_10_net_[15] , \_10_net_[14] , \_10_net_[13] , \_10_net_[12] ,
         \_10_net_[11] , \_10_net_[10] , \_10_net_[9] , \_10_net_[8] ,
         \_10_net_[7] , \_10_net_[6] , \_12_net_[31] , \_12_net_[30] ,
         \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] ,
         \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] ,
         \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] ,
         \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] ,
         \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] ,
         \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , \_14_net_[31] ,
         \_14_net_[30] , \_14_net_[29] , \_14_net_[28] , \_14_net_[27] ,
         \_14_net_[26] , \_14_net_[25] , \_14_net_[24] , \_14_net_[23] ,
         \_14_net_[22] , \_14_net_[21] , \_14_net_[20] , \_14_net_[19] ,
         \_14_net_[18] , \_14_net_[17] , \_14_net_[16] , \_14_net_[15] ,
         \_14_net_[14] , \_14_net_[13] , \_14_net_[12] , \_14_net_[11] ,
         \_14_net_[10] , \_14_net_[9] , \_14_net_[8] , \_16_net_[31] ,
         \_16_net_[30] , \_16_net_[29] , \_16_net_[28] , \_16_net_[27] ,
         \_16_net_[26] , \_16_net_[25] , \_16_net_[24] , \_16_net_[23] ,
         \_16_net_[22] , \_16_net_[21] , \_16_net_[20] , \_16_net_[19] ,
         \_16_net_[18] , \_16_net_[17] , \_16_net_[16] , \_16_net_[15] ,
         \_16_net_[14] , \_16_net_[13] , \_16_net_[12] , \_16_net_[11] ,
         \_16_net_[10] , \_16_net_[9] , \_18_net_[31] , \_18_net_[30] ,
         \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] ,
         \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] ,
         \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] ,
         \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] ,
         \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] ,
         \_20_net_[31] , \_20_net_[30] , \_20_net_[29] , \_20_net_[28] ,
         \_20_net_[27] , \_20_net_[26] , \_20_net_[25] , \_20_net_[24] ,
         \_20_net_[23] , \_20_net_[22] , \_20_net_[21] , \_20_net_[20] ,
         \_20_net_[19] , \_20_net_[18] , \_20_net_[17] , \_20_net_[16] ,
         \_20_net_[15] , \_20_net_[14] , \_20_net_[13] , \_20_net_[12] ,
         \_20_net_[11] , \_22_net_[31] , \_22_net_[30] , \_22_net_[29] ,
         \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , \_22_net_[25] ,
         \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , \_22_net_[21] ,
         \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , \_22_net_[17] ,
         \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , \_22_net_[13] ,
         \_22_net_[12] , \_24_net_[31] , \_24_net_[30] , \_24_net_[29] ,
         \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , \_24_net_[25] ,
         \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , \_24_net_[21] ,
         \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , \_24_net_[17] ,
         \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , \_24_net_[13] ,
         \_26_net_[31] , \_26_net_[30] , \_26_net_[29] , \_26_net_[28] ,
         \_26_net_[27] , \_26_net_[26] , \_26_net_[25] , \_26_net_[24] ,
         \_26_net_[23] , \_26_net_[22] , \_26_net_[21] , \_26_net_[20] ,
         \_26_net_[19] , \_26_net_[18] , \_26_net_[17] , \_26_net_[16] ,
         \_26_net_[15] , \_26_net_[14] , \_28_net_[31] , \_28_net_[30] ,
         \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] ,
         \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] ,
         \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] ,
         \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , \_30_net_[31] ,
         \_30_net_[30] , \_30_net_[29] , \_30_net_[28] , \_30_net_[27] ,
         \_30_net_[26] , \_30_net_[25] , \_30_net_[24] , \_30_net_[23] ,
         \_30_net_[22] , \_30_net_[21] , \_30_net_[20] , \_30_net_[19] ,
         \_30_net_[18] , \_30_net_[17] , \_30_net_[16] , \_32_net_[31] ,
         \_32_net_[30] , \_32_net_[29] , \_32_net_[28] , \_32_net_[27] ,
         \_32_net_[26] , \_32_net_[25] , \_32_net_[24] , \_32_net_[23] ,
         \_32_net_[22] , \_32_net_[21] , \_32_net_[20] , \_32_net_[19] ,
         \_32_net_[18] , \_32_net_[17] , \_34_net_[31] , \_34_net_[30] ,
         \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] ,
         \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] ,
         \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] ,
         \_36_net_[31] , \_36_net_[30] , \_36_net_[29] , \_36_net_[28] ,
         \_36_net_[27] , \_36_net_[26] , \_36_net_[25] , \_36_net_[24] ,
         \_36_net_[23] , \_36_net_[22] , \_36_net_[21] , \_36_net_[20] ,
         \_36_net_[19] , \_38_net_[31] , \_38_net_[30] , \_38_net_[29] ,
         \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , \_38_net_[25] ,
         \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , \_38_net_[21] ,
         \_38_net_[20] , \_40_net_[31] , \_40_net_[30] , \_40_net_[29] ,
         \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , \_40_net_[25] ,
         \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , \_40_net_[21] ,
         \_42_net_[31] , \_42_net_[30] , \_42_net_[29] , \_42_net_[28] ,
         \_42_net_[27] , \_42_net_[26] , \_42_net_[25] , \_42_net_[24] ,
         \_42_net_[23] , \_42_net_[22] , \_44_net_[31] , \_44_net_[30] ,
         \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] ,
         \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , \_46_net_[31] ,
         \_46_net_[30] , \_46_net_[29] , \_46_net_[28] , \_46_net_[27] ,
         \_46_net_[26] , \_46_net_[25] , \_46_net_[24] , \_48_net_[31] ,
         \_48_net_[30] , \_48_net_[29] , \_48_net_[28] , \_48_net_[27] ,
         \_48_net_[26] , \_48_net_[25] , \_50_net_[31] , \_50_net_[30] ,
         \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] ,
         \_52_net_[31] , \_52_net_[30] , \_52_net_[29] , \_52_net_[28] ,
         \_52_net_[27] , \_54_net_[31] , \_54_net_[30] , \_54_net_[29] ,
         \_54_net_[28] , \_56_net_[31] , \_56_net_[30] , \_56_net_[29] ,
         \_58_net_[31] , \_58_net_[30] , \_60_net_[31] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  ADD_N32_93 \FAINST[1].ADD_  ( .A({\_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .S({
        \w[2][31] , \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , 
        \w[2][25] , \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , 
        \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , 
        \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , 
        \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , 
        \w[2][1] , SYNOPSYS_UNCONNECTED__0}) );
  ADD_N32_92 \FAINST[2].ADD_  ( .A({\_2_net_[31] , \_2_net_[30] , 
        \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , \_2_net_[26] , 
        \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , \_2_net_[22] , 
        \_2_net_[21] , \_2_net_[20] , \_2_net_[19] , \_2_net_[18] , 
        \_2_net_[17] , \_2_net_[16] , \_2_net_[15] , \_2_net_[14] , 
        \_2_net_[13] , \_2_net_[12] , \_2_net_[11] , \_2_net_[10] , 
        \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , \_2_net_[5] , 
        \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , 1'b0, 1'b0}), .B({\w[2][31] , 
        \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] , 
        \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , \w[2][19] , 
        \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , \w[2][13] , 
        \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , \w[2][7] , 
        \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , \w[2][1] , 1'b0}), .CI(1'b0), .S({\w[3][31] , \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , 
        \w[3][26] , \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , 
        \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , 
        \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , 
        \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , 
        \w[3][2] , \w[3][1] , SYNOPSYS_UNCONNECTED__1}) );
  ADD_N32_91 \FAINST[3].ADD_  ( .A({\_4_net_[31] , \_4_net_[30] , 
        \_4_net_[29] , \_4_net_[28] , \_4_net_[27] , \_4_net_[26] , 
        \_4_net_[25] , \_4_net_[24] , \_4_net_[23] , \_4_net_[22] , 
        \_4_net_[21] , \_4_net_[20] , \_4_net_[19] , \_4_net_[18] , 
        \_4_net_[17] , \_4_net_[16] , \_4_net_[15] , \_4_net_[14] , 
        \_4_net_[13] , \_4_net_[12] , \_4_net_[11] , \_4_net_[10] , 
        \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] , \_4_net_[5] , 
        \_4_net_[4] , \_4_net_[3] , 1'b0, 1'b0, 1'b0}), .B({\w[3][31] , 
        \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] , \w[3][25] , 
        \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , \w[3][20] , \w[3][19] , 
        \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , \w[3][14] , \w[3][13] , 
        \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , 
        \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , 1'b0}), .CI(1'b0), .S({\w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] , 
        \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] , \w[4][21] , 
        \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] , \w[4][16] , \w[4][15] , 
        \w[4][14] , \w[4][13] , \w[4][12] , \w[4][11] , \w[4][10] , \w[4][9] , 
        \w[4][8] , \w[4][7] , \w[4][6] , \w[4][5] , \w[4][4] , \w[4][3] , 
        \w[4][2] , \w[4][1] , SYNOPSYS_UNCONNECTED__2}) );
  ADD_N32_90 \FAINST[4].ADD_  ( .A({\_6_net_[31] , \_6_net_[30] , 
        \_6_net_[29] , \_6_net_[28] , \_6_net_[27] , \_6_net_[26] , 
        \_6_net_[25] , \_6_net_[24] , \_6_net_[23] , \_6_net_[22] , 
        \_6_net_[21] , \_6_net_[20] , \_6_net_[19] , \_6_net_[18] , 
        \_6_net_[17] , \_6_net_[16] , \_6_net_[15] , \_6_net_[14] , 
        \_6_net_[13] , \_6_net_[12] , \_6_net_[11] , \_6_net_[10] , 
        \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] , \_6_net_[5] , 
        \_6_net_[4] , 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[4][31] , \w[4][30] , 
        \w[4][29] , \w[4][28] , \w[4][27] , \w[4][26] , \w[4][25] , \w[4][24] , 
        \w[4][23] , \w[4][22] , \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , 
        \w[4][17] , \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] , 
        \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] , 
        \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , 1'b0}), .CI(
        1'b0), .S({\w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] , \w[5][27] , 
        \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , \w[5][22] , \w[5][21] , 
        \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , \w[5][16] , \w[5][15] , 
        \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , 
        \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , 
        \w[5][2] , \w[5][1] , SYNOPSYS_UNCONNECTED__3}) );
  ADD_N32_89 \FAINST[5].ADD_  ( .A({\_8_net_[31] , \_8_net_[30] , 
        \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] , 
        \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] , 
        \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] , 
        \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] , 
        \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] , 
        \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[5][31] , \w[5][30] , \w[5][29] , 
        \w[5][28] , \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , 
        \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , 
        \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , 
        \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , 
        \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] , 1'b0}), .CI(1'b0), .S({
        \w[6][31] , \w[6][30] , \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , 
        \w[6][25] , \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] , 
        \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] , \w[6][14] , 
        \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] , \w[6][8] , 
        \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] , \w[6][2] , 
        \w[6][1] , SYNOPSYS_UNCONNECTED__4}) );
  ADD_N32_88 \FAINST[6].ADD_  ( .A({\_10_net_[31] , \_10_net_[30] , 
        \_10_net_[29] , \_10_net_[28] , \_10_net_[27] , \_10_net_[26] , 
        \_10_net_[25] , \_10_net_[24] , \_10_net_[23] , \_10_net_[22] , 
        \_10_net_[21] , \_10_net_[20] , \_10_net_[19] , \_10_net_[18] , 
        \_10_net_[17] , \_10_net_[16] , \_10_net_[15] , \_10_net_[14] , 
        \_10_net_[13] , \_10_net_[12] , \_10_net_[11] , \_10_net_[10] , 
        \_10_net_[9] , \_10_net_[8] , \_10_net_[7] , \_10_net_[6] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[6][31] , \w[6][30] , \w[6][29] , 
        \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] , \w[6][24] , \w[6][23] , 
        \w[6][22] , \w[6][21] , \w[6][20] , \w[6][19] , \w[6][18] , \w[6][17] , 
        \w[6][16] , \w[6][15] , \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , 
        \w[6][10] , \w[6][9] , \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , 
        \w[6][4] , \w[6][3] , \w[6][2] , \w[6][1] , 1'b0}), .CI(1'b0), .S({
        \w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] , 
        \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] , \w[7][20] , 
        \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , \w[7][15] , \w[7][14] , 
        \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , \w[7][9] , \w[7][8] , 
        \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , \w[7][3] , \w[7][2] , 
        \w[7][1] , SYNOPSYS_UNCONNECTED__5}) );
  ADD_N32_87 \FAINST[7].ADD_  ( .A({\_12_net_[31] , \_12_net_[30] , 
        \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] , 
        \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] , 
        \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] , 
        \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] , 
        \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] , 
        \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , 
        \w[7][27] , \w[7][26] , \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , 
        \w[7][21] , \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , 
        \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , 
        \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , 
        \w[7][3] , \w[7][2] , \w[7][1] , 1'b0}), .CI(1'b0), .S({\w[8][31] , 
        \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , \w[8][26] , \w[8][25] , 
        \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , \w[8][20] , \w[8][19] , 
        \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , 
        \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , 
        \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , 
        SYNOPSYS_UNCONNECTED__6}) );
  ADD_N32_86 \FAINST[8].ADD_  ( .A({\_14_net_[31] , \_14_net_[30] , 
        \_14_net_[29] , \_14_net_[28] , \_14_net_[27] , \_14_net_[26] , 
        \_14_net_[25] , \_14_net_[24] , \_14_net_[23] , \_14_net_[22] , 
        \_14_net_[21] , \_14_net_[20] , \_14_net_[19] , \_14_net_[18] , 
        \_14_net_[17] , \_14_net_[16] , \_14_net_[15] , \_14_net_[14] , 
        \_14_net_[13] , \_14_net_[12] , \_14_net_[11] , \_14_net_[10] , 
        \_14_net_[9] , \_14_net_[8] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , 
        \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , 
        \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , 
        \w[8][14] , \w[8][13] , \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , 
        \w[8][8] , \w[8][7] , \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , 
        \w[8][2] , \w[8][1] , 1'b0}), .CI(1'b0), .S({\w[9][31] , \w[9][30] , 
        \w[9][29] , \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] , 
        \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] , \w[9][18] , 
        \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] , \w[9][13] , \w[9][12] , 
        \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] , \w[9][7] , \w[9][6] , 
        \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] , \w[9][1] , 
        SYNOPSYS_UNCONNECTED__7}) );
  ADD_N32_85 \FAINST[9].ADD_  ( .A({\_16_net_[31] , \_16_net_[30] , 
        \_16_net_[29] , \_16_net_[28] , \_16_net_[27] , \_16_net_[26] , 
        \_16_net_[25] , \_16_net_[24] , \_16_net_[23] , \_16_net_[22] , 
        \_16_net_[21] , \_16_net_[20] , \_16_net_[19] , \_16_net_[18] , 
        \_16_net_[17] , \_16_net_[16] , \_16_net_[15] , \_16_net_[14] , 
        \_16_net_[13] , \_16_net_[12] , \_16_net_[11] , \_16_net_[10] , 
        \_16_net_[9] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[9][31] , \w[9][30] , \w[9][29] , \w[9][28] , \w[9][27] , 
        \w[9][26] , \w[9][25] , \w[9][24] , \w[9][23] , \w[9][22] , \w[9][21] , 
        \w[9][20] , \w[9][19] , \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , 
        \w[9][14] , \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , 
        \w[9][8] , \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , 
        \w[9][2] , \w[9][1] , 1'b0}), .CI(1'b0), .S({\w[10][31] , \w[10][30] , 
        \w[10][29] , \w[10][28] , \w[10][27] , \w[10][26] , \w[10][25] , 
        \w[10][24] , \w[10][23] , \w[10][22] , \w[10][21] , \w[10][20] , 
        \w[10][19] , \w[10][18] , \w[10][17] , \w[10][16] , \w[10][15] , 
        \w[10][14] , \w[10][13] , \w[10][12] , \w[10][11] , \w[10][10] , 
        \w[10][9] , \w[10][8] , \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , 
        \w[10][3] , \w[10][2] , \w[10][1] , SYNOPSYS_UNCONNECTED__8}) );
  ADD_N32_84 \FAINST[10].ADD_  ( .A({\_18_net_[31] , \_18_net_[30] , 
        \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] , 
        \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] , 
        \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] , 
        \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] , 
        \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] , \w[10][27] , 
        \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] , \w[10][22] , 
        \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] , \w[10][17] , 
        \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] , \w[10][12] , 
        \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] , \w[10][7] , 
        \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] , \w[10][2] , \w[10][1] , 
        1'b0}), .CI(1'b0), .S({\w[11][31] , \w[11][30] , \w[11][29] , 
        \w[11][28] , \w[11][27] , \w[11][26] , \w[11][25] , \w[11][24] , 
        \w[11][23] , \w[11][22] , \w[11][21] , \w[11][20] , \w[11][19] , 
        \w[11][18] , \w[11][17] , \w[11][16] , \w[11][15] , \w[11][14] , 
        \w[11][13] , \w[11][12] , \w[11][11] , \w[11][10] , \w[11][9] , 
        \w[11][8] , \w[11][7] , \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , 
        \w[11][2] , \w[11][1] , SYNOPSYS_UNCONNECTED__9}) );
  ADD_N32_83 \FAINST[11].ADD_  ( .A({\_20_net_[31] , \_20_net_[30] , 
        \_20_net_[29] , \_20_net_[28] , \_20_net_[27] , \_20_net_[26] , 
        \_20_net_[25] , \_20_net_[24] , \_20_net_[23] , \_20_net_[22] , 
        \_20_net_[21] , \_20_net_[20] , \_20_net_[19] , \_20_net_[18] , 
        \_20_net_[17] , \_20_net_[16] , \_20_net_[15] , \_20_net_[14] , 
        \_20_net_[13] , \_20_net_[12] , \_20_net_[11] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[11][31] , 
        \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] , \w[11][26] , 
        \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] , \w[11][21] , 
        \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] , \w[11][16] , 
        \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] , \w[11][11] , 
        \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] , \w[11][6] , 
        \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] , \w[11][1] , 1'b0}), 
        .CI(1'b0), .S({\w[12][31] , \w[12][30] , \w[12][29] , \w[12][28] , 
        \w[12][27] , \w[12][26] , \w[12][25] , \w[12][24] , \w[12][23] , 
        \w[12][22] , \w[12][21] , \w[12][20] , \w[12][19] , \w[12][18] , 
        \w[12][17] , \w[12][16] , \w[12][15] , \w[12][14] , \w[12][13] , 
        \w[12][12] , \w[12][11] , \w[12][10] , \w[12][9] , \w[12][8] , 
        \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , 
        \w[12][1] , SYNOPSYS_UNCONNECTED__10}) );
  ADD_N32_82 \FAINST[12].ADD_  ( .A({\_22_net_[31] , \_22_net_[30] , 
        \_22_net_[29] , \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , 
        \_22_net_[25] , \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , 
        \_22_net_[21] , \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , 
        \_22_net_[17] , \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , 
        \_22_net_[13] , \_22_net_[12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[12][31] , \w[12][30] , 
        \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] , \w[12][25] , 
        \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] , \w[12][20] , 
        \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] , \w[12][15] , 
        \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] , \w[12][10] , 
        \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , 
        \w[12][3] , \w[12][2] , \w[12][1] , 1'b0}), .CI(1'b0), .S({\w[13][31] , 
        \w[13][30] , \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , 
        \w[13][25] , \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , 
        \w[13][20] , \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , 
        \w[13][15] , \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , 
        \w[13][10] , \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , 
        \w[13][5] , \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , 
        SYNOPSYS_UNCONNECTED__11}) );
  ADD_N32_81 \FAINST[13].ADD_  ( .A({\_24_net_[31] , \_24_net_[30] , 
        \_24_net_[29] , \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , 
        \_24_net_[25] , \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , 
        \_24_net_[21] , \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , 
        \_24_net_[17] , \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , 
        \_24_net_[13] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[13][31] , \w[13][30] , \w[13][29] , 
        \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] , \w[13][24] , 
        \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] , \w[13][19] , 
        \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] , \w[13][14] , 
        \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] , \w[13][9] , 
        \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] , \w[13][4] , \w[13][3] , 
        \w[13][2] , \w[13][1] , 1'b0}), .CI(1'b0), .S({\w[14][31] , 
        \w[14][30] , \w[14][29] , \w[14][28] , \w[14][27] , \w[14][26] , 
        \w[14][25] , \w[14][24] , \w[14][23] , \w[14][22] , \w[14][21] , 
        \w[14][20] , \w[14][19] , \w[14][18] , \w[14][17] , \w[14][16] , 
        \w[14][15] , \w[14][14] , \w[14][13] , \w[14][12] , \w[14][11] , 
        \w[14][10] , \w[14][9] , \w[14][8] , \w[14][7] , \w[14][6] , 
        \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , \w[14][1] , 
        SYNOPSYS_UNCONNECTED__12}) );
  ADD_N32_80 \FAINST[14].ADD_  ( .A({\_26_net_[31] , \_26_net_[30] , 
        \_26_net_[29] , \_26_net_[28] , \_26_net_[27] , \_26_net_[26] , 
        \_26_net_[25] , \_26_net_[24] , \_26_net_[23] , \_26_net_[22] , 
        \_26_net_[21] , \_26_net_[20] , \_26_net_[19] , \_26_net_[18] , 
        \_26_net_[17] , \_26_net_[16] , \_26_net_[15] , \_26_net_[14] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[14][31] , \w[14][30] , \w[14][29] , \w[14][28] , 
        \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] , \w[14][23] , 
        \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] , \w[14][18] , 
        \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] , \w[14][13] , 
        \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] , \w[14][8] , 
        \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , 
        \w[14][1] , 1'b0}), .CI(1'b0), .S({\w[15][31] , \w[15][30] , 
        \w[15][29] , \w[15][28] , \w[15][27] , \w[15][26] , \w[15][25] , 
        \w[15][24] , \w[15][23] , \w[15][22] , \w[15][21] , \w[15][20] , 
        \w[15][19] , \w[15][18] , \w[15][17] , \w[15][16] , \w[15][15] , 
        \w[15][14] , \w[15][13] , \w[15][12] , \w[15][11] , \w[15][10] , 
        \w[15][9] , \w[15][8] , \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , 
        \w[15][3] , \w[15][2] , \w[15][1] , SYNOPSYS_UNCONNECTED__13}) );
  ADD_N32_79 \FAINST[15].ADD_  ( .A({\_28_net_[31] , \_28_net_[30] , 
        \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] , 
        \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] , 
        \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] , 
        \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] , \w[15][27] , 
        \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] , \w[15][22] , 
        \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] , \w[15][17] , 
        \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] , \w[15][12] , 
        \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] , \w[15][7] , 
        \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] , \w[15][2] , \w[15][1] , 
        1'b0}), .CI(1'b0), .S({\w[16][31] , \w[16][30] , \w[16][29] , 
        \w[16][28] , \w[16][27] , \w[16][26] , \w[16][25] , \w[16][24] , 
        \w[16][23] , \w[16][22] , \w[16][21] , \w[16][20] , \w[16][19] , 
        \w[16][18] , \w[16][17] , \w[16][16] , \w[16][15] , \w[16][14] , 
        \w[16][13] , \w[16][12] , \w[16][11] , \w[16][10] , \w[16][9] , 
        \w[16][8] , \w[16][7] , \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , 
        \w[16][2] , \w[16][1] , SYNOPSYS_UNCONNECTED__14}) );
  ADD_N32_78 \FAINST[16].ADD_  ( .A({\_30_net_[31] , \_30_net_[30] , 
        \_30_net_[29] , \_30_net_[28] , \_30_net_[27] , \_30_net_[26] , 
        \_30_net_[25] , \_30_net_[24] , \_30_net_[23] , \_30_net_[22] , 
        \_30_net_[21] , \_30_net_[20] , \_30_net_[19] , \_30_net_[18] , 
        \_30_net_[17] , \_30_net_[16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] , 
        \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] , 
        \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] , 
        \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] , 
        \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] , 
        \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] , \w[16][1] , 
        1'b0}), .CI(1'b0), .S({\w[17][31] , \w[17][30] , \w[17][29] , 
        \w[17][28] , \w[17][27] , \w[17][26] , \w[17][25] , \w[17][24] , 
        \w[17][23] , \w[17][22] , \w[17][21] , \w[17][20] , \w[17][19] , 
        \w[17][18] , \w[17][17] , \w[17][16] , \w[17][15] , \w[17][14] , 
        \w[17][13] , \w[17][12] , \w[17][11] , \w[17][10] , \w[17][9] , 
        \w[17][8] , \w[17][7] , \w[17][6] , \w[17][5] , \w[17][4] , \w[17][3] , 
        \w[17][2] , \w[17][1] , SYNOPSYS_UNCONNECTED__15}) );
  ADD_N32_77 \FAINST[17].ADD_  ( .A({\_32_net_[31] , \_32_net_[30] , 
        \_32_net_[29] , \_32_net_[28] , \_32_net_[27] , \_32_net_[26] , 
        \_32_net_[25] , \_32_net_[24] , \_32_net_[23] , \_32_net_[22] , 
        \_32_net_[21] , \_32_net_[20] , \_32_net_[19] , \_32_net_[18] , 
        \_32_net_[17] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[17][31] , 
        \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] , 
        \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] , 
        \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] , 
        \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] , 
        \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] , 
        \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] , 1'b0}), 
        .CI(1'b0), .S({\w[18][31] , \w[18][30] , \w[18][29] , \w[18][28] , 
        \w[18][27] , \w[18][26] , \w[18][25] , \w[18][24] , \w[18][23] , 
        \w[18][22] , \w[18][21] , \w[18][20] , \w[18][19] , \w[18][18] , 
        \w[18][17] , \w[18][16] , \w[18][15] , \w[18][14] , \w[18][13] , 
        \w[18][12] , \w[18][11] , \w[18][10] , \w[18][9] , \w[18][8] , 
        \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , \w[18][3] , \w[18][2] , 
        \w[18][1] , SYNOPSYS_UNCONNECTED__16}) );
  ADD_N32_76 \FAINST[18].ADD_  ( .A({\_34_net_[31] , \_34_net_[30] , 
        \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] , 
        \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] , 
        \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[18][31] , \w[18][30] , 
        \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] , 
        \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] , 
        \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] , 
        \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] , 
        \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , 
        \w[18][3] , \w[18][2] , \w[18][1] , 1'b0}), .CI(1'b0), .S({\w[19][31] , 
        \w[19][30] , \w[19][29] , \w[19][28] , \w[19][27] , \w[19][26] , 
        \w[19][25] , \w[19][24] , \w[19][23] , \w[19][22] , \w[19][21] , 
        \w[19][20] , \w[19][19] , \w[19][18] , \w[19][17] , \w[19][16] , 
        \w[19][15] , \w[19][14] , \w[19][13] , \w[19][12] , \w[19][11] , 
        \w[19][10] , \w[19][9] , \w[19][8] , \w[19][7] , \w[19][6] , 
        \w[19][5] , \w[19][4] , \w[19][3] , \w[19][2] , \w[19][1] , 
        SYNOPSYS_UNCONNECTED__17}) );
  ADD_N32_75 \FAINST[19].ADD_  ( .A({\_36_net_[31] , \_36_net_[30] , 
        \_36_net_[29] , \_36_net_[28] , \_36_net_[27] , \_36_net_[26] , 
        \_36_net_[25] , \_36_net_[24] , \_36_net_[23] , \_36_net_[22] , 
        \_36_net_[21] , \_36_net_[20] , \_36_net_[19] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[19][31] , \w[19][30] , \w[19][29] , 
        \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] , 
        \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] , 
        \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] , 
        \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] , 
        \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] , \w[19][3] , 
        \w[19][2] , \w[19][1] , 1'b0}), .CI(1'b0), .S({\w[20][31] , 
        \w[20][30] , \w[20][29] , \w[20][28] , \w[20][27] , \w[20][26] , 
        \w[20][25] , \w[20][24] , \w[20][23] , \w[20][22] , \w[20][21] , 
        \w[20][20] , \w[20][19] , \w[20][18] , \w[20][17] , \w[20][16] , 
        \w[20][15] , \w[20][14] , \w[20][13] , \w[20][12] , \w[20][11] , 
        \w[20][10] , \w[20][9] , \w[20][8] , \w[20][7] , \w[20][6] , 
        \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , \w[20][1] , 
        SYNOPSYS_UNCONNECTED__18}) );
  ADD_N32_74 \FAINST[20].ADD_  ( .A({\_38_net_[31] , \_38_net_[30] , 
        \_38_net_[29] , \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , 
        \_38_net_[25] , \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , 
        \_38_net_[21] , \_38_net_[20] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({\w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] , 
        \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] , 
        \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] , 
        \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] , 
        \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] , 
        \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , 
        \w[20][1] , 1'b0}), .CI(1'b0), .S({\w[21][31] , \w[21][30] , 
        \w[21][29] , \w[21][28] , \w[21][27] , \w[21][26] , \w[21][25] , 
        \w[21][24] , \w[21][23] , \w[21][22] , \w[21][21] , \w[21][20] , 
        \w[21][19] , \w[21][18] , \w[21][17] , \w[21][16] , \w[21][15] , 
        \w[21][14] , \w[21][13] , \w[21][12] , \w[21][11] , \w[21][10] , 
        \w[21][9] , \w[21][8] , \w[21][7] , \w[21][6] , \w[21][5] , \w[21][4] , 
        \w[21][3] , \w[21][2] , \w[21][1] , SYNOPSYS_UNCONNECTED__19}) );
  ADD_N32_73 \FAINST[21].ADD_  ( .A({\_40_net_[31] , \_40_net_[30] , 
        \_40_net_[29] , \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , 
        \_40_net_[25] , \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , 
        \_40_net_[21] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] , 
        \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] , 
        \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] , 
        \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] , 
        \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] , 
        \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] , \w[21][1] , 
        1'b0}), .CI(1'b0), .S({\w[22][31] , \w[22][30] , \w[22][29] , 
        \w[22][28] , \w[22][27] , \w[22][26] , \w[22][25] , \w[22][24] , 
        \w[22][23] , \w[22][22] , \w[22][21] , \w[22][20] , \w[22][19] , 
        \w[22][18] , \w[22][17] , \w[22][16] , \w[22][15] , \w[22][14] , 
        \w[22][13] , \w[22][12] , \w[22][11] , \w[22][10] , \w[22][9] , 
        \w[22][8] , \w[22][7] , \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , 
        \w[22][2] , \w[22][1] , SYNOPSYS_UNCONNECTED__20}) );
  ADD_N32_72 \FAINST[22].ADD_  ( .A({\_42_net_[31] , \_42_net_[30] , 
        \_42_net_[29] , \_42_net_[28] , \_42_net_[27] , \_42_net_[26] , 
        \_42_net_[25] , \_42_net_[24] , \_42_net_[23] , \_42_net_[22] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[22][31] , \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , 
        \w[22][26] , \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , 
        \w[22][21] , \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , 
        \w[22][16] , \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , 
        \w[22][11] , \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , 
        \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] , 
        1'b0}), .CI(1'b0), .S({\w[23][31] , \w[23][30] , \w[23][29] , 
        \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] , \w[23][24] , 
        \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] , \w[23][19] , 
        \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] , \w[23][14] , 
        \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] , \w[23][9] , 
        \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] , \w[23][4] , \w[23][3] , 
        \w[23][2] , \w[23][1] , SYNOPSYS_UNCONNECTED__21}) );
  ADD_N32_71 \FAINST[23].ADD_  ( .A({\_44_net_[31] , \_44_net_[30] , 
        \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] , 
        \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[23][31] , 
        \w[23][30] , \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , 
        \w[23][25] , \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , 
        \w[23][20] , \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , 
        \w[23][15] , \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , 
        \w[23][10] , \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , 
        \w[23][5] , \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , 1'b0}), 
        .CI(1'b0), .S({\w[24][31] , \w[24][30] , \w[24][29] , \w[24][28] , 
        \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] , \w[24][23] , 
        \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] , \w[24][18] , 
        \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] , \w[24][13] , 
        \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] , \w[24][8] , 
        \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , \w[24][3] , \w[24][2] , 
        \w[24][1] , SYNOPSYS_UNCONNECTED__22}) );
  ADD_N32_70 \FAINST[24].ADD_  ( .A({\_46_net_[31] , \_46_net_[30] , 
        \_46_net_[29] , \_46_net_[28] , \_46_net_[27] , \_46_net_[26] , 
        \_46_net_[25] , \_46_net_[24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[24][31] , \w[24][30] , 
        \w[24][29] , \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , 
        \w[24][24] , \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , 
        \w[24][19] , \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , 
        \w[24][14] , \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , 
        \w[24][9] , \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , 
        \w[24][3] , \w[24][2] , \w[24][1] , 1'b0}), .CI(1'b0), .S({\w[25][31] , 
        \w[25][30] , \w[25][29] , \w[25][28] , \w[25][27] , \w[25][26] , 
        \w[25][25] , \w[25][24] , \w[25][23] , \w[25][22] , \w[25][21] , 
        \w[25][20] , \w[25][19] , \w[25][18] , \w[25][17] , \w[25][16] , 
        \w[25][15] , \w[25][14] , \w[25][13] , \w[25][12] , \w[25][11] , 
        \w[25][10] , \w[25][9] , \w[25][8] , \w[25][7] , \w[25][6] , 
        \w[25][5] , \w[25][4] , \w[25][3] , \w[25][2] , \w[25][1] , 
        SYNOPSYS_UNCONNECTED__23}) );
  ADD_N32_69 \FAINST[25].ADD_  ( .A({\_48_net_[31] , \_48_net_[30] , 
        \_48_net_[29] , \_48_net_[28] , \_48_net_[27] , \_48_net_[26] , 
        \_48_net_[25] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[25][31] , \w[25][30] , \w[25][29] , 
        \w[25][28] , \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , 
        \w[25][23] , \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , 
        \w[25][18] , \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , 
        \w[25][13] , \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , 
        \w[25][8] , \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] , 
        \w[25][2] , \w[25][1] , 1'b0}), .CI(1'b0), .S({\w[26][31] , 
        \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] , \w[26][26] , 
        \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] , \w[26][21] , 
        \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] , \w[26][16] , 
        \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] , \w[26][11] , 
        \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] , \w[26][6] , 
        \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , \w[26][1] , 
        SYNOPSYS_UNCONNECTED__24}) );
  ADD_N32_68 \FAINST[26].ADD_  ( .A({\_50_net_[31] , \_50_net_[30] , 
        \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , 
        \w[26][27] , \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , 
        \w[26][22] , \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , 
        \w[26][17] , \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , 
        \w[26][12] , \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , 
        \w[26][7] , \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , 
        \w[26][1] , 1'b0}), .CI(1'b0), .S({\w[27][31] , \w[27][30] , 
        \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] , \w[27][25] , 
        \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] , \w[27][20] , 
        \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] , \w[27][15] , 
        \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] , \w[27][10] , 
        \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] , \w[27][5] , \w[27][4] , 
        \w[27][3] , \w[27][2] , \w[27][1] , SYNOPSYS_UNCONNECTED__25}) );
  ADD_N32_67 \FAINST[27].ADD_  ( .A({\_52_net_[31] , \_52_net_[30] , 
        \_52_net_[29] , \_52_net_[28] , \_52_net_[27] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[27][31] , \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , 
        \w[27][26] , \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , 
        \w[27][21] , \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , 
        \w[27][16] , \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , 
        \w[27][11] , \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , 
        \w[27][6] , \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] , 
        1'b0}), .CI(1'b0), .S({\w[28][31] , \w[28][30] , \w[28][29] , 
        \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] , \w[28][24] , 
        \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] , \w[28][19] , 
        \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] , \w[28][14] , 
        \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] , \w[28][9] , 
        \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , 
        \w[28][2] , \w[28][1] , SYNOPSYS_UNCONNECTED__26}) );
  ADD_N32_66 \FAINST[28].ADD_  ( .A({\_54_net_[31] , \_54_net_[30] , 
        \_54_net_[29] , \_54_net_[28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[28][31] , \w[28][30] , \w[28][29] , \w[28][28] , \w[28][27] , 
        \w[28][26] , \w[28][25] , \w[28][24] , \w[28][23] , \w[28][22] , 
        \w[28][21] , \w[28][20] , \w[28][19] , \w[28][18] , \w[28][17] , 
        \w[28][16] , \w[28][15] , \w[28][14] , \w[28][13] , \w[28][12] , 
        \w[28][11] , \w[28][10] , \w[28][9] , \w[28][8] , \w[28][7] , 
        \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , 
        1'b0}), .CI(1'b0), .S({\w[29][31] , \w[29][30] , \w[29][29] , 
        \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] , 
        \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] , 
        \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] , 
        \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] , 
        \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] , \w[29][3] , 
        \w[29][2] , \w[29][1] , SYNOPSYS_UNCONNECTED__27}) );
  ADD_N32_65 \FAINST[29].ADD_  ( .A({\_56_net_[31] , \_56_net_[30] , 
        \_56_net_[29] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[29][31] , 
        \w[29][30] , \w[29][29] , \w[29][28] , \w[29][27] , \w[29][26] , 
        \w[29][25] , \w[29][24] , \w[29][23] , \w[29][22] , \w[29][21] , 
        \w[29][20] , \w[29][19] , \w[29][18] , \w[29][17] , \w[29][16] , 
        \w[29][15] , \w[29][14] , \w[29][13] , \w[29][12] , \w[29][11] , 
        \w[29][10] , \w[29][9] , \w[29][8] , \w[29][7] , \w[29][6] , 
        \w[29][5] , \w[29][4] , \w[29][3] , \w[29][2] , \w[29][1] , 1'b0}), 
        .CI(1'b0), .S({\w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] , 
        \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] , 
        \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] , 
        \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] , 
        \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] , 
        \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] , \w[30][2] , 
        \w[30][1] , SYNOPSYS_UNCONNECTED__28}) );
  ADD_N32_64 \FAINST[30].ADD_  ( .A({\_58_net_[31] , \_58_net_[30] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[30][31] , \w[30][30] , 
        \w[30][29] , \w[30][28] , \w[30][27] , \w[30][26] , \w[30][25] , 
        \w[30][24] , \w[30][23] , \w[30][22] , \w[30][21] , \w[30][20] , 
        \w[30][19] , \w[30][18] , \w[30][17] , \w[30][16] , \w[30][15] , 
        \w[30][14] , \w[30][13] , \w[30][12] , \w[30][11] , \w[30][10] , 
        \w[30][9] , \w[30][8] , \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , 
        \w[30][3] , \w[30][2] , \w[30][1] , 1'b0}), .CI(1'b0), .S({\w[31][31] , 
        \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] , \w[31][26] , 
        \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] , \w[31][21] , 
        \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] , \w[31][16] , 
        \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] , \w[31][11] , 
        \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] , \w[31][6] , 
        \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] , \w[31][1] , 
        SYNOPSYS_UNCONNECTED__29}) );
  ADD_N32_63 \FAINST[31].ADD_  ( .A({\_60_net_[31] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[31][31] , \w[31][30] , \w[31][29] , 
        \w[31][28] , \w[31][27] , \w[31][26] , \w[31][25] , \w[31][24] , 
        \w[31][23] , \w[31][22] , \w[31][21] , \w[31][20] , \w[31][19] , 
        \w[31][18] , \w[31][17] , \w[31][16] , \w[31][15] , \w[31][14] , 
        \w[31][13] , \w[31][12] , \w[31][11] , \w[31][10] , \w[31][9] , 
        \w[31][8] , \w[31][7] , \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , 
        \w[31][2] , \w[31][1] , 1'b0}), .CI(1'b0), .S({O[31:1], 
        SYNOPSYS_UNCONNECTED__30}) );
  AND U2 ( .A(A[5]), .B(B[4]), .Z(\_8_net_[9] ) );
  AND U3 ( .A(A[5]), .B(B[3]), .Z(\_8_net_[8] ) );
  AND U4 ( .A(A[5]), .B(B[2]), .Z(\_8_net_[7] ) );
  AND U5 ( .A(A[5]), .B(B[1]), .Z(\_8_net_[6] ) );
  AND U6 ( .A(A[5]), .B(B[0]), .Z(\_8_net_[5] ) );
  AND U7 ( .A(A[5]), .B(B[26]), .Z(\_8_net_[31] ) );
  AND U8 ( .A(A[5]), .B(B[25]), .Z(\_8_net_[30] ) );
  AND U9 ( .A(A[5]), .B(B[24]), .Z(\_8_net_[29] ) );
  AND U10 ( .A(A[5]), .B(B[23]), .Z(\_8_net_[28] ) );
  AND U11 ( .A(A[5]), .B(B[22]), .Z(\_8_net_[27] ) );
  AND U12 ( .A(A[5]), .B(B[21]), .Z(\_8_net_[26] ) );
  AND U13 ( .A(A[5]), .B(B[20]), .Z(\_8_net_[25] ) );
  AND U14 ( .A(A[5]), .B(B[19]), .Z(\_8_net_[24] ) );
  AND U15 ( .A(A[5]), .B(B[18]), .Z(\_8_net_[23] ) );
  AND U16 ( .A(A[5]), .B(B[17]), .Z(\_8_net_[22] ) );
  AND U17 ( .A(A[5]), .B(B[16]), .Z(\_8_net_[21] ) );
  AND U18 ( .A(A[5]), .B(B[15]), .Z(\_8_net_[20] ) );
  AND U19 ( .A(A[5]), .B(B[14]), .Z(\_8_net_[19] ) );
  AND U20 ( .A(A[5]), .B(B[13]), .Z(\_8_net_[18] ) );
  AND U21 ( .A(A[5]), .B(B[12]), .Z(\_8_net_[17] ) );
  AND U22 ( .A(A[5]), .B(B[11]), .Z(\_8_net_[16] ) );
  AND U23 ( .A(A[5]), .B(B[10]), .Z(\_8_net_[15] ) );
  AND U24 ( .A(A[5]), .B(B[9]), .Z(\_8_net_[14] ) );
  AND U25 ( .A(A[5]), .B(B[8]), .Z(\_8_net_[13] ) );
  AND U26 ( .A(A[5]), .B(B[7]), .Z(\_8_net_[12] ) );
  AND U27 ( .A(A[5]), .B(B[6]), .Z(\_8_net_[11] ) );
  AND U28 ( .A(A[5]), .B(B[5]), .Z(\_8_net_[10] ) );
  AND U29 ( .A(B[5]), .B(A[4]), .Z(\_6_net_[9] ) );
  AND U30 ( .A(B[4]), .B(A[4]), .Z(\_6_net_[8] ) );
  AND U31 ( .A(B[3]), .B(A[4]), .Z(\_6_net_[7] ) );
  AND U32 ( .A(B[2]), .B(A[4]), .Z(\_6_net_[6] ) );
  AND U33 ( .A(B[1]), .B(A[4]), .Z(\_6_net_[5] ) );
  AND U34 ( .A(B[0]), .B(A[4]), .Z(\_6_net_[4] ) );
  AND U35 ( .A(A[4]), .B(B[27]), .Z(\_6_net_[31] ) );
  AND U36 ( .A(B[26]), .B(A[4]), .Z(\_6_net_[30] ) );
  AND U37 ( .A(B[25]), .B(A[4]), .Z(\_6_net_[29] ) );
  AND U38 ( .A(B[24]), .B(A[4]), .Z(\_6_net_[28] ) );
  AND U39 ( .A(B[23]), .B(A[4]), .Z(\_6_net_[27] ) );
  AND U40 ( .A(B[22]), .B(A[4]), .Z(\_6_net_[26] ) );
  AND U41 ( .A(B[21]), .B(A[4]), .Z(\_6_net_[25] ) );
  AND U42 ( .A(B[20]), .B(A[4]), .Z(\_6_net_[24] ) );
  AND U43 ( .A(B[19]), .B(A[4]), .Z(\_6_net_[23] ) );
  AND U44 ( .A(B[18]), .B(A[4]), .Z(\_6_net_[22] ) );
  AND U45 ( .A(B[17]), .B(A[4]), .Z(\_6_net_[21] ) );
  AND U46 ( .A(B[16]), .B(A[4]), .Z(\_6_net_[20] ) );
  AND U47 ( .A(B[15]), .B(A[4]), .Z(\_6_net_[19] ) );
  AND U48 ( .A(B[14]), .B(A[4]), .Z(\_6_net_[18] ) );
  AND U49 ( .A(B[13]), .B(A[4]), .Z(\_6_net_[17] ) );
  AND U50 ( .A(B[12]), .B(A[4]), .Z(\_6_net_[16] ) );
  AND U51 ( .A(B[11]), .B(A[4]), .Z(\_6_net_[15] ) );
  AND U52 ( .A(B[10]), .B(A[4]), .Z(\_6_net_[14] ) );
  AND U53 ( .A(B[9]), .B(A[4]), .Z(\_6_net_[13] ) );
  AND U54 ( .A(B[8]), .B(A[4]), .Z(\_6_net_[12] ) );
  AND U55 ( .A(B[7]), .B(A[4]), .Z(\_6_net_[11] ) );
  AND U56 ( .A(B[6]), .B(A[4]), .Z(\_6_net_[10] ) );
  AND U57 ( .A(A[31]), .B(B[0]), .Z(\_60_net_[31] ) );
  AND U58 ( .A(B[1]), .B(A[30]), .Z(\_58_net_[31] ) );
  AND U59 ( .A(A[30]), .B(B[0]), .Z(\_58_net_[30] ) );
  AND U60 ( .A(B[2]), .B(A[29]), .Z(\_56_net_[31] ) );
  AND U61 ( .A(B[1]), .B(A[29]), .Z(\_56_net_[30] ) );
  AND U62 ( .A(A[29]), .B(B[0]), .Z(\_56_net_[29] ) );
  AND U63 ( .A(B[3]), .B(A[28]), .Z(\_54_net_[31] ) );
  AND U64 ( .A(B[2]), .B(A[28]), .Z(\_54_net_[30] ) );
  AND U65 ( .A(B[1]), .B(A[28]), .Z(\_54_net_[29] ) );
  AND U66 ( .A(A[28]), .B(B[0]), .Z(\_54_net_[28] ) );
  AND U67 ( .A(B[4]), .B(A[27]), .Z(\_52_net_[31] ) );
  AND U68 ( .A(B[3]), .B(A[27]), .Z(\_52_net_[30] ) );
  AND U69 ( .A(B[2]), .B(A[27]), .Z(\_52_net_[29] ) );
  AND U70 ( .A(B[1]), .B(A[27]), .Z(\_52_net_[28] ) );
  AND U71 ( .A(A[27]), .B(B[0]), .Z(\_52_net_[27] ) );
  AND U72 ( .A(B[5]), .B(A[26]), .Z(\_50_net_[31] ) );
  AND U73 ( .A(B[4]), .B(A[26]), .Z(\_50_net_[30] ) );
  AND U74 ( .A(B[3]), .B(A[26]), .Z(\_50_net_[29] ) );
  AND U75 ( .A(B[2]), .B(A[26]), .Z(\_50_net_[28] ) );
  AND U76 ( .A(B[1]), .B(A[26]), .Z(\_50_net_[27] ) );
  AND U77 ( .A(A[26]), .B(B[0]), .Z(\_50_net_[26] ) );
  AND U78 ( .A(B[6]), .B(A[3]), .Z(\_4_net_[9] ) );
  AND U79 ( .A(B[5]), .B(A[3]), .Z(\_4_net_[8] ) );
  AND U80 ( .A(B[4]), .B(A[3]), .Z(\_4_net_[7] ) );
  AND U81 ( .A(B[3]), .B(A[3]), .Z(\_4_net_[6] ) );
  AND U82 ( .A(B[2]), .B(A[3]), .Z(\_4_net_[5] ) );
  AND U83 ( .A(B[1]), .B(A[3]), .Z(\_4_net_[4] ) );
  AND U84 ( .A(B[0]), .B(A[3]), .Z(\_4_net_[3] ) );
  AND U85 ( .A(A[3]), .B(B[28]), .Z(\_4_net_[31] ) );
  AND U86 ( .A(B[27]), .B(A[3]), .Z(\_4_net_[30] ) );
  AND U87 ( .A(B[26]), .B(A[3]), .Z(\_4_net_[29] ) );
  AND U88 ( .A(B[25]), .B(A[3]), .Z(\_4_net_[28] ) );
  AND U89 ( .A(B[24]), .B(A[3]), .Z(\_4_net_[27] ) );
  AND U90 ( .A(B[23]), .B(A[3]), .Z(\_4_net_[26] ) );
  AND U91 ( .A(B[22]), .B(A[3]), .Z(\_4_net_[25] ) );
  AND U92 ( .A(B[21]), .B(A[3]), .Z(\_4_net_[24] ) );
  AND U93 ( .A(B[20]), .B(A[3]), .Z(\_4_net_[23] ) );
  AND U94 ( .A(B[19]), .B(A[3]), .Z(\_4_net_[22] ) );
  AND U95 ( .A(B[18]), .B(A[3]), .Z(\_4_net_[21] ) );
  AND U96 ( .A(B[17]), .B(A[3]), .Z(\_4_net_[20] ) );
  AND U97 ( .A(B[16]), .B(A[3]), .Z(\_4_net_[19] ) );
  AND U98 ( .A(B[15]), .B(A[3]), .Z(\_4_net_[18] ) );
  AND U99 ( .A(B[14]), .B(A[3]), .Z(\_4_net_[17] ) );
  AND U100 ( .A(B[13]), .B(A[3]), .Z(\_4_net_[16] ) );
  AND U101 ( .A(B[12]), .B(A[3]), .Z(\_4_net_[15] ) );
  AND U102 ( .A(B[11]), .B(A[3]), .Z(\_4_net_[14] ) );
  AND U103 ( .A(B[10]), .B(A[3]), .Z(\_4_net_[13] ) );
  AND U104 ( .A(B[9]), .B(A[3]), .Z(\_4_net_[12] ) );
  AND U105 ( .A(B[8]), .B(A[3]), .Z(\_4_net_[11] ) );
  AND U106 ( .A(B[7]), .B(A[3]), .Z(\_4_net_[10] ) );
  AND U107 ( .A(B[6]), .B(A[25]), .Z(\_48_net_[31] ) );
  AND U108 ( .A(B[5]), .B(A[25]), .Z(\_48_net_[30] ) );
  AND U109 ( .A(B[4]), .B(A[25]), .Z(\_48_net_[29] ) );
  AND U110 ( .A(B[3]), .B(A[25]), .Z(\_48_net_[28] ) );
  AND U111 ( .A(B[2]), .B(A[25]), .Z(\_48_net_[27] ) );
  AND U112 ( .A(B[1]), .B(A[25]), .Z(\_48_net_[26] ) );
  AND U113 ( .A(A[25]), .B(B[0]), .Z(\_48_net_[25] ) );
  AND U114 ( .A(B[7]), .B(A[24]), .Z(\_46_net_[31] ) );
  AND U115 ( .A(B[6]), .B(A[24]), .Z(\_46_net_[30] ) );
  AND U116 ( .A(B[5]), .B(A[24]), .Z(\_46_net_[29] ) );
  AND U117 ( .A(B[4]), .B(A[24]), .Z(\_46_net_[28] ) );
  AND U118 ( .A(B[3]), .B(A[24]), .Z(\_46_net_[27] ) );
  AND U119 ( .A(B[2]), .B(A[24]), .Z(\_46_net_[26] ) );
  AND U120 ( .A(B[1]), .B(A[24]), .Z(\_46_net_[25] ) );
  AND U121 ( .A(A[24]), .B(B[0]), .Z(\_46_net_[24] ) );
  AND U122 ( .A(B[8]), .B(A[23]), .Z(\_44_net_[31] ) );
  AND U123 ( .A(B[7]), .B(A[23]), .Z(\_44_net_[30] ) );
  AND U124 ( .A(B[6]), .B(A[23]), .Z(\_44_net_[29] ) );
  AND U125 ( .A(B[5]), .B(A[23]), .Z(\_44_net_[28] ) );
  AND U126 ( .A(B[4]), .B(A[23]), .Z(\_44_net_[27] ) );
  AND U127 ( .A(B[3]), .B(A[23]), .Z(\_44_net_[26] ) );
  AND U128 ( .A(B[2]), .B(A[23]), .Z(\_44_net_[25] ) );
  AND U129 ( .A(B[1]), .B(A[23]), .Z(\_44_net_[24] ) );
  AND U130 ( .A(A[23]), .B(B[0]), .Z(\_44_net_[23] ) );
  AND U131 ( .A(B[9]), .B(A[22]), .Z(\_42_net_[31] ) );
  AND U132 ( .A(B[8]), .B(A[22]), .Z(\_42_net_[30] ) );
  AND U133 ( .A(B[7]), .B(A[22]), .Z(\_42_net_[29] ) );
  AND U134 ( .A(B[6]), .B(A[22]), .Z(\_42_net_[28] ) );
  AND U135 ( .A(B[5]), .B(A[22]), .Z(\_42_net_[27] ) );
  AND U136 ( .A(B[4]), .B(A[22]), .Z(\_42_net_[26] ) );
  AND U137 ( .A(B[3]), .B(A[22]), .Z(\_42_net_[25] ) );
  AND U138 ( .A(B[2]), .B(A[22]), .Z(\_42_net_[24] ) );
  AND U139 ( .A(B[1]), .B(A[22]), .Z(\_42_net_[23] ) );
  AND U140 ( .A(A[22]), .B(B[0]), .Z(\_42_net_[22] ) );
  AND U141 ( .A(B[10]), .B(A[21]), .Z(\_40_net_[31] ) );
  AND U142 ( .A(B[9]), .B(A[21]), .Z(\_40_net_[30] ) );
  AND U143 ( .A(B[8]), .B(A[21]), .Z(\_40_net_[29] ) );
  AND U144 ( .A(B[7]), .B(A[21]), .Z(\_40_net_[28] ) );
  AND U145 ( .A(B[6]), .B(A[21]), .Z(\_40_net_[27] ) );
  AND U146 ( .A(B[5]), .B(A[21]), .Z(\_40_net_[26] ) );
  AND U147 ( .A(B[4]), .B(A[21]), .Z(\_40_net_[25] ) );
  AND U148 ( .A(B[3]), .B(A[21]), .Z(\_40_net_[24] ) );
  AND U149 ( .A(B[2]), .B(A[21]), .Z(\_40_net_[23] ) );
  AND U150 ( .A(B[1]), .B(A[21]), .Z(\_40_net_[22] ) );
  AND U151 ( .A(A[21]), .B(B[0]), .Z(\_40_net_[21] ) );
  AND U152 ( .A(B[11]), .B(A[20]), .Z(\_38_net_[31] ) );
  AND U153 ( .A(B[10]), .B(A[20]), .Z(\_38_net_[30] ) );
  AND U154 ( .A(B[9]), .B(A[20]), .Z(\_38_net_[29] ) );
  AND U155 ( .A(B[8]), .B(A[20]), .Z(\_38_net_[28] ) );
  AND U156 ( .A(B[7]), .B(A[20]), .Z(\_38_net_[27] ) );
  AND U157 ( .A(B[6]), .B(A[20]), .Z(\_38_net_[26] ) );
  AND U158 ( .A(B[5]), .B(A[20]), .Z(\_38_net_[25] ) );
  AND U159 ( .A(B[4]), .B(A[20]), .Z(\_38_net_[24] ) );
  AND U160 ( .A(B[3]), .B(A[20]), .Z(\_38_net_[23] ) );
  AND U161 ( .A(B[2]), .B(A[20]), .Z(\_38_net_[22] ) );
  AND U162 ( .A(B[1]), .B(A[20]), .Z(\_38_net_[21] ) );
  AND U163 ( .A(A[20]), .B(B[0]), .Z(\_38_net_[20] ) );
  AND U164 ( .A(B[12]), .B(A[19]), .Z(\_36_net_[31] ) );
  AND U165 ( .A(B[11]), .B(A[19]), .Z(\_36_net_[30] ) );
  AND U166 ( .A(B[10]), .B(A[19]), .Z(\_36_net_[29] ) );
  AND U167 ( .A(B[9]), .B(A[19]), .Z(\_36_net_[28] ) );
  AND U168 ( .A(B[8]), .B(A[19]), .Z(\_36_net_[27] ) );
  AND U169 ( .A(B[7]), .B(A[19]), .Z(\_36_net_[26] ) );
  AND U170 ( .A(B[6]), .B(A[19]), .Z(\_36_net_[25] ) );
  AND U171 ( .A(B[5]), .B(A[19]), .Z(\_36_net_[24] ) );
  AND U172 ( .A(B[4]), .B(A[19]), .Z(\_36_net_[23] ) );
  AND U173 ( .A(B[3]), .B(A[19]), .Z(\_36_net_[22] ) );
  AND U174 ( .A(B[2]), .B(A[19]), .Z(\_36_net_[21] ) );
  AND U175 ( .A(B[1]), .B(A[19]), .Z(\_36_net_[20] ) );
  AND U176 ( .A(A[19]), .B(B[0]), .Z(\_36_net_[19] ) );
  AND U177 ( .A(B[13]), .B(A[18]), .Z(\_34_net_[31] ) );
  AND U178 ( .A(B[12]), .B(A[18]), .Z(\_34_net_[30] ) );
  AND U179 ( .A(B[11]), .B(A[18]), .Z(\_34_net_[29] ) );
  AND U180 ( .A(B[10]), .B(A[18]), .Z(\_34_net_[28] ) );
  AND U181 ( .A(B[9]), .B(A[18]), .Z(\_34_net_[27] ) );
  AND U182 ( .A(B[8]), .B(A[18]), .Z(\_34_net_[26] ) );
  AND U183 ( .A(B[7]), .B(A[18]), .Z(\_34_net_[25] ) );
  AND U184 ( .A(B[6]), .B(A[18]), .Z(\_34_net_[24] ) );
  AND U185 ( .A(B[5]), .B(A[18]), .Z(\_34_net_[23] ) );
  AND U186 ( .A(B[4]), .B(A[18]), .Z(\_34_net_[22] ) );
  AND U187 ( .A(B[3]), .B(A[18]), .Z(\_34_net_[21] ) );
  AND U188 ( .A(B[2]), .B(A[18]), .Z(\_34_net_[20] ) );
  AND U189 ( .A(B[1]), .B(A[18]), .Z(\_34_net_[19] ) );
  AND U190 ( .A(A[18]), .B(B[0]), .Z(\_34_net_[18] ) );
  AND U191 ( .A(B[14]), .B(A[17]), .Z(\_32_net_[31] ) );
  AND U192 ( .A(B[13]), .B(A[17]), .Z(\_32_net_[30] ) );
  AND U193 ( .A(B[12]), .B(A[17]), .Z(\_32_net_[29] ) );
  AND U194 ( .A(B[11]), .B(A[17]), .Z(\_32_net_[28] ) );
  AND U195 ( .A(B[10]), .B(A[17]), .Z(\_32_net_[27] ) );
  AND U196 ( .A(B[9]), .B(A[17]), .Z(\_32_net_[26] ) );
  AND U197 ( .A(B[8]), .B(A[17]), .Z(\_32_net_[25] ) );
  AND U198 ( .A(B[7]), .B(A[17]), .Z(\_32_net_[24] ) );
  AND U199 ( .A(B[6]), .B(A[17]), .Z(\_32_net_[23] ) );
  AND U200 ( .A(B[5]), .B(A[17]), .Z(\_32_net_[22] ) );
  AND U201 ( .A(B[4]), .B(A[17]), .Z(\_32_net_[21] ) );
  AND U202 ( .A(B[3]), .B(A[17]), .Z(\_32_net_[20] ) );
  AND U203 ( .A(B[2]), .B(A[17]), .Z(\_32_net_[19] ) );
  AND U204 ( .A(B[1]), .B(A[17]), .Z(\_32_net_[18] ) );
  AND U205 ( .A(A[17]), .B(B[0]), .Z(\_32_net_[17] ) );
  AND U206 ( .A(B[15]), .B(A[16]), .Z(\_30_net_[31] ) );
  AND U207 ( .A(B[14]), .B(A[16]), .Z(\_30_net_[30] ) );
  AND U208 ( .A(B[13]), .B(A[16]), .Z(\_30_net_[29] ) );
  AND U209 ( .A(B[12]), .B(A[16]), .Z(\_30_net_[28] ) );
  AND U210 ( .A(B[11]), .B(A[16]), .Z(\_30_net_[27] ) );
  AND U211 ( .A(B[10]), .B(A[16]), .Z(\_30_net_[26] ) );
  AND U212 ( .A(B[9]), .B(A[16]), .Z(\_30_net_[25] ) );
  AND U213 ( .A(B[8]), .B(A[16]), .Z(\_30_net_[24] ) );
  AND U214 ( .A(B[7]), .B(A[16]), .Z(\_30_net_[23] ) );
  AND U215 ( .A(B[6]), .B(A[16]), .Z(\_30_net_[22] ) );
  AND U216 ( .A(B[5]), .B(A[16]), .Z(\_30_net_[21] ) );
  AND U217 ( .A(B[4]), .B(A[16]), .Z(\_30_net_[20] ) );
  AND U218 ( .A(B[3]), .B(A[16]), .Z(\_30_net_[19] ) );
  AND U219 ( .A(B[2]), .B(A[16]), .Z(\_30_net_[18] ) );
  AND U220 ( .A(B[1]), .B(A[16]), .Z(\_30_net_[17] ) );
  AND U221 ( .A(A[16]), .B(B[0]), .Z(\_30_net_[16] ) );
  AND U222 ( .A(B[7]), .B(A[2]), .Z(\_2_net_[9] ) );
  AND U223 ( .A(B[6]), .B(A[2]), .Z(\_2_net_[8] ) );
  AND U224 ( .A(B[5]), .B(A[2]), .Z(\_2_net_[7] ) );
  AND U225 ( .A(B[4]), .B(A[2]), .Z(\_2_net_[6] ) );
  AND U226 ( .A(B[3]), .B(A[2]), .Z(\_2_net_[5] ) );
  AND U227 ( .A(B[2]), .B(A[2]), .Z(\_2_net_[4] ) );
  AND U228 ( .A(B[1]), .B(A[2]), .Z(\_2_net_[3] ) );
  AND U229 ( .A(A[2]), .B(B[29]), .Z(\_2_net_[31] ) );
  AND U230 ( .A(B[28]), .B(A[2]), .Z(\_2_net_[30] ) );
  AND U231 ( .A(B[0]), .B(A[2]), .Z(\_2_net_[2] ) );
  AND U232 ( .A(B[27]), .B(A[2]), .Z(\_2_net_[29] ) );
  AND U233 ( .A(B[26]), .B(A[2]), .Z(\_2_net_[28] ) );
  AND U234 ( .A(B[25]), .B(A[2]), .Z(\_2_net_[27] ) );
  AND U235 ( .A(B[24]), .B(A[2]), .Z(\_2_net_[26] ) );
  AND U236 ( .A(B[23]), .B(A[2]), .Z(\_2_net_[25] ) );
  AND U237 ( .A(B[22]), .B(A[2]), .Z(\_2_net_[24] ) );
  AND U238 ( .A(B[21]), .B(A[2]), .Z(\_2_net_[23] ) );
  AND U239 ( .A(B[20]), .B(A[2]), .Z(\_2_net_[22] ) );
  AND U240 ( .A(B[19]), .B(A[2]), .Z(\_2_net_[21] ) );
  AND U241 ( .A(B[18]), .B(A[2]), .Z(\_2_net_[20] ) );
  AND U242 ( .A(B[17]), .B(A[2]), .Z(\_2_net_[19] ) );
  AND U243 ( .A(B[16]), .B(A[2]), .Z(\_2_net_[18] ) );
  AND U244 ( .A(B[15]), .B(A[2]), .Z(\_2_net_[17] ) );
  AND U245 ( .A(B[14]), .B(A[2]), .Z(\_2_net_[16] ) );
  AND U246 ( .A(B[13]), .B(A[2]), .Z(\_2_net_[15] ) );
  AND U247 ( .A(B[12]), .B(A[2]), .Z(\_2_net_[14] ) );
  AND U248 ( .A(B[11]), .B(A[2]), .Z(\_2_net_[13] ) );
  AND U249 ( .A(B[10]), .B(A[2]), .Z(\_2_net_[12] ) );
  AND U250 ( .A(B[9]), .B(A[2]), .Z(\_2_net_[11] ) );
  AND U251 ( .A(B[8]), .B(A[2]), .Z(\_2_net_[10] ) );
  AND U252 ( .A(B[16]), .B(A[15]), .Z(\_28_net_[31] ) );
  AND U253 ( .A(B[15]), .B(A[15]), .Z(\_28_net_[30] ) );
  AND U254 ( .A(B[14]), .B(A[15]), .Z(\_28_net_[29] ) );
  AND U255 ( .A(B[13]), .B(A[15]), .Z(\_28_net_[28] ) );
  AND U256 ( .A(B[12]), .B(A[15]), .Z(\_28_net_[27] ) );
  AND U257 ( .A(B[11]), .B(A[15]), .Z(\_28_net_[26] ) );
  AND U258 ( .A(B[10]), .B(A[15]), .Z(\_28_net_[25] ) );
  AND U259 ( .A(B[9]), .B(A[15]), .Z(\_28_net_[24] ) );
  AND U260 ( .A(B[8]), .B(A[15]), .Z(\_28_net_[23] ) );
  AND U261 ( .A(B[7]), .B(A[15]), .Z(\_28_net_[22] ) );
  AND U262 ( .A(B[6]), .B(A[15]), .Z(\_28_net_[21] ) );
  AND U263 ( .A(B[5]), .B(A[15]), .Z(\_28_net_[20] ) );
  AND U264 ( .A(B[4]), .B(A[15]), .Z(\_28_net_[19] ) );
  AND U265 ( .A(B[3]), .B(A[15]), .Z(\_28_net_[18] ) );
  AND U266 ( .A(B[2]), .B(A[15]), .Z(\_28_net_[17] ) );
  AND U267 ( .A(B[1]), .B(A[15]), .Z(\_28_net_[16] ) );
  AND U268 ( .A(A[15]), .B(B[0]), .Z(\_28_net_[15] ) );
  AND U269 ( .A(B[17]), .B(A[14]), .Z(\_26_net_[31] ) );
  AND U270 ( .A(B[16]), .B(A[14]), .Z(\_26_net_[30] ) );
  AND U271 ( .A(B[15]), .B(A[14]), .Z(\_26_net_[29] ) );
  AND U272 ( .A(B[14]), .B(A[14]), .Z(\_26_net_[28] ) );
  AND U273 ( .A(B[13]), .B(A[14]), .Z(\_26_net_[27] ) );
  AND U274 ( .A(B[12]), .B(A[14]), .Z(\_26_net_[26] ) );
  AND U275 ( .A(B[11]), .B(A[14]), .Z(\_26_net_[25] ) );
  AND U276 ( .A(B[10]), .B(A[14]), .Z(\_26_net_[24] ) );
  AND U277 ( .A(B[9]), .B(A[14]), .Z(\_26_net_[23] ) );
  AND U278 ( .A(B[8]), .B(A[14]), .Z(\_26_net_[22] ) );
  AND U279 ( .A(B[7]), .B(A[14]), .Z(\_26_net_[21] ) );
  AND U280 ( .A(B[6]), .B(A[14]), .Z(\_26_net_[20] ) );
  AND U281 ( .A(B[5]), .B(A[14]), .Z(\_26_net_[19] ) );
  AND U282 ( .A(B[4]), .B(A[14]), .Z(\_26_net_[18] ) );
  AND U283 ( .A(B[3]), .B(A[14]), .Z(\_26_net_[17] ) );
  AND U284 ( .A(B[2]), .B(A[14]), .Z(\_26_net_[16] ) );
  AND U285 ( .A(B[1]), .B(A[14]), .Z(\_26_net_[15] ) );
  AND U286 ( .A(A[14]), .B(B[0]), .Z(\_26_net_[14] ) );
  AND U287 ( .A(B[18]), .B(A[13]), .Z(\_24_net_[31] ) );
  AND U288 ( .A(B[17]), .B(A[13]), .Z(\_24_net_[30] ) );
  AND U289 ( .A(B[16]), .B(A[13]), .Z(\_24_net_[29] ) );
  AND U290 ( .A(B[15]), .B(A[13]), .Z(\_24_net_[28] ) );
  AND U291 ( .A(B[14]), .B(A[13]), .Z(\_24_net_[27] ) );
  AND U292 ( .A(B[13]), .B(A[13]), .Z(\_24_net_[26] ) );
  AND U293 ( .A(B[12]), .B(A[13]), .Z(\_24_net_[25] ) );
  AND U294 ( .A(B[11]), .B(A[13]), .Z(\_24_net_[24] ) );
  AND U295 ( .A(B[10]), .B(A[13]), .Z(\_24_net_[23] ) );
  AND U296 ( .A(B[9]), .B(A[13]), .Z(\_24_net_[22] ) );
  AND U297 ( .A(B[8]), .B(A[13]), .Z(\_24_net_[21] ) );
  AND U298 ( .A(B[7]), .B(A[13]), .Z(\_24_net_[20] ) );
  AND U299 ( .A(B[6]), .B(A[13]), .Z(\_24_net_[19] ) );
  AND U300 ( .A(B[5]), .B(A[13]), .Z(\_24_net_[18] ) );
  AND U301 ( .A(B[4]), .B(A[13]), .Z(\_24_net_[17] ) );
  AND U302 ( .A(B[3]), .B(A[13]), .Z(\_24_net_[16] ) );
  AND U303 ( .A(B[2]), .B(A[13]), .Z(\_24_net_[15] ) );
  AND U304 ( .A(B[1]), .B(A[13]), .Z(\_24_net_[14] ) );
  AND U305 ( .A(A[13]), .B(B[0]), .Z(\_24_net_[13] ) );
  AND U306 ( .A(B[19]), .B(A[12]), .Z(\_22_net_[31] ) );
  AND U307 ( .A(B[18]), .B(A[12]), .Z(\_22_net_[30] ) );
  AND U308 ( .A(B[17]), .B(A[12]), .Z(\_22_net_[29] ) );
  AND U309 ( .A(B[16]), .B(A[12]), .Z(\_22_net_[28] ) );
  AND U310 ( .A(B[15]), .B(A[12]), .Z(\_22_net_[27] ) );
  AND U311 ( .A(B[14]), .B(A[12]), .Z(\_22_net_[26] ) );
  AND U312 ( .A(B[13]), .B(A[12]), .Z(\_22_net_[25] ) );
  AND U313 ( .A(B[12]), .B(A[12]), .Z(\_22_net_[24] ) );
  AND U314 ( .A(B[11]), .B(A[12]), .Z(\_22_net_[23] ) );
  AND U315 ( .A(B[10]), .B(A[12]), .Z(\_22_net_[22] ) );
  AND U316 ( .A(B[9]), .B(A[12]), .Z(\_22_net_[21] ) );
  AND U317 ( .A(B[8]), .B(A[12]), .Z(\_22_net_[20] ) );
  AND U318 ( .A(B[7]), .B(A[12]), .Z(\_22_net_[19] ) );
  AND U319 ( .A(B[6]), .B(A[12]), .Z(\_22_net_[18] ) );
  AND U320 ( .A(B[5]), .B(A[12]), .Z(\_22_net_[17] ) );
  AND U321 ( .A(B[4]), .B(A[12]), .Z(\_22_net_[16] ) );
  AND U322 ( .A(B[3]), .B(A[12]), .Z(\_22_net_[15] ) );
  AND U323 ( .A(B[2]), .B(A[12]), .Z(\_22_net_[14] ) );
  AND U324 ( .A(B[1]), .B(A[12]), .Z(\_22_net_[13] ) );
  AND U325 ( .A(A[12]), .B(B[0]), .Z(\_22_net_[12] ) );
  AND U326 ( .A(B[20]), .B(A[11]), .Z(\_20_net_[31] ) );
  AND U327 ( .A(B[19]), .B(A[11]), .Z(\_20_net_[30] ) );
  AND U328 ( .A(B[18]), .B(A[11]), .Z(\_20_net_[29] ) );
  AND U329 ( .A(B[17]), .B(A[11]), .Z(\_20_net_[28] ) );
  AND U330 ( .A(B[16]), .B(A[11]), .Z(\_20_net_[27] ) );
  AND U331 ( .A(B[15]), .B(A[11]), .Z(\_20_net_[26] ) );
  AND U332 ( .A(B[14]), .B(A[11]), .Z(\_20_net_[25] ) );
  AND U333 ( .A(B[13]), .B(A[11]), .Z(\_20_net_[24] ) );
  AND U334 ( .A(B[12]), .B(A[11]), .Z(\_20_net_[23] ) );
  AND U335 ( .A(B[11]), .B(A[11]), .Z(\_20_net_[22] ) );
  AND U336 ( .A(B[10]), .B(A[11]), .Z(\_20_net_[21] ) );
  AND U337 ( .A(B[9]), .B(A[11]), .Z(\_20_net_[20] ) );
  AND U338 ( .A(B[8]), .B(A[11]), .Z(\_20_net_[19] ) );
  AND U339 ( .A(B[7]), .B(A[11]), .Z(\_20_net_[18] ) );
  AND U340 ( .A(B[6]), .B(A[11]), .Z(\_20_net_[17] ) );
  AND U341 ( .A(B[5]), .B(A[11]), .Z(\_20_net_[16] ) );
  AND U342 ( .A(B[4]), .B(A[11]), .Z(\_20_net_[15] ) );
  AND U343 ( .A(B[3]), .B(A[11]), .Z(\_20_net_[14] ) );
  AND U344 ( .A(B[2]), .B(A[11]), .Z(\_20_net_[13] ) );
  AND U345 ( .A(B[1]), .B(A[11]), .Z(\_20_net_[12] ) );
  AND U346 ( .A(A[11]), .B(B[0]), .Z(\_20_net_[11] ) );
  AND U347 ( .A(B[21]), .B(A[10]), .Z(\_18_net_[31] ) );
  AND U348 ( .A(B[20]), .B(A[10]), .Z(\_18_net_[30] ) );
  AND U349 ( .A(B[19]), .B(A[10]), .Z(\_18_net_[29] ) );
  AND U350 ( .A(B[18]), .B(A[10]), .Z(\_18_net_[28] ) );
  AND U351 ( .A(B[17]), .B(A[10]), .Z(\_18_net_[27] ) );
  AND U352 ( .A(B[16]), .B(A[10]), .Z(\_18_net_[26] ) );
  AND U353 ( .A(B[15]), .B(A[10]), .Z(\_18_net_[25] ) );
  AND U354 ( .A(B[14]), .B(A[10]), .Z(\_18_net_[24] ) );
  AND U355 ( .A(B[13]), .B(A[10]), .Z(\_18_net_[23] ) );
  AND U356 ( .A(B[12]), .B(A[10]), .Z(\_18_net_[22] ) );
  AND U357 ( .A(B[11]), .B(A[10]), .Z(\_18_net_[21] ) );
  AND U358 ( .A(B[10]), .B(A[10]), .Z(\_18_net_[20] ) );
  AND U359 ( .A(B[9]), .B(A[10]), .Z(\_18_net_[19] ) );
  AND U360 ( .A(B[8]), .B(A[10]), .Z(\_18_net_[18] ) );
  AND U361 ( .A(B[7]), .B(A[10]), .Z(\_18_net_[17] ) );
  AND U362 ( .A(B[6]), .B(A[10]), .Z(\_18_net_[16] ) );
  AND U363 ( .A(B[5]), .B(A[10]), .Z(\_18_net_[15] ) );
  AND U364 ( .A(B[4]), .B(A[10]), .Z(\_18_net_[14] ) );
  AND U365 ( .A(B[3]), .B(A[10]), .Z(\_18_net_[13] ) );
  AND U366 ( .A(B[2]), .B(A[10]), .Z(\_18_net_[12] ) );
  AND U367 ( .A(B[1]), .B(A[10]), .Z(\_18_net_[11] ) );
  AND U368 ( .A(A[10]), .B(B[0]), .Z(\_18_net_[10] ) );
  AND U369 ( .A(B[0]), .B(A[9]), .Z(\_16_net_[9] ) );
  AND U370 ( .A(B[22]), .B(A[9]), .Z(\_16_net_[31] ) );
  AND U371 ( .A(B[21]), .B(A[9]), .Z(\_16_net_[30] ) );
  AND U372 ( .A(B[20]), .B(A[9]), .Z(\_16_net_[29] ) );
  AND U373 ( .A(B[19]), .B(A[9]), .Z(\_16_net_[28] ) );
  AND U374 ( .A(B[18]), .B(A[9]), .Z(\_16_net_[27] ) );
  AND U375 ( .A(B[17]), .B(A[9]), .Z(\_16_net_[26] ) );
  AND U376 ( .A(B[16]), .B(A[9]), .Z(\_16_net_[25] ) );
  AND U377 ( .A(B[15]), .B(A[9]), .Z(\_16_net_[24] ) );
  AND U378 ( .A(B[14]), .B(A[9]), .Z(\_16_net_[23] ) );
  AND U379 ( .A(B[13]), .B(A[9]), .Z(\_16_net_[22] ) );
  AND U380 ( .A(B[12]), .B(A[9]), .Z(\_16_net_[21] ) );
  AND U381 ( .A(B[11]), .B(A[9]), .Z(\_16_net_[20] ) );
  AND U382 ( .A(B[10]), .B(A[9]), .Z(\_16_net_[19] ) );
  AND U383 ( .A(B[9]), .B(A[9]), .Z(\_16_net_[18] ) );
  AND U384 ( .A(B[8]), .B(A[9]), .Z(\_16_net_[17] ) );
  AND U385 ( .A(B[7]), .B(A[9]), .Z(\_16_net_[16] ) );
  AND U386 ( .A(B[6]), .B(A[9]), .Z(\_16_net_[15] ) );
  AND U387 ( .A(B[5]), .B(A[9]), .Z(\_16_net_[14] ) );
  AND U388 ( .A(B[4]), .B(A[9]), .Z(\_16_net_[13] ) );
  AND U389 ( .A(B[3]), .B(A[9]), .Z(\_16_net_[12] ) );
  AND U390 ( .A(B[2]), .B(A[9]), .Z(\_16_net_[11] ) );
  AND U391 ( .A(A[9]), .B(B[1]), .Z(\_16_net_[10] ) );
  AND U392 ( .A(B[1]), .B(A[8]), .Z(\_14_net_[9] ) );
  AND U393 ( .A(B[0]), .B(A[8]), .Z(\_14_net_[8] ) );
  AND U394 ( .A(B[23]), .B(A[8]), .Z(\_14_net_[31] ) );
  AND U395 ( .A(B[22]), .B(A[8]), .Z(\_14_net_[30] ) );
  AND U396 ( .A(B[21]), .B(A[8]), .Z(\_14_net_[29] ) );
  AND U397 ( .A(B[20]), .B(A[8]), .Z(\_14_net_[28] ) );
  AND U398 ( .A(B[19]), .B(A[8]), .Z(\_14_net_[27] ) );
  AND U399 ( .A(B[18]), .B(A[8]), .Z(\_14_net_[26] ) );
  AND U400 ( .A(B[17]), .B(A[8]), .Z(\_14_net_[25] ) );
  AND U401 ( .A(B[16]), .B(A[8]), .Z(\_14_net_[24] ) );
  AND U402 ( .A(B[15]), .B(A[8]), .Z(\_14_net_[23] ) );
  AND U403 ( .A(B[14]), .B(A[8]), .Z(\_14_net_[22] ) );
  AND U404 ( .A(B[13]), .B(A[8]), .Z(\_14_net_[21] ) );
  AND U405 ( .A(B[12]), .B(A[8]), .Z(\_14_net_[20] ) );
  AND U406 ( .A(B[11]), .B(A[8]), .Z(\_14_net_[19] ) );
  AND U407 ( .A(B[10]), .B(A[8]), .Z(\_14_net_[18] ) );
  AND U408 ( .A(B[9]), .B(A[8]), .Z(\_14_net_[17] ) );
  AND U409 ( .A(B[8]), .B(A[8]), .Z(\_14_net_[16] ) );
  AND U410 ( .A(B[7]), .B(A[8]), .Z(\_14_net_[15] ) );
  AND U411 ( .A(B[6]), .B(A[8]), .Z(\_14_net_[14] ) );
  AND U412 ( .A(B[5]), .B(A[8]), .Z(\_14_net_[13] ) );
  AND U413 ( .A(B[4]), .B(A[8]), .Z(\_14_net_[12] ) );
  AND U414 ( .A(B[3]), .B(A[8]), .Z(\_14_net_[11] ) );
  AND U415 ( .A(A[8]), .B(B[2]), .Z(\_14_net_[10] ) );
  AND U416 ( .A(B[2]), .B(A[7]), .Z(\_12_net_[9] ) );
  AND U417 ( .A(B[1]), .B(A[7]), .Z(\_12_net_[8] ) );
  AND U418 ( .A(B[0]), .B(A[7]), .Z(\_12_net_[7] ) );
  AND U419 ( .A(B[24]), .B(A[7]), .Z(\_12_net_[31] ) );
  AND U420 ( .A(B[23]), .B(A[7]), .Z(\_12_net_[30] ) );
  AND U421 ( .A(B[22]), .B(A[7]), .Z(\_12_net_[29] ) );
  AND U422 ( .A(B[21]), .B(A[7]), .Z(\_12_net_[28] ) );
  AND U423 ( .A(B[20]), .B(A[7]), .Z(\_12_net_[27] ) );
  AND U424 ( .A(B[19]), .B(A[7]), .Z(\_12_net_[26] ) );
  AND U425 ( .A(B[18]), .B(A[7]), .Z(\_12_net_[25] ) );
  AND U426 ( .A(B[17]), .B(A[7]), .Z(\_12_net_[24] ) );
  AND U427 ( .A(B[16]), .B(A[7]), .Z(\_12_net_[23] ) );
  AND U428 ( .A(B[15]), .B(A[7]), .Z(\_12_net_[22] ) );
  AND U429 ( .A(B[14]), .B(A[7]), .Z(\_12_net_[21] ) );
  AND U430 ( .A(B[13]), .B(A[7]), .Z(\_12_net_[20] ) );
  AND U431 ( .A(B[12]), .B(A[7]), .Z(\_12_net_[19] ) );
  AND U432 ( .A(B[11]), .B(A[7]), .Z(\_12_net_[18] ) );
  AND U433 ( .A(B[10]), .B(A[7]), .Z(\_12_net_[17] ) );
  AND U434 ( .A(B[9]), .B(A[7]), .Z(\_12_net_[16] ) );
  AND U435 ( .A(B[8]), .B(A[7]), .Z(\_12_net_[15] ) );
  AND U436 ( .A(B[7]), .B(A[7]), .Z(\_12_net_[14] ) );
  AND U437 ( .A(B[6]), .B(A[7]), .Z(\_12_net_[13] ) );
  AND U438 ( .A(B[5]), .B(A[7]), .Z(\_12_net_[12] ) );
  AND U439 ( .A(B[4]), .B(A[7]), .Z(\_12_net_[11] ) );
  AND U440 ( .A(A[7]), .B(B[3]), .Z(\_12_net_[10] ) );
  AND U441 ( .A(B[3]), .B(A[6]), .Z(\_10_net_[9] ) );
  AND U442 ( .A(B[2]), .B(A[6]), .Z(\_10_net_[8] ) );
  AND U443 ( .A(B[1]), .B(A[6]), .Z(\_10_net_[7] ) );
  AND U444 ( .A(B[0]), .B(A[6]), .Z(\_10_net_[6] ) );
  AND U445 ( .A(B[25]), .B(A[6]), .Z(\_10_net_[31] ) );
  AND U446 ( .A(B[24]), .B(A[6]), .Z(\_10_net_[30] ) );
  AND U447 ( .A(B[23]), .B(A[6]), .Z(\_10_net_[29] ) );
  AND U448 ( .A(B[22]), .B(A[6]), .Z(\_10_net_[28] ) );
  AND U449 ( .A(B[21]), .B(A[6]), .Z(\_10_net_[27] ) );
  AND U450 ( .A(B[20]), .B(A[6]), .Z(\_10_net_[26] ) );
  AND U451 ( .A(B[19]), .B(A[6]), .Z(\_10_net_[25] ) );
  AND U452 ( .A(B[18]), .B(A[6]), .Z(\_10_net_[24] ) );
  AND U453 ( .A(B[17]), .B(A[6]), .Z(\_10_net_[23] ) );
  AND U454 ( .A(B[16]), .B(A[6]), .Z(\_10_net_[22] ) );
  AND U455 ( .A(B[15]), .B(A[6]), .Z(\_10_net_[21] ) );
  AND U456 ( .A(B[14]), .B(A[6]), .Z(\_10_net_[20] ) );
  AND U457 ( .A(B[13]), .B(A[6]), .Z(\_10_net_[19] ) );
  AND U458 ( .A(B[12]), .B(A[6]), .Z(\_10_net_[18] ) );
  AND U459 ( .A(B[11]), .B(A[6]), .Z(\_10_net_[17] ) );
  AND U460 ( .A(B[10]), .B(A[6]), .Z(\_10_net_[16] ) );
  AND U461 ( .A(B[9]), .B(A[6]), .Z(\_10_net_[15] ) );
  AND U462 ( .A(B[8]), .B(A[6]), .Z(\_10_net_[14] ) );
  AND U463 ( .A(B[7]), .B(A[6]), .Z(\_10_net_[13] ) );
  AND U464 ( .A(B[6]), .B(A[6]), .Z(\_10_net_[12] ) );
  AND U465 ( .A(B[5]), .B(A[6]), .Z(\_10_net_[11] ) );
  AND U466 ( .A(A[6]), .B(B[4]), .Z(\_10_net_[10] ) );
  AND U467 ( .A(B[8]), .B(A[1]), .Z(\_0_net_[9] ) );
  AND U468 ( .A(B[7]), .B(A[1]), .Z(\_0_net_[8] ) );
  AND U469 ( .A(B[6]), .B(A[1]), .Z(\_0_net_[7] ) );
  AND U470 ( .A(B[5]), .B(A[1]), .Z(\_0_net_[6] ) );
  AND U471 ( .A(B[4]), .B(A[1]), .Z(\_0_net_[5] ) );
  AND U472 ( .A(B[3]), .B(A[1]), .Z(\_0_net_[4] ) );
  AND U473 ( .A(B[2]), .B(A[1]), .Z(\_0_net_[3] ) );
  AND U474 ( .A(B[30]), .B(A[1]), .Z(\_0_net_[31] ) );
  AND U475 ( .A(B[29]), .B(A[1]), .Z(\_0_net_[30] ) );
  AND U476 ( .A(B[1]), .B(A[1]), .Z(\_0_net_[2] ) );
  AND U477 ( .A(B[28]), .B(A[1]), .Z(\_0_net_[29] ) );
  AND U478 ( .A(B[27]), .B(A[1]), .Z(\_0_net_[28] ) );
  AND U479 ( .A(B[26]), .B(A[1]), .Z(\_0_net_[27] ) );
  AND U480 ( .A(B[25]), .B(A[1]), .Z(\_0_net_[26] ) );
  AND U481 ( .A(B[24]), .B(A[1]), .Z(\_0_net_[25] ) );
  AND U482 ( .A(B[23]), .B(A[1]), .Z(\_0_net_[24] ) );
  AND U483 ( .A(B[22]), .B(A[1]), .Z(\_0_net_[23] ) );
  AND U484 ( .A(B[21]), .B(A[1]), .Z(\_0_net_[22] ) );
  AND U485 ( .A(B[20]), .B(A[1]), .Z(\_0_net_[21] ) );
  AND U486 ( .A(B[19]), .B(A[1]), .Z(\_0_net_[20] ) );
  AND U487 ( .A(B[0]), .B(A[1]), .Z(\_0_net_[1] ) );
  AND U488 ( .A(B[18]), .B(A[1]), .Z(\_0_net_[19] ) );
  AND U489 ( .A(B[17]), .B(A[1]), .Z(\_0_net_[18] ) );
  AND U490 ( .A(B[16]), .B(A[1]), .Z(\_0_net_[17] ) );
  AND U491 ( .A(B[15]), .B(A[1]), .Z(\_0_net_[16] ) );
  AND U492 ( .A(B[14]), .B(A[1]), .Z(\_0_net_[15] ) );
  AND U493 ( .A(B[13]), .B(A[1]), .Z(\_0_net_[14] ) );
  AND U494 ( .A(B[12]), .B(A[1]), .Z(\_0_net_[13] ) );
  AND U495 ( .A(B[11]), .B(A[1]), .Z(\_0_net_[12] ) );
  AND U496 ( .A(B[10]), .B(A[1]), .Z(\_0_net_[11] ) );
  AND U497 ( .A(A[1]), .B(B[9]), .Z(\_0_net_[10] ) );
endmodule


module FA_3041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N32_0 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3071 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_3070 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_3069 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_3068 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_3067 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_3066 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3065 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3064 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3063 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3062 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3061 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3060 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3059 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3058 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3057 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3056 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3055 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3054 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3053 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3052 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3051 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3050 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3049 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3048 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3047 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3046 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3045 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3044 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3043 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3042 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3041 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_2 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_4 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_6 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_7 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_8 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_9 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_10 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_11 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_12 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_13 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_14 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_15 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_16 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_17 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_18 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_19 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_20 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_21 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_22 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_23 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_24 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_25 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_26 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_27 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_28 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_29 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_30 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_31 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_1 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_31 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_30 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_29 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_28 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_27 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_26 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_25 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_24 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_23 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_22 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_21 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_20 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_19 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_18 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_17 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_16 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_15 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_14 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_13 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_12 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_11 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_10 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_9 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_8 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_7 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_6 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_5 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_4 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_3 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_2 \FAINST[30].FA_  ( .A(1'b0), .B(B[30]), .CI(1'b0), .S(S[30]) );
  FA_1 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(1'b0), .S(S[31]) );
endmodule


module FA_33 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_34 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_35 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_36 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_37 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_38 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_39 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_40 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_41 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_42 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_43 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_44 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_45 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_46 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_47 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_48 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_49 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_50 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_51 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_52 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_53 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_54 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_55 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_56 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_57 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_58 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_59 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_60 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_61 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_62 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_63 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_2 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;
  wire   \C[31] ;

  FA_63 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_62 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_61 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_60 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_59 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_58 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_57 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_56 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_55 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_54 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_53 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_52 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_51 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_50 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_49 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_48 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_47 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_46 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_45 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_44 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_43 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_42 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_41 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_40 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_39 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_38 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_37 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_36 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_35 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_34 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(1'b0), .S(S[30]), .CO(
        \C[31] ) );
  FA_33 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(\C[31] ), .S(S[31]) );
endmodule


module FA_65 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_66 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_67 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_68 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_69 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_70 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_71 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_72 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_73 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_74 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_75 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_76 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_77 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_78 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_79 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_80 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_81 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_82 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_83 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_84 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_85 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_86 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_87 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_88 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_89 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_90 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_91 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_92 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_93 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_94 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_95 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_3 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_95 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_94 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_93 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_92 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_91 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_90 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_89 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_88 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_87 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_86 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_85 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_84 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_83 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_82 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_81 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_80 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_79 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_78 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_77 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_76 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_75 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_74 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_73 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_72 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_71 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_70 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_69 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_68 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_67 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(1'b0), .S(S[29]), .CO(
        C[30]) );
  FA_66 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_65 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_97 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_98 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_99 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_4 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_127 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_126 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_125 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_124 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_123 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_122 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_121 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_120 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_119 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_118 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_117 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_116 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_115 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_114 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_113 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_112 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_111 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_110 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_109 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_108 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_107 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_106 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_105 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_104 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_103 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_102 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_101 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_100 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(1'b0), .S(S[28]), .CO(
        C[29]) );
  FA_99 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_98 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_97 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_5 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_159 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_158 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_157 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_156 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_155 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_154 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_153 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_152 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_151 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_150 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_149 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_148 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_147 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_146 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_145 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_144 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_143 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_142 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_141 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_140 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_139 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_138 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_137 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_136 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_135 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_134 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_133 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(1'b0), .S(S[27]), .CO(
        C[28]) );
  FA_132 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_131 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_130 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_129 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_6 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_191 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_190 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_189 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_188 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_187 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_186 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_185 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_184 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_183 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_182 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_181 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_180 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_179 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_178 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_177 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_176 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_175 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_174 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_173 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_172 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_171 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_170 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_169 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_168 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_167 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_166 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(1'b0), .S(S[26]), .CO(
        C[27]) );
  FA_165 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_164 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_163 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_162 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_161 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_7 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_223 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_222 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_221 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_220 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_219 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_218 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_217 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_216 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_215 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_214 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_213 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_212 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_211 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_210 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_209 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_208 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_207 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_206 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_205 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_204 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_203 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_202 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_201 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_200 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_199 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(1'b0), .S(S[25]), .CO(
        C[26]) );
  FA_198 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_197 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_196 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_195 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_194 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_193 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_8 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_255 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_254 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_253 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_252 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_251 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_250 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_249 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_248 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_247 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_246 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_245 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_244 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_243 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_242 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_241 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_240 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_239 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_238 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_237 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_236 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_235 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_234 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_233 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_232 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(1'b0), .S(S[24]), .CO(
        C[25]) );
  FA_231 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_230 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_229 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_228 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_227 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_226 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_225 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_9 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_287 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_286 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_285 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_284 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_283 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_282 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_281 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_280 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_279 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_278 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_277 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_276 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_275 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_274 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_273 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_272 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_271 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_270 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_269 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_268 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_267 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_266 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_265 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(1'b0), .S(S[23]), .CO(
        C[24]) );
  FA_264 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_263 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_262 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_261 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_260 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_259 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_258 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_257 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_10 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_319 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_318 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_317 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_316 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_315 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_314 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_313 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_312 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_311 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_310 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_309 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_308 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_307 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_306 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_305 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_304 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_303 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_302 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_301 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_300 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_299 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_298 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(1'b0), .S(S[22]), .CO(
        C[23]) );
  FA_297 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_296 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_295 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_294 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_293 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_292 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_291 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_290 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_289 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_11 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_351 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_350 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_349 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_348 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_347 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_346 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_345 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_344 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_343 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_342 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_341 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_340 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_339 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_338 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_337 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_336 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_335 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_334 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_333 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_332 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_331 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(1'b0), .S(S[21]), .CO(
        C[22]) );
  FA_330 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_329 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_328 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_327 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_326 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_325 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_324 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_323 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_322 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_321 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_12 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_383 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_382 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_381 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_380 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_379 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_378 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_377 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_376 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_375 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_374 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_373 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_372 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_371 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_370 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_369 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_368 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_367 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_366 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_365 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_364 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(1'b0), .S(S[20]), .CO(
        C[21]) );
  FA_363 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_362 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_361 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_360 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_359 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_358 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_357 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_356 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_355 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_354 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_353 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_13 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_415 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_414 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_413 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_412 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_411 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_410 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_409 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_408 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_407 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_406 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_405 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_404 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_403 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_402 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_401 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_400 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_399 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_398 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_397 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(1'b0), .S(S[19]), .CO(
        C[20]) );
  FA_396 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_395 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_394 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_393 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_392 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_391 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_390 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_389 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_388 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_387 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_386 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_385 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_14 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_447 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_446 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_445 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_444 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_443 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_442 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_441 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_440 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_439 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_438 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_437 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_436 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_435 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_434 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_433 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_432 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_431 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_430 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(1'b0), .S(S[18]), .CO(
        C[19]) );
  FA_429 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_428 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_427 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_426 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_425 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_424 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_423 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_422 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_421 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_420 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_419 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_418 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_417 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_15 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_479 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_478 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_477 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_476 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_475 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_474 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_473 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_472 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_471 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_470 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_469 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_468 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_467 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_466 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_465 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_464 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_463 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(1'b0), .S(S[17]), .CO(
        C[18]) );
  FA_462 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_461 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_460 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_459 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_458 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_457 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_456 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_455 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_454 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_453 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_452 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_451 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_450 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_449 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_16 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_511 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_510 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_509 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_508 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_507 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_506 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_505 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_504 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_503 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_502 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_501 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_500 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_499 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_498 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_497 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_496 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(1'b0), .S(S[16]), .CO(
        C[17]) );
  FA_495 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_494 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_493 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_492 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_491 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_490 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_489 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_488 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_487 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_486 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_485 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_484 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_483 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_482 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_481 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_17 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_543 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_542 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_541 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_540 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_539 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_538 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_537 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_536 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_535 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_534 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_533 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_532 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_531 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_530 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_529 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(1'b0), .S(S[15]), .CO(
        C[16]) );
  FA_528 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_527 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_526 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_525 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_524 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_523 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_522 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_521 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_520 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_519 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_518 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_517 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_516 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_515 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_514 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_513 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_18 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_575 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_574 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_573 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_572 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_571 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_570 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_569 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_568 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_567 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_566 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_565 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_564 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_563 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_562 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(1'b0), .S(S[14]), .CO(
        C[15]) );
  FA_561 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_560 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_559 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_558 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_557 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_556 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_555 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_554 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_553 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_552 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_551 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_550 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_549 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_548 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_547 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_546 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_545 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_19 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_607 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_606 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_605 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_604 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_603 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_602 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_601 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_600 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_599 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_598 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_597 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_596 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_595 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(1'b0), .S(S[13]), .CO(
        C[14]) );
  FA_594 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_593 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_592 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_591 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_590 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_589 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_588 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_587 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_586 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_585 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_584 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_583 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_582 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_581 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_580 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_579 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_578 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_577 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_20 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_639 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_638 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_637 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_636 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_635 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_634 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_633 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_632 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_631 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_630 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_629 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_628 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(1'b0), .S(S[12]), .CO(
        C[13]) );
  FA_627 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_626 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_625 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_624 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_623 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_622 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_621 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_620 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_619 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_618 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_617 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_616 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_615 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_614 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_613 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_612 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_611 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_610 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_609 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_21 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_671 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_670 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_669 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_668 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_667 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_666 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_665 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_664 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_663 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_662 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_661 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(1'b0), .S(S[11]), .CO(
        C[12]) );
  FA_660 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_659 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_658 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_657 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_656 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_655 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_654 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_653 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_652 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_651 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_650 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_649 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_648 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_647 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_646 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_645 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_644 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_643 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_642 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_641 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_22 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_703 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_702 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_701 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_700 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_699 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_698 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_697 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_696 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_695 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_694 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(1'b0), .S(S[10]), .CO(
        C[11]) );
  FA_693 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_692 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_691 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_690 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_689 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_688 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_687 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_686 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_685 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_684 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_683 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_682 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_681 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_680 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_679 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_678 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_677 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_676 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_675 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_674 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_673 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_23 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_735 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_734 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_733 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_732 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_731 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_730 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_729 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_728 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_727 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(1'b0), .S(S[9]), .CO(C[10])
         );
  FA_726 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_725 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_724 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_723 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_722 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_721 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_720 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_719 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_718 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_717 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_716 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_715 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_714 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_713 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_712 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_711 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_710 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_709 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_708 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_707 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_706 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_705 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_24 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_767 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_766 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_765 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_764 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_763 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_762 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_761 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_760 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(1'b0), .S(S[8]), .CO(C[9])
         );
  FA_759 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10])
         );
  FA_758 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_757 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_756 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_755 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_754 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_753 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_752 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_751 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_750 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_749 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_748 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_747 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_746 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_745 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_744 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_743 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_742 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_741 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_740 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_739 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_738 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_737 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_25 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_799 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_798 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_797 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_796 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_795 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_794 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_793 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(1'b0), .S(S[7]), .CO(C[8])
         );
  FA_792 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_791 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10])
         );
  FA_790 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_789 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_788 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_787 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_786 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_785 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_784 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_783 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_782 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_781 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_780 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_779 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_778 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_777 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_776 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_775 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_774 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_773 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_772 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_771 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_770 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_769 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_26 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_831 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_830 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_829 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_828 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_827 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_826 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(1'b0), .S(S[6]), .CO(C[7])
         );
  FA_825 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_824 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_823 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10])
         );
  FA_822 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_821 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_820 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_819 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_818 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_817 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_816 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_815 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_814 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_813 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_812 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_811 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_810 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_809 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_808 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_807 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_806 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_805 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_804 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_803 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_802 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_801 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_27 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_863 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_862 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_861 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_860 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_859 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(1'b0), .S(S[5]), .CO(C[6])
         );
  FA_858 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_857 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_856 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_855 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10])
         );
  FA_854 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_853 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_852 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_851 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_850 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_849 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_848 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_847 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_846 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_845 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_844 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_843 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_842 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_841 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_840 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_839 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_838 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_837 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_836 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_835 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_834 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_833 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_28 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_895 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_894 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_893 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_892 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(1'b0), .S(S[4]), .CO(C[5])
         );
  FA_891 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_890 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_889 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_888 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_887 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10])
         );
  FA_886 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_885 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_884 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_883 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_882 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_881 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_880 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_879 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_878 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_877 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_876 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_875 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_874 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_873 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_872 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_871 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_870 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_869 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_868 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_867 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_866 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_865 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_29 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_927 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_926 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_925 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(1'b0), .S(S[3]), .CO(C[4])
         );
  FA_924 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_923 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_922 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_921 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_920 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_919 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10])
         );
  FA_918 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_917 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_916 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_915 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_914 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_913 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_912 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_911 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_910 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_909 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_908 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_907 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_906 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_905 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_904 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_903 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_902 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_901 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_900 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_899 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_898 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_897 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_30 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_959 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_958 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(1'b0), .S(S[2]), .CO(C[3])
         );
  FA_957 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_956 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_955 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_954 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_953 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_952 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_951 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10])
         );
  FA_950 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_949 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_948 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_947 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_946 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_945 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_944 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_943 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_942 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_941 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_940 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_939 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_938 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_937 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_936 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_935 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_934 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_933 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_932 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_931 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_930 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_929 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module ADD_N32_31 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_991 \FAINST[1].FA_  ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(S[1]) );
  FA_990 \FAINST[2].FA_  ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(S[2]) );
  FA_989 \FAINST[3].FA_  ( .A(A[3]), .B(1'b0), .CI(1'b0), .S(S[3]) );
  FA_988 \FAINST[4].FA_  ( .A(A[4]), .B(1'b0), .CI(1'b0), .S(S[4]) );
  FA_987 \FAINST[5].FA_  ( .A(A[5]), .B(1'b0), .CI(1'b0), .S(S[5]) );
  FA_986 \FAINST[6].FA_  ( .A(A[6]), .B(1'b0), .CI(1'b0), .S(S[6]) );
  FA_985 \FAINST[7].FA_  ( .A(A[7]), .B(1'b0), .CI(1'b0), .S(S[7]) );
  FA_984 \FAINST[8].FA_  ( .A(A[8]), .B(1'b0), .CI(1'b0), .S(S[8]) );
  FA_983 \FAINST[9].FA_  ( .A(A[9]), .B(1'b0), .CI(1'b0), .S(S[9]) );
  FA_982 \FAINST[10].FA_  ( .A(A[10]), .B(1'b0), .CI(1'b0), .S(S[10]) );
  FA_981 \FAINST[11].FA_  ( .A(A[11]), .B(1'b0), .CI(1'b0), .S(S[11]) );
  FA_980 \FAINST[12].FA_  ( .A(A[12]), .B(1'b0), .CI(1'b0), .S(S[12]) );
  FA_979 \FAINST[13].FA_  ( .A(A[13]), .B(1'b0), .CI(1'b0), .S(S[13]) );
  FA_978 \FAINST[14].FA_  ( .A(A[14]), .B(1'b0), .CI(1'b0), .S(S[14]) );
  FA_977 \FAINST[15].FA_  ( .A(A[15]), .B(1'b0), .CI(1'b0), .S(S[15]) );
  FA_976 \FAINST[16].FA_  ( .A(A[16]), .B(1'b0), .CI(1'b0), .S(S[16]) );
  FA_975 \FAINST[17].FA_  ( .A(A[17]), .B(1'b0), .CI(1'b0), .S(S[17]) );
  FA_974 \FAINST[18].FA_  ( .A(A[18]), .B(1'b0), .CI(1'b0), .S(S[18]) );
  FA_973 \FAINST[19].FA_  ( .A(A[19]), .B(1'b0), .CI(1'b0), .S(S[19]) );
  FA_972 \FAINST[20].FA_  ( .A(A[20]), .B(1'b0), .CI(1'b0), .S(S[20]) );
  FA_971 \FAINST[21].FA_  ( .A(A[21]), .B(1'b0), .CI(1'b0), .S(S[21]) );
  FA_970 \FAINST[22].FA_  ( .A(A[22]), .B(1'b0), .CI(1'b0), .S(S[22]) );
  FA_969 \FAINST[23].FA_  ( .A(A[23]), .B(1'b0), .CI(1'b0), .S(S[23]) );
  FA_968 \FAINST[24].FA_  ( .A(A[24]), .B(1'b0), .CI(1'b0), .S(S[24]) );
  FA_967 \FAINST[25].FA_  ( .A(A[25]), .B(1'b0), .CI(1'b0), .S(S[25]) );
  FA_966 \FAINST[26].FA_  ( .A(A[26]), .B(1'b0), .CI(1'b0), .S(S[26]) );
  FA_965 \FAINST[27].FA_  ( .A(A[27]), .B(1'b0), .CI(1'b0), .S(S[27]) );
  FA_964 \FAINST[28].FA_  ( .A(A[28]), .B(1'b0), .CI(1'b0), .S(S[28]) );
  FA_963 \FAINST[29].FA_  ( .A(A[29]), .B(1'b0), .CI(1'b0), .S(S[29]) );
  FA_962 \FAINST[30].FA_  ( .A(A[30]), .B(1'b0), .CI(1'b0), .S(S[30]) );
  FA_961 \FAINST[31].FA_  ( .A(A[31]), .B(1'b0), .CI(1'b0), .S(S[31]) );
endmodule


module MULT_N32_1 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   \w[31][31] , \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] ,
         \w[31][26] , \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] ,
         \w[31][21] , \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] ,
         \w[31][16] , \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] ,
         \w[31][11] , \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] ,
         \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] ,
         \w[31][1] , \w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] ,
         \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] ,
         \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] ,
         \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] ,
         \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] ,
         \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] ,
         \w[30][2] , \w[30][1] , \w[29][31] , \w[29][30] , \w[29][29] ,
         \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] ,
         \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] ,
         \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] ,
         \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] ,
         \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] ,
         \w[29][3] , \w[29][2] , \w[29][1] , \w[28][31] , \w[28][30] ,
         \w[28][29] , \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] ,
         \w[28][24] , \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] ,
         \w[28][19] , \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] ,
         \w[28][14] , \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] ,
         \w[28][9] , \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] ,
         \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , \w[27][31] ,
         \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] ,
         \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] ,
         \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] ,
         \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] ,
         \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] ,
         \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] ,
         \w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] ,
         \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] ,
         \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] ,
         \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] ,
         \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] ,
         \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] ,
         \w[26][1] , \w[25][31] , \w[25][30] , \w[25][29] , \w[25][28] ,
         \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , \w[25][23] ,
         \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , \w[25][18] ,
         \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , \w[25][13] ,
         \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , \w[25][8] ,
         \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] ,
         \w[25][2] , \w[25][1] , \w[24][31] , \w[24][30] , \w[24][29] ,
         \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] ,
         \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] ,
         \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] ,
         \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] ,
         \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] ,
         \w[24][3] , \w[24][2] , \w[24][1] , \w[23][31] , \w[23][30] ,
         \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] ,
         \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] ,
         \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] ,
         \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] ,
         \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] ,
         \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , \w[22][31] ,
         \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , \w[22][26] ,
         \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , \w[22][21] ,
         \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , \w[22][16] ,
         \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , \w[22][11] ,
         \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , \w[22][6] ,
         \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] ,
         \w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] ,
         \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] ,
         \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] ,
         \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] ,
         \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] ,
         \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] ,
         \w[21][1] , \w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] ,
         \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] ,
         \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] ,
         \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] ,
         \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] ,
         \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] ,
         \w[20][2] , \w[20][1] , \w[19][31] , \w[19][30] , \w[19][29] ,
         \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] ,
         \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] ,
         \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] ,
         \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] ,
         \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] ,
         \w[19][3] , \w[19][2] , \w[19][1] , \w[18][31] , \w[18][30] ,
         \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] ,
         \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] ,
         \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] ,
         \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] ,
         \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] ,
         \w[18][4] , \w[18][3] , \w[18][2] , \w[18][1] , \w[17][31] ,
         \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] ,
         \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] ,
         \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] ,
         \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] ,
         \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] ,
         \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] ,
         \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] ,
         \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] ,
         \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] ,
         \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] ,
         \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] ,
         \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] ,
         \w[16][1] , \w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] ,
         \w[15][27] , \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] ,
         \w[15][22] , \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] ,
         \w[15][17] , \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] ,
         \w[15][12] , \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] ,
         \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] ,
         \w[15][2] , \w[15][1] , \w[14][31] , \w[14][30] , \w[14][29] ,
         \w[14][28] , \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] ,
         \w[14][23] , \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] ,
         \w[14][18] , \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] ,
         \w[14][13] , \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] ,
         \w[14][8] , \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] ,
         \w[14][3] , \w[14][2] , \w[14][1] , \w[13][31] , \w[13][30] ,
         \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] ,
         \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] ,
         \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] ,
         \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] ,
         \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] ,
         \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , \w[12][31] ,
         \w[12][30] , \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] ,
         \w[12][25] , \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] ,
         \w[12][20] , \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] ,
         \w[12][15] , \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] ,
         \w[12][10] , \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] ,
         \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , \w[12][1] ,
         \w[11][31] , \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] ,
         \w[11][26] , \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] ,
         \w[11][21] , \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] ,
         \w[11][16] , \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] ,
         \w[11][11] , \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] ,
         \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] ,
         \w[11][1] , \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] ,
         \w[10][27] , \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] ,
         \w[10][22] , \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] ,
         \w[10][17] , \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] ,
         \w[10][12] , \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] ,
         \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] ,
         \w[10][2] , \w[10][1] , \w[9][31] , \w[9][30] , \w[9][29] ,
         \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] ,
         \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] ,
         \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] ,
         \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] ,
         \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] ,
         \w[9][1] , \w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] ,
         \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] ,
         \w[8][21] , \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] ,
         \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , \w[8][12] ,
         \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , \w[8][6] ,
         \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , \w[7][31] ,
         \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] ,
         \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] ,
         \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] ,
         \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] ,
         \w[7][10] , \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] ,
         \w[7][4] , \w[7][3] , \w[7][2] , \w[7][1] , \w[6][31] , \w[6][30] ,
         \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] ,
         \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] ,
         \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] ,
         \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] ,
         \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] ,
         \w[6][2] , \w[6][1] , \w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] ,
         \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] ,
         \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] ,
         \w[5][17] , \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] ,
         \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] ,
         \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] ,
         \w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] ,
         \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] ,
         \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] ,
         \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] ,
         \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] ,
         \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , \w[3][31] ,
         \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] ,
         \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] ,
         \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] ,
         \w[3][15] , \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] ,
         \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] ,
         \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , \w[2][31] , \w[2][30] ,
         \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] ,
         \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] ,
         \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] ,
         \w[2][14] , \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] ,
         \w[2][8] , \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] ,
         \w[2][2] , \w[2][1] , \_0_net_[31] , \_0_net_[30] , \_0_net_[29] ,
         \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , \_0_net_[25] ,
         \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , \_0_net_[21] ,
         \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , \_0_net_[17] ,
         \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , \_0_net_[13] ,
         \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , \_0_net_[9] ,
         \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] ,
         \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_2_net_[31] ,
         \_2_net_[30] , \_2_net_[29] , \_2_net_[28] , \_2_net_[27] ,
         \_2_net_[26] , \_2_net_[25] , \_2_net_[24] , \_2_net_[23] ,
         \_2_net_[22] , \_2_net_[21] , \_2_net_[20] , \_2_net_[19] ,
         \_2_net_[18] , \_2_net_[17] , \_2_net_[16] , \_2_net_[15] ,
         \_2_net_[14] , \_2_net_[13] , \_2_net_[12] , \_2_net_[11] ,
         \_2_net_[10] , \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] ,
         \_2_net_[5] , \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , \_4_net_[31] ,
         \_4_net_[30] , \_4_net_[29] , \_4_net_[28] , \_4_net_[27] ,
         \_4_net_[26] , \_4_net_[25] , \_4_net_[24] , \_4_net_[23] ,
         \_4_net_[22] , \_4_net_[21] , \_4_net_[20] , \_4_net_[19] ,
         \_4_net_[18] , \_4_net_[17] , \_4_net_[16] , \_4_net_[15] ,
         \_4_net_[14] , \_4_net_[13] , \_4_net_[12] , \_4_net_[11] ,
         \_4_net_[10] , \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] ,
         \_4_net_[5] , \_4_net_[4] , \_4_net_[3] , \_6_net_[31] ,
         \_6_net_[30] , \_6_net_[29] , \_6_net_[28] , \_6_net_[27] ,
         \_6_net_[26] , \_6_net_[25] , \_6_net_[24] , \_6_net_[23] ,
         \_6_net_[22] , \_6_net_[21] , \_6_net_[20] , \_6_net_[19] ,
         \_6_net_[18] , \_6_net_[17] , \_6_net_[16] , \_6_net_[15] ,
         \_6_net_[14] , \_6_net_[13] , \_6_net_[12] , \_6_net_[11] ,
         \_6_net_[10] , \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] ,
         \_6_net_[5] , \_6_net_[4] , \_8_net_[31] , \_8_net_[30] ,
         \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] ,
         \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] ,
         \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] ,
         \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] ,
         \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] ,
         \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] ,
         \_10_net_[31] , \_10_net_[30] , \_10_net_[29] , \_10_net_[28] ,
         \_10_net_[27] , \_10_net_[26] , \_10_net_[25] , \_10_net_[24] ,
         \_10_net_[23] , \_10_net_[22] , \_10_net_[21] , \_10_net_[20] ,
         \_10_net_[19] , \_10_net_[18] , \_10_net_[17] , \_10_net_[16] ,
         \_10_net_[15] , \_10_net_[14] , \_10_net_[13] , \_10_net_[12] ,
         \_10_net_[11] , \_10_net_[10] , \_10_net_[9] , \_10_net_[8] ,
         \_10_net_[7] , \_10_net_[6] , \_12_net_[31] , \_12_net_[30] ,
         \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] ,
         \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] ,
         \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] ,
         \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] ,
         \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] ,
         \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , \_14_net_[31] ,
         \_14_net_[30] , \_14_net_[29] , \_14_net_[28] , \_14_net_[27] ,
         \_14_net_[26] , \_14_net_[25] , \_14_net_[24] , \_14_net_[23] ,
         \_14_net_[22] , \_14_net_[21] , \_14_net_[20] , \_14_net_[19] ,
         \_14_net_[18] , \_14_net_[17] , \_14_net_[16] , \_14_net_[15] ,
         \_14_net_[14] , \_14_net_[13] , \_14_net_[12] , \_14_net_[11] ,
         \_14_net_[10] , \_14_net_[9] , \_14_net_[8] , \_16_net_[31] ,
         \_16_net_[30] , \_16_net_[29] , \_16_net_[28] , \_16_net_[27] ,
         \_16_net_[26] , \_16_net_[25] , \_16_net_[24] , \_16_net_[23] ,
         \_16_net_[22] , \_16_net_[21] , \_16_net_[20] , \_16_net_[19] ,
         \_16_net_[18] , \_16_net_[17] , \_16_net_[16] , \_16_net_[15] ,
         \_16_net_[14] , \_16_net_[13] , \_16_net_[12] , \_16_net_[11] ,
         \_16_net_[10] , \_16_net_[9] , \_18_net_[31] , \_18_net_[30] ,
         \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] ,
         \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] ,
         \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] ,
         \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] ,
         \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] ,
         \_20_net_[31] , \_20_net_[30] , \_20_net_[29] , \_20_net_[28] ,
         \_20_net_[27] , \_20_net_[26] , \_20_net_[25] , \_20_net_[24] ,
         \_20_net_[23] , \_20_net_[22] , \_20_net_[21] , \_20_net_[20] ,
         \_20_net_[19] , \_20_net_[18] , \_20_net_[17] , \_20_net_[16] ,
         \_20_net_[15] , \_20_net_[14] , \_20_net_[13] , \_20_net_[12] ,
         \_20_net_[11] , \_22_net_[31] , \_22_net_[30] , \_22_net_[29] ,
         \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , \_22_net_[25] ,
         \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , \_22_net_[21] ,
         \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , \_22_net_[17] ,
         \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , \_22_net_[13] ,
         \_22_net_[12] , \_24_net_[31] , \_24_net_[30] , \_24_net_[29] ,
         \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , \_24_net_[25] ,
         \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , \_24_net_[21] ,
         \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , \_24_net_[17] ,
         \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , \_24_net_[13] ,
         \_26_net_[31] , \_26_net_[30] , \_26_net_[29] , \_26_net_[28] ,
         \_26_net_[27] , \_26_net_[26] , \_26_net_[25] , \_26_net_[24] ,
         \_26_net_[23] , \_26_net_[22] , \_26_net_[21] , \_26_net_[20] ,
         \_26_net_[19] , \_26_net_[18] , \_26_net_[17] , \_26_net_[16] ,
         \_26_net_[15] , \_26_net_[14] , \_28_net_[31] , \_28_net_[30] ,
         \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] ,
         \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] ,
         \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] ,
         \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , \_30_net_[31] ,
         \_30_net_[30] , \_30_net_[29] , \_30_net_[28] , \_30_net_[27] ,
         \_30_net_[26] , \_30_net_[25] , \_30_net_[24] , \_30_net_[23] ,
         \_30_net_[22] , \_30_net_[21] , \_30_net_[20] , \_30_net_[19] ,
         \_30_net_[18] , \_30_net_[17] , \_30_net_[16] , \_32_net_[31] ,
         \_32_net_[30] , \_32_net_[29] , \_32_net_[28] , \_32_net_[27] ,
         \_32_net_[26] , \_32_net_[25] , \_32_net_[24] , \_32_net_[23] ,
         \_32_net_[22] , \_32_net_[21] , \_32_net_[20] , \_32_net_[19] ,
         \_32_net_[18] , \_32_net_[17] , \_34_net_[31] , \_34_net_[30] ,
         \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] ,
         \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] ,
         \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] ,
         \_36_net_[31] , \_36_net_[30] , \_36_net_[29] , \_36_net_[28] ,
         \_36_net_[27] , \_36_net_[26] , \_36_net_[25] , \_36_net_[24] ,
         \_36_net_[23] , \_36_net_[22] , \_36_net_[21] , \_36_net_[20] ,
         \_36_net_[19] , \_38_net_[31] , \_38_net_[30] , \_38_net_[29] ,
         \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , \_38_net_[25] ,
         \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , \_38_net_[21] ,
         \_38_net_[20] , \_40_net_[31] , \_40_net_[30] , \_40_net_[29] ,
         \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , \_40_net_[25] ,
         \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , \_40_net_[21] ,
         \_42_net_[31] , \_42_net_[30] , \_42_net_[29] , \_42_net_[28] ,
         \_42_net_[27] , \_42_net_[26] , \_42_net_[25] , \_42_net_[24] ,
         \_42_net_[23] , \_42_net_[22] , \_44_net_[31] , \_44_net_[30] ,
         \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] ,
         \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , \_46_net_[31] ,
         \_46_net_[30] , \_46_net_[29] , \_46_net_[28] , \_46_net_[27] ,
         \_46_net_[26] , \_46_net_[25] , \_46_net_[24] , \_48_net_[31] ,
         \_48_net_[30] , \_48_net_[29] , \_48_net_[28] , \_48_net_[27] ,
         \_48_net_[26] , \_48_net_[25] , \_50_net_[31] , \_50_net_[30] ,
         \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] ,
         \_52_net_[31] , \_52_net_[30] , \_52_net_[29] , \_52_net_[28] ,
         \_52_net_[27] , \_54_net_[31] , \_54_net_[30] , \_54_net_[29] ,
         \_54_net_[28] , \_56_net_[31] , \_56_net_[30] , \_56_net_[29] ,
         \_58_net_[31] , \_58_net_[30] , \_60_net_[31] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  ADD_N32_31 \FAINST[1].ADD_  ( .A({\_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .S({
        \w[2][31] , \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , 
        \w[2][25] , \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , 
        \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , 
        \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , 
        \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , 
        \w[2][1] , SYNOPSYS_UNCONNECTED__0}) );
  ADD_N32_30 \FAINST[2].ADD_  ( .A({\_2_net_[31] , \_2_net_[30] , 
        \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , \_2_net_[26] , 
        \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , \_2_net_[22] , 
        \_2_net_[21] , \_2_net_[20] , \_2_net_[19] , \_2_net_[18] , 
        \_2_net_[17] , \_2_net_[16] , \_2_net_[15] , \_2_net_[14] , 
        \_2_net_[13] , \_2_net_[12] , \_2_net_[11] , \_2_net_[10] , 
        \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , \_2_net_[5] , 
        \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , 1'b0, 1'b0}), .B({\w[2][31] , 
        \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] , 
        \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , \w[2][19] , 
        \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , \w[2][13] , 
        \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , \w[2][7] , 
        \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , \w[2][1] , 1'b0}), .CI(1'b0), .S({\w[3][31] , \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , 
        \w[3][26] , \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , 
        \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , 
        \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , 
        \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , 
        \w[3][2] , \w[3][1] , SYNOPSYS_UNCONNECTED__1}) );
  ADD_N32_29 \FAINST[3].ADD_  ( .A({\_4_net_[31] , \_4_net_[30] , 
        \_4_net_[29] , \_4_net_[28] , \_4_net_[27] , \_4_net_[26] , 
        \_4_net_[25] , \_4_net_[24] , \_4_net_[23] , \_4_net_[22] , 
        \_4_net_[21] , \_4_net_[20] , \_4_net_[19] , \_4_net_[18] , 
        \_4_net_[17] , \_4_net_[16] , \_4_net_[15] , \_4_net_[14] , 
        \_4_net_[13] , \_4_net_[12] , \_4_net_[11] , \_4_net_[10] , 
        \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] , \_4_net_[5] , 
        \_4_net_[4] , \_4_net_[3] , 1'b0, 1'b0, 1'b0}), .B({\w[3][31] , 
        \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] , \w[3][25] , 
        \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , \w[3][20] , \w[3][19] , 
        \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , \w[3][14] , \w[3][13] , 
        \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , 
        \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , 1'b0}), .CI(1'b0), .S({\w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] , 
        \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] , \w[4][21] , 
        \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] , \w[4][16] , \w[4][15] , 
        \w[4][14] , \w[4][13] , \w[4][12] , \w[4][11] , \w[4][10] , \w[4][9] , 
        \w[4][8] , \w[4][7] , \w[4][6] , \w[4][5] , \w[4][4] , \w[4][3] , 
        \w[4][2] , \w[4][1] , SYNOPSYS_UNCONNECTED__2}) );
  ADD_N32_28 \FAINST[4].ADD_  ( .A({\_6_net_[31] , \_6_net_[30] , 
        \_6_net_[29] , \_6_net_[28] , \_6_net_[27] , \_6_net_[26] , 
        \_6_net_[25] , \_6_net_[24] , \_6_net_[23] , \_6_net_[22] , 
        \_6_net_[21] , \_6_net_[20] , \_6_net_[19] , \_6_net_[18] , 
        \_6_net_[17] , \_6_net_[16] , \_6_net_[15] , \_6_net_[14] , 
        \_6_net_[13] , \_6_net_[12] , \_6_net_[11] , \_6_net_[10] , 
        \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] , \_6_net_[5] , 
        \_6_net_[4] , 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[4][31] , \w[4][30] , 
        \w[4][29] , \w[4][28] , \w[4][27] , \w[4][26] , \w[4][25] , \w[4][24] , 
        \w[4][23] , \w[4][22] , \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , 
        \w[4][17] , \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] , 
        \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] , 
        \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , 1'b0}), .CI(
        1'b0), .S({\w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] , \w[5][27] , 
        \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , \w[5][22] , \w[5][21] , 
        \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , \w[5][16] , \w[5][15] , 
        \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , 
        \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , 
        \w[5][2] , \w[5][1] , SYNOPSYS_UNCONNECTED__3}) );
  ADD_N32_27 \FAINST[5].ADD_  ( .A({\_8_net_[31] , \_8_net_[30] , 
        \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] , 
        \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] , 
        \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] , 
        \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] , 
        \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] , 
        \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[5][31] , \w[5][30] , \w[5][29] , 
        \w[5][28] , \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , 
        \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , 
        \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , 
        \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , 
        \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] , 1'b0}), .CI(1'b0), .S({
        \w[6][31] , \w[6][30] , \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , 
        \w[6][25] , \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] , 
        \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] , \w[6][14] , 
        \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] , \w[6][8] , 
        \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] , \w[6][2] , 
        \w[6][1] , SYNOPSYS_UNCONNECTED__4}) );
  ADD_N32_26 \FAINST[6].ADD_  ( .A({\_10_net_[31] , \_10_net_[30] , 
        \_10_net_[29] , \_10_net_[28] , \_10_net_[27] , \_10_net_[26] , 
        \_10_net_[25] , \_10_net_[24] , \_10_net_[23] , \_10_net_[22] , 
        \_10_net_[21] , \_10_net_[20] , \_10_net_[19] , \_10_net_[18] , 
        \_10_net_[17] , \_10_net_[16] , \_10_net_[15] , \_10_net_[14] , 
        \_10_net_[13] , \_10_net_[12] , \_10_net_[11] , \_10_net_[10] , 
        \_10_net_[9] , \_10_net_[8] , \_10_net_[7] , \_10_net_[6] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[6][31] , \w[6][30] , \w[6][29] , 
        \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] , \w[6][24] , \w[6][23] , 
        \w[6][22] , \w[6][21] , \w[6][20] , \w[6][19] , \w[6][18] , \w[6][17] , 
        \w[6][16] , \w[6][15] , \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , 
        \w[6][10] , \w[6][9] , \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , 
        \w[6][4] , \w[6][3] , \w[6][2] , \w[6][1] , 1'b0}), .CI(1'b0), .S({
        \w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] , 
        \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] , \w[7][20] , 
        \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , \w[7][15] , \w[7][14] , 
        \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , \w[7][9] , \w[7][8] , 
        \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , \w[7][3] , \w[7][2] , 
        \w[7][1] , SYNOPSYS_UNCONNECTED__5}) );
  ADD_N32_25 \FAINST[7].ADD_  ( .A({\_12_net_[31] , \_12_net_[30] , 
        \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] , 
        \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] , 
        \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] , 
        \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] , 
        \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] , 
        \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , 
        \w[7][27] , \w[7][26] , \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , 
        \w[7][21] , \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , 
        \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , 
        \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , 
        \w[7][3] , \w[7][2] , \w[7][1] , 1'b0}), .CI(1'b0), .S({\w[8][31] , 
        \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , \w[8][26] , \w[8][25] , 
        \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , \w[8][20] , \w[8][19] , 
        \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , 
        \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , 
        \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , 
        SYNOPSYS_UNCONNECTED__6}) );
  ADD_N32_24 \FAINST[8].ADD_  ( .A({\_14_net_[31] , \_14_net_[30] , 
        \_14_net_[29] , \_14_net_[28] , \_14_net_[27] , \_14_net_[26] , 
        \_14_net_[25] , \_14_net_[24] , \_14_net_[23] , \_14_net_[22] , 
        \_14_net_[21] , \_14_net_[20] , \_14_net_[19] , \_14_net_[18] , 
        \_14_net_[17] , \_14_net_[16] , \_14_net_[15] , \_14_net_[14] , 
        \_14_net_[13] , \_14_net_[12] , \_14_net_[11] , \_14_net_[10] , 
        \_14_net_[9] , \_14_net_[8] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , 
        \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , 
        \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , 
        \w[8][14] , \w[8][13] , \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , 
        \w[8][8] , \w[8][7] , \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , 
        \w[8][2] , \w[8][1] , 1'b0}), .CI(1'b0), .S({\w[9][31] , \w[9][30] , 
        \w[9][29] , \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] , 
        \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] , \w[9][18] , 
        \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] , \w[9][13] , \w[9][12] , 
        \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] , \w[9][7] , \w[9][6] , 
        \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] , \w[9][1] , 
        SYNOPSYS_UNCONNECTED__7}) );
  ADD_N32_23 \FAINST[9].ADD_  ( .A({\_16_net_[31] , \_16_net_[30] , 
        \_16_net_[29] , \_16_net_[28] , \_16_net_[27] , \_16_net_[26] , 
        \_16_net_[25] , \_16_net_[24] , \_16_net_[23] , \_16_net_[22] , 
        \_16_net_[21] , \_16_net_[20] , \_16_net_[19] , \_16_net_[18] , 
        \_16_net_[17] , \_16_net_[16] , \_16_net_[15] , \_16_net_[14] , 
        \_16_net_[13] , \_16_net_[12] , \_16_net_[11] , \_16_net_[10] , 
        \_16_net_[9] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[9][31] , \w[9][30] , \w[9][29] , \w[9][28] , \w[9][27] , 
        \w[9][26] , \w[9][25] , \w[9][24] , \w[9][23] , \w[9][22] , \w[9][21] , 
        \w[9][20] , \w[9][19] , \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , 
        \w[9][14] , \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , 
        \w[9][8] , \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , 
        \w[9][2] , \w[9][1] , 1'b0}), .CI(1'b0), .S({\w[10][31] , \w[10][30] , 
        \w[10][29] , \w[10][28] , \w[10][27] , \w[10][26] , \w[10][25] , 
        \w[10][24] , \w[10][23] , \w[10][22] , \w[10][21] , \w[10][20] , 
        \w[10][19] , \w[10][18] , \w[10][17] , \w[10][16] , \w[10][15] , 
        \w[10][14] , \w[10][13] , \w[10][12] , \w[10][11] , \w[10][10] , 
        \w[10][9] , \w[10][8] , \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , 
        \w[10][3] , \w[10][2] , \w[10][1] , SYNOPSYS_UNCONNECTED__8}) );
  ADD_N32_22 \FAINST[10].ADD_  ( .A({\_18_net_[31] , \_18_net_[30] , 
        \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] , 
        \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] , 
        \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] , 
        \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] , 
        \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] , \w[10][27] , 
        \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] , \w[10][22] , 
        \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] , \w[10][17] , 
        \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] , \w[10][12] , 
        \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] , \w[10][7] , 
        \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] , \w[10][2] , \w[10][1] , 
        1'b0}), .CI(1'b0), .S({\w[11][31] , \w[11][30] , \w[11][29] , 
        \w[11][28] , \w[11][27] , \w[11][26] , \w[11][25] , \w[11][24] , 
        \w[11][23] , \w[11][22] , \w[11][21] , \w[11][20] , \w[11][19] , 
        \w[11][18] , \w[11][17] , \w[11][16] , \w[11][15] , \w[11][14] , 
        \w[11][13] , \w[11][12] , \w[11][11] , \w[11][10] , \w[11][9] , 
        \w[11][8] , \w[11][7] , \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , 
        \w[11][2] , \w[11][1] , SYNOPSYS_UNCONNECTED__9}) );
  ADD_N32_21 \FAINST[11].ADD_  ( .A({\_20_net_[31] , \_20_net_[30] , 
        \_20_net_[29] , \_20_net_[28] , \_20_net_[27] , \_20_net_[26] , 
        \_20_net_[25] , \_20_net_[24] , \_20_net_[23] , \_20_net_[22] , 
        \_20_net_[21] , \_20_net_[20] , \_20_net_[19] , \_20_net_[18] , 
        \_20_net_[17] , \_20_net_[16] , \_20_net_[15] , \_20_net_[14] , 
        \_20_net_[13] , \_20_net_[12] , \_20_net_[11] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[11][31] , 
        \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] , \w[11][26] , 
        \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] , \w[11][21] , 
        \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] , \w[11][16] , 
        \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] , \w[11][11] , 
        \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] , \w[11][6] , 
        \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] , \w[11][1] , 1'b0}), 
        .CI(1'b0), .S({\w[12][31] , \w[12][30] , \w[12][29] , \w[12][28] , 
        \w[12][27] , \w[12][26] , \w[12][25] , \w[12][24] , \w[12][23] , 
        \w[12][22] , \w[12][21] , \w[12][20] , \w[12][19] , \w[12][18] , 
        \w[12][17] , \w[12][16] , \w[12][15] , \w[12][14] , \w[12][13] , 
        \w[12][12] , \w[12][11] , \w[12][10] , \w[12][9] , \w[12][8] , 
        \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , 
        \w[12][1] , SYNOPSYS_UNCONNECTED__10}) );
  ADD_N32_20 \FAINST[12].ADD_  ( .A({\_22_net_[31] , \_22_net_[30] , 
        \_22_net_[29] , \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , 
        \_22_net_[25] , \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , 
        \_22_net_[21] , \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , 
        \_22_net_[17] , \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , 
        \_22_net_[13] , \_22_net_[12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[12][31] , \w[12][30] , 
        \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] , \w[12][25] , 
        \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] , \w[12][20] , 
        \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] , \w[12][15] , 
        \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] , \w[12][10] , 
        \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , 
        \w[12][3] , \w[12][2] , \w[12][1] , 1'b0}), .CI(1'b0), .S({\w[13][31] , 
        \w[13][30] , \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , 
        \w[13][25] , \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , 
        \w[13][20] , \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , 
        \w[13][15] , \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , 
        \w[13][10] , \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , 
        \w[13][5] , \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , 
        SYNOPSYS_UNCONNECTED__11}) );
  ADD_N32_19 \FAINST[13].ADD_  ( .A({\_24_net_[31] , \_24_net_[30] , 
        \_24_net_[29] , \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , 
        \_24_net_[25] , \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , 
        \_24_net_[21] , \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , 
        \_24_net_[17] , \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , 
        \_24_net_[13] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[13][31] , \w[13][30] , \w[13][29] , 
        \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] , \w[13][24] , 
        \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] , \w[13][19] , 
        \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] , \w[13][14] , 
        \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] , \w[13][9] , 
        \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] , \w[13][4] , \w[13][3] , 
        \w[13][2] , \w[13][1] , 1'b0}), .CI(1'b0), .S({\w[14][31] , 
        \w[14][30] , \w[14][29] , \w[14][28] , \w[14][27] , \w[14][26] , 
        \w[14][25] , \w[14][24] , \w[14][23] , \w[14][22] , \w[14][21] , 
        \w[14][20] , \w[14][19] , \w[14][18] , \w[14][17] , \w[14][16] , 
        \w[14][15] , \w[14][14] , \w[14][13] , \w[14][12] , \w[14][11] , 
        \w[14][10] , \w[14][9] , \w[14][8] , \w[14][7] , \w[14][6] , 
        \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , \w[14][1] , 
        SYNOPSYS_UNCONNECTED__12}) );
  ADD_N32_18 \FAINST[14].ADD_  ( .A({\_26_net_[31] , \_26_net_[30] , 
        \_26_net_[29] , \_26_net_[28] , \_26_net_[27] , \_26_net_[26] , 
        \_26_net_[25] , \_26_net_[24] , \_26_net_[23] , \_26_net_[22] , 
        \_26_net_[21] , \_26_net_[20] , \_26_net_[19] , \_26_net_[18] , 
        \_26_net_[17] , \_26_net_[16] , \_26_net_[15] , \_26_net_[14] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[14][31] , \w[14][30] , \w[14][29] , \w[14][28] , 
        \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] , \w[14][23] , 
        \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] , \w[14][18] , 
        \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] , \w[14][13] , 
        \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] , \w[14][8] , 
        \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , 
        \w[14][1] , 1'b0}), .CI(1'b0), .S({\w[15][31] , \w[15][30] , 
        \w[15][29] , \w[15][28] , \w[15][27] , \w[15][26] , \w[15][25] , 
        \w[15][24] , \w[15][23] , \w[15][22] , \w[15][21] , \w[15][20] , 
        \w[15][19] , \w[15][18] , \w[15][17] , \w[15][16] , \w[15][15] , 
        \w[15][14] , \w[15][13] , \w[15][12] , \w[15][11] , \w[15][10] , 
        \w[15][9] , \w[15][8] , \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , 
        \w[15][3] , \w[15][2] , \w[15][1] , SYNOPSYS_UNCONNECTED__13}) );
  ADD_N32_17 \FAINST[15].ADD_  ( .A({\_28_net_[31] , \_28_net_[30] , 
        \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] , 
        \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] , 
        \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] , 
        \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] , \w[15][27] , 
        \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] , \w[15][22] , 
        \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] , \w[15][17] , 
        \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] , \w[15][12] , 
        \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] , \w[15][7] , 
        \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] , \w[15][2] , \w[15][1] , 
        1'b0}), .CI(1'b0), .S({\w[16][31] , \w[16][30] , \w[16][29] , 
        \w[16][28] , \w[16][27] , \w[16][26] , \w[16][25] , \w[16][24] , 
        \w[16][23] , \w[16][22] , \w[16][21] , \w[16][20] , \w[16][19] , 
        \w[16][18] , \w[16][17] , \w[16][16] , \w[16][15] , \w[16][14] , 
        \w[16][13] , \w[16][12] , \w[16][11] , \w[16][10] , \w[16][9] , 
        \w[16][8] , \w[16][7] , \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , 
        \w[16][2] , \w[16][1] , SYNOPSYS_UNCONNECTED__14}) );
  ADD_N32_16 \FAINST[16].ADD_  ( .A({\_30_net_[31] , \_30_net_[30] , 
        \_30_net_[29] , \_30_net_[28] , \_30_net_[27] , \_30_net_[26] , 
        \_30_net_[25] , \_30_net_[24] , \_30_net_[23] , \_30_net_[22] , 
        \_30_net_[21] , \_30_net_[20] , \_30_net_[19] , \_30_net_[18] , 
        \_30_net_[17] , \_30_net_[16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] , 
        \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] , 
        \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] , 
        \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] , 
        \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] , 
        \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] , \w[16][1] , 
        1'b0}), .CI(1'b0), .S({\w[17][31] , \w[17][30] , \w[17][29] , 
        \w[17][28] , \w[17][27] , \w[17][26] , \w[17][25] , \w[17][24] , 
        \w[17][23] , \w[17][22] , \w[17][21] , \w[17][20] , \w[17][19] , 
        \w[17][18] , \w[17][17] , \w[17][16] , \w[17][15] , \w[17][14] , 
        \w[17][13] , \w[17][12] , \w[17][11] , \w[17][10] , \w[17][9] , 
        \w[17][8] , \w[17][7] , \w[17][6] , \w[17][5] , \w[17][4] , \w[17][3] , 
        \w[17][2] , \w[17][1] , SYNOPSYS_UNCONNECTED__15}) );
  ADD_N32_15 \FAINST[17].ADD_  ( .A({\_32_net_[31] , \_32_net_[30] , 
        \_32_net_[29] , \_32_net_[28] , \_32_net_[27] , \_32_net_[26] , 
        \_32_net_[25] , \_32_net_[24] , \_32_net_[23] , \_32_net_[22] , 
        \_32_net_[21] , \_32_net_[20] , \_32_net_[19] , \_32_net_[18] , 
        \_32_net_[17] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[17][31] , 
        \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] , 
        \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] , 
        \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] , 
        \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] , 
        \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] , 
        \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] , 1'b0}), 
        .CI(1'b0), .S({\w[18][31] , \w[18][30] , \w[18][29] , \w[18][28] , 
        \w[18][27] , \w[18][26] , \w[18][25] , \w[18][24] , \w[18][23] , 
        \w[18][22] , \w[18][21] , \w[18][20] , \w[18][19] , \w[18][18] , 
        \w[18][17] , \w[18][16] , \w[18][15] , \w[18][14] , \w[18][13] , 
        \w[18][12] , \w[18][11] , \w[18][10] , \w[18][9] , \w[18][8] , 
        \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , \w[18][3] , \w[18][2] , 
        \w[18][1] , SYNOPSYS_UNCONNECTED__16}) );
  ADD_N32_14 \FAINST[18].ADD_  ( .A({\_34_net_[31] , \_34_net_[30] , 
        \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] , 
        \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] , 
        \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[18][31] , \w[18][30] , 
        \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] , 
        \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] , 
        \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] , 
        \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] , 
        \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , 
        \w[18][3] , \w[18][2] , \w[18][1] , 1'b0}), .CI(1'b0), .S({\w[19][31] , 
        \w[19][30] , \w[19][29] , \w[19][28] , \w[19][27] , \w[19][26] , 
        \w[19][25] , \w[19][24] , \w[19][23] , \w[19][22] , \w[19][21] , 
        \w[19][20] , \w[19][19] , \w[19][18] , \w[19][17] , \w[19][16] , 
        \w[19][15] , \w[19][14] , \w[19][13] , \w[19][12] , \w[19][11] , 
        \w[19][10] , \w[19][9] , \w[19][8] , \w[19][7] , \w[19][6] , 
        \w[19][5] , \w[19][4] , \w[19][3] , \w[19][2] , \w[19][1] , 
        SYNOPSYS_UNCONNECTED__17}) );
  ADD_N32_13 \FAINST[19].ADD_  ( .A({\_36_net_[31] , \_36_net_[30] , 
        \_36_net_[29] , \_36_net_[28] , \_36_net_[27] , \_36_net_[26] , 
        \_36_net_[25] , \_36_net_[24] , \_36_net_[23] , \_36_net_[22] , 
        \_36_net_[21] , \_36_net_[20] , \_36_net_[19] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[19][31] , \w[19][30] , \w[19][29] , 
        \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] , 
        \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] , 
        \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] , 
        \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] , 
        \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] , \w[19][3] , 
        \w[19][2] , \w[19][1] , 1'b0}), .CI(1'b0), .S({\w[20][31] , 
        \w[20][30] , \w[20][29] , \w[20][28] , \w[20][27] , \w[20][26] , 
        \w[20][25] , \w[20][24] , \w[20][23] , \w[20][22] , \w[20][21] , 
        \w[20][20] , \w[20][19] , \w[20][18] , \w[20][17] , \w[20][16] , 
        \w[20][15] , \w[20][14] , \w[20][13] , \w[20][12] , \w[20][11] , 
        \w[20][10] , \w[20][9] , \w[20][8] , \w[20][7] , \w[20][6] , 
        \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , \w[20][1] , 
        SYNOPSYS_UNCONNECTED__18}) );
  ADD_N32_12 \FAINST[20].ADD_  ( .A({\_38_net_[31] , \_38_net_[30] , 
        \_38_net_[29] , \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , 
        \_38_net_[25] , \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , 
        \_38_net_[21] , \_38_net_[20] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({\w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] , 
        \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] , 
        \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] , 
        \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] , 
        \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] , 
        \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , 
        \w[20][1] , 1'b0}), .CI(1'b0), .S({\w[21][31] , \w[21][30] , 
        \w[21][29] , \w[21][28] , \w[21][27] , \w[21][26] , \w[21][25] , 
        \w[21][24] , \w[21][23] , \w[21][22] , \w[21][21] , \w[21][20] , 
        \w[21][19] , \w[21][18] , \w[21][17] , \w[21][16] , \w[21][15] , 
        \w[21][14] , \w[21][13] , \w[21][12] , \w[21][11] , \w[21][10] , 
        \w[21][9] , \w[21][8] , \w[21][7] , \w[21][6] , \w[21][5] , \w[21][4] , 
        \w[21][3] , \w[21][2] , \w[21][1] , SYNOPSYS_UNCONNECTED__19}) );
  ADD_N32_11 \FAINST[21].ADD_  ( .A({\_40_net_[31] , \_40_net_[30] , 
        \_40_net_[29] , \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , 
        \_40_net_[25] , \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , 
        \_40_net_[21] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] , 
        \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] , 
        \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] , 
        \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] , 
        \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] , 
        \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] , \w[21][1] , 
        1'b0}), .CI(1'b0), .S({\w[22][31] , \w[22][30] , \w[22][29] , 
        \w[22][28] , \w[22][27] , \w[22][26] , \w[22][25] , \w[22][24] , 
        \w[22][23] , \w[22][22] , \w[22][21] , \w[22][20] , \w[22][19] , 
        \w[22][18] , \w[22][17] , \w[22][16] , \w[22][15] , \w[22][14] , 
        \w[22][13] , \w[22][12] , \w[22][11] , \w[22][10] , \w[22][9] , 
        \w[22][8] , \w[22][7] , \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , 
        \w[22][2] , \w[22][1] , SYNOPSYS_UNCONNECTED__20}) );
  ADD_N32_10 \FAINST[22].ADD_  ( .A({\_42_net_[31] , \_42_net_[30] , 
        \_42_net_[29] , \_42_net_[28] , \_42_net_[27] , \_42_net_[26] , 
        \_42_net_[25] , \_42_net_[24] , \_42_net_[23] , \_42_net_[22] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[22][31] , \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , 
        \w[22][26] , \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , 
        \w[22][21] , \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , 
        \w[22][16] , \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , 
        \w[22][11] , \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , 
        \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] , 
        1'b0}), .CI(1'b0), .S({\w[23][31] , \w[23][30] , \w[23][29] , 
        \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] , \w[23][24] , 
        \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] , \w[23][19] , 
        \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] , \w[23][14] , 
        \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] , \w[23][9] , 
        \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] , \w[23][4] , \w[23][3] , 
        \w[23][2] , \w[23][1] , SYNOPSYS_UNCONNECTED__21}) );
  ADD_N32_9 \FAINST[23].ADD_  ( .A({\_44_net_[31] , \_44_net_[30] , 
        \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] , 
        \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[23][31] , 
        \w[23][30] , \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , 
        \w[23][25] , \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , 
        \w[23][20] , \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , 
        \w[23][15] , \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , 
        \w[23][10] , \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , 
        \w[23][5] , \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , 1'b0}), 
        .CI(1'b0), .S({\w[24][31] , \w[24][30] , \w[24][29] , \w[24][28] , 
        \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] , \w[24][23] , 
        \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] , \w[24][18] , 
        \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] , \w[24][13] , 
        \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] , \w[24][8] , 
        \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , \w[24][3] , \w[24][2] , 
        \w[24][1] , SYNOPSYS_UNCONNECTED__22}) );
  ADD_N32_8 \FAINST[24].ADD_  ( .A({\_46_net_[31] , \_46_net_[30] , 
        \_46_net_[29] , \_46_net_[28] , \_46_net_[27] , \_46_net_[26] , 
        \_46_net_[25] , \_46_net_[24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[24][31] , \w[24][30] , 
        \w[24][29] , \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , 
        \w[24][24] , \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , 
        \w[24][19] , \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , 
        \w[24][14] , \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , 
        \w[24][9] , \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , 
        \w[24][3] , \w[24][2] , \w[24][1] , 1'b0}), .CI(1'b0), .S({\w[25][31] , 
        \w[25][30] , \w[25][29] , \w[25][28] , \w[25][27] , \w[25][26] , 
        \w[25][25] , \w[25][24] , \w[25][23] , \w[25][22] , \w[25][21] , 
        \w[25][20] , \w[25][19] , \w[25][18] , \w[25][17] , \w[25][16] , 
        \w[25][15] , \w[25][14] , \w[25][13] , \w[25][12] , \w[25][11] , 
        \w[25][10] , \w[25][9] , \w[25][8] , \w[25][7] , \w[25][6] , 
        \w[25][5] , \w[25][4] , \w[25][3] , \w[25][2] , \w[25][1] , 
        SYNOPSYS_UNCONNECTED__23}) );
  ADD_N32_7 \FAINST[25].ADD_  ( .A({\_48_net_[31] , \_48_net_[30] , 
        \_48_net_[29] , \_48_net_[28] , \_48_net_[27] , \_48_net_[26] , 
        \_48_net_[25] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[25][31] , \w[25][30] , \w[25][29] , 
        \w[25][28] , \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , 
        \w[25][23] , \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , 
        \w[25][18] , \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , 
        \w[25][13] , \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , 
        \w[25][8] , \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] , 
        \w[25][2] , \w[25][1] , 1'b0}), .CI(1'b0), .S({\w[26][31] , 
        \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] , \w[26][26] , 
        \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] , \w[26][21] , 
        \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] , \w[26][16] , 
        \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] , \w[26][11] , 
        \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] , \w[26][6] , 
        \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , \w[26][1] , 
        SYNOPSYS_UNCONNECTED__24}) );
  ADD_N32_6 \FAINST[26].ADD_  ( .A({\_50_net_[31] , \_50_net_[30] , 
        \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , 
        \w[26][27] , \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , 
        \w[26][22] , \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , 
        \w[26][17] , \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , 
        \w[26][12] , \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , 
        \w[26][7] , \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , 
        \w[26][1] , 1'b0}), .CI(1'b0), .S({\w[27][31] , \w[27][30] , 
        \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] , \w[27][25] , 
        \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] , \w[27][20] , 
        \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] , \w[27][15] , 
        \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] , \w[27][10] , 
        \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] , \w[27][5] , \w[27][4] , 
        \w[27][3] , \w[27][2] , \w[27][1] , SYNOPSYS_UNCONNECTED__25}) );
  ADD_N32_5 \FAINST[27].ADD_  ( .A({\_52_net_[31] , \_52_net_[30] , 
        \_52_net_[29] , \_52_net_[28] , \_52_net_[27] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[27][31] , \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , 
        \w[27][26] , \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , 
        \w[27][21] , \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , 
        \w[27][16] , \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , 
        \w[27][11] , \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , 
        \w[27][6] , \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] , 
        1'b0}), .CI(1'b0), .S({\w[28][31] , \w[28][30] , \w[28][29] , 
        \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] , \w[28][24] , 
        \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] , \w[28][19] , 
        \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] , \w[28][14] , 
        \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] , \w[28][9] , 
        \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , 
        \w[28][2] , \w[28][1] , SYNOPSYS_UNCONNECTED__26}) );
  ADD_N32_4 \FAINST[28].ADD_  ( .A({\_54_net_[31] , \_54_net_[30] , 
        \_54_net_[29] , \_54_net_[28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[28][31] , \w[28][30] , \w[28][29] , \w[28][28] , \w[28][27] , 
        \w[28][26] , \w[28][25] , \w[28][24] , \w[28][23] , \w[28][22] , 
        \w[28][21] , \w[28][20] , \w[28][19] , \w[28][18] , \w[28][17] , 
        \w[28][16] , \w[28][15] , \w[28][14] , \w[28][13] , \w[28][12] , 
        \w[28][11] , \w[28][10] , \w[28][9] , \w[28][8] , \w[28][7] , 
        \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , 
        1'b0}), .CI(1'b0), .S({\w[29][31] , \w[29][30] , \w[29][29] , 
        \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] , 
        \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] , 
        \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] , 
        \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] , 
        \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] , \w[29][3] , 
        \w[29][2] , \w[29][1] , SYNOPSYS_UNCONNECTED__27}) );
  ADD_N32_3 \FAINST[29].ADD_  ( .A({\_56_net_[31] , \_56_net_[30] , 
        \_56_net_[29] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[29][31] , 
        \w[29][30] , \w[29][29] , \w[29][28] , \w[29][27] , \w[29][26] , 
        \w[29][25] , \w[29][24] , \w[29][23] , \w[29][22] , \w[29][21] , 
        \w[29][20] , \w[29][19] , \w[29][18] , \w[29][17] , \w[29][16] , 
        \w[29][15] , \w[29][14] , \w[29][13] , \w[29][12] , \w[29][11] , 
        \w[29][10] , \w[29][9] , \w[29][8] , \w[29][7] , \w[29][6] , 
        \w[29][5] , \w[29][4] , \w[29][3] , \w[29][2] , \w[29][1] , 1'b0}), 
        .CI(1'b0), .S({\w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] , 
        \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] , 
        \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] , 
        \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] , 
        \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] , 
        \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] , \w[30][2] , 
        \w[30][1] , SYNOPSYS_UNCONNECTED__28}) );
  ADD_N32_2 \FAINST[30].ADD_  ( .A({\_58_net_[31] , \_58_net_[30] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[30][31] , \w[30][30] , \w[30][29] , 
        \w[30][28] , \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , 
        \w[30][23] , \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , 
        \w[30][18] , \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , 
        \w[30][13] , \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , 
        \w[30][8] , \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] , 
        \w[30][2] , \w[30][1] , 1'b0}), .CI(1'b0), .S({\w[31][31] , 
        \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] , \w[31][26] , 
        \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] , \w[31][21] , 
        \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] , \w[31][16] , 
        \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] , \w[31][11] , 
        \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] , \w[31][6] , 
        \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] , \w[31][1] , 
        SYNOPSYS_UNCONNECTED__29}) );
  ADD_N32_1 \FAINST[31].ADD_  ( .A({\_60_net_[31] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[31][31] , \w[31][30] , \w[31][29] , 
        \w[31][28] , \w[31][27] , \w[31][26] , \w[31][25] , \w[31][24] , 
        \w[31][23] , \w[31][22] , \w[31][21] , \w[31][20] , \w[31][19] , 
        \w[31][18] , \w[31][17] , \w[31][16] , \w[31][15] , \w[31][14] , 
        \w[31][13] , \w[31][12] , \w[31][11] , \w[31][10] , \w[31][9] , 
        \w[31][8] , \w[31][7] , \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , 
        \w[31][2] , \w[31][1] , 1'b0}), .CI(1'b0), .S({O[31:1], 
        SYNOPSYS_UNCONNECTED__30}) );
  AND U2 ( .A(A[5]), .B(B[4]), .Z(\_8_net_[9] ) );
  AND U3 ( .A(A[5]), .B(B[3]), .Z(\_8_net_[8] ) );
  AND U4 ( .A(A[5]), .B(B[2]), .Z(\_8_net_[7] ) );
  AND U5 ( .A(A[5]), .B(B[1]), .Z(\_8_net_[6] ) );
  AND U6 ( .A(A[5]), .B(B[0]), .Z(\_8_net_[5] ) );
  AND U7 ( .A(A[5]), .B(B[26]), .Z(\_8_net_[31] ) );
  AND U8 ( .A(A[5]), .B(B[25]), .Z(\_8_net_[30] ) );
  AND U9 ( .A(A[5]), .B(B[24]), .Z(\_8_net_[29] ) );
  AND U10 ( .A(A[5]), .B(B[23]), .Z(\_8_net_[28] ) );
  AND U11 ( .A(A[5]), .B(B[22]), .Z(\_8_net_[27] ) );
  AND U12 ( .A(A[5]), .B(B[21]), .Z(\_8_net_[26] ) );
  AND U13 ( .A(A[5]), .B(B[20]), .Z(\_8_net_[25] ) );
  AND U14 ( .A(A[5]), .B(B[19]), .Z(\_8_net_[24] ) );
  AND U15 ( .A(A[5]), .B(B[18]), .Z(\_8_net_[23] ) );
  AND U16 ( .A(A[5]), .B(B[17]), .Z(\_8_net_[22] ) );
  AND U17 ( .A(A[5]), .B(B[16]), .Z(\_8_net_[21] ) );
  AND U18 ( .A(A[5]), .B(B[15]), .Z(\_8_net_[20] ) );
  AND U19 ( .A(A[5]), .B(B[14]), .Z(\_8_net_[19] ) );
  AND U20 ( .A(A[5]), .B(B[13]), .Z(\_8_net_[18] ) );
  AND U21 ( .A(A[5]), .B(B[12]), .Z(\_8_net_[17] ) );
  AND U22 ( .A(A[5]), .B(B[11]), .Z(\_8_net_[16] ) );
  AND U23 ( .A(A[5]), .B(B[10]), .Z(\_8_net_[15] ) );
  AND U24 ( .A(A[5]), .B(B[9]), .Z(\_8_net_[14] ) );
  AND U25 ( .A(A[5]), .B(B[8]), .Z(\_8_net_[13] ) );
  AND U26 ( .A(A[5]), .B(B[7]), .Z(\_8_net_[12] ) );
  AND U27 ( .A(A[5]), .B(B[6]), .Z(\_8_net_[11] ) );
  AND U28 ( .A(A[5]), .B(B[5]), .Z(\_8_net_[10] ) );
  AND U29 ( .A(B[5]), .B(A[4]), .Z(\_6_net_[9] ) );
  AND U30 ( .A(B[4]), .B(A[4]), .Z(\_6_net_[8] ) );
  AND U31 ( .A(B[3]), .B(A[4]), .Z(\_6_net_[7] ) );
  AND U32 ( .A(B[2]), .B(A[4]), .Z(\_6_net_[6] ) );
  AND U33 ( .A(B[1]), .B(A[4]), .Z(\_6_net_[5] ) );
  AND U34 ( .A(B[0]), .B(A[4]), .Z(\_6_net_[4] ) );
  AND U35 ( .A(A[4]), .B(B[27]), .Z(\_6_net_[31] ) );
  AND U36 ( .A(B[26]), .B(A[4]), .Z(\_6_net_[30] ) );
  AND U37 ( .A(B[25]), .B(A[4]), .Z(\_6_net_[29] ) );
  AND U38 ( .A(B[24]), .B(A[4]), .Z(\_6_net_[28] ) );
  AND U39 ( .A(B[23]), .B(A[4]), .Z(\_6_net_[27] ) );
  AND U40 ( .A(B[22]), .B(A[4]), .Z(\_6_net_[26] ) );
  AND U41 ( .A(B[21]), .B(A[4]), .Z(\_6_net_[25] ) );
  AND U42 ( .A(B[20]), .B(A[4]), .Z(\_6_net_[24] ) );
  AND U43 ( .A(B[19]), .B(A[4]), .Z(\_6_net_[23] ) );
  AND U44 ( .A(B[18]), .B(A[4]), .Z(\_6_net_[22] ) );
  AND U45 ( .A(B[17]), .B(A[4]), .Z(\_6_net_[21] ) );
  AND U46 ( .A(B[16]), .B(A[4]), .Z(\_6_net_[20] ) );
  AND U47 ( .A(B[15]), .B(A[4]), .Z(\_6_net_[19] ) );
  AND U48 ( .A(B[14]), .B(A[4]), .Z(\_6_net_[18] ) );
  AND U49 ( .A(B[13]), .B(A[4]), .Z(\_6_net_[17] ) );
  AND U50 ( .A(B[12]), .B(A[4]), .Z(\_6_net_[16] ) );
  AND U51 ( .A(B[11]), .B(A[4]), .Z(\_6_net_[15] ) );
  AND U52 ( .A(B[10]), .B(A[4]), .Z(\_6_net_[14] ) );
  AND U53 ( .A(B[9]), .B(A[4]), .Z(\_6_net_[13] ) );
  AND U54 ( .A(B[8]), .B(A[4]), .Z(\_6_net_[12] ) );
  AND U55 ( .A(B[7]), .B(A[4]), .Z(\_6_net_[11] ) );
  AND U56 ( .A(B[6]), .B(A[4]), .Z(\_6_net_[10] ) );
  AND U57 ( .A(A[31]), .B(B[0]), .Z(\_60_net_[31] ) );
  AND U58 ( .A(B[1]), .B(A[30]), .Z(\_58_net_[31] ) );
  AND U59 ( .A(A[30]), .B(B[0]), .Z(\_58_net_[30] ) );
  AND U60 ( .A(B[2]), .B(A[29]), .Z(\_56_net_[31] ) );
  AND U61 ( .A(B[1]), .B(A[29]), .Z(\_56_net_[30] ) );
  AND U62 ( .A(A[29]), .B(B[0]), .Z(\_56_net_[29] ) );
  AND U63 ( .A(B[3]), .B(A[28]), .Z(\_54_net_[31] ) );
  AND U64 ( .A(B[2]), .B(A[28]), .Z(\_54_net_[30] ) );
  AND U65 ( .A(B[1]), .B(A[28]), .Z(\_54_net_[29] ) );
  AND U66 ( .A(A[28]), .B(B[0]), .Z(\_54_net_[28] ) );
  AND U67 ( .A(B[4]), .B(A[27]), .Z(\_52_net_[31] ) );
  AND U68 ( .A(B[3]), .B(A[27]), .Z(\_52_net_[30] ) );
  AND U69 ( .A(B[2]), .B(A[27]), .Z(\_52_net_[29] ) );
  AND U70 ( .A(B[1]), .B(A[27]), .Z(\_52_net_[28] ) );
  AND U71 ( .A(A[27]), .B(B[0]), .Z(\_52_net_[27] ) );
  AND U72 ( .A(B[5]), .B(A[26]), .Z(\_50_net_[31] ) );
  AND U73 ( .A(B[4]), .B(A[26]), .Z(\_50_net_[30] ) );
  AND U74 ( .A(B[3]), .B(A[26]), .Z(\_50_net_[29] ) );
  AND U75 ( .A(B[2]), .B(A[26]), .Z(\_50_net_[28] ) );
  AND U76 ( .A(B[1]), .B(A[26]), .Z(\_50_net_[27] ) );
  AND U77 ( .A(A[26]), .B(B[0]), .Z(\_50_net_[26] ) );
  AND U78 ( .A(B[6]), .B(A[3]), .Z(\_4_net_[9] ) );
  AND U79 ( .A(B[5]), .B(A[3]), .Z(\_4_net_[8] ) );
  AND U80 ( .A(B[4]), .B(A[3]), .Z(\_4_net_[7] ) );
  AND U81 ( .A(B[3]), .B(A[3]), .Z(\_4_net_[6] ) );
  AND U82 ( .A(B[2]), .B(A[3]), .Z(\_4_net_[5] ) );
  AND U83 ( .A(B[1]), .B(A[3]), .Z(\_4_net_[4] ) );
  AND U84 ( .A(B[0]), .B(A[3]), .Z(\_4_net_[3] ) );
  AND U85 ( .A(A[3]), .B(B[28]), .Z(\_4_net_[31] ) );
  AND U86 ( .A(B[27]), .B(A[3]), .Z(\_4_net_[30] ) );
  AND U87 ( .A(B[26]), .B(A[3]), .Z(\_4_net_[29] ) );
  AND U88 ( .A(B[25]), .B(A[3]), .Z(\_4_net_[28] ) );
  AND U89 ( .A(B[24]), .B(A[3]), .Z(\_4_net_[27] ) );
  AND U90 ( .A(B[23]), .B(A[3]), .Z(\_4_net_[26] ) );
  AND U91 ( .A(B[22]), .B(A[3]), .Z(\_4_net_[25] ) );
  AND U92 ( .A(B[21]), .B(A[3]), .Z(\_4_net_[24] ) );
  AND U93 ( .A(B[20]), .B(A[3]), .Z(\_4_net_[23] ) );
  AND U94 ( .A(B[19]), .B(A[3]), .Z(\_4_net_[22] ) );
  AND U95 ( .A(B[18]), .B(A[3]), .Z(\_4_net_[21] ) );
  AND U96 ( .A(B[17]), .B(A[3]), .Z(\_4_net_[20] ) );
  AND U97 ( .A(B[16]), .B(A[3]), .Z(\_4_net_[19] ) );
  AND U98 ( .A(B[15]), .B(A[3]), .Z(\_4_net_[18] ) );
  AND U99 ( .A(B[14]), .B(A[3]), .Z(\_4_net_[17] ) );
  AND U100 ( .A(B[13]), .B(A[3]), .Z(\_4_net_[16] ) );
  AND U101 ( .A(B[12]), .B(A[3]), .Z(\_4_net_[15] ) );
  AND U102 ( .A(B[11]), .B(A[3]), .Z(\_4_net_[14] ) );
  AND U103 ( .A(B[10]), .B(A[3]), .Z(\_4_net_[13] ) );
  AND U104 ( .A(B[9]), .B(A[3]), .Z(\_4_net_[12] ) );
  AND U105 ( .A(B[8]), .B(A[3]), .Z(\_4_net_[11] ) );
  AND U106 ( .A(B[7]), .B(A[3]), .Z(\_4_net_[10] ) );
  AND U107 ( .A(B[6]), .B(A[25]), .Z(\_48_net_[31] ) );
  AND U108 ( .A(B[5]), .B(A[25]), .Z(\_48_net_[30] ) );
  AND U109 ( .A(B[4]), .B(A[25]), .Z(\_48_net_[29] ) );
  AND U110 ( .A(B[3]), .B(A[25]), .Z(\_48_net_[28] ) );
  AND U111 ( .A(B[2]), .B(A[25]), .Z(\_48_net_[27] ) );
  AND U112 ( .A(B[1]), .B(A[25]), .Z(\_48_net_[26] ) );
  AND U113 ( .A(A[25]), .B(B[0]), .Z(\_48_net_[25] ) );
  AND U114 ( .A(B[7]), .B(A[24]), .Z(\_46_net_[31] ) );
  AND U115 ( .A(B[6]), .B(A[24]), .Z(\_46_net_[30] ) );
  AND U116 ( .A(B[5]), .B(A[24]), .Z(\_46_net_[29] ) );
  AND U117 ( .A(B[4]), .B(A[24]), .Z(\_46_net_[28] ) );
  AND U118 ( .A(B[3]), .B(A[24]), .Z(\_46_net_[27] ) );
  AND U119 ( .A(B[2]), .B(A[24]), .Z(\_46_net_[26] ) );
  AND U120 ( .A(B[1]), .B(A[24]), .Z(\_46_net_[25] ) );
  AND U121 ( .A(A[24]), .B(B[0]), .Z(\_46_net_[24] ) );
  AND U122 ( .A(B[8]), .B(A[23]), .Z(\_44_net_[31] ) );
  AND U123 ( .A(B[7]), .B(A[23]), .Z(\_44_net_[30] ) );
  AND U124 ( .A(B[6]), .B(A[23]), .Z(\_44_net_[29] ) );
  AND U125 ( .A(B[5]), .B(A[23]), .Z(\_44_net_[28] ) );
  AND U126 ( .A(B[4]), .B(A[23]), .Z(\_44_net_[27] ) );
  AND U127 ( .A(B[3]), .B(A[23]), .Z(\_44_net_[26] ) );
  AND U128 ( .A(B[2]), .B(A[23]), .Z(\_44_net_[25] ) );
  AND U129 ( .A(B[1]), .B(A[23]), .Z(\_44_net_[24] ) );
  AND U130 ( .A(A[23]), .B(B[0]), .Z(\_44_net_[23] ) );
  AND U131 ( .A(B[9]), .B(A[22]), .Z(\_42_net_[31] ) );
  AND U132 ( .A(B[8]), .B(A[22]), .Z(\_42_net_[30] ) );
  AND U133 ( .A(B[7]), .B(A[22]), .Z(\_42_net_[29] ) );
  AND U134 ( .A(B[6]), .B(A[22]), .Z(\_42_net_[28] ) );
  AND U135 ( .A(B[5]), .B(A[22]), .Z(\_42_net_[27] ) );
  AND U136 ( .A(B[4]), .B(A[22]), .Z(\_42_net_[26] ) );
  AND U137 ( .A(B[3]), .B(A[22]), .Z(\_42_net_[25] ) );
  AND U138 ( .A(B[2]), .B(A[22]), .Z(\_42_net_[24] ) );
  AND U139 ( .A(B[1]), .B(A[22]), .Z(\_42_net_[23] ) );
  AND U140 ( .A(A[22]), .B(B[0]), .Z(\_42_net_[22] ) );
  AND U141 ( .A(B[10]), .B(A[21]), .Z(\_40_net_[31] ) );
  AND U142 ( .A(B[9]), .B(A[21]), .Z(\_40_net_[30] ) );
  AND U143 ( .A(B[8]), .B(A[21]), .Z(\_40_net_[29] ) );
  AND U144 ( .A(B[7]), .B(A[21]), .Z(\_40_net_[28] ) );
  AND U145 ( .A(B[6]), .B(A[21]), .Z(\_40_net_[27] ) );
  AND U146 ( .A(B[5]), .B(A[21]), .Z(\_40_net_[26] ) );
  AND U147 ( .A(B[4]), .B(A[21]), .Z(\_40_net_[25] ) );
  AND U148 ( .A(B[3]), .B(A[21]), .Z(\_40_net_[24] ) );
  AND U149 ( .A(B[2]), .B(A[21]), .Z(\_40_net_[23] ) );
  AND U150 ( .A(B[1]), .B(A[21]), .Z(\_40_net_[22] ) );
  AND U151 ( .A(A[21]), .B(B[0]), .Z(\_40_net_[21] ) );
  AND U152 ( .A(B[11]), .B(A[20]), .Z(\_38_net_[31] ) );
  AND U153 ( .A(B[10]), .B(A[20]), .Z(\_38_net_[30] ) );
  AND U154 ( .A(B[9]), .B(A[20]), .Z(\_38_net_[29] ) );
  AND U155 ( .A(B[8]), .B(A[20]), .Z(\_38_net_[28] ) );
  AND U156 ( .A(B[7]), .B(A[20]), .Z(\_38_net_[27] ) );
  AND U157 ( .A(B[6]), .B(A[20]), .Z(\_38_net_[26] ) );
  AND U158 ( .A(B[5]), .B(A[20]), .Z(\_38_net_[25] ) );
  AND U159 ( .A(B[4]), .B(A[20]), .Z(\_38_net_[24] ) );
  AND U160 ( .A(B[3]), .B(A[20]), .Z(\_38_net_[23] ) );
  AND U161 ( .A(B[2]), .B(A[20]), .Z(\_38_net_[22] ) );
  AND U162 ( .A(B[1]), .B(A[20]), .Z(\_38_net_[21] ) );
  AND U163 ( .A(A[20]), .B(B[0]), .Z(\_38_net_[20] ) );
  AND U164 ( .A(B[12]), .B(A[19]), .Z(\_36_net_[31] ) );
  AND U165 ( .A(B[11]), .B(A[19]), .Z(\_36_net_[30] ) );
  AND U166 ( .A(B[10]), .B(A[19]), .Z(\_36_net_[29] ) );
  AND U167 ( .A(B[9]), .B(A[19]), .Z(\_36_net_[28] ) );
  AND U168 ( .A(B[8]), .B(A[19]), .Z(\_36_net_[27] ) );
  AND U169 ( .A(B[7]), .B(A[19]), .Z(\_36_net_[26] ) );
  AND U170 ( .A(B[6]), .B(A[19]), .Z(\_36_net_[25] ) );
  AND U171 ( .A(B[5]), .B(A[19]), .Z(\_36_net_[24] ) );
  AND U172 ( .A(B[4]), .B(A[19]), .Z(\_36_net_[23] ) );
  AND U173 ( .A(B[3]), .B(A[19]), .Z(\_36_net_[22] ) );
  AND U174 ( .A(B[2]), .B(A[19]), .Z(\_36_net_[21] ) );
  AND U175 ( .A(B[1]), .B(A[19]), .Z(\_36_net_[20] ) );
  AND U176 ( .A(A[19]), .B(B[0]), .Z(\_36_net_[19] ) );
  AND U177 ( .A(B[13]), .B(A[18]), .Z(\_34_net_[31] ) );
  AND U178 ( .A(B[12]), .B(A[18]), .Z(\_34_net_[30] ) );
  AND U179 ( .A(B[11]), .B(A[18]), .Z(\_34_net_[29] ) );
  AND U180 ( .A(B[10]), .B(A[18]), .Z(\_34_net_[28] ) );
  AND U181 ( .A(B[9]), .B(A[18]), .Z(\_34_net_[27] ) );
  AND U182 ( .A(B[8]), .B(A[18]), .Z(\_34_net_[26] ) );
  AND U183 ( .A(B[7]), .B(A[18]), .Z(\_34_net_[25] ) );
  AND U184 ( .A(B[6]), .B(A[18]), .Z(\_34_net_[24] ) );
  AND U185 ( .A(B[5]), .B(A[18]), .Z(\_34_net_[23] ) );
  AND U186 ( .A(B[4]), .B(A[18]), .Z(\_34_net_[22] ) );
  AND U187 ( .A(B[3]), .B(A[18]), .Z(\_34_net_[21] ) );
  AND U188 ( .A(B[2]), .B(A[18]), .Z(\_34_net_[20] ) );
  AND U189 ( .A(B[1]), .B(A[18]), .Z(\_34_net_[19] ) );
  AND U190 ( .A(A[18]), .B(B[0]), .Z(\_34_net_[18] ) );
  AND U191 ( .A(B[14]), .B(A[17]), .Z(\_32_net_[31] ) );
  AND U192 ( .A(B[13]), .B(A[17]), .Z(\_32_net_[30] ) );
  AND U193 ( .A(B[12]), .B(A[17]), .Z(\_32_net_[29] ) );
  AND U194 ( .A(B[11]), .B(A[17]), .Z(\_32_net_[28] ) );
  AND U195 ( .A(B[10]), .B(A[17]), .Z(\_32_net_[27] ) );
  AND U196 ( .A(B[9]), .B(A[17]), .Z(\_32_net_[26] ) );
  AND U197 ( .A(B[8]), .B(A[17]), .Z(\_32_net_[25] ) );
  AND U198 ( .A(B[7]), .B(A[17]), .Z(\_32_net_[24] ) );
  AND U199 ( .A(B[6]), .B(A[17]), .Z(\_32_net_[23] ) );
  AND U200 ( .A(B[5]), .B(A[17]), .Z(\_32_net_[22] ) );
  AND U201 ( .A(B[4]), .B(A[17]), .Z(\_32_net_[21] ) );
  AND U202 ( .A(B[3]), .B(A[17]), .Z(\_32_net_[20] ) );
  AND U203 ( .A(B[2]), .B(A[17]), .Z(\_32_net_[19] ) );
  AND U204 ( .A(B[1]), .B(A[17]), .Z(\_32_net_[18] ) );
  AND U205 ( .A(A[17]), .B(B[0]), .Z(\_32_net_[17] ) );
  AND U206 ( .A(B[15]), .B(A[16]), .Z(\_30_net_[31] ) );
  AND U207 ( .A(B[14]), .B(A[16]), .Z(\_30_net_[30] ) );
  AND U208 ( .A(B[13]), .B(A[16]), .Z(\_30_net_[29] ) );
  AND U209 ( .A(B[12]), .B(A[16]), .Z(\_30_net_[28] ) );
  AND U210 ( .A(B[11]), .B(A[16]), .Z(\_30_net_[27] ) );
  AND U211 ( .A(B[10]), .B(A[16]), .Z(\_30_net_[26] ) );
  AND U212 ( .A(B[9]), .B(A[16]), .Z(\_30_net_[25] ) );
  AND U213 ( .A(B[8]), .B(A[16]), .Z(\_30_net_[24] ) );
  AND U214 ( .A(B[7]), .B(A[16]), .Z(\_30_net_[23] ) );
  AND U215 ( .A(B[6]), .B(A[16]), .Z(\_30_net_[22] ) );
  AND U216 ( .A(B[5]), .B(A[16]), .Z(\_30_net_[21] ) );
  AND U217 ( .A(B[4]), .B(A[16]), .Z(\_30_net_[20] ) );
  AND U218 ( .A(B[3]), .B(A[16]), .Z(\_30_net_[19] ) );
  AND U219 ( .A(B[2]), .B(A[16]), .Z(\_30_net_[18] ) );
  AND U220 ( .A(B[1]), .B(A[16]), .Z(\_30_net_[17] ) );
  AND U221 ( .A(A[16]), .B(B[0]), .Z(\_30_net_[16] ) );
  AND U222 ( .A(B[7]), .B(A[2]), .Z(\_2_net_[9] ) );
  AND U223 ( .A(B[6]), .B(A[2]), .Z(\_2_net_[8] ) );
  AND U224 ( .A(B[5]), .B(A[2]), .Z(\_2_net_[7] ) );
  AND U225 ( .A(B[4]), .B(A[2]), .Z(\_2_net_[6] ) );
  AND U226 ( .A(B[3]), .B(A[2]), .Z(\_2_net_[5] ) );
  AND U227 ( .A(B[2]), .B(A[2]), .Z(\_2_net_[4] ) );
  AND U228 ( .A(B[1]), .B(A[2]), .Z(\_2_net_[3] ) );
  AND U229 ( .A(A[2]), .B(B[29]), .Z(\_2_net_[31] ) );
  AND U230 ( .A(B[28]), .B(A[2]), .Z(\_2_net_[30] ) );
  AND U231 ( .A(B[0]), .B(A[2]), .Z(\_2_net_[2] ) );
  AND U232 ( .A(B[27]), .B(A[2]), .Z(\_2_net_[29] ) );
  AND U233 ( .A(B[26]), .B(A[2]), .Z(\_2_net_[28] ) );
  AND U234 ( .A(B[25]), .B(A[2]), .Z(\_2_net_[27] ) );
  AND U235 ( .A(B[24]), .B(A[2]), .Z(\_2_net_[26] ) );
  AND U236 ( .A(B[23]), .B(A[2]), .Z(\_2_net_[25] ) );
  AND U237 ( .A(B[22]), .B(A[2]), .Z(\_2_net_[24] ) );
  AND U238 ( .A(B[21]), .B(A[2]), .Z(\_2_net_[23] ) );
  AND U239 ( .A(B[20]), .B(A[2]), .Z(\_2_net_[22] ) );
  AND U240 ( .A(B[19]), .B(A[2]), .Z(\_2_net_[21] ) );
  AND U241 ( .A(B[18]), .B(A[2]), .Z(\_2_net_[20] ) );
  AND U242 ( .A(B[17]), .B(A[2]), .Z(\_2_net_[19] ) );
  AND U243 ( .A(B[16]), .B(A[2]), .Z(\_2_net_[18] ) );
  AND U244 ( .A(B[15]), .B(A[2]), .Z(\_2_net_[17] ) );
  AND U245 ( .A(B[14]), .B(A[2]), .Z(\_2_net_[16] ) );
  AND U246 ( .A(B[13]), .B(A[2]), .Z(\_2_net_[15] ) );
  AND U247 ( .A(B[12]), .B(A[2]), .Z(\_2_net_[14] ) );
  AND U248 ( .A(B[11]), .B(A[2]), .Z(\_2_net_[13] ) );
  AND U249 ( .A(B[10]), .B(A[2]), .Z(\_2_net_[12] ) );
  AND U250 ( .A(B[9]), .B(A[2]), .Z(\_2_net_[11] ) );
  AND U251 ( .A(B[8]), .B(A[2]), .Z(\_2_net_[10] ) );
  AND U252 ( .A(B[16]), .B(A[15]), .Z(\_28_net_[31] ) );
  AND U253 ( .A(B[15]), .B(A[15]), .Z(\_28_net_[30] ) );
  AND U254 ( .A(B[14]), .B(A[15]), .Z(\_28_net_[29] ) );
  AND U255 ( .A(B[13]), .B(A[15]), .Z(\_28_net_[28] ) );
  AND U256 ( .A(B[12]), .B(A[15]), .Z(\_28_net_[27] ) );
  AND U257 ( .A(B[11]), .B(A[15]), .Z(\_28_net_[26] ) );
  AND U258 ( .A(B[10]), .B(A[15]), .Z(\_28_net_[25] ) );
  AND U259 ( .A(B[9]), .B(A[15]), .Z(\_28_net_[24] ) );
  AND U260 ( .A(B[8]), .B(A[15]), .Z(\_28_net_[23] ) );
  AND U261 ( .A(B[7]), .B(A[15]), .Z(\_28_net_[22] ) );
  AND U262 ( .A(B[6]), .B(A[15]), .Z(\_28_net_[21] ) );
  AND U263 ( .A(B[5]), .B(A[15]), .Z(\_28_net_[20] ) );
  AND U264 ( .A(B[4]), .B(A[15]), .Z(\_28_net_[19] ) );
  AND U265 ( .A(B[3]), .B(A[15]), .Z(\_28_net_[18] ) );
  AND U266 ( .A(B[2]), .B(A[15]), .Z(\_28_net_[17] ) );
  AND U267 ( .A(B[1]), .B(A[15]), .Z(\_28_net_[16] ) );
  AND U268 ( .A(A[15]), .B(B[0]), .Z(\_28_net_[15] ) );
  AND U269 ( .A(B[17]), .B(A[14]), .Z(\_26_net_[31] ) );
  AND U270 ( .A(B[16]), .B(A[14]), .Z(\_26_net_[30] ) );
  AND U271 ( .A(B[15]), .B(A[14]), .Z(\_26_net_[29] ) );
  AND U272 ( .A(B[14]), .B(A[14]), .Z(\_26_net_[28] ) );
  AND U273 ( .A(B[13]), .B(A[14]), .Z(\_26_net_[27] ) );
  AND U274 ( .A(B[12]), .B(A[14]), .Z(\_26_net_[26] ) );
  AND U275 ( .A(B[11]), .B(A[14]), .Z(\_26_net_[25] ) );
  AND U276 ( .A(B[10]), .B(A[14]), .Z(\_26_net_[24] ) );
  AND U277 ( .A(B[9]), .B(A[14]), .Z(\_26_net_[23] ) );
  AND U278 ( .A(B[8]), .B(A[14]), .Z(\_26_net_[22] ) );
  AND U279 ( .A(B[7]), .B(A[14]), .Z(\_26_net_[21] ) );
  AND U280 ( .A(B[6]), .B(A[14]), .Z(\_26_net_[20] ) );
  AND U281 ( .A(B[5]), .B(A[14]), .Z(\_26_net_[19] ) );
  AND U282 ( .A(B[4]), .B(A[14]), .Z(\_26_net_[18] ) );
  AND U283 ( .A(B[3]), .B(A[14]), .Z(\_26_net_[17] ) );
  AND U284 ( .A(B[2]), .B(A[14]), .Z(\_26_net_[16] ) );
  AND U285 ( .A(B[1]), .B(A[14]), .Z(\_26_net_[15] ) );
  AND U286 ( .A(A[14]), .B(B[0]), .Z(\_26_net_[14] ) );
  AND U287 ( .A(B[18]), .B(A[13]), .Z(\_24_net_[31] ) );
  AND U288 ( .A(B[17]), .B(A[13]), .Z(\_24_net_[30] ) );
  AND U289 ( .A(B[16]), .B(A[13]), .Z(\_24_net_[29] ) );
  AND U290 ( .A(B[15]), .B(A[13]), .Z(\_24_net_[28] ) );
  AND U291 ( .A(B[14]), .B(A[13]), .Z(\_24_net_[27] ) );
  AND U292 ( .A(B[13]), .B(A[13]), .Z(\_24_net_[26] ) );
  AND U293 ( .A(B[12]), .B(A[13]), .Z(\_24_net_[25] ) );
  AND U294 ( .A(B[11]), .B(A[13]), .Z(\_24_net_[24] ) );
  AND U295 ( .A(B[10]), .B(A[13]), .Z(\_24_net_[23] ) );
  AND U296 ( .A(B[9]), .B(A[13]), .Z(\_24_net_[22] ) );
  AND U297 ( .A(B[8]), .B(A[13]), .Z(\_24_net_[21] ) );
  AND U298 ( .A(B[7]), .B(A[13]), .Z(\_24_net_[20] ) );
  AND U299 ( .A(B[6]), .B(A[13]), .Z(\_24_net_[19] ) );
  AND U300 ( .A(B[5]), .B(A[13]), .Z(\_24_net_[18] ) );
  AND U301 ( .A(B[4]), .B(A[13]), .Z(\_24_net_[17] ) );
  AND U302 ( .A(B[3]), .B(A[13]), .Z(\_24_net_[16] ) );
  AND U303 ( .A(B[2]), .B(A[13]), .Z(\_24_net_[15] ) );
  AND U304 ( .A(B[1]), .B(A[13]), .Z(\_24_net_[14] ) );
  AND U305 ( .A(A[13]), .B(B[0]), .Z(\_24_net_[13] ) );
  AND U306 ( .A(B[19]), .B(A[12]), .Z(\_22_net_[31] ) );
  AND U307 ( .A(B[18]), .B(A[12]), .Z(\_22_net_[30] ) );
  AND U308 ( .A(B[17]), .B(A[12]), .Z(\_22_net_[29] ) );
  AND U309 ( .A(B[16]), .B(A[12]), .Z(\_22_net_[28] ) );
  AND U310 ( .A(B[15]), .B(A[12]), .Z(\_22_net_[27] ) );
  AND U311 ( .A(B[14]), .B(A[12]), .Z(\_22_net_[26] ) );
  AND U312 ( .A(B[13]), .B(A[12]), .Z(\_22_net_[25] ) );
  AND U313 ( .A(B[12]), .B(A[12]), .Z(\_22_net_[24] ) );
  AND U314 ( .A(B[11]), .B(A[12]), .Z(\_22_net_[23] ) );
  AND U315 ( .A(B[10]), .B(A[12]), .Z(\_22_net_[22] ) );
  AND U316 ( .A(B[9]), .B(A[12]), .Z(\_22_net_[21] ) );
  AND U317 ( .A(B[8]), .B(A[12]), .Z(\_22_net_[20] ) );
  AND U318 ( .A(B[7]), .B(A[12]), .Z(\_22_net_[19] ) );
  AND U319 ( .A(B[6]), .B(A[12]), .Z(\_22_net_[18] ) );
  AND U320 ( .A(B[5]), .B(A[12]), .Z(\_22_net_[17] ) );
  AND U321 ( .A(B[4]), .B(A[12]), .Z(\_22_net_[16] ) );
  AND U322 ( .A(B[3]), .B(A[12]), .Z(\_22_net_[15] ) );
  AND U323 ( .A(B[2]), .B(A[12]), .Z(\_22_net_[14] ) );
  AND U324 ( .A(B[1]), .B(A[12]), .Z(\_22_net_[13] ) );
  AND U325 ( .A(A[12]), .B(B[0]), .Z(\_22_net_[12] ) );
  AND U326 ( .A(B[20]), .B(A[11]), .Z(\_20_net_[31] ) );
  AND U327 ( .A(B[19]), .B(A[11]), .Z(\_20_net_[30] ) );
  AND U328 ( .A(B[18]), .B(A[11]), .Z(\_20_net_[29] ) );
  AND U329 ( .A(B[17]), .B(A[11]), .Z(\_20_net_[28] ) );
  AND U330 ( .A(B[16]), .B(A[11]), .Z(\_20_net_[27] ) );
  AND U331 ( .A(B[15]), .B(A[11]), .Z(\_20_net_[26] ) );
  AND U332 ( .A(B[14]), .B(A[11]), .Z(\_20_net_[25] ) );
  AND U333 ( .A(B[13]), .B(A[11]), .Z(\_20_net_[24] ) );
  AND U334 ( .A(B[12]), .B(A[11]), .Z(\_20_net_[23] ) );
  AND U335 ( .A(B[11]), .B(A[11]), .Z(\_20_net_[22] ) );
  AND U336 ( .A(B[10]), .B(A[11]), .Z(\_20_net_[21] ) );
  AND U337 ( .A(B[9]), .B(A[11]), .Z(\_20_net_[20] ) );
  AND U338 ( .A(B[8]), .B(A[11]), .Z(\_20_net_[19] ) );
  AND U339 ( .A(B[7]), .B(A[11]), .Z(\_20_net_[18] ) );
  AND U340 ( .A(B[6]), .B(A[11]), .Z(\_20_net_[17] ) );
  AND U341 ( .A(B[5]), .B(A[11]), .Z(\_20_net_[16] ) );
  AND U342 ( .A(B[4]), .B(A[11]), .Z(\_20_net_[15] ) );
  AND U343 ( .A(B[3]), .B(A[11]), .Z(\_20_net_[14] ) );
  AND U344 ( .A(B[2]), .B(A[11]), .Z(\_20_net_[13] ) );
  AND U345 ( .A(B[1]), .B(A[11]), .Z(\_20_net_[12] ) );
  AND U346 ( .A(A[11]), .B(B[0]), .Z(\_20_net_[11] ) );
  AND U347 ( .A(B[21]), .B(A[10]), .Z(\_18_net_[31] ) );
  AND U348 ( .A(B[20]), .B(A[10]), .Z(\_18_net_[30] ) );
  AND U349 ( .A(B[19]), .B(A[10]), .Z(\_18_net_[29] ) );
  AND U350 ( .A(B[18]), .B(A[10]), .Z(\_18_net_[28] ) );
  AND U351 ( .A(B[17]), .B(A[10]), .Z(\_18_net_[27] ) );
  AND U352 ( .A(B[16]), .B(A[10]), .Z(\_18_net_[26] ) );
  AND U353 ( .A(B[15]), .B(A[10]), .Z(\_18_net_[25] ) );
  AND U354 ( .A(B[14]), .B(A[10]), .Z(\_18_net_[24] ) );
  AND U355 ( .A(B[13]), .B(A[10]), .Z(\_18_net_[23] ) );
  AND U356 ( .A(B[12]), .B(A[10]), .Z(\_18_net_[22] ) );
  AND U357 ( .A(B[11]), .B(A[10]), .Z(\_18_net_[21] ) );
  AND U358 ( .A(B[10]), .B(A[10]), .Z(\_18_net_[20] ) );
  AND U359 ( .A(B[9]), .B(A[10]), .Z(\_18_net_[19] ) );
  AND U360 ( .A(B[8]), .B(A[10]), .Z(\_18_net_[18] ) );
  AND U361 ( .A(B[7]), .B(A[10]), .Z(\_18_net_[17] ) );
  AND U362 ( .A(B[6]), .B(A[10]), .Z(\_18_net_[16] ) );
  AND U363 ( .A(B[5]), .B(A[10]), .Z(\_18_net_[15] ) );
  AND U364 ( .A(B[4]), .B(A[10]), .Z(\_18_net_[14] ) );
  AND U365 ( .A(B[3]), .B(A[10]), .Z(\_18_net_[13] ) );
  AND U366 ( .A(B[2]), .B(A[10]), .Z(\_18_net_[12] ) );
  AND U367 ( .A(B[1]), .B(A[10]), .Z(\_18_net_[11] ) );
  AND U368 ( .A(A[10]), .B(B[0]), .Z(\_18_net_[10] ) );
  AND U369 ( .A(B[0]), .B(A[9]), .Z(\_16_net_[9] ) );
  AND U370 ( .A(B[22]), .B(A[9]), .Z(\_16_net_[31] ) );
  AND U371 ( .A(B[21]), .B(A[9]), .Z(\_16_net_[30] ) );
  AND U372 ( .A(B[20]), .B(A[9]), .Z(\_16_net_[29] ) );
  AND U373 ( .A(B[19]), .B(A[9]), .Z(\_16_net_[28] ) );
  AND U374 ( .A(B[18]), .B(A[9]), .Z(\_16_net_[27] ) );
  AND U375 ( .A(B[17]), .B(A[9]), .Z(\_16_net_[26] ) );
  AND U376 ( .A(B[16]), .B(A[9]), .Z(\_16_net_[25] ) );
  AND U377 ( .A(B[15]), .B(A[9]), .Z(\_16_net_[24] ) );
  AND U378 ( .A(B[14]), .B(A[9]), .Z(\_16_net_[23] ) );
  AND U379 ( .A(B[13]), .B(A[9]), .Z(\_16_net_[22] ) );
  AND U380 ( .A(B[12]), .B(A[9]), .Z(\_16_net_[21] ) );
  AND U381 ( .A(B[11]), .B(A[9]), .Z(\_16_net_[20] ) );
  AND U382 ( .A(B[10]), .B(A[9]), .Z(\_16_net_[19] ) );
  AND U383 ( .A(B[9]), .B(A[9]), .Z(\_16_net_[18] ) );
  AND U384 ( .A(B[8]), .B(A[9]), .Z(\_16_net_[17] ) );
  AND U385 ( .A(B[7]), .B(A[9]), .Z(\_16_net_[16] ) );
  AND U386 ( .A(B[6]), .B(A[9]), .Z(\_16_net_[15] ) );
  AND U387 ( .A(B[5]), .B(A[9]), .Z(\_16_net_[14] ) );
  AND U388 ( .A(B[4]), .B(A[9]), .Z(\_16_net_[13] ) );
  AND U389 ( .A(B[3]), .B(A[9]), .Z(\_16_net_[12] ) );
  AND U390 ( .A(B[2]), .B(A[9]), .Z(\_16_net_[11] ) );
  AND U391 ( .A(A[9]), .B(B[1]), .Z(\_16_net_[10] ) );
  AND U392 ( .A(B[1]), .B(A[8]), .Z(\_14_net_[9] ) );
  AND U393 ( .A(B[0]), .B(A[8]), .Z(\_14_net_[8] ) );
  AND U394 ( .A(B[23]), .B(A[8]), .Z(\_14_net_[31] ) );
  AND U395 ( .A(B[22]), .B(A[8]), .Z(\_14_net_[30] ) );
  AND U396 ( .A(B[21]), .B(A[8]), .Z(\_14_net_[29] ) );
  AND U397 ( .A(B[20]), .B(A[8]), .Z(\_14_net_[28] ) );
  AND U398 ( .A(B[19]), .B(A[8]), .Z(\_14_net_[27] ) );
  AND U399 ( .A(B[18]), .B(A[8]), .Z(\_14_net_[26] ) );
  AND U400 ( .A(B[17]), .B(A[8]), .Z(\_14_net_[25] ) );
  AND U401 ( .A(B[16]), .B(A[8]), .Z(\_14_net_[24] ) );
  AND U402 ( .A(B[15]), .B(A[8]), .Z(\_14_net_[23] ) );
  AND U403 ( .A(B[14]), .B(A[8]), .Z(\_14_net_[22] ) );
  AND U404 ( .A(B[13]), .B(A[8]), .Z(\_14_net_[21] ) );
  AND U405 ( .A(B[12]), .B(A[8]), .Z(\_14_net_[20] ) );
  AND U406 ( .A(B[11]), .B(A[8]), .Z(\_14_net_[19] ) );
  AND U407 ( .A(B[10]), .B(A[8]), .Z(\_14_net_[18] ) );
  AND U408 ( .A(B[9]), .B(A[8]), .Z(\_14_net_[17] ) );
  AND U409 ( .A(B[8]), .B(A[8]), .Z(\_14_net_[16] ) );
  AND U410 ( .A(B[7]), .B(A[8]), .Z(\_14_net_[15] ) );
  AND U411 ( .A(B[6]), .B(A[8]), .Z(\_14_net_[14] ) );
  AND U412 ( .A(B[5]), .B(A[8]), .Z(\_14_net_[13] ) );
  AND U413 ( .A(B[4]), .B(A[8]), .Z(\_14_net_[12] ) );
  AND U414 ( .A(B[3]), .B(A[8]), .Z(\_14_net_[11] ) );
  AND U415 ( .A(A[8]), .B(B[2]), .Z(\_14_net_[10] ) );
  AND U416 ( .A(B[2]), .B(A[7]), .Z(\_12_net_[9] ) );
  AND U417 ( .A(B[1]), .B(A[7]), .Z(\_12_net_[8] ) );
  AND U418 ( .A(B[0]), .B(A[7]), .Z(\_12_net_[7] ) );
  AND U419 ( .A(B[24]), .B(A[7]), .Z(\_12_net_[31] ) );
  AND U420 ( .A(B[23]), .B(A[7]), .Z(\_12_net_[30] ) );
  AND U421 ( .A(B[22]), .B(A[7]), .Z(\_12_net_[29] ) );
  AND U422 ( .A(B[21]), .B(A[7]), .Z(\_12_net_[28] ) );
  AND U423 ( .A(B[20]), .B(A[7]), .Z(\_12_net_[27] ) );
  AND U424 ( .A(B[19]), .B(A[7]), .Z(\_12_net_[26] ) );
  AND U425 ( .A(B[18]), .B(A[7]), .Z(\_12_net_[25] ) );
  AND U426 ( .A(B[17]), .B(A[7]), .Z(\_12_net_[24] ) );
  AND U427 ( .A(B[16]), .B(A[7]), .Z(\_12_net_[23] ) );
  AND U428 ( .A(B[15]), .B(A[7]), .Z(\_12_net_[22] ) );
  AND U429 ( .A(B[14]), .B(A[7]), .Z(\_12_net_[21] ) );
  AND U430 ( .A(B[13]), .B(A[7]), .Z(\_12_net_[20] ) );
  AND U431 ( .A(B[12]), .B(A[7]), .Z(\_12_net_[19] ) );
  AND U432 ( .A(B[11]), .B(A[7]), .Z(\_12_net_[18] ) );
  AND U433 ( .A(B[10]), .B(A[7]), .Z(\_12_net_[17] ) );
  AND U434 ( .A(B[9]), .B(A[7]), .Z(\_12_net_[16] ) );
  AND U435 ( .A(B[8]), .B(A[7]), .Z(\_12_net_[15] ) );
  AND U436 ( .A(B[7]), .B(A[7]), .Z(\_12_net_[14] ) );
  AND U437 ( .A(B[6]), .B(A[7]), .Z(\_12_net_[13] ) );
  AND U438 ( .A(B[5]), .B(A[7]), .Z(\_12_net_[12] ) );
  AND U439 ( .A(B[4]), .B(A[7]), .Z(\_12_net_[11] ) );
  AND U440 ( .A(A[7]), .B(B[3]), .Z(\_12_net_[10] ) );
  AND U441 ( .A(B[3]), .B(A[6]), .Z(\_10_net_[9] ) );
  AND U442 ( .A(B[2]), .B(A[6]), .Z(\_10_net_[8] ) );
  AND U443 ( .A(B[1]), .B(A[6]), .Z(\_10_net_[7] ) );
  AND U444 ( .A(B[0]), .B(A[6]), .Z(\_10_net_[6] ) );
  AND U445 ( .A(B[25]), .B(A[6]), .Z(\_10_net_[31] ) );
  AND U446 ( .A(B[24]), .B(A[6]), .Z(\_10_net_[30] ) );
  AND U447 ( .A(B[23]), .B(A[6]), .Z(\_10_net_[29] ) );
  AND U448 ( .A(B[22]), .B(A[6]), .Z(\_10_net_[28] ) );
  AND U449 ( .A(B[21]), .B(A[6]), .Z(\_10_net_[27] ) );
  AND U450 ( .A(B[20]), .B(A[6]), .Z(\_10_net_[26] ) );
  AND U451 ( .A(B[19]), .B(A[6]), .Z(\_10_net_[25] ) );
  AND U452 ( .A(B[18]), .B(A[6]), .Z(\_10_net_[24] ) );
  AND U453 ( .A(B[17]), .B(A[6]), .Z(\_10_net_[23] ) );
  AND U454 ( .A(B[16]), .B(A[6]), .Z(\_10_net_[22] ) );
  AND U455 ( .A(B[15]), .B(A[6]), .Z(\_10_net_[21] ) );
  AND U456 ( .A(B[14]), .B(A[6]), .Z(\_10_net_[20] ) );
  AND U457 ( .A(B[13]), .B(A[6]), .Z(\_10_net_[19] ) );
  AND U458 ( .A(B[12]), .B(A[6]), .Z(\_10_net_[18] ) );
  AND U459 ( .A(B[11]), .B(A[6]), .Z(\_10_net_[17] ) );
  AND U460 ( .A(B[10]), .B(A[6]), .Z(\_10_net_[16] ) );
  AND U461 ( .A(B[9]), .B(A[6]), .Z(\_10_net_[15] ) );
  AND U462 ( .A(B[8]), .B(A[6]), .Z(\_10_net_[14] ) );
  AND U463 ( .A(B[7]), .B(A[6]), .Z(\_10_net_[13] ) );
  AND U464 ( .A(B[6]), .B(A[6]), .Z(\_10_net_[12] ) );
  AND U465 ( .A(B[5]), .B(A[6]), .Z(\_10_net_[11] ) );
  AND U466 ( .A(A[6]), .B(B[4]), .Z(\_10_net_[10] ) );
  AND U467 ( .A(B[8]), .B(A[1]), .Z(\_0_net_[9] ) );
  AND U468 ( .A(B[7]), .B(A[1]), .Z(\_0_net_[8] ) );
  AND U469 ( .A(B[6]), .B(A[1]), .Z(\_0_net_[7] ) );
  AND U470 ( .A(B[5]), .B(A[1]), .Z(\_0_net_[6] ) );
  AND U471 ( .A(B[4]), .B(A[1]), .Z(\_0_net_[5] ) );
  AND U472 ( .A(B[3]), .B(A[1]), .Z(\_0_net_[4] ) );
  AND U473 ( .A(B[2]), .B(A[1]), .Z(\_0_net_[3] ) );
  AND U474 ( .A(B[30]), .B(A[1]), .Z(\_0_net_[31] ) );
  AND U475 ( .A(B[29]), .B(A[1]), .Z(\_0_net_[30] ) );
  AND U476 ( .A(B[1]), .B(A[1]), .Z(\_0_net_[2] ) );
  AND U477 ( .A(B[28]), .B(A[1]), .Z(\_0_net_[29] ) );
  AND U478 ( .A(B[27]), .B(A[1]), .Z(\_0_net_[28] ) );
  AND U479 ( .A(B[26]), .B(A[1]), .Z(\_0_net_[27] ) );
  AND U480 ( .A(B[25]), .B(A[1]), .Z(\_0_net_[26] ) );
  AND U481 ( .A(B[24]), .B(A[1]), .Z(\_0_net_[25] ) );
  AND U482 ( .A(B[23]), .B(A[1]), .Z(\_0_net_[24] ) );
  AND U483 ( .A(B[22]), .B(A[1]), .Z(\_0_net_[23] ) );
  AND U484 ( .A(B[21]), .B(A[1]), .Z(\_0_net_[22] ) );
  AND U485 ( .A(B[20]), .B(A[1]), .Z(\_0_net_[21] ) );
  AND U486 ( .A(B[19]), .B(A[1]), .Z(\_0_net_[20] ) );
  AND U487 ( .A(B[0]), .B(A[1]), .Z(\_0_net_[1] ) );
  AND U488 ( .A(B[18]), .B(A[1]), .Z(\_0_net_[19] ) );
  AND U489 ( .A(B[17]), .B(A[1]), .Z(\_0_net_[18] ) );
  AND U490 ( .A(B[16]), .B(A[1]), .Z(\_0_net_[17] ) );
  AND U491 ( .A(B[15]), .B(A[1]), .Z(\_0_net_[16] ) );
  AND U492 ( .A(B[14]), .B(A[1]), .Z(\_0_net_[15] ) );
  AND U493 ( .A(B[13]), .B(A[1]), .Z(\_0_net_[14] ) );
  AND U494 ( .A(B[12]), .B(A[1]), .Z(\_0_net_[13] ) );
  AND U495 ( .A(B[11]), .B(A[1]), .Z(\_0_net_[12] ) );
  AND U496 ( .A(B[10]), .B(A[1]), .Z(\_0_net_[11] ) );
  AND U497 ( .A(A[1]), .B(B[9]), .Z(\_0_net_[10] ) );
endmodule


module FA_993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_32 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_1023 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1022 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1021 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1020 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1019 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1018 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1017 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1016 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1015 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1014 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1013 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1012 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1011 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1010 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1009 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1008 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1007 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1006 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1005 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1004 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1003 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1002 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1001 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1000 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_999 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_998 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_997 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_996 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_995 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_994 \FAINST[30].FA_  ( .A(1'b0), .B(B[30]), .CI(1'b0), .S(S[30]) );
  FA_993 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(1'b0), .S(S[31]) );
endmodule


module FA_1025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_33 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;
  wire   \C[31] ;

  FA_1055 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1054 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1053 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1052 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1051 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1050 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1049 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1048 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1047 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1046 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1045 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1044 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1043 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1042 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1041 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1040 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1039 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1038 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1037 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1036 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1035 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1034 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1033 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1032 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1031 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_1030 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_1029 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_1028 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_1027 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_1026 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(1'b0), .S(S[30]), .CO(
        \C[31] ) );
  FA_1025 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(\C[31] ), .S(S[31]) );
endmodule


module FA_1057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_34 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1087 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1086 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1085 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1084 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1083 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1082 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1081 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1080 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1079 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1078 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1077 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1076 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1075 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1074 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1073 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1072 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1071 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1070 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1069 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1068 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1067 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1066 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1065 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1064 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1063 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_1062 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_1061 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_1060 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_1059 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(1'b0), .S(S[29]), .CO(
        C[30]) );
  FA_1058 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1057 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_35 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1119 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1118 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1117 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1116 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1115 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1114 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1113 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1112 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1111 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1110 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1109 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1108 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1107 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1106 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1105 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1104 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1103 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1102 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1101 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1100 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1099 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1098 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1097 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1096 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1095 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_1094 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_1093 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_1092 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(1'b0), .S(S[28]), .CO(
        C[29]) );
  FA_1091 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1090 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1089 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_36 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1151 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1150 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1149 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1148 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1147 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1146 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1145 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1144 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1143 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1142 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1141 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1140 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1139 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1138 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1137 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1136 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1135 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1134 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1133 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1132 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1131 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1130 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1129 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1128 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1127 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_1126 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_1125 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(1'b0), .S(S[27]), .CO(
        C[28]) );
  FA_1124 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1123 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1122 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1121 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_37 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1183 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1182 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1181 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1180 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1179 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1178 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1177 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1176 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1175 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1174 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1173 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1172 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1171 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1170 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1169 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1168 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1167 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1166 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1165 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1164 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1163 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1162 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1161 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1160 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1159 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_1158 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(1'b0), .S(S[26]), .CO(
        C[27]) );
  FA_1157 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1156 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1155 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1154 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1153 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_38 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1215 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1214 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1213 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1212 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1211 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1210 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1209 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1208 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1207 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1206 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1205 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1204 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1203 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1202 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1201 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1200 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1199 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1198 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1197 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1196 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1195 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1194 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1193 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1192 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1191 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(1'b0), .S(S[25]), .CO(
        C[26]) );
  FA_1190 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1189 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1188 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1187 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1186 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1185 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_39 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1247 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1246 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1245 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1244 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1243 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1242 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1241 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1240 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1239 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1238 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1237 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1236 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1235 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1234 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1233 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1232 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1231 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1230 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1229 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1228 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1227 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1226 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1225 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1224 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(1'b0), .S(S[24]), .CO(
        C[25]) );
  FA_1223 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1222 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1221 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1220 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1219 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1218 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1217 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_40 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1279 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1278 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1277 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1276 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1275 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1274 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1273 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1272 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1271 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1270 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1269 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1268 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1267 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1266 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1265 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1264 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1263 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1262 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1261 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1260 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1259 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1258 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1257 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(1'b0), .S(S[23]), .CO(
        C[24]) );
  FA_1256 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1255 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1254 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1253 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1252 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1251 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1250 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1249 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_41 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1311 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1310 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1309 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1308 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1307 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1306 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1305 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1304 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1303 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1302 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1301 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1300 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1299 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1298 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1297 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1296 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1295 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1294 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1293 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1292 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1291 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1290 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(1'b0), .S(S[22]), .CO(
        C[23]) );
  FA_1289 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1288 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1287 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1286 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1285 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1284 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1283 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1282 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1281 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_42 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1343 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1342 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1341 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1340 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1339 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1338 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1337 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1336 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1335 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1334 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1333 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1332 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1331 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1330 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1329 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1328 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1327 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1326 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1325 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1324 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1323 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(1'b0), .S(S[21]), .CO(
        C[22]) );
  FA_1322 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1321 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1320 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1319 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1318 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1317 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1316 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1315 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1314 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1313 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_43 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1375 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1374 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1373 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1372 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1371 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1370 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1369 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1368 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1367 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1366 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1365 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1364 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1363 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1362 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1361 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1360 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1359 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1358 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1357 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1356 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(1'b0), .S(S[20]), .CO(
        C[21]) );
  FA_1355 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1354 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1353 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1352 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1351 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1350 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1349 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1348 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1347 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1346 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1345 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_44 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1407 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1406 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1405 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1404 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1403 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1402 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1401 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1400 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1399 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1398 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1397 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1396 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1395 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1394 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1393 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1392 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1391 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1390 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1389 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(1'b0), .S(S[19]), .CO(
        C[20]) );
  FA_1388 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1387 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1386 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1385 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1384 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1383 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1382 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1381 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1380 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1379 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1378 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1377 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_45 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1439 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1438 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1437 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1436 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1435 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1434 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1433 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1432 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1431 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1430 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1429 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1428 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1427 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1426 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1425 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1424 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1423 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1422 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(1'b0), .S(S[18]), .CO(
        C[19]) );
  FA_1421 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1420 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1419 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1418 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1417 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1416 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1415 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1414 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1413 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1412 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1411 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1410 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1409 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_46 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1471 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1470 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1469 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1468 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1467 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1466 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1465 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1464 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1463 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1462 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1461 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1460 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1459 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1458 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1457 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1456 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1455 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(1'b0), .S(S[17]), .CO(
        C[18]) );
  FA_1454 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1453 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1452 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1451 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1450 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1449 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1448 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1447 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1446 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1445 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1444 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1443 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1442 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1441 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_47 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1503 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1502 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1501 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1500 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1499 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1498 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1497 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1496 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1495 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1494 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1493 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1492 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1491 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1490 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1489 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1488 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(1'b0), .S(S[16]), .CO(
        C[17]) );
  FA_1487 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1486 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1485 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1484 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1483 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1482 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1481 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1480 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1479 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1478 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1477 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1476 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1475 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1474 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1473 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_48 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1535 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1534 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1533 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1532 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1531 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1530 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1529 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1528 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1527 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1526 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1525 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1524 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1523 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1522 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1521 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(1'b0), .S(S[15]), .CO(
        C[16]) );
  FA_1520 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1519 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1518 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1517 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1516 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1515 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1514 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1513 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1512 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1511 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1510 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1509 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1508 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1507 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1506 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1505 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_49 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1567 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1566 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1565 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1564 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1563 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1562 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1561 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1560 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1559 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1558 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1557 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1556 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1555 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1554 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(1'b0), .S(S[14]), .CO(
        C[15]) );
  FA_1553 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1552 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1551 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1550 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1549 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1548 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1547 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1546 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1545 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1544 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1543 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1542 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1541 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1540 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1539 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1538 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1537 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_50 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1599 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1598 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1597 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1596 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1595 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1594 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1593 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1592 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1591 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1590 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1589 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1588 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1587 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(1'b0), .S(S[13]), .CO(
        C[14]) );
  FA_1586 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1585 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1584 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1583 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1582 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1581 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1580 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1579 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1578 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1577 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1576 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1575 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1574 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1573 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1572 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1571 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1570 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1569 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_51 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1631 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1630 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1629 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1628 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1627 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1626 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1625 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1624 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1623 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1622 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1621 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1620 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(1'b0), .S(S[12]), .CO(
        C[13]) );
  FA_1619 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1618 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1617 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1616 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1615 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1614 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1613 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1612 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1611 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1610 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1609 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1608 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1607 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1606 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1605 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1604 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1603 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1602 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1601 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_52 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1663 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1662 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1661 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1660 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1659 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1658 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1657 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1656 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1655 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1654 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1653 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(1'b0), .S(S[11]), .CO(
        C[12]) );
  FA_1652 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1651 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1650 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1649 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1648 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1647 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1646 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1645 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1644 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1643 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1642 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1641 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1640 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1639 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1638 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1637 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1636 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1635 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1634 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1633 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_53 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1695 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1694 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1693 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1692 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1691 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1690 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1689 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1688 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1687 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1686 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(1'b0), .S(S[10]), .CO(
        C[11]) );
  FA_1685 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1684 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1683 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1682 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1681 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1680 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1679 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1678 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1677 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1676 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1675 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1674 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1673 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1672 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1671 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1670 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1669 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1668 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1667 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1666 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1665 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_54 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1727 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1726 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1725 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1724 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1723 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1722 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1721 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1720 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1719 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(1'b0), .S(S[9]), .CO(C[10]) );
  FA_1718 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1717 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1716 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1715 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1714 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1713 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1712 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1711 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1710 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1709 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1708 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1707 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1706 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1705 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1704 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1703 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1702 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1701 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1700 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1699 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1698 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1697 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_55 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1759 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1758 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1757 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1756 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1755 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1754 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1753 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1752 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(1'b0), .S(S[8]), .CO(C[9])
         );
  FA_1751 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1750 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1749 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1748 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1747 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1746 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1745 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1744 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1743 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1742 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1741 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1740 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1739 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1738 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1737 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1736 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1735 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1734 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1733 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1732 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1731 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1730 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1729 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_56 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1791 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1790 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1789 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1788 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1787 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1786 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1785 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(1'b0), .S(S[7]), .CO(C[8])
         );
  FA_1784 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1783 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1782 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1781 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1780 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1779 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1778 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1777 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1776 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1775 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1774 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1773 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1772 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1771 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1770 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1769 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1768 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1767 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1766 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1765 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1764 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1763 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1762 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1761 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_57 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1823 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1822 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1821 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1820 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1819 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1818 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(1'b0), .S(S[6]), .CO(C[7])
         );
  FA_1817 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_1816 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1815 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1814 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1813 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1812 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1811 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1810 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1809 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1808 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1807 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1806 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1805 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1804 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1803 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1802 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1801 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1800 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1799 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1798 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1797 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1796 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1795 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1794 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1793 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_58 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1855 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1854 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1853 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1852 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1851 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(1'b0), .S(S[5]), .CO(C[6])
         );
  FA_1850 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_1849 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_1848 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1847 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1846 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1845 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1844 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1843 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1842 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1841 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1840 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1839 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1838 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1837 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1836 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1835 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1834 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1833 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1832 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1831 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1830 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1829 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1828 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1827 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1826 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1825 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_59 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1887 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1886 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1885 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1884 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(1'b0), .S(S[4]), .CO(C[5])
         );
  FA_1883 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_1882 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_1881 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_1880 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1879 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1878 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1877 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1876 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1875 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1874 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1873 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1872 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1871 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1870 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1869 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1868 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1867 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1866 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1865 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1864 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1863 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1862 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1861 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1860 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1859 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1858 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1857 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_60 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1919 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1918 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1917 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(1'b0), .S(S[3]), .CO(C[4])
         );
  FA_1916 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_1915 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_1914 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_1913 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_1912 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1911 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1910 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1909 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1908 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1907 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1906 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1905 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1904 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1903 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1902 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1901 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1900 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1899 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1898 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1897 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1896 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1895 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1894 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1893 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1892 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1891 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1890 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1889 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_61 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1951 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1950 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(1'b0), .S(S[2]), .CO(C[3])
         );
  FA_1949 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_1948 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_1947 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_1946 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_1945 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_1944 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1943 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1942 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1941 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1940 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1939 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1938 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1937 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1936 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1935 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1934 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1933 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1932 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1931 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1930 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1929 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1928 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1927 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1926 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1925 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1924 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1923 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1922 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1921 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module ADD_N32_62 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_1983 \FAINST[1].FA_  ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(S[1]) );
  FA_1982 \FAINST[2].FA_  ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(S[2]) );
  FA_1981 \FAINST[3].FA_  ( .A(A[3]), .B(1'b0), .CI(1'b0), .S(S[3]) );
  FA_1980 \FAINST[4].FA_  ( .A(A[4]), .B(1'b0), .CI(1'b0), .S(S[4]) );
  FA_1979 \FAINST[5].FA_  ( .A(A[5]), .B(1'b0), .CI(1'b0), .S(S[5]) );
  FA_1978 \FAINST[6].FA_  ( .A(A[6]), .B(1'b0), .CI(1'b0), .S(S[6]) );
  FA_1977 \FAINST[7].FA_  ( .A(A[7]), .B(1'b0), .CI(1'b0), .S(S[7]) );
  FA_1976 \FAINST[8].FA_  ( .A(A[8]), .B(1'b0), .CI(1'b0), .S(S[8]) );
  FA_1975 \FAINST[9].FA_  ( .A(A[9]), .B(1'b0), .CI(1'b0), .S(S[9]) );
  FA_1974 \FAINST[10].FA_  ( .A(A[10]), .B(1'b0), .CI(1'b0), .S(S[10]) );
  FA_1973 \FAINST[11].FA_  ( .A(A[11]), .B(1'b0), .CI(1'b0), .S(S[11]) );
  FA_1972 \FAINST[12].FA_  ( .A(A[12]), .B(1'b0), .CI(1'b0), .S(S[12]) );
  FA_1971 \FAINST[13].FA_  ( .A(A[13]), .B(1'b0), .CI(1'b0), .S(S[13]) );
  FA_1970 \FAINST[14].FA_  ( .A(A[14]), .B(1'b0), .CI(1'b0), .S(S[14]) );
  FA_1969 \FAINST[15].FA_  ( .A(A[15]), .B(1'b0), .CI(1'b0), .S(S[15]) );
  FA_1968 \FAINST[16].FA_  ( .A(A[16]), .B(1'b0), .CI(1'b0), .S(S[16]) );
  FA_1967 \FAINST[17].FA_  ( .A(A[17]), .B(1'b0), .CI(1'b0), .S(S[17]) );
  FA_1966 \FAINST[18].FA_  ( .A(A[18]), .B(1'b0), .CI(1'b0), .S(S[18]) );
  FA_1965 \FAINST[19].FA_  ( .A(A[19]), .B(1'b0), .CI(1'b0), .S(S[19]) );
  FA_1964 \FAINST[20].FA_  ( .A(A[20]), .B(1'b0), .CI(1'b0), .S(S[20]) );
  FA_1963 \FAINST[21].FA_  ( .A(A[21]), .B(1'b0), .CI(1'b0), .S(S[21]) );
  FA_1962 \FAINST[22].FA_  ( .A(A[22]), .B(1'b0), .CI(1'b0), .S(S[22]) );
  FA_1961 \FAINST[23].FA_  ( .A(A[23]), .B(1'b0), .CI(1'b0), .S(S[23]) );
  FA_1960 \FAINST[24].FA_  ( .A(A[24]), .B(1'b0), .CI(1'b0), .S(S[24]) );
  FA_1959 \FAINST[25].FA_  ( .A(A[25]), .B(1'b0), .CI(1'b0), .S(S[25]) );
  FA_1958 \FAINST[26].FA_  ( .A(A[26]), .B(1'b0), .CI(1'b0), .S(S[26]) );
  FA_1957 \FAINST[27].FA_  ( .A(A[27]), .B(1'b0), .CI(1'b0), .S(S[27]) );
  FA_1956 \FAINST[28].FA_  ( .A(A[28]), .B(1'b0), .CI(1'b0), .S(S[28]) );
  FA_1955 \FAINST[29].FA_  ( .A(A[29]), .B(1'b0), .CI(1'b0), .S(S[29]) );
  FA_1954 \FAINST[30].FA_  ( .A(A[30]), .B(1'b0), .CI(1'b0), .S(S[30]) );
  FA_1953 \FAINST[31].FA_  ( .A(A[31]), .B(1'b0), .CI(1'b0), .S(S[31]) );
endmodule


module MULT_N32_2 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   \w[31][31] , \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] ,
         \w[31][26] , \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] ,
         \w[31][21] , \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] ,
         \w[31][16] , \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] ,
         \w[31][11] , \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] ,
         \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] ,
         \w[31][1] , \w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] ,
         \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] ,
         \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] ,
         \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] ,
         \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] ,
         \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] ,
         \w[30][2] , \w[30][1] , \w[29][31] , \w[29][30] , \w[29][29] ,
         \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] ,
         \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] ,
         \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] ,
         \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] ,
         \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] ,
         \w[29][3] , \w[29][2] , \w[29][1] , \w[28][31] , \w[28][30] ,
         \w[28][29] , \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] ,
         \w[28][24] , \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] ,
         \w[28][19] , \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] ,
         \w[28][14] , \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] ,
         \w[28][9] , \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] ,
         \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , \w[27][31] ,
         \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] ,
         \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] ,
         \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] ,
         \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] ,
         \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] ,
         \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] ,
         \w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] ,
         \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] ,
         \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] ,
         \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] ,
         \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] ,
         \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] ,
         \w[26][1] , \w[25][31] , \w[25][30] , \w[25][29] , \w[25][28] ,
         \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , \w[25][23] ,
         \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , \w[25][18] ,
         \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , \w[25][13] ,
         \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , \w[25][8] ,
         \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] ,
         \w[25][2] , \w[25][1] , \w[24][31] , \w[24][30] , \w[24][29] ,
         \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] ,
         \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] ,
         \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] ,
         \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] ,
         \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] ,
         \w[24][3] , \w[24][2] , \w[24][1] , \w[23][31] , \w[23][30] ,
         \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] ,
         \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] ,
         \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] ,
         \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] ,
         \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] ,
         \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , \w[22][31] ,
         \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , \w[22][26] ,
         \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , \w[22][21] ,
         \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , \w[22][16] ,
         \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , \w[22][11] ,
         \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , \w[22][6] ,
         \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] ,
         \w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] ,
         \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] ,
         \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] ,
         \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] ,
         \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] ,
         \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] ,
         \w[21][1] , \w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] ,
         \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] ,
         \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] ,
         \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] ,
         \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] ,
         \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] ,
         \w[20][2] , \w[20][1] , \w[19][31] , \w[19][30] , \w[19][29] ,
         \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] ,
         \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] ,
         \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] ,
         \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] ,
         \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] ,
         \w[19][3] , \w[19][2] , \w[19][1] , \w[18][31] , \w[18][30] ,
         \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] ,
         \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] ,
         \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] ,
         \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] ,
         \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] ,
         \w[18][4] , \w[18][3] , \w[18][2] , \w[18][1] , \w[17][31] ,
         \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] ,
         \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] ,
         \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] ,
         \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] ,
         \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] ,
         \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] ,
         \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] ,
         \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] ,
         \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] ,
         \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] ,
         \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] ,
         \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] ,
         \w[16][1] , \w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] ,
         \w[15][27] , \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] ,
         \w[15][22] , \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] ,
         \w[15][17] , \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] ,
         \w[15][12] , \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] ,
         \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] ,
         \w[15][2] , \w[15][1] , \w[14][31] , \w[14][30] , \w[14][29] ,
         \w[14][28] , \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] ,
         \w[14][23] , \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] ,
         \w[14][18] , \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] ,
         \w[14][13] , \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] ,
         \w[14][8] , \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] ,
         \w[14][3] , \w[14][2] , \w[14][1] , \w[13][31] , \w[13][30] ,
         \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] ,
         \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] ,
         \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] ,
         \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] ,
         \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] ,
         \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , \w[12][31] ,
         \w[12][30] , \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] ,
         \w[12][25] , \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] ,
         \w[12][20] , \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] ,
         \w[12][15] , \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] ,
         \w[12][10] , \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] ,
         \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , \w[12][1] ,
         \w[11][31] , \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] ,
         \w[11][26] , \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] ,
         \w[11][21] , \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] ,
         \w[11][16] , \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] ,
         \w[11][11] , \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] ,
         \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] ,
         \w[11][1] , \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] ,
         \w[10][27] , \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] ,
         \w[10][22] , \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] ,
         \w[10][17] , \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] ,
         \w[10][12] , \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] ,
         \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] ,
         \w[10][2] , \w[10][1] , \w[9][31] , \w[9][30] , \w[9][29] ,
         \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] ,
         \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] ,
         \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] ,
         \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] ,
         \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] ,
         \w[9][1] , \w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] ,
         \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] ,
         \w[8][21] , \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] ,
         \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , \w[8][12] ,
         \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , \w[8][6] ,
         \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , \w[7][31] ,
         \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] ,
         \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] ,
         \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] ,
         \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] ,
         \w[7][10] , \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] ,
         \w[7][4] , \w[7][3] , \w[7][2] , \w[7][1] , \w[6][31] , \w[6][30] ,
         \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] ,
         \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] ,
         \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] ,
         \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] ,
         \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] ,
         \w[6][2] , \w[6][1] , \w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] ,
         \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] ,
         \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] ,
         \w[5][17] , \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] ,
         \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] ,
         \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] ,
         \w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] ,
         \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] ,
         \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] ,
         \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] ,
         \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] ,
         \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , \w[3][31] ,
         \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] ,
         \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] ,
         \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] ,
         \w[3][15] , \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] ,
         \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] ,
         \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , \w[2][31] , \w[2][30] ,
         \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] ,
         \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] ,
         \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] ,
         \w[2][14] , \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] ,
         \w[2][8] , \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] ,
         \w[2][2] , \w[2][1] , \_0_net_[31] , \_0_net_[30] , \_0_net_[29] ,
         \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , \_0_net_[25] ,
         \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , \_0_net_[21] ,
         \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , \_0_net_[17] ,
         \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , \_0_net_[13] ,
         \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , \_0_net_[9] ,
         \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] ,
         \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_2_net_[31] ,
         \_2_net_[30] , \_2_net_[29] , \_2_net_[28] , \_2_net_[27] ,
         \_2_net_[26] , \_2_net_[25] , \_2_net_[24] , \_2_net_[23] ,
         \_2_net_[22] , \_2_net_[21] , \_2_net_[20] , \_2_net_[19] ,
         \_2_net_[18] , \_2_net_[17] , \_2_net_[16] , \_2_net_[15] ,
         \_2_net_[14] , \_2_net_[13] , \_2_net_[12] , \_2_net_[11] ,
         \_2_net_[10] , \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] ,
         \_2_net_[5] , \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , \_4_net_[31] ,
         \_4_net_[30] , \_4_net_[29] , \_4_net_[28] , \_4_net_[27] ,
         \_4_net_[26] , \_4_net_[25] , \_4_net_[24] , \_4_net_[23] ,
         \_4_net_[22] , \_4_net_[21] , \_4_net_[20] , \_4_net_[19] ,
         \_4_net_[18] , \_4_net_[17] , \_4_net_[16] , \_4_net_[15] ,
         \_4_net_[14] , \_4_net_[13] , \_4_net_[12] , \_4_net_[11] ,
         \_4_net_[10] , \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] ,
         \_4_net_[5] , \_4_net_[4] , \_4_net_[3] , \_6_net_[31] ,
         \_6_net_[30] , \_6_net_[29] , \_6_net_[28] , \_6_net_[27] ,
         \_6_net_[26] , \_6_net_[25] , \_6_net_[24] , \_6_net_[23] ,
         \_6_net_[22] , \_6_net_[21] , \_6_net_[20] , \_6_net_[19] ,
         \_6_net_[18] , \_6_net_[17] , \_6_net_[16] , \_6_net_[15] ,
         \_6_net_[14] , \_6_net_[13] , \_6_net_[12] , \_6_net_[11] ,
         \_6_net_[10] , \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] ,
         \_6_net_[5] , \_6_net_[4] , \_8_net_[31] , \_8_net_[30] ,
         \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] ,
         \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] ,
         \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] ,
         \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] ,
         \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] ,
         \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] ,
         \_10_net_[31] , \_10_net_[30] , \_10_net_[29] , \_10_net_[28] ,
         \_10_net_[27] , \_10_net_[26] , \_10_net_[25] , \_10_net_[24] ,
         \_10_net_[23] , \_10_net_[22] , \_10_net_[21] , \_10_net_[20] ,
         \_10_net_[19] , \_10_net_[18] , \_10_net_[17] , \_10_net_[16] ,
         \_10_net_[15] , \_10_net_[14] , \_10_net_[13] , \_10_net_[12] ,
         \_10_net_[11] , \_10_net_[10] , \_10_net_[9] , \_10_net_[8] ,
         \_10_net_[7] , \_10_net_[6] , \_12_net_[31] , \_12_net_[30] ,
         \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] ,
         \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] ,
         \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] ,
         \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] ,
         \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] ,
         \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , \_14_net_[31] ,
         \_14_net_[30] , \_14_net_[29] , \_14_net_[28] , \_14_net_[27] ,
         \_14_net_[26] , \_14_net_[25] , \_14_net_[24] , \_14_net_[23] ,
         \_14_net_[22] , \_14_net_[21] , \_14_net_[20] , \_14_net_[19] ,
         \_14_net_[18] , \_14_net_[17] , \_14_net_[16] , \_14_net_[15] ,
         \_14_net_[14] , \_14_net_[13] , \_14_net_[12] , \_14_net_[11] ,
         \_14_net_[10] , \_14_net_[9] , \_14_net_[8] , \_16_net_[31] ,
         \_16_net_[30] , \_16_net_[29] , \_16_net_[28] , \_16_net_[27] ,
         \_16_net_[26] , \_16_net_[25] , \_16_net_[24] , \_16_net_[23] ,
         \_16_net_[22] , \_16_net_[21] , \_16_net_[20] , \_16_net_[19] ,
         \_16_net_[18] , \_16_net_[17] , \_16_net_[16] , \_16_net_[15] ,
         \_16_net_[14] , \_16_net_[13] , \_16_net_[12] , \_16_net_[11] ,
         \_16_net_[10] , \_16_net_[9] , \_18_net_[31] , \_18_net_[30] ,
         \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] ,
         \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] ,
         \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] ,
         \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] ,
         \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] ,
         \_20_net_[31] , \_20_net_[30] , \_20_net_[29] , \_20_net_[28] ,
         \_20_net_[27] , \_20_net_[26] , \_20_net_[25] , \_20_net_[24] ,
         \_20_net_[23] , \_20_net_[22] , \_20_net_[21] , \_20_net_[20] ,
         \_20_net_[19] , \_20_net_[18] , \_20_net_[17] , \_20_net_[16] ,
         \_20_net_[15] , \_20_net_[14] , \_20_net_[13] , \_20_net_[12] ,
         \_20_net_[11] , \_22_net_[31] , \_22_net_[30] , \_22_net_[29] ,
         \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , \_22_net_[25] ,
         \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , \_22_net_[21] ,
         \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , \_22_net_[17] ,
         \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , \_22_net_[13] ,
         \_22_net_[12] , \_24_net_[31] , \_24_net_[30] , \_24_net_[29] ,
         \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , \_24_net_[25] ,
         \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , \_24_net_[21] ,
         \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , \_24_net_[17] ,
         \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , \_24_net_[13] ,
         \_26_net_[31] , \_26_net_[30] , \_26_net_[29] , \_26_net_[28] ,
         \_26_net_[27] , \_26_net_[26] , \_26_net_[25] , \_26_net_[24] ,
         \_26_net_[23] , \_26_net_[22] , \_26_net_[21] , \_26_net_[20] ,
         \_26_net_[19] , \_26_net_[18] , \_26_net_[17] , \_26_net_[16] ,
         \_26_net_[15] , \_26_net_[14] , \_28_net_[31] , \_28_net_[30] ,
         \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] ,
         \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] ,
         \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] ,
         \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , \_30_net_[31] ,
         \_30_net_[30] , \_30_net_[29] , \_30_net_[28] , \_30_net_[27] ,
         \_30_net_[26] , \_30_net_[25] , \_30_net_[24] , \_30_net_[23] ,
         \_30_net_[22] , \_30_net_[21] , \_30_net_[20] , \_30_net_[19] ,
         \_30_net_[18] , \_30_net_[17] , \_30_net_[16] , \_32_net_[31] ,
         \_32_net_[30] , \_32_net_[29] , \_32_net_[28] , \_32_net_[27] ,
         \_32_net_[26] , \_32_net_[25] , \_32_net_[24] , \_32_net_[23] ,
         \_32_net_[22] , \_32_net_[21] , \_32_net_[20] , \_32_net_[19] ,
         \_32_net_[18] , \_32_net_[17] , \_34_net_[31] , \_34_net_[30] ,
         \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] ,
         \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] ,
         \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] ,
         \_36_net_[31] , \_36_net_[30] , \_36_net_[29] , \_36_net_[28] ,
         \_36_net_[27] , \_36_net_[26] , \_36_net_[25] , \_36_net_[24] ,
         \_36_net_[23] , \_36_net_[22] , \_36_net_[21] , \_36_net_[20] ,
         \_36_net_[19] , \_38_net_[31] , \_38_net_[30] , \_38_net_[29] ,
         \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , \_38_net_[25] ,
         \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , \_38_net_[21] ,
         \_38_net_[20] , \_40_net_[31] , \_40_net_[30] , \_40_net_[29] ,
         \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , \_40_net_[25] ,
         \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , \_40_net_[21] ,
         \_42_net_[31] , \_42_net_[30] , \_42_net_[29] , \_42_net_[28] ,
         \_42_net_[27] , \_42_net_[26] , \_42_net_[25] , \_42_net_[24] ,
         \_42_net_[23] , \_42_net_[22] , \_44_net_[31] , \_44_net_[30] ,
         \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] ,
         \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , \_46_net_[31] ,
         \_46_net_[30] , \_46_net_[29] , \_46_net_[28] , \_46_net_[27] ,
         \_46_net_[26] , \_46_net_[25] , \_46_net_[24] , \_48_net_[31] ,
         \_48_net_[30] , \_48_net_[29] , \_48_net_[28] , \_48_net_[27] ,
         \_48_net_[26] , \_48_net_[25] , \_50_net_[31] , \_50_net_[30] ,
         \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] ,
         \_52_net_[31] , \_52_net_[30] , \_52_net_[29] , \_52_net_[28] ,
         \_52_net_[27] , \_54_net_[31] , \_54_net_[30] , \_54_net_[29] ,
         \_54_net_[28] , \_56_net_[31] , \_56_net_[30] , \_56_net_[29] ,
         \_58_net_[31] , \_58_net_[30] , \_60_net_[31] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  ADD_N32_62 \FAINST[1].ADD_  ( .A({\_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .S({
        \w[2][31] , \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , 
        \w[2][25] , \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , 
        \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , 
        \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , 
        \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , 
        \w[2][1] , SYNOPSYS_UNCONNECTED__0}) );
  ADD_N32_61 \FAINST[2].ADD_  ( .A({\_2_net_[31] , \_2_net_[30] , 
        \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , \_2_net_[26] , 
        \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , \_2_net_[22] , 
        \_2_net_[21] , \_2_net_[20] , \_2_net_[19] , \_2_net_[18] , 
        \_2_net_[17] , \_2_net_[16] , \_2_net_[15] , \_2_net_[14] , 
        \_2_net_[13] , \_2_net_[12] , \_2_net_[11] , \_2_net_[10] , 
        \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , \_2_net_[5] , 
        \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , 1'b0, 1'b0}), .B({\w[2][31] , 
        \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] , 
        \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , \w[2][19] , 
        \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , \w[2][13] , 
        \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , \w[2][7] , 
        \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , \w[2][1] , 1'b0}), .CI(1'b0), .S({\w[3][31] , \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , 
        \w[3][26] , \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , 
        \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , 
        \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , 
        \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , 
        \w[3][2] , \w[3][1] , SYNOPSYS_UNCONNECTED__1}) );
  ADD_N32_60 \FAINST[3].ADD_  ( .A({\_4_net_[31] , \_4_net_[30] , 
        \_4_net_[29] , \_4_net_[28] , \_4_net_[27] , \_4_net_[26] , 
        \_4_net_[25] , \_4_net_[24] , \_4_net_[23] , \_4_net_[22] , 
        \_4_net_[21] , \_4_net_[20] , \_4_net_[19] , \_4_net_[18] , 
        \_4_net_[17] , \_4_net_[16] , \_4_net_[15] , \_4_net_[14] , 
        \_4_net_[13] , \_4_net_[12] , \_4_net_[11] , \_4_net_[10] , 
        \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] , \_4_net_[5] , 
        \_4_net_[4] , \_4_net_[3] , 1'b0, 1'b0, 1'b0}), .B({\w[3][31] , 
        \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] , \w[3][25] , 
        \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , \w[3][20] , \w[3][19] , 
        \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , \w[3][14] , \w[3][13] , 
        \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , 
        \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , 1'b0}), .CI(1'b0), .S({\w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] , 
        \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] , \w[4][21] , 
        \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] , \w[4][16] , \w[4][15] , 
        \w[4][14] , \w[4][13] , \w[4][12] , \w[4][11] , \w[4][10] , \w[4][9] , 
        \w[4][8] , \w[4][7] , \w[4][6] , \w[4][5] , \w[4][4] , \w[4][3] , 
        \w[4][2] , \w[4][1] , SYNOPSYS_UNCONNECTED__2}) );
  ADD_N32_59 \FAINST[4].ADD_  ( .A({\_6_net_[31] , \_6_net_[30] , 
        \_6_net_[29] , \_6_net_[28] , \_6_net_[27] , \_6_net_[26] , 
        \_6_net_[25] , \_6_net_[24] , \_6_net_[23] , \_6_net_[22] , 
        \_6_net_[21] , \_6_net_[20] , \_6_net_[19] , \_6_net_[18] , 
        \_6_net_[17] , \_6_net_[16] , \_6_net_[15] , \_6_net_[14] , 
        \_6_net_[13] , \_6_net_[12] , \_6_net_[11] , \_6_net_[10] , 
        \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] , \_6_net_[5] , 
        \_6_net_[4] , 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[4][31] , \w[4][30] , 
        \w[4][29] , \w[4][28] , \w[4][27] , \w[4][26] , \w[4][25] , \w[4][24] , 
        \w[4][23] , \w[4][22] , \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , 
        \w[4][17] , \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] , 
        \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] , 
        \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , 1'b0}), .CI(
        1'b0), .S({\w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] , \w[5][27] , 
        \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , \w[5][22] , \w[5][21] , 
        \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , \w[5][16] , \w[5][15] , 
        \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , 
        \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , 
        \w[5][2] , \w[5][1] , SYNOPSYS_UNCONNECTED__3}) );
  ADD_N32_58 \FAINST[5].ADD_  ( .A({\_8_net_[31] , \_8_net_[30] , 
        \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] , 
        \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] , 
        \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] , 
        \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] , 
        \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] , 
        \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[5][31] , \w[5][30] , \w[5][29] , 
        \w[5][28] , \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , 
        \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , 
        \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , 
        \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , 
        \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] , 1'b0}), .CI(1'b0), .S({
        \w[6][31] , \w[6][30] , \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , 
        \w[6][25] , \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] , 
        \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] , \w[6][14] , 
        \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] , \w[6][8] , 
        \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] , \w[6][2] , 
        \w[6][1] , SYNOPSYS_UNCONNECTED__4}) );
  ADD_N32_57 \FAINST[6].ADD_  ( .A({\_10_net_[31] , \_10_net_[30] , 
        \_10_net_[29] , \_10_net_[28] , \_10_net_[27] , \_10_net_[26] , 
        \_10_net_[25] , \_10_net_[24] , \_10_net_[23] , \_10_net_[22] , 
        \_10_net_[21] , \_10_net_[20] , \_10_net_[19] , \_10_net_[18] , 
        \_10_net_[17] , \_10_net_[16] , \_10_net_[15] , \_10_net_[14] , 
        \_10_net_[13] , \_10_net_[12] , \_10_net_[11] , \_10_net_[10] , 
        \_10_net_[9] , \_10_net_[8] , \_10_net_[7] , \_10_net_[6] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[6][31] , \w[6][30] , \w[6][29] , 
        \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] , \w[6][24] , \w[6][23] , 
        \w[6][22] , \w[6][21] , \w[6][20] , \w[6][19] , \w[6][18] , \w[6][17] , 
        \w[6][16] , \w[6][15] , \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , 
        \w[6][10] , \w[6][9] , \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , 
        \w[6][4] , \w[6][3] , \w[6][2] , \w[6][1] , 1'b0}), .CI(1'b0), .S({
        \w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] , 
        \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] , \w[7][20] , 
        \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , \w[7][15] , \w[7][14] , 
        \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , \w[7][9] , \w[7][8] , 
        \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , \w[7][3] , \w[7][2] , 
        \w[7][1] , SYNOPSYS_UNCONNECTED__5}) );
  ADD_N32_56 \FAINST[7].ADD_  ( .A({\_12_net_[31] , \_12_net_[30] , 
        \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] , 
        \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] , 
        \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] , 
        \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] , 
        \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] , 
        \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , 
        \w[7][27] , \w[7][26] , \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , 
        \w[7][21] , \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , 
        \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , 
        \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , 
        \w[7][3] , \w[7][2] , \w[7][1] , 1'b0}), .CI(1'b0), .S({\w[8][31] , 
        \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , \w[8][26] , \w[8][25] , 
        \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , \w[8][20] , \w[8][19] , 
        \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , 
        \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , 
        \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , 
        SYNOPSYS_UNCONNECTED__6}) );
  ADD_N32_55 \FAINST[8].ADD_  ( .A({\_14_net_[31] , \_14_net_[30] , 
        \_14_net_[29] , \_14_net_[28] , \_14_net_[27] , \_14_net_[26] , 
        \_14_net_[25] , \_14_net_[24] , \_14_net_[23] , \_14_net_[22] , 
        \_14_net_[21] , \_14_net_[20] , \_14_net_[19] , \_14_net_[18] , 
        \_14_net_[17] , \_14_net_[16] , \_14_net_[15] , \_14_net_[14] , 
        \_14_net_[13] , \_14_net_[12] , \_14_net_[11] , \_14_net_[10] , 
        \_14_net_[9] , \_14_net_[8] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , 
        \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , 
        \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , 
        \w[8][14] , \w[8][13] , \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , 
        \w[8][8] , \w[8][7] , \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , 
        \w[8][2] , \w[8][1] , 1'b0}), .CI(1'b0), .S({\w[9][31] , \w[9][30] , 
        \w[9][29] , \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] , 
        \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] , \w[9][18] , 
        \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] , \w[9][13] , \w[9][12] , 
        \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] , \w[9][7] , \w[9][6] , 
        \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] , \w[9][1] , 
        SYNOPSYS_UNCONNECTED__7}) );
  ADD_N32_54 \FAINST[9].ADD_  ( .A({\_16_net_[31] , \_16_net_[30] , 
        \_16_net_[29] , \_16_net_[28] , \_16_net_[27] , \_16_net_[26] , 
        \_16_net_[25] , \_16_net_[24] , \_16_net_[23] , \_16_net_[22] , 
        \_16_net_[21] , \_16_net_[20] , \_16_net_[19] , \_16_net_[18] , 
        \_16_net_[17] , \_16_net_[16] , \_16_net_[15] , \_16_net_[14] , 
        \_16_net_[13] , \_16_net_[12] , \_16_net_[11] , \_16_net_[10] , 
        \_16_net_[9] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[9][31] , \w[9][30] , \w[9][29] , \w[9][28] , \w[9][27] , 
        \w[9][26] , \w[9][25] , \w[9][24] , \w[9][23] , \w[9][22] , \w[9][21] , 
        \w[9][20] , \w[9][19] , \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , 
        \w[9][14] , \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , 
        \w[9][8] , \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , 
        \w[9][2] , \w[9][1] , 1'b0}), .CI(1'b0), .S({\w[10][31] , \w[10][30] , 
        \w[10][29] , \w[10][28] , \w[10][27] , \w[10][26] , \w[10][25] , 
        \w[10][24] , \w[10][23] , \w[10][22] , \w[10][21] , \w[10][20] , 
        \w[10][19] , \w[10][18] , \w[10][17] , \w[10][16] , \w[10][15] , 
        \w[10][14] , \w[10][13] , \w[10][12] , \w[10][11] , \w[10][10] , 
        \w[10][9] , \w[10][8] , \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , 
        \w[10][3] , \w[10][2] , \w[10][1] , SYNOPSYS_UNCONNECTED__8}) );
  ADD_N32_53 \FAINST[10].ADD_  ( .A({\_18_net_[31] , \_18_net_[30] , 
        \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] , 
        \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] , 
        \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] , 
        \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] , 
        \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] , \w[10][27] , 
        \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] , \w[10][22] , 
        \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] , \w[10][17] , 
        \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] , \w[10][12] , 
        \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] , \w[10][7] , 
        \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] , \w[10][2] , \w[10][1] , 
        1'b0}), .CI(1'b0), .S({\w[11][31] , \w[11][30] , \w[11][29] , 
        \w[11][28] , \w[11][27] , \w[11][26] , \w[11][25] , \w[11][24] , 
        \w[11][23] , \w[11][22] , \w[11][21] , \w[11][20] , \w[11][19] , 
        \w[11][18] , \w[11][17] , \w[11][16] , \w[11][15] , \w[11][14] , 
        \w[11][13] , \w[11][12] , \w[11][11] , \w[11][10] , \w[11][9] , 
        \w[11][8] , \w[11][7] , \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , 
        \w[11][2] , \w[11][1] , SYNOPSYS_UNCONNECTED__9}) );
  ADD_N32_52 \FAINST[11].ADD_  ( .A({\_20_net_[31] , \_20_net_[30] , 
        \_20_net_[29] , \_20_net_[28] , \_20_net_[27] , \_20_net_[26] , 
        \_20_net_[25] , \_20_net_[24] , \_20_net_[23] , \_20_net_[22] , 
        \_20_net_[21] , \_20_net_[20] , \_20_net_[19] , \_20_net_[18] , 
        \_20_net_[17] , \_20_net_[16] , \_20_net_[15] , \_20_net_[14] , 
        \_20_net_[13] , \_20_net_[12] , \_20_net_[11] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[11][31] , 
        \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] , \w[11][26] , 
        \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] , \w[11][21] , 
        \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] , \w[11][16] , 
        \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] , \w[11][11] , 
        \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] , \w[11][6] , 
        \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] , \w[11][1] , 1'b0}), 
        .CI(1'b0), .S({\w[12][31] , \w[12][30] , \w[12][29] , \w[12][28] , 
        \w[12][27] , \w[12][26] , \w[12][25] , \w[12][24] , \w[12][23] , 
        \w[12][22] , \w[12][21] , \w[12][20] , \w[12][19] , \w[12][18] , 
        \w[12][17] , \w[12][16] , \w[12][15] , \w[12][14] , \w[12][13] , 
        \w[12][12] , \w[12][11] , \w[12][10] , \w[12][9] , \w[12][8] , 
        \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , 
        \w[12][1] , SYNOPSYS_UNCONNECTED__10}) );
  ADD_N32_51 \FAINST[12].ADD_  ( .A({\_22_net_[31] , \_22_net_[30] , 
        \_22_net_[29] , \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , 
        \_22_net_[25] , \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , 
        \_22_net_[21] , \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , 
        \_22_net_[17] , \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , 
        \_22_net_[13] , \_22_net_[12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[12][31] , \w[12][30] , 
        \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] , \w[12][25] , 
        \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] , \w[12][20] , 
        \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] , \w[12][15] , 
        \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] , \w[12][10] , 
        \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , 
        \w[12][3] , \w[12][2] , \w[12][1] , 1'b0}), .CI(1'b0), .S({\w[13][31] , 
        \w[13][30] , \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , 
        \w[13][25] , \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , 
        \w[13][20] , \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , 
        \w[13][15] , \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , 
        \w[13][10] , \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , 
        \w[13][5] , \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , 
        SYNOPSYS_UNCONNECTED__11}) );
  ADD_N32_50 \FAINST[13].ADD_  ( .A({\_24_net_[31] , \_24_net_[30] , 
        \_24_net_[29] , \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , 
        \_24_net_[25] , \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , 
        \_24_net_[21] , \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , 
        \_24_net_[17] , \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , 
        \_24_net_[13] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[13][31] , \w[13][30] , \w[13][29] , 
        \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] , \w[13][24] , 
        \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] , \w[13][19] , 
        \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] , \w[13][14] , 
        \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] , \w[13][9] , 
        \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] , \w[13][4] , \w[13][3] , 
        \w[13][2] , \w[13][1] , 1'b0}), .CI(1'b0), .S({\w[14][31] , 
        \w[14][30] , \w[14][29] , \w[14][28] , \w[14][27] , \w[14][26] , 
        \w[14][25] , \w[14][24] , \w[14][23] , \w[14][22] , \w[14][21] , 
        \w[14][20] , \w[14][19] , \w[14][18] , \w[14][17] , \w[14][16] , 
        \w[14][15] , \w[14][14] , \w[14][13] , \w[14][12] , \w[14][11] , 
        \w[14][10] , \w[14][9] , \w[14][8] , \w[14][7] , \w[14][6] , 
        \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , \w[14][1] , 
        SYNOPSYS_UNCONNECTED__12}) );
  ADD_N32_49 \FAINST[14].ADD_  ( .A({\_26_net_[31] , \_26_net_[30] , 
        \_26_net_[29] , \_26_net_[28] , \_26_net_[27] , \_26_net_[26] , 
        \_26_net_[25] , \_26_net_[24] , \_26_net_[23] , \_26_net_[22] , 
        \_26_net_[21] , \_26_net_[20] , \_26_net_[19] , \_26_net_[18] , 
        \_26_net_[17] , \_26_net_[16] , \_26_net_[15] , \_26_net_[14] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[14][31] , \w[14][30] , \w[14][29] , \w[14][28] , 
        \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] , \w[14][23] , 
        \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] , \w[14][18] , 
        \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] , \w[14][13] , 
        \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] , \w[14][8] , 
        \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , 
        \w[14][1] , 1'b0}), .CI(1'b0), .S({\w[15][31] , \w[15][30] , 
        \w[15][29] , \w[15][28] , \w[15][27] , \w[15][26] , \w[15][25] , 
        \w[15][24] , \w[15][23] , \w[15][22] , \w[15][21] , \w[15][20] , 
        \w[15][19] , \w[15][18] , \w[15][17] , \w[15][16] , \w[15][15] , 
        \w[15][14] , \w[15][13] , \w[15][12] , \w[15][11] , \w[15][10] , 
        \w[15][9] , \w[15][8] , \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , 
        \w[15][3] , \w[15][2] , \w[15][1] , SYNOPSYS_UNCONNECTED__13}) );
  ADD_N32_48 \FAINST[15].ADD_  ( .A({\_28_net_[31] , \_28_net_[30] , 
        \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] , 
        \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] , 
        \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] , 
        \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] , \w[15][27] , 
        \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] , \w[15][22] , 
        \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] , \w[15][17] , 
        \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] , \w[15][12] , 
        \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] , \w[15][7] , 
        \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] , \w[15][2] , \w[15][1] , 
        1'b0}), .CI(1'b0), .S({\w[16][31] , \w[16][30] , \w[16][29] , 
        \w[16][28] , \w[16][27] , \w[16][26] , \w[16][25] , \w[16][24] , 
        \w[16][23] , \w[16][22] , \w[16][21] , \w[16][20] , \w[16][19] , 
        \w[16][18] , \w[16][17] , \w[16][16] , \w[16][15] , \w[16][14] , 
        \w[16][13] , \w[16][12] , \w[16][11] , \w[16][10] , \w[16][9] , 
        \w[16][8] , \w[16][7] , \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , 
        \w[16][2] , \w[16][1] , SYNOPSYS_UNCONNECTED__14}) );
  ADD_N32_47 \FAINST[16].ADD_  ( .A({\_30_net_[31] , \_30_net_[30] , 
        \_30_net_[29] , \_30_net_[28] , \_30_net_[27] , \_30_net_[26] , 
        \_30_net_[25] , \_30_net_[24] , \_30_net_[23] , \_30_net_[22] , 
        \_30_net_[21] , \_30_net_[20] , \_30_net_[19] , \_30_net_[18] , 
        \_30_net_[17] , \_30_net_[16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] , 
        \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] , 
        \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] , 
        \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] , 
        \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] , 
        \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] , \w[16][1] , 
        1'b0}), .CI(1'b0), .S({\w[17][31] , \w[17][30] , \w[17][29] , 
        \w[17][28] , \w[17][27] , \w[17][26] , \w[17][25] , \w[17][24] , 
        \w[17][23] , \w[17][22] , \w[17][21] , \w[17][20] , \w[17][19] , 
        \w[17][18] , \w[17][17] , \w[17][16] , \w[17][15] , \w[17][14] , 
        \w[17][13] , \w[17][12] , \w[17][11] , \w[17][10] , \w[17][9] , 
        \w[17][8] , \w[17][7] , \w[17][6] , \w[17][5] , \w[17][4] , \w[17][3] , 
        \w[17][2] , \w[17][1] , SYNOPSYS_UNCONNECTED__15}) );
  ADD_N32_46 \FAINST[17].ADD_  ( .A({\_32_net_[31] , \_32_net_[30] , 
        \_32_net_[29] , \_32_net_[28] , \_32_net_[27] , \_32_net_[26] , 
        \_32_net_[25] , \_32_net_[24] , \_32_net_[23] , \_32_net_[22] , 
        \_32_net_[21] , \_32_net_[20] , \_32_net_[19] , \_32_net_[18] , 
        \_32_net_[17] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[17][31] , 
        \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] , 
        \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] , 
        \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] , 
        \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] , 
        \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] , 
        \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] , 1'b0}), 
        .CI(1'b0), .S({\w[18][31] , \w[18][30] , \w[18][29] , \w[18][28] , 
        \w[18][27] , \w[18][26] , \w[18][25] , \w[18][24] , \w[18][23] , 
        \w[18][22] , \w[18][21] , \w[18][20] , \w[18][19] , \w[18][18] , 
        \w[18][17] , \w[18][16] , \w[18][15] , \w[18][14] , \w[18][13] , 
        \w[18][12] , \w[18][11] , \w[18][10] , \w[18][9] , \w[18][8] , 
        \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , \w[18][3] , \w[18][2] , 
        \w[18][1] , SYNOPSYS_UNCONNECTED__16}) );
  ADD_N32_45 \FAINST[18].ADD_  ( .A({\_34_net_[31] , \_34_net_[30] , 
        \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] , 
        \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] , 
        \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[18][31] , \w[18][30] , 
        \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] , 
        \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] , 
        \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] , 
        \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] , 
        \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , 
        \w[18][3] , \w[18][2] , \w[18][1] , 1'b0}), .CI(1'b0), .S({\w[19][31] , 
        \w[19][30] , \w[19][29] , \w[19][28] , \w[19][27] , \w[19][26] , 
        \w[19][25] , \w[19][24] , \w[19][23] , \w[19][22] , \w[19][21] , 
        \w[19][20] , \w[19][19] , \w[19][18] , \w[19][17] , \w[19][16] , 
        \w[19][15] , \w[19][14] , \w[19][13] , \w[19][12] , \w[19][11] , 
        \w[19][10] , \w[19][9] , \w[19][8] , \w[19][7] , \w[19][6] , 
        \w[19][5] , \w[19][4] , \w[19][3] , \w[19][2] , \w[19][1] , 
        SYNOPSYS_UNCONNECTED__17}) );
  ADD_N32_44 \FAINST[19].ADD_  ( .A({\_36_net_[31] , \_36_net_[30] , 
        \_36_net_[29] , \_36_net_[28] , \_36_net_[27] , \_36_net_[26] , 
        \_36_net_[25] , \_36_net_[24] , \_36_net_[23] , \_36_net_[22] , 
        \_36_net_[21] , \_36_net_[20] , \_36_net_[19] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[19][31] , \w[19][30] , \w[19][29] , 
        \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] , 
        \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] , 
        \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] , 
        \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] , 
        \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] , \w[19][3] , 
        \w[19][2] , \w[19][1] , 1'b0}), .CI(1'b0), .S({\w[20][31] , 
        \w[20][30] , \w[20][29] , \w[20][28] , \w[20][27] , \w[20][26] , 
        \w[20][25] , \w[20][24] , \w[20][23] , \w[20][22] , \w[20][21] , 
        \w[20][20] , \w[20][19] , \w[20][18] , \w[20][17] , \w[20][16] , 
        \w[20][15] , \w[20][14] , \w[20][13] , \w[20][12] , \w[20][11] , 
        \w[20][10] , \w[20][9] , \w[20][8] , \w[20][7] , \w[20][6] , 
        \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , \w[20][1] , 
        SYNOPSYS_UNCONNECTED__18}) );
  ADD_N32_43 \FAINST[20].ADD_  ( .A({\_38_net_[31] , \_38_net_[30] , 
        \_38_net_[29] , \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , 
        \_38_net_[25] , \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , 
        \_38_net_[21] , \_38_net_[20] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({\w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] , 
        \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] , 
        \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] , 
        \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] , 
        \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] , 
        \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , 
        \w[20][1] , 1'b0}), .CI(1'b0), .S({\w[21][31] , \w[21][30] , 
        \w[21][29] , \w[21][28] , \w[21][27] , \w[21][26] , \w[21][25] , 
        \w[21][24] , \w[21][23] , \w[21][22] , \w[21][21] , \w[21][20] , 
        \w[21][19] , \w[21][18] , \w[21][17] , \w[21][16] , \w[21][15] , 
        \w[21][14] , \w[21][13] , \w[21][12] , \w[21][11] , \w[21][10] , 
        \w[21][9] , \w[21][8] , \w[21][7] , \w[21][6] , \w[21][5] , \w[21][4] , 
        \w[21][3] , \w[21][2] , \w[21][1] , SYNOPSYS_UNCONNECTED__19}) );
  ADD_N32_42 \FAINST[21].ADD_  ( .A({\_40_net_[31] , \_40_net_[30] , 
        \_40_net_[29] , \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , 
        \_40_net_[25] , \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , 
        \_40_net_[21] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] , 
        \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] , 
        \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] , 
        \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] , 
        \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] , 
        \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] , \w[21][1] , 
        1'b0}), .CI(1'b0), .S({\w[22][31] , \w[22][30] , \w[22][29] , 
        \w[22][28] , \w[22][27] , \w[22][26] , \w[22][25] , \w[22][24] , 
        \w[22][23] , \w[22][22] , \w[22][21] , \w[22][20] , \w[22][19] , 
        \w[22][18] , \w[22][17] , \w[22][16] , \w[22][15] , \w[22][14] , 
        \w[22][13] , \w[22][12] , \w[22][11] , \w[22][10] , \w[22][9] , 
        \w[22][8] , \w[22][7] , \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , 
        \w[22][2] , \w[22][1] , SYNOPSYS_UNCONNECTED__20}) );
  ADD_N32_41 \FAINST[22].ADD_  ( .A({\_42_net_[31] , \_42_net_[30] , 
        \_42_net_[29] , \_42_net_[28] , \_42_net_[27] , \_42_net_[26] , 
        \_42_net_[25] , \_42_net_[24] , \_42_net_[23] , \_42_net_[22] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[22][31] , \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , 
        \w[22][26] , \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , 
        \w[22][21] , \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , 
        \w[22][16] , \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , 
        \w[22][11] , \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , 
        \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] , 
        1'b0}), .CI(1'b0), .S({\w[23][31] , \w[23][30] , \w[23][29] , 
        \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] , \w[23][24] , 
        \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] , \w[23][19] , 
        \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] , \w[23][14] , 
        \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] , \w[23][9] , 
        \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] , \w[23][4] , \w[23][3] , 
        \w[23][2] , \w[23][1] , SYNOPSYS_UNCONNECTED__21}) );
  ADD_N32_40 \FAINST[23].ADD_  ( .A({\_44_net_[31] , \_44_net_[30] , 
        \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] , 
        \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[23][31] , 
        \w[23][30] , \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , 
        \w[23][25] , \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , 
        \w[23][20] , \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , 
        \w[23][15] , \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , 
        \w[23][10] , \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , 
        \w[23][5] , \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , 1'b0}), 
        .CI(1'b0), .S({\w[24][31] , \w[24][30] , \w[24][29] , \w[24][28] , 
        \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] , \w[24][23] , 
        \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] , \w[24][18] , 
        \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] , \w[24][13] , 
        \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] , \w[24][8] , 
        \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , \w[24][3] , \w[24][2] , 
        \w[24][1] , SYNOPSYS_UNCONNECTED__22}) );
  ADD_N32_39 \FAINST[24].ADD_  ( .A({\_46_net_[31] , \_46_net_[30] , 
        \_46_net_[29] , \_46_net_[28] , \_46_net_[27] , \_46_net_[26] , 
        \_46_net_[25] , \_46_net_[24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[24][31] , \w[24][30] , 
        \w[24][29] , \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , 
        \w[24][24] , \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , 
        \w[24][19] , \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , 
        \w[24][14] , \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , 
        \w[24][9] , \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , 
        \w[24][3] , \w[24][2] , \w[24][1] , 1'b0}), .CI(1'b0), .S({\w[25][31] , 
        \w[25][30] , \w[25][29] , \w[25][28] , \w[25][27] , \w[25][26] , 
        \w[25][25] , \w[25][24] , \w[25][23] , \w[25][22] , \w[25][21] , 
        \w[25][20] , \w[25][19] , \w[25][18] , \w[25][17] , \w[25][16] , 
        \w[25][15] , \w[25][14] , \w[25][13] , \w[25][12] , \w[25][11] , 
        \w[25][10] , \w[25][9] , \w[25][8] , \w[25][7] , \w[25][6] , 
        \w[25][5] , \w[25][4] , \w[25][3] , \w[25][2] , \w[25][1] , 
        SYNOPSYS_UNCONNECTED__23}) );
  ADD_N32_38 \FAINST[25].ADD_  ( .A({\_48_net_[31] , \_48_net_[30] , 
        \_48_net_[29] , \_48_net_[28] , \_48_net_[27] , \_48_net_[26] , 
        \_48_net_[25] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[25][31] , \w[25][30] , \w[25][29] , 
        \w[25][28] , \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , 
        \w[25][23] , \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , 
        \w[25][18] , \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , 
        \w[25][13] , \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , 
        \w[25][8] , \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] , 
        \w[25][2] , \w[25][1] , 1'b0}), .CI(1'b0), .S({\w[26][31] , 
        \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] , \w[26][26] , 
        \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] , \w[26][21] , 
        \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] , \w[26][16] , 
        \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] , \w[26][11] , 
        \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] , \w[26][6] , 
        \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , \w[26][1] , 
        SYNOPSYS_UNCONNECTED__24}) );
  ADD_N32_37 \FAINST[26].ADD_  ( .A({\_50_net_[31] , \_50_net_[30] , 
        \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , 
        \w[26][27] , \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , 
        \w[26][22] , \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , 
        \w[26][17] , \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , 
        \w[26][12] , \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , 
        \w[26][7] , \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , 
        \w[26][1] , 1'b0}), .CI(1'b0), .S({\w[27][31] , \w[27][30] , 
        \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] , \w[27][25] , 
        \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] , \w[27][20] , 
        \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] , \w[27][15] , 
        \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] , \w[27][10] , 
        \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] , \w[27][5] , \w[27][4] , 
        \w[27][3] , \w[27][2] , \w[27][1] , SYNOPSYS_UNCONNECTED__25}) );
  ADD_N32_36 \FAINST[27].ADD_  ( .A({\_52_net_[31] , \_52_net_[30] , 
        \_52_net_[29] , \_52_net_[28] , \_52_net_[27] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[27][31] , \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , 
        \w[27][26] , \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , 
        \w[27][21] , \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , 
        \w[27][16] , \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , 
        \w[27][11] , \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , 
        \w[27][6] , \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] , 
        1'b0}), .CI(1'b0), .S({\w[28][31] , \w[28][30] , \w[28][29] , 
        \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] , \w[28][24] , 
        \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] , \w[28][19] , 
        \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] , \w[28][14] , 
        \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] , \w[28][9] , 
        \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , 
        \w[28][2] , \w[28][1] , SYNOPSYS_UNCONNECTED__26}) );
  ADD_N32_35 \FAINST[28].ADD_  ( .A({\_54_net_[31] , \_54_net_[30] , 
        \_54_net_[29] , \_54_net_[28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[28][31] , \w[28][30] , \w[28][29] , \w[28][28] , \w[28][27] , 
        \w[28][26] , \w[28][25] , \w[28][24] , \w[28][23] , \w[28][22] , 
        \w[28][21] , \w[28][20] , \w[28][19] , \w[28][18] , \w[28][17] , 
        \w[28][16] , \w[28][15] , \w[28][14] , \w[28][13] , \w[28][12] , 
        \w[28][11] , \w[28][10] , \w[28][9] , \w[28][8] , \w[28][7] , 
        \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , 
        1'b0}), .CI(1'b0), .S({\w[29][31] , \w[29][30] , \w[29][29] , 
        \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] , 
        \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] , 
        \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] , 
        \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] , 
        \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] , \w[29][3] , 
        \w[29][2] , \w[29][1] , SYNOPSYS_UNCONNECTED__27}) );
  ADD_N32_34 \FAINST[29].ADD_  ( .A({\_56_net_[31] , \_56_net_[30] , 
        \_56_net_[29] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[29][31] , 
        \w[29][30] , \w[29][29] , \w[29][28] , \w[29][27] , \w[29][26] , 
        \w[29][25] , \w[29][24] , \w[29][23] , \w[29][22] , \w[29][21] , 
        \w[29][20] , \w[29][19] , \w[29][18] , \w[29][17] , \w[29][16] , 
        \w[29][15] , \w[29][14] , \w[29][13] , \w[29][12] , \w[29][11] , 
        \w[29][10] , \w[29][9] , \w[29][8] , \w[29][7] , \w[29][6] , 
        \w[29][5] , \w[29][4] , \w[29][3] , \w[29][2] , \w[29][1] , 1'b0}), 
        .CI(1'b0), .S({\w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] , 
        \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] , 
        \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] , 
        \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] , 
        \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] , 
        \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] , \w[30][2] , 
        \w[30][1] , SYNOPSYS_UNCONNECTED__28}) );
  ADD_N32_33 \FAINST[30].ADD_  ( .A({\_58_net_[31] , \_58_net_[30] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[30][31] , \w[30][30] , 
        \w[30][29] , \w[30][28] , \w[30][27] , \w[30][26] , \w[30][25] , 
        \w[30][24] , \w[30][23] , \w[30][22] , \w[30][21] , \w[30][20] , 
        \w[30][19] , \w[30][18] , \w[30][17] , \w[30][16] , \w[30][15] , 
        \w[30][14] , \w[30][13] , \w[30][12] , \w[30][11] , \w[30][10] , 
        \w[30][9] , \w[30][8] , \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , 
        \w[30][3] , \w[30][2] , \w[30][1] , 1'b0}), .CI(1'b0), .S({\w[31][31] , 
        \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] , \w[31][26] , 
        \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] , \w[31][21] , 
        \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] , \w[31][16] , 
        \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] , \w[31][11] , 
        \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] , \w[31][6] , 
        \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] , \w[31][1] , 
        SYNOPSYS_UNCONNECTED__29}) );
  ADD_N32_32 \FAINST[31].ADD_  ( .A({\_60_net_[31] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[31][31] , \w[31][30] , \w[31][29] , 
        \w[31][28] , \w[31][27] , \w[31][26] , \w[31][25] , \w[31][24] , 
        \w[31][23] , \w[31][22] , \w[31][21] , \w[31][20] , \w[31][19] , 
        \w[31][18] , \w[31][17] , \w[31][16] , \w[31][15] , \w[31][14] , 
        \w[31][13] , \w[31][12] , \w[31][11] , \w[31][10] , \w[31][9] , 
        \w[31][8] , \w[31][7] , \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , 
        \w[31][2] , \w[31][1] , 1'b0}), .CI(1'b0), .S({O[31:1], 
        SYNOPSYS_UNCONNECTED__30}) );
  AND U2 ( .A(A[5]), .B(B[4]), .Z(\_8_net_[9] ) );
  AND U3 ( .A(A[5]), .B(B[3]), .Z(\_8_net_[8] ) );
  AND U4 ( .A(A[5]), .B(B[2]), .Z(\_8_net_[7] ) );
  AND U5 ( .A(A[5]), .B(B[1]), .Z(\_8_net_[6] ) );
  AND U6 ( .A(A[5]), .B(B[0]), .Z(\_8_net_[5] ) );
  AND U7 ( .A(A[5]), .B(B[26]), .Z(\_8_net_[31] ) );
  AND U8 ( .A(A[5]), .B(B[25]), .Z(\_8_net_[30] ) );
  AND U9 ( .A(A[5]), .B(B[24]), .Z(\_8_net_[29] ) );
  AND U10 ( .A(A[5]), .B(B[23]), .Z(\_8_net_[28] ) );
  AND U11 ( .A(A[5]), .B(B[22]), .Z(\_8_net_[27] ) );
  AND U12 ( .A(A[5]), .B(B[21]), .Z(\_8_net_[26] ) );
  AND U13 ( .A(A[5]), .B(B[20]), .Z(\_8_net_[25] ) );
  AND U14 ( .A(A[5]), .B(B[19]), .Z(\_8_net_[24] ) );
  AND U15 ( .A(A[5]), .B(B[18]), .Z(\_8_net_[23] ) );
  AND U16 ( .A(A[5]), .B(B[17]), .Z(\_8_net_[22] ) );
  AND U17 ( .A(A[5]), .B(B[16]), .Z(\_8_net_[21] ) );
  AND U18 ( .A(A[5]), .B(B[15]), .Z(\_8_net_[20] ) );
  AND U19 ( .A(A[5]), .B(B[14]), .Z(\_8_net_[19] ) );
  AND U20 ( .A(A[5]), .B(B[13]), .Z(\_8_net_[18] ) );
  AND U21 ( .A(A[5]), .B(B[12]), .Z(\_8_net_[17] ) );
  AND U22 ( .A(A[5]), .B(B[11]), .Z(\_8_net_[16] ) );
  AND U23 ( .A(A[5]), .B(B[10]), .Z(\_8_net_[15] ) );
  AND U24 ( .A(A[5]), .B(B[9]), .Z(\_8_net_[14] ) );
  AND U25 ( .A(A[5]), .B(B[8]), .Z(\_8_net_[13] ) );
  AND U26 ( .A(A[5]), .B(B[7]), .Z(\_8_net_[12] ) );
  AND U27 ( .A(A[5]), .B(B[6]), .Z(\_8_net_[11] ) );
  AND U28 ( .A(A[5]), .B(B[5]), .Z(\_8_net_[10] ) );
  AND U29 ( .A(B[5]), .B(A[4]), .Z(\_6_net_[9] ) );
  AND U30 ( .A(B[4]), .B(A[4]), .Z(\_6_net_[8] ) );
  AND U31 ( .A(B[3]), .B(A[4]), .Z(\_6_net_[7] ) );
  AND U32 ( .A(B[2]), .B(A[4]), .Z(\_6_net_[6] ) );
  AND U33 ( .A(B[1]), .B(A[4]), .Z(\_6_net_[5] ) );
  AND U34 ( .A(B[0]), .B(A[4]), .Z(\_6_net_[4] ) );
  AND U35 ( .A(A[4]), .B(B[27]), .Z(\_6_net_[31] ) );
  AND U36 ( .A(B[26]), .B(A[4]), .Z(\_6_net_[30] ) );
  AND U37 ( .A(B[25]), .B(A[4]), .Z(\_6_net_[29] ) );
  AND U38 ( .A(B[24]), .B(A[4]), .Z(\_6_net_[28] ) );
  AND U39 ( .A(B[23]), .B(A[4]), .Z(\_6_net_[27] ) );
  AND U40 ( .A(B[22]), .B(A[4]), .Z(\_6_net_[26] ) );
  AND U41 ( .A(B[21]), .B(A[4]), .Z(\_6_net_[25] ) );
  AND U42 ( .A(B[20]), .B(A[4]), .Z(\_6_net_[24] ) );
  AND U43 ( .A(B[19]), .B(A[4]), .Z(\_6_net_[23] ) );
  AND U44 ( .A(B[18]), .B(A[4]), .Z(\_6_net_[22] ) );
  AND U45 ( .A(B[17]), .B(A[4]), .Z(\_6_net_[21] ) );
  AND U46 ( .A(B[16]), .B(A[4]), .Z(\_6_net_[20] ) );
  AND U47 ( .A(B[15]), .B(A[4]), .Z(\_6_net_[19] ) );
  AND U48 ( .A(B[14]), .B(A[4]), .Z(\_6_net_[18] ) );
  AND U49 ( .A(B[13]), .B(A[4]), .Z(\_6_net_[17] ) );
  AND U50 ( .A(B[12]), .B(A[4]), .Z(\_6_net_[16] ) );
  AND U51 ( .A(B[11]), .B(A[4]), .Z(\_6_net_[15] ) );
  AND U52 ( .A(B[10]), .B(A[4]), .Z(\_6_net_[14] ) );
  AND U53 ( .A(B[9]), .B(A[4]), .Z(\_6_net_[13] ) );
  AND U54 ( .A(B[8]), .B(A[4]), .Z(\_6_net_[12] ) );
  AND U55 ( .A(B[7]), .B(A[4]), .Z(\_6_net_[11] ) );
  AND U56 ( .A(B[6]), .B(A[4]), .Z(\_6_net_[10] ) );
  AND U57 ( .A(A[31]), .B(B[0]), .Z(\_60_net_[31] ) );
  AND U58 ( .A(B[1]), .B(A[30]), .Z(\_58_net_[31] ) );
  AND U59 ( .A(A[30]), .B(B[0]), .Z(\_58_net_[30] ) );
  AND U60 ( .A(B[2]), .B(A[29]), .Z(\_56_net_[31] ) );
  AND U61 ( .A(B[1]), .B(A[29]), .Z(\_56_net_[30] ) );
  AND U62 ( .A(A[29]), .B(B[0]), .Z(\_56_net_[29] ) );
  AND U63 ( .A(B[3]), .B(A[28]), .Z(\_54_net_[31] ) );
  AND U64 ( .A(B[2]), .B(A[28]), .Z(\_54_net_[30] ) );
  AND U65 ( .A(B[1]), .B(A[28]), .Z(\_54_net_[29] ) );
  AND U66 ( .A(A[28]), .B(B[0]), .Z(\_54_net_[28] ) );
  AND U67 ( .A(B[4]), .B(A[27]), .Z(\_52_net_[31] ) );
  AND U68 ( .A(B[3]), .B(A[27]), .Z(\_52_net_[30] ) );
  AND U69 ( .A(B[2]), .B(A[27]), .Z(\_52_net_[29] ) );
  AND U70 ( .A(B[1]), .B(A[27]), .Z(\_52_net_[28] ) );
  AND U71 ( .A(A[27]), .B(B[0]), .Z(\_52_net_[27] ) );
  AND U72 ( .A(B[5]), .B(A[26]), .Z(\_50_net_[31] ) );
  AND U73 ( .A(B[4]), .B(A[26]), .Z(\_50_net_[30] ) );
  AND U74 ( .A(B[3]), .B(A[26]), .Z(\_50_net_[29] ) );
  AND U75 ( .A(B[2]), .B(A[26]), .Z(\_50_net_[28] ) );
  AND U76 ( .A(B[1]), .B(A[26]), .Z(\_50_net_[27] ) );
  AND U77 ( .A(A[26]), .B(B[0]), .Z(\_50_net_[26] ) );
  AND U78 ( .A(B[6]), .B(A[3]), .Z(\_4_net_[9] ) );
  AND U79 ( .A(B[5]), .B(A[3]), .Z(\_4_net_[8] ) );
  AND U80 ( .A(B[4]), .B(A[3]), .Z(\_4_net_[7] ) );
  AND U81 ( .A(B[3]), .B(A[3]), .Z(\_4_net_[6] ) );
  AND U82 ( .A(B[2]), .B(A[3]), .Z(\_4_net_[5] ) );
  AND U83 ( .A(B[1]), .B(A[3]), .Z(\_4_net_[4] ) );
  AND U84 ( .A(B[0]), .B(A[3]), .Z(\_4_net_[3] ) );
  AND U85 ( .A(A[3]), .B(B[28]), .Z(\_4_net_[31] ) );
  AND U86 ( .A(B[27]), .B(A[3]), .Z(\_4_net_[30] ) );
  AND U87 ( .A(B[26]), .B(A[3]), .Z(\_4_net_[29] ) );
  AND U88 ( .A(B[25]), .B(A[3]), .Z(\_4_net_[28] ) );
  AND U89 ( .A(B[24]), .B(A[3]), .Z(\_4_net_[27] ) );
  AND U90 ( .A(B[23]), .B(A[3]), .Z(\_4_net_[26] ) );
  AND U91 ( .A(B[22]), .B(A[3]), .Z(\_4_net_[25] ) );
  AND U92 ( .A(B[21]), .B(A[3]), .Z(\_4_net_[24] ) );
  AND U93 ( .A(B[20]), .B(A[3]), .Z(\_4_net_[23] ) );
  AND U94 ( .A(B[19]), .B(A[3]), .Z(\_4_net_[22] ) );
  AND U95 ( .A(B[18]), .B(A[3]), .Z(\_4_net_[21] ) );
  AND U96 ( .A(B[17]), .B(A[3]), .Z(\_4_net_[20] ) );
  AND U97 ( .A(B[16]), .B(A[3]), .Z(\_4_net_[19] ) );
  AND U98 ( .A(B[15]), .B(A[3]), .Z(\_4_net_[18] ) );
  AND U99 ( .A(B[14]), .B(A[3]), .Z(\_4_net_[17] ) );
  AND U100 ( .A(B[13]), .B(A[3]), .Z(\_4_net_[16] ) );
  AND U101 ( .A(B[12]), .B(A[3]), .Z(\_4_net_[15] ) );
  AND U102 ( .A(B[11]), .B(A[3]), .Z(\_4_net_[14] ) );
  AND U103 ( .A(B[10]), .B(A[3]), .Z(\_4_net_[13] ) );
  AND U104 ( .A(B[9]), .B(A[3]), .Z(\_4_net_[12] ) );
  AND U105 ( .A(B[8]), .B(A[3]), .Z(\_4_net_[11] ) );
  AND U106 ( .A(B[7]), .B(A[3]), .Z(\_4_net_[10] ) );
  AND U107 ( .A(B[6]), .B(A[25]), .Z(\_48_net_[31] ) );
  AND U108 ( .A(B[5]), .B(A[25]), .Z(\_48_net_[30] ) );
  AND U109 ( .A(B[4]), .B(A[25]), .Z(\_48_net_[29] ) );
  AND U110 ( .A(B[3]), .B(A[25]), .Z(\_48_net_[28] ) );
  AND U111 ( .A(B[2]), .B(A[25]), .Z(\_48_net_[27] ) );
  AND U112 ( .A(B[1]), .B(A[25]), .Z(\_48_net_[26] ) );
  AND U113 ( .A(A[25]), .B(B[0]), .Z(\_48_net_[25] ) );
  AND U114 ( .A(B[7]), .B(A[24]), .Z(\_46_net_[31] ) );
  AND U115 ( .A(B[6]), .B(A[24]), .Z(\_46_net_[30] ) );
  AND U116 ( .A(B[5]), .B(A[24]), .Z(\_46_net_[29] ) );
  AND U117 ( .A(B[4]), .B(A[24]), .Z(\_46_net_[28] ) );
  AND U118 ( .A(B[3]), .B(A[24]), .Z(\_46_net_[27] ) );
  AND U119 ( .A(B[2]), .B(A[24]), .Z(\_46_net_[26] ) );
  AND U120 ( .A(B[1]), .B(A[24]), .Z(\_46_net_[25] ) );
  AND U121 ( .A(A[24]), .B(B[0]), .Z(\_46_net_[24] ) );
  AND U122 ( .A(B[8]), .B(A[23]), .Z(\_44_net_[31] ) );
  AND U123 ( .A(B[7]), .B(A[23]), .Z(\_44_net_[30] ) );
  AND U124 ( .A(B[6]), .B(A[23]), .Z(\_44_net_[29] ) );
  AND U125 ( .A(B[5]), .B(A[23]), .Z(\_44_net_[28] ) );
  AND U126 ( .A(B[4]), .B(A[23]), .Z(\_44_net_[27] ) );
  AND U127 ( .A(B[3]), .B(A[23]), .Z(\_44_net_[26] ) );
  AND U128 ( .A(B[2]), .B(A[23]), .Z(\_44_net_[25] ) );
  AND U129 ( .A(B[1]), .B(A[23]), .Z(\_44_net_[24] ) );
  AND U130 ( .A(A[23]), .B(B[0]), .Z(\_44_net_[23] ) );
  AND U131 ( .A(B[9]), .B(A[22]), .Z(\_42_net_[31] ) );
  AND U132 ( .A(B[8]), .B(A[22]), .Z(\_42_net_[30] ) );
  AND U133 ( .A(B[7]), .B(A[22]), .Z(\_42_net_[29] ) );
  AND U134 ( .A(B[6]), .B(A[22]), .Z(\_42_net_[28] ) );
  AND U135 ( .A(B[5]), .B(A[22]), .Z(\_42_net_[27] ) );
  AND U136 ( .A(B[4]), .B(A[22]), .Z(\_42_net_[26] ) );
  AND U137 ( .A(B[3]), .B(A[22]), .Z(\_42_net_[25] ) );
  AND U138 ( .A(B[2]), .B(A[22]), .Z(\_42_net_[24] ) );
  AND U139 ( .A(B[1]), .B(A[22]), .Z(\_42_net_[23] ) );
  AND U140 ( .A(A[22]), .B(B[0]), .Z(\_42_net_[22] ) );
  AND U141 ( .A(B[10]), .B(A[21]), .Z(\_40_net_[31] ) );
  AND U142 ( .A(B[9]), .B(A[21]), .Z(\_40_net_[30] ) );
  AND U143 ( .A(B[8]), .B(A[21]), .Z(\_40_net_[29] ) );
  AND U144 ( .A(B[7]), .B(A[21]), .Z(\_40_net_[28] ) );
  AND U145 ( .A(B[6]), .B(A[21]), .Z(\_40_net_[27] ) );
  AND U146 ( .A(B[5]), .B(A[21]), .Z(\_40_net_[26] ) );
  AND U147 ( .A(B[4]), .B(A[21]), .Z(\_40_net_[25] ) );
  AND U148 ( .A(B[3]), .B(A[21]), .Z(\_40_net_[24] ) );
  AND U149 ( .A(B[2]), .B(A[21]), .Z(\_40_net_[23] ) );
  AND U150 ( .A(B[1]), .B(A[21]), .Z(\_40_net_[22] ) );
  AND U151 ( .A(A[21]), .B(B[0]), .Z(\_40_net_[21] ) );
  AND U152 ( .A(B[11]), .B(A[20]), .Z(\_38_net_[31] ) );
  AND U153 ( .A(B[10]), .B(A[20]), .Z(\_38_net_[30] ) );
  AND U154 ( .A(B[9]), .B(A[20]), .Z(\_38_net_[29] ) );
  AND U155 ( .A(B[8]), .B(A[20]), .Z(\_38_net_[28] ) );
  AND U156 ( .A(B[7]), .B(A[20]), .Z(\_38_net_[27] ) );
  AND U157 ( .A(B[6]), .B(A[20]), .Z(\_38_net_[26] ) );
  AND U158 ( .A(B[5]), .B(A[20]), .Z(\_38_net_[25] ) );
  AND U159 ( .A(B[4]), .B(A[20]), .Z(\_38_net_[24] ) );
  AND U160 ( .A(B[3]), .B(A[20]), .Z(\_38_net_[23] ) );
  AND U161 ( .A(B[2]), .B(A[20]), .Z(\_38_net_[22] ) );
  AND U162 ( .A(B[1]), .B(A[20]), .Z(\_38_net_[21] ) );
  AND U163 ( .A(A[20]), .B(B[0]), .Z(\_38_net_[20] ) );
  AND U164 ( .A(B[12]), .B(A[19]), .Z(\_36_net_[31] ) );
  AND U165 ( .A(B[11]), .B(A[19]), .Z(\_36_net_[30] ) );
  AND U166 ( .A(B[10]), .B(A[19]), .Z(\_36_net_[29] ) );
  AND U167 ( .A(B[9]), .B(A[19]), .Z(\_36_net_[28] ) );
  AND U168 ( .A(B[8]), .B(A[19]), .Z(\_36_net_[27] ) );
  AND U169 ( .A(B[7]), .B(A[19]), .Z(\_36_net_[26] ) );
  AND U170 ( .A(B[6]), .B(A[19]), .Z(\_36_net_[25] ) );
  AND U171 ( .A(B[5]), .B(A[19]), .Z(\_36_net_[24] ) );
  AND U172 ( .A(B[4]), .B(A[19]), .Z(\_36_net_[23] ) );
  AND U173 ( .A(B[3]), .B(A[19]), .Z(\_36_net_[22] ) );
  AND U174 ( .A(B[2]), .B(A[19]), .Z(\_36_net_[21] ) );
  AND U175 ( .A(B[1]), .B(A[19]), .Z(\_36_net_[20] ) );
  AND U176 ( .A(A[19]), .B(B[0]), .Z(\_36_net_[19] ) );
  AND U177 ( .A(B[13]), .B(A[18]), .Z(\_34_net_[31] ) );
  AND U178 ( .A(B[12]), .B(A[18]), .Z(\_34_net_[30] ) );
  AND U179 ( .A(B[11]), .B(A[18]), .Z(\_34_net_[29] ) );
  AND U180 ( .A(B[10]), .B(A[18]), .Z(\_34_net_[28] ) );
  AND U181 ( .A(B[9]), .B(A[18]), .Z(\_34_net_[27] ) );
  AND U182 ( .A(B[8]), .B(A[18]), .Z(\_34_net_[26] ) );
  AND U183 ( .A(B[7]), .B(A[18]), .Z(\_34_net_[25] ) );
  AND U184 ( .A(B[6]), .B(A[18]), .Z(\_34_net_[24] ) );
  AND U185 ( .A(B[5]), .B(A[18]), .Z(\_34_net_[23] ) );
  AND U186 ( .A(B[4]), .B(A[18]), .Z(\_34_net_[22] ) );
  AND U187 ( .A(B[3]), .B(A[18]), .Z(\_34_net_[21] ) );
  AND U188 ( .A(B[2]), .B(A[18]), .Z(\_34_net_[20] ) );
  AND U189 ( .A(B[1]), .B(A[18]), .Z(\_34_net_[19] ) );
  AND U190 ( .A(A[18]), .B(B[0]), .Z(\_34_net_[18] ) );
  AND U191 ( .A(B[14]), .B(A[17]), .Z(\_32_net_[31] ) );
  AND U192 ( .A(B[13]), .B(A[17]), .Z(\_32_net_[30] ) );
  AND U193 ( .A(B[12]), .B(A[17]), .Z(\_32_net_[29] ) );
  AND U194 ( .A(B[11]), .B(A[17]), .Z(\_32_net_[28] ) );
  AND U195 ( .A(B[10]), .B(A[17]), .Z(\_32_net_[27] ) );
  AND U196 ( .A(B[9]), .B(A[17]), .Z(\_32_net_[26] ) );
  AND U197 ( .A(B[8]), .B(A[17]), .Z(\_32_net_[25] ) );
  AND U198 ( .A(B[7]), .B(A[17]), .Z(\_32_net_[24] ) );
  AND U199 ( .A(B[6]), .B(A[17]), .Z(\_32_net_[23] ) );
  AND U200 ( .A(B[5]), .B(A[17]), .Z(\_32_net_[22] ) );
  AND U201 ( .A(B[4]), .B(A[17]), .Z(\_32_net_[21] ) );
  AND U202 ( .A(B[3]), .B(A[17]), .Z(\_32_net_[20] ) );
  AND U203 ( .A(B[2]), .B(A[17]), .Z(\_32_net_[19] ) );
  AND U204 ( .A(B[1]), .B(A[17]), .Z(\_32_net_[18] ) );
  AND U205 ( .A(A[17]), .B(B[0]), .Z(\_32_net_[17] ) );
  AND U206 ( .A(B[15]), .B(A[16]), .Z(\_30_net_[31] ) );
  AND U207 ( .A(B[14]), .B(A[16]), .Z(\_30_net_[30] ) );
  AND U208 ( .A(B[13]), .B(A[16]), .Z(\_30_net_[29] ) );
  AND U209 ( .A(B[12]), .B(A[16]), .Z(\_30_net_[28] ) );
  AND U210 ( .A(B[11]), .B(A[16]), .Z(\_30_net_[27] ) );
  AND U211 ( .A(B[10]), .B(A[16]), .Z(\_30_net_[26] ) );
  AND U212 ( .A(B[9]), .B(A[16]), .Z(\_30_net_[25] ) );
  AND U213 ( .A(B[8]), .B(A[16]), .Z(\_30_net_[24] ) );
  AND U214 ( .A(B[7]), .B(A[16]), .Z(\_30_net_[23] ) );
  AND U215 ( .A(B[6]), .B(A[16]), .Z(\_30_net_[22] ) );
  AND U216 ( .A(B[5]), .B(A[16]), .Z(\_30_net_[21] ) );
  AND U217 ( .A(B[4]), .B(A[16]), .Z(\_30_net_[20] ) );
  AND U218 ( .A(B[3]), .B(A[16]), .Z(\_30_net_[19] ) );
  AND U219 ( .A(B[2]), .B(A[16]), .Z(\_30_net_[18] ) );
  AND U220 ( .A(B[1]), .B(A[16]), .Z(\_30_net_[17] ) );
  AND U221 ( .A(A[16]), .B(B[0]), .Z(\_30_net_[16] ) );
  AND U222 ( .A(B[7]), .B(A[2]), .Z(\_2_net_[9] ) );
  AND U223 ( .A(B[6]), .B(A[2]), .Z(\_2_net_[8] ) );
  AND U224 ( .A(B[5]), .B(A[2]), .Z(\_2_net_[7] ) );
  AND U225 ( .A(B[4]), .B(A[2]), .Z(\_2_net_[6] ) );
  AND U226 ( .A(B[3]), .B(A[2]), .Z(\_2_net_[5] ) );
  AND U227 ( .A(B[2]), .B(A[2]), .Z(\_2_net_[4] ) );
  AND U228 ( .A(B[1]), .B(A[2]), .Z(\_2_net_[3] ) );
  AND U229 ( .A(A[2]), .B(B[29]), .Z(\_2_net_[31] ) );
  AND U230 ( .A(B[28]), .B(A[2]), .Z(\_2_net_[30] ) );
  AND U231 ( .A(B[0]), .B(A[2]), .Z(\_2_net_[2] ) );
  AND U232 ( .A(B[27]), .B(A[2]), .Z(\_2_net_[29] ) );
  AND U233 ( .A(B[26]), .B(A[2]), .Z(\_2_net_[28] ) );
  AND U234 ( .A(B[25]), .B(A[2]), .Z(\_2_net_[27] ) );
  AND U235 ( .A(B[24]), .B(A[2]), .Z(\_2_net_[26] ) );
  AND U236 ( .A(B[23]), .B(A[2]), .Z(\_2_net_[25] ) );
  AND U237 ( .A(B[22]), .B(A[2]), .Z(\_2_net_[24] ) );
  AND U238 ( .A(B[21]), .B(A[2]), .Z(\_2_net_[23] ) );
  AND U239 ( .A(B[20]), .B(A[2]), .Z(\_2_net_[22] ) );
  AND U240 ( .A(B[19]), .B(A[2]), .Z(\_2_net_[21] ) );
  AND U241 ( .A(B[18]), .B(A[2]), .Z(\_2_net_[20] ) );
  AND U242 ( .A(B[17]), .B(A[2]), .Z(\_2_net_[19] ) );
  AND U243 ( .A(B[16]), .B(A[2]), .Z(\_2_net_[18] ) );
  AND U244 ( .A(B[15]), .B(A[2]), .Z(\_2_net_[17] ) );
  AND U245 ( .A(B[14]), .B(A[2]), .Z(\_2_net_[16] ) );
  AND U246 ( .A(B[13]), .B(A[2]), .Z(\_2_net_[15] ) );
  AND U247 ( .A(B[12]), .B(A[2]), .Z(\_2_net_[14] ) );
  AND U248 ( .A(B[11]), .B(A[2]), .Z(\_2_net_[13] ) );
  AND U249 ( .A(B[10]), .B(A[2]), .Z(\_2_net_[12] ) );
  AND U250 ( .A(B[9]), .B(A[2]), .Z(\_2_net_[11] ) );
  AND U251 ( .A(B[8]), .B(A[2]), .Z(\_2_net_[10] ) );
  AND U252 ( .A(B[16]), .B(A[15]), .Z(\_28_net_[31] ) );
  AND U253 ( .A(B[15]), .B(A[15]), .Z(\_28_net_[30] ) );
  AND U254 ( .A(B[14]), .B(A[15]), .Z(\_28_net_[29] ) );
  AND U255 ( .A(B[13]), .B(A[15]), .Z(\_28_net_[28] ) );
  AND U256 ( .A(B[12]), .B(A[15]), .Z(\_28_net_[27] ) );
  AND U257 ( .A(B[11]), .B(A[15]), .Z(\_28_net_[26] ) );
  AND U258 ( .A(B[10]), .B(A[15]), .Z(\_28_net_[25] ) );
  AND U259 ( .A(B[9]), .B(A[15]), .Z(\_28_net_[24] ) );
  AND U260 ( .A(B[8]), .B(A[15]), .Z(\_28_net_[23] ) );
  AND U261 ( .A(B[7]), .B(A[15]), .Z(\_28_net_[22] ) );
  AND U262 ( .A(B[6]), .B(A[15]), .Z(\_28_net_[21] ) );
  AND U263 ( .A(B[5]), .B(A[15]), .Z(\_28_net_[20] ) );
  AND U264 ( .A(B[4]), .B(A[15]), .Z(\_28_net_[19] ) );
  AND U265 ( .A(B[3]), .B(A[15]), .Z(\_28_net_[18] ) );
  AND U266 ( .A(B[2]), .B(A[15]), .Z(\_28_net_[17] ) );
  AND U267 ( .A(B[1]), .B(A[15]), .Z(\_28_net_[16] ) );
  AND U268 ( .A(A[15]), .B(B[0]), .Z(\_28_net_[15] ) );
  AND U269 ( .A(B[17]), .B(A[14]), .Z(\_26_net_[31] ) );
  AND U270 ( .A(B[16]), .B(A[14]), .Z(\_26_net_[30] ) );
  AND U271 ( .A(B[15]), .B(A[14]), .Z(\_26_net_[29] ) );
  AND U272 ( .A(B[14]), .B(A[14]), .Z(\_26_net_[28] ) );
  AND U273 ( .A(B[13]), .B(A[14]), .Z(\_26_net_[27] ) );
  AND U274 ( .A(B[12]), .B(A[14]), .Z(\_26_net_[26] ) );
  AND U275 ( .A(B[11]), .B(A[14]), .Z(\_26_net_[25] ) );
  AND U276 ( .A(B[10]), .B(A[14]), .Z(\_26_net_[24] ) );
  AND U277 ( .A(B[9]), .B(A[14]), .Z(\_26_net_[23] ) );
  AND U278 ( .A(B[8]), .B(A[14]), .Z(\_26_net_[22] ) );
  AND U279 ( .A(B[7]), .B(A[14]), .Z(\_26_net_[21] ) );
  AND U280 ( .A(B[6]), .B(A[14]), .Z(\_26_net_[20] ) );
  AND U281 ( .A(B[5]), .B(A[14]), .Z(\_26_net_[19] ) );
  AND U282 ( .A(B[4]), .B(A[14]), .Z(\_26_net_[18] ) );
  AND U283 ( .A(B[3]), .B(A[14]), .Z(\_26_net_[17] ) );
  AND U284 ( .A(B[2]), .B(A[14]), .Z(\_26_net_[16] ) );
  AND U285 ( .A(B[1]), .B(A[14]), .Z(\_26_net_[15] ) );
  AND U286 ( .A(A[14]), .B(B[0]), .Z(\_26_net_[14] ) );
  AND U287 ( .A(B[18]), .B(A[13]), .Z(\_24_net_[31] ) );
  AND U288 ( .A(B[17]), .B(A[13]), .Z(\_24_net_[30] ) );
  AND U289 ( .A(B[16]), .B(A[13]), .Z(\_24_net_[29] ) );
  AND U290 ( .A(B[15]), .B(A[13]), .Z(\_24_net_[28] ) );
  AND U291 ( .A(B[14]), .B(A[13]), .Z(\_24_net_[27] ) );
  AND U292 ( .A(B[13]), .B(A[13]), .Z(\_24_net_[26] ) );
  AND U293 ( .A(B[12]), .B(A[13]), .Z(\_24_net_[25] ) );
  AND U294 ( .A(B[11]), .B(A[13]), .Z(\_24_net_[24] ) );
  AND U295 ( .A(B[10]), .B(A[13]), .Z(\_24_net_[23] ) );
  AND U296 ( .A(B[9]), .B(A[13]), .Z(\_24_net_[22] ) );
  AND U297 ( .A(B[8]), .B(A[13]), .Z(\_24_net_[21] ) );
  AND U298 ( .A(B[7]), .B(A[13]), .Z(\_24_net_[20] ) );
  AND U299 ( .A(B[6]), .B(A[13]), .Z(\_24_net_[19] ) );
  AND U300 ( .A(B[5]), .B(A[13]), .Z(\_24_net_[18] ) );
  AND U301 ( .A(B[4]), .B(A[13]), .Z(\_24_net_[17] ) );
  AND U302 ( .A(B[3]), .B(A[13]), .Z(\_24_net_[16] ) );
  AND U303 ( .A(B[2]), .B(A[13]), .Z(\_24_net_[15] ) );
  AND U304 ( .A(B[1]), .B(A[13]), .Z(\_24_net_[14] ) );
  AND U305 ( .A(A[13]), .B(B[0]), .Z(\_24_net_[13] ) );
  AND U306 ( .A(B[19]), .B(A[12]), .Z(\_22_net_[31] ) );
  AND U307 ( .A(B[18]), .B(A[12]), .Z(\_22_net_[30] ) );
  AND U308 ( .A(B[17]), .B(A[12]), .Z(\_22_net_[29] ) );
  AND U309 ( .A(B[16]), .B(A[12]), .Z(\_22_net_[28] ) );
  AND U310 ( .A(B[15]), .B(A[12]), .Z(\_22_net_[27] ) );
  AND U311 ( .A(B[14]), .B(A[12]), .Z(\_22_net_[26] ) );
  AND U312 ( .A(B[13]), .B(A[12]), .Z(\_22_net_[25] ) );
  AND U313 ( .A(B[12]), .B(A[12]), .Z(\_22_net_[24] ) );
  AND U314 ( .A(B[11]), .B(A[12]), .Z(\_22_net_[23] ) );
  AND U315 ( .A(B[10]), .B(A[12]), .Z(\_22_net_[22] ) );
  AND U316 ( .A(B[9]), .B(A[12]), .Z(\_22_net_[21] ) );
  AND U317 ( .A(B[8]), .B(A[12]), .Z(\_22_net_[20] ) );
  AND U318 ( .A(B[7]), .B(A[12]), .Z(\_22_net_[19] ) );
  AND U319 ( .A(B[6]), .B(A[12]), .Z(\_22_net_[18] ) );
  AND U320 ( .A(B[5]), .B(A[12]), .Z(\_22_net_[17] ) );
  AND U321 ( .A(B[4]), .B(A[12]), .Z(\_22_net_[16] ) );
  AND U322 ( .A(B[3]), .B(A[12]), .Z(\_22_net_[15] ) );
  AND U323 ( .A(B[2]), .B(A[12]), .Z(\_22_net_[14] ) );
  AND U324 ( .A(B[1]), .B(A[12]), .Z(\_22_net_[13] ) );
  AND U325 ( .A(A[12]), .B(B[0]), .Z(\_22_net_[12] ) );
  AND U326 ( .A(B[20]), .B(A[11]), .Z(\_20_net_[31] ) );
  AND U327 ( .A(B[19]), .B(A[11]), .Z(\_20_net_[30] ) );
  AND U328 ( .A(B[18]), .B(A[11]), .Z(\_20_net_[29] ) );
  AND U329 ( .A(B[17]), .B(A[11]), .Z(\_20_net_[28] ) );
  AND U330 ( .A(B[16]), .B(A[11]), .Z(\_20_net_[27] ) );
  AND U331 ( .A(B[15]), .B(A[11]), .Z(\_20_net_[26] ) );
  AND U332 ( .A(B[14]), .B(A[11]), .Z(\_20_net_[25] ) );
  AND U333 ( .A(B[13]), .B(A[11]), .Z(\_20_net_[24] ) );
  AND U334 ( .A(B[12]), .B(A[11]), .Z(\_20_net_[23] ) );
  AND U335 ( .A(B[11]), .B(A[11]), .Z(\_20_net_[22] ) );
  AND U336 ( .A(B[10]), .B(A[11]), .Z(\_20_net_[21] ) );
  AND U337 ( .A(B[9]), .B(A[11]), .Z(\_20_net_[20] ) );
  AND U338 ( .A(B[8]), .B(A[11]), .Z(\_20_net_[19] ) );
  AND U339 ( .A(B[7]), .B(A[11]), .Z(\_20_net_[18] ) );
  AND U340 ( .A(B[6]), .B(A[11]), .Z(\_20_net_[17] ) );
  AND U341 ( .A(B[5]), .B(A[11]), .Z(\_20_net_[16] ) );
  AND U342 ( .A(B[4]), .B(A[11]), .Z(\_20_net_[15] ) );
  AND U343 ( .A(B[3]), .B(A[11]), .Z(\_20_net_[14] ) );
  AND U344 ( .A(B[2]), .B(A[11]), .Z(\_20_net_[13] ) );
  AND U345 ( .A(B[1]), .B(A[11]), .Z(\_20_net_[12] ) );
  AND U346 ( .A(A[11]), .B(B[0]), .Z(\_20_net_[11] ) );
  AND U347 ( .A(B[21]), .B(A[10]), .Z(\_18_net_[31] ) );
  AND U348 ( .A(B[20]), .B(A[10]), .Z(\_18_net_[30] ) );
  AND U349 ( .A(B[19]), .B(A[10]), .Z(\_18_net_[29] ) );
  AND U350 ( .A(B[18]), .B(A[10]), .Z(\_18_net_[28] ) );
  AND U351 ( .A(B[17]), .B(A[10]), .Z(\_18_net_[27] ) );
  AND U352 ( .A(B[16]), .B(A[10]), .Z(\_18_net_[26] ) );
  AND U353 ( .A(B[15]), .B(A[10]), .Z(\_18_net_[25] ) );
  AND U354 ( .A(B[14]), .B(A[10]), .Z(\_18_net_[24] ) );
  AND U355 ( .A(B[13]), .B(A[10]), .Z(\_18_net_[23] ) );
  AND U356 ( .A(B[12]), .B(A[10]), .Z(\_18_net_[22] ) );
  AND U357 ( .A(B[11]), .B(A[10]), .Z(\_18_net_[21] ) );
  AND U358 ( .A(B[10]), .B(A[10]), .Z(\_18_net_[20] ) );
  AND U359 ( .A(B[9]), .B(A[10]), .Z(\_18_net_[19] ) );
  AND U360 ( .A(B[8]), .B(A[10]), .Z(\_18_net_[18] ) );
  AND U361 ( .A(B[7]), .B(A[10]), .Z(\_18_net_[17] ) );
  AND U362 ( .A(B[6]), .B(A[10]), .Z(\_18_net_[16] ) );
  AND U363 ( .A(B[5]), .B(A[10]), .Z(\_18_net_[15] ) );
  AND U364 ( .A(B[4]), .B(A[10]), .Z(\_18_net_[14] ) );
  AND U365 ( .A(B[3]), .B(A[10]), .Z(\_18_net_[13] ) );
  AND U366 ( .A(B[2]), .B(A[10]), .Z(\_18_net_[12] ) );
  AND U367 ( .A(B[1]), .B(A[10]), .Z(\_18_net_[11] ) );
  AND U368 ( .A(A[10]), .B(B[0]), .Z(\_18_net_[10] ) );
  AND U369 ( .A(B[0]), .B(A[9]), .Z(\_16_net_[9] ) );
  AND U370 ( .A(B[22]), .B(A[9]), .Z(\_16_net_[31] ) );
  AND U371 ( .A(B[21]), .B(A[9]), .Z(\_16_net_[30] ) );
  AND U372 ( .A(B[20]), .B(A[9]), .Z(\_16_net_[29] ) );
  AND U373 ( .A(B[19]), .B(A[9]), .Z(\_16_net_[28] ) );
  AND U374 ( .A(B[18]), .B(A[9]), .Z(\_16_net_[27] ) );
  AND U375 ( .A(B[17]), .B(A[9]), .Z(\_16_net_[26] ) );
  AND U376 ( .A(B[16]), .B(A[9]), .Z(\_16_net_[25] ) );
  AND U377 ( .A(B[15]), .B(A[9]), .Z(\_16_net_[24] ) );
  AND U378 ( .A(B[14]), .B(A[9]), .Z(\_16_net_[23] ) );
  AND U379 ( .A(B[13]), .B(A[9]), .Z(\_16_net_[22] ) );
  AND U380 ( .A(B[12]), .B(A[9]), .Z(\_16_net_[21] ) );
  AND U381 ( .A(B[11]), .B(A[9]), .Z(\_16_net_[20] ) );
  AND U382 ( .A(B[10]), .B(A[9]), .Z(\_16_net_[19] ) );
  AND U383 ( .A(B[9]), .B(A[9]), .Z(\_16_net_[18] ) );
  AND U384 ( .A(B[8]), .B(A[9]), .Z(\_16_net_[17] ) );
  AND U385 ( .A(B[7]), .B(A[9]), .Z(\_16_net_[16] ) );
  AND U386 ( .A(B[6]), .B(A[9]), .Z(\_16_net_[15] ) );
  AND U387 ( .A(B[5]), .B(A[9]), .Z(\_16_net_[14] ) );
  AND U388 ( .A(B[4]), .B(A[9]), .Z(\_16_net_[13] ) );
  AND U389 ( .A(B[3]), .B(A[9]), .Z(\_16_net_[12] ) );
  AND U390 ( .A(B[2]), .B(A[9]), .Z(\_16_net_[11] ) );
  AND U391 ( .A(A[9]), .B(B[1]), .Z(\_16_net_[10] ) );
  AND U392 ( .A(B[1]), .B(A[8]), .Z(\_14_net_[9] ) );
  AND U393 ( .A(B[0]), .B(A[8]), .Z(\_14_net_[8] ) );
  AND U394 ( .A(B[23]), .B(A[8]), .Z(\_14_net_[31] ) );
  AND U395 ( .A(B[22]), .B(A[8]), .Z(\_14_net_[30] ) );
  AND U396 ( .A(B[21]), .B(A[8]), .Z(\_14_net_[29] ) );
  AND U397 ( .A(B[20]), .B(A[8]), .Z(\_14_net_[28] ) );
  AND U398 ( .A(B[19]), .B(A[8]), .Z(\_14_net_[27] ) );
  AND U399 ( .A(B[18]), .B(A[8]), .Z(\_14_net_[26] ) );
  AND U400 ( .A(B[17]), .B(A[8]), .Z(\_14_net_[25] ) );
  AND U401 ( .A(B[16]), .B(A[8]), .Z(\_14_net_[24] ) );
  AND U402 ( .A(B[15]), .B(A[8]), .Z(\_14_net_[23] ) );
  AND U403 ( .A(B[14]), .B(A[8]), .Z(\_14_net_[22] ) );
  AND U404 ( .A(B[13]), .B(A[8]), .Z(\_14_net_[21] ) );
  AND U405 ( .A(B[12]), .B(A[8]), .Z(\_14_net_[20] ) );
  AND U406 ( .A(B[11]), .B(A[8]), .Z(\_14_net_[19] ) );
  AND U407 ( .A(B[10]), .B(A[8]), .Z(\_14_net_[18] ) );
  AND U408 ( .A(B[9]), .B(A[8]), .Z(\_14_net_[17] ) );
  AND U409 ( .A(B[8]), .B(A[8]), .Z(\_14_net_[16] ) );
  AND U410 ( .A(B[7]), .B(A[8]), .Z(\_14_net_[15] ) );
  AND U411 ( .A(B[6]), .B(A[8]), .Z(\_14_net_[14] ) );
  AND U412 ( .A(B[5]), .B(A[8]), .Z(\_14_net_[13] ) );
  AND U413 ( .A(B[4]), .B(A[8]), .Z(\_14_net_[12] ) );
  AND U414 ( .A(B[3]), .B(A[8]), .Z(\_14_net_[11] ) );
  AND U415 ( .A(A[8]), .B(B[2]), .Z(\_14_net_[10] ) );
  AND U416 ( .A(B[2]), .B(A[7]), .Z(\_12_net_[9] ) );
  AND U417 ( .A(B[1]), .B(A[7]), .Z(\_12_net_[8] ) );
  AND U418 ( .A(B[0]), .B(A[7]), .Z(\_12_net_[7] ) );
  AND U419 ( .A(B[24]), .B(A[7]), .Z(\_12_net_[31] ) );
  AND U420 ( .A(B[23]), .B(A[7]), .Z(\_12_net_[30] ) );
  AND U421 ( .A(B[22]), .B(A[7]), .Z(\_12_net_[29] ) );
  AND U422 ( .A(B[21]), .B(A[7]), .Z(\_12_net_[28] ) );
  AND U423 ( .A(B[20]), .B(A[7]), .Z(\_12_net_[27] ) );
  AND U424 ( .A(B[19]), .B(A[7]), .Z(\_12_net_[26] ) );
  AND U425 ( .A(B[18]), .B(A[7]), .Z(\_12_net_[25] ) );
  AND U426 ( .A(B[17]), .B(A[7]), .Z(\_12_net_[24] ) );
  AND U427 ( .A(B[16]), .B(A[7]), .Z(\_12_net_[23] ) );
  AND U428 ( .A(B[15]), .B(A[7]), .Z(\_12_net_[22] ) );
  AND U429 ( .A(B[14]), .B(A[7]), .Z(\_12_net_[21] ) );
  AND U430 ( .A(B[13]), .B(A[7]), .Z(\_12_net_[20] ) );
  AND U431 ( .A(B[12]), .B(A[7]), .Z(\_12_net_[19] ) );
  AND U432 ( .A(B[11]), .B(A[7]), .Z(\_12_net_[18] ) );
  AND U433 ( .A(B[10]), .B(A[7]), .Z(\_12_net_[17] ) );
  AND U434 ( .A(B[9]), .B(A[7]), .Z(\_12_net_[16] ) );
  AND U435 ( .A(B[8]), .B(A[7]), .Z(\_12_net_[15] ) );
  AND U436 ( .A(B[7]), .B(A[7]), .Z(\_12_net_[14] ) );
  AND U437 ( .A(B[6]), .B(A[7]), .Z(\_12_net_[13] ) );
  AND U438 ( .A(B[5]), .B(A[7]), .Z(\_12_net_[12] ) );
  AND U439 ( .A(B[4]), .B(A[7]), .Z(\_12_net_[11] ) );
  AND U440 ( .A(A[7]), .B(B[3]), .Z(\_12_net_[10] ) );
  AND U441 ( .A(B[3]), .B(A[6]), .Z(\_10_net_[9] ) );
  AND U442 ( .A(B[2]), .B(A[6]), .Z(\_10_net_[8] ) );
  AND U443 ( .A(B[1]), .B(A[6]), .Z(\_10_net_[7] ) );
  AND U444 ( .A(B[0]), .B(A[6]), .Z(\_10_net_[6] ) );
  AND U445 ( .A(B[25]), .B(A[6]), .Z(\_10_net_[31] ) );
  AND U446 ( .A(B[24]), .B(A[6]), .Z(\_10_net_[30] ) );
  AND U447 ( .A(B[23]), .B(A[6]), .Z(\_10_net_[29] ) );
  AND U448 ( .A(B[22]), .B(A[6]), .Z(\_10_net_[28] ) );
  AND U449 ( .A(B[21]), .B(A[6]), .Z(\_10_net_[27] ) );
  AND U450 ( .A(B[20]), .B(A[6]), .Z(\_10_net_[26] ) );
  AND U451 ( .A(B[19]), .B(A[6]), .Z(\_10_net_[25] ) );
  AND U452 ( .A(B[18]), .B(A[6]), .Z(\_10_net_[24] ) );
  AND U453 ( .A(B[17]), .B(A[6]), .Z(\_10_net_[23] ) );
  AND U454 ( .A(B[16]), .B(A[6]), .Z(\_10_net_[22] ) );
  AND U455 ( .A(B[15]), .B(A[6]), .Z(\_10_net_[21] ) );
  AND U456 ( .A(B[14]), .B(A[6]), .Z(\_10_net_[20] ) );
  AND U457 ( .A(B[13]), .B(A[6]), .Z(\_10_net_[19] ) );
  AND U458 ( .A(B[12]), .B(A[6]), .Z(\_10_net_[18] ) );
  AND U459 ( .A(B[11]), .B(A[6]), .Z(\_10_net_[17] ) );
  AND U460 ( .A(B[10]), .B(A[6]), .Z(\_10_net_[16] ) );
  AND U461 ( .A(B[9]), .B(A[6]), .Z(\_10_net_[15] ) );
  AND U462 ( .A(B[8]), .B(A[6]), .Z(\_10_net_[14] ) );
  AND U463 ( .A(B[7]), .B(A[6]), .Z(\_10_net_[13] ) );
  AND U464 ( .A(B[6]), .B(A[6]), .Z(\_10_net_[12] ) );
  AND U465 ( .A(B[5]), .B(A[6]), .Z(\_10_net_[11] ) );
  AND U466 ( .A(A[6]), .B(B[4]), .Z(\_10_net_[10] ) );
  AND U467 ( .A(B[8]), .B(A[1]), .Z(\_0_net_[9] ) );
  AND U468 ( .A(B[7]), .B(A[1]), .Z(\_0_net_[8] ) );
  AND U469 ( .A(B[6]), .B(A[1]), .Z(\_0_net_[7] ) );
  AND U470 ( .A(B[5]), .B(A[1]), .Z(\_0_net_[6] ) );
  AND U471 ( .A(B[4]), .B(A[1]), .Z(\_0_net_[5] ) );
  AND U472 ( .A(B[3]), .B(A[1]), .Z(\_0_net_[4] ) );
  AND U473 ( .A(B[2]), .B(A[1]), .Z(\_0_net_[3] ) );
  AND U474 ( .A(B[30]), .B(A[1]), .Z(\_0_net_[31] ) );
  AND U475 ( .A(B[29]), .B(A[1]), .Z(\_0_net_[30] ) );
  AND U476 ( .A(B[1]), .B(A[1]), .Z(\_0_net_[2] ) );
  AND U477 ( .A(B[28]), .B(A[1]), .Z(\_0_net_[29] ) );
  AND U478 ( .A(B[27]), .B(A[1]), .Z(\_0_net_[28] ) );
  AND U479 ( .A(B[26]), .B(A[1]), .Z(\_0_net_[27] ) );
  AND U480 ( .A(B[25]), .B(A[1]), .Z(\_0_net_[26] ) );
  AND U481 ( .A(B[24]), .B(A[1]), .Z(\_0_net_[25] ) );
  AND U482 ( .A(B[23]), .B(A[1]), .Z(\_0_net_[24] ) );
  AND U483 ( .A(B[22]), .B(A[1]), .Z(\_0_net_[23] ) );
  AND U484 ( .A(B[21]), .B(A[1]), .Z(\_0_net_[22] ) );
  AND U485 ( .A(B[20]), .B(A[1]), .Z(\_0_net_[21] ) );
  AND U486 ( .A(B[19]), .B(A[1]), .Z(\_0_net_[20] ) );
  AND U487 ( .A(B[0]), .B(A[1]), .Z(\_0_net_[1] ) );
  AND U488 ( .A(B[18]), .B(A[1]), .Z(\_0_net_[19] ) );
  AND U489 ( .A(B[17]), .B(A[1]), .Z(\_0_net_[18] ) );
  AND U490 ( .A(B[16]), .B(A[1]), .Z(\_0_net_[17] ) );
  AND U491 ( .A(B[15]), .B(A[1]), .Z(\_0_net_[16] ) );
  AND U492 ( .A(B[14]), .B(A[1]), .Z(\_0_net_[15] ) );
  AND U493 ( .A(B[13]), .B(A[1]), .Z(\_0_net_[14] ) );
  AND U494 ( .A(B[12]), .B(A[1]), .Z(\_0_net_[13] ) );
  AND U495 ( .A(B[11]), .B(A[1]), .Z(\_0_net_[12] ) );
  AND U496 ( .A(B[10]), .B(A[1]), .Z(\_0_net_[11] ) );
  AND U497 ( .A(A[1]), .B(B[9]), .Z(\_0_net_[10] ) );
endmodule


module FA_2977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_2978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N32_94 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3007 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_3006 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_3005 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_3004 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_3003 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_3002 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3001 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3000 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_2999 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_2998 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2997 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2996 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2995 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2994 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2993 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2992 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2991 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2990 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2989 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2988 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2987 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2986 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2985 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2984 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2983 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2982 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2981 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2980 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2979 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2978 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2977 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N32_95 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3039 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_3038 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_3037 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_3036 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_3035 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_3034 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3033 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3032 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3031 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3030 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3029 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3028 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3027 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3026 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3025 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3024 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3023 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3022 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3021 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3020 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3019 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3018 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3017 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3016 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3015 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3014 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3013 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3012 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3011 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3010 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3009 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module matrixMult_N_M_2_N3_M32 ( clk, rst, x, y, o );
  input [95:0] x;
  input [95:0] y;
  output [31:0] o;
  input clk, rst;
  wire   \xyi[2][31] , \xyi[2][30] , \xyi[2][29] , \xyi[2][28] , \xyi[2][27] ,
         \xyi[2][26] , \xyi[2][25] , \xyi[2][24] , \xyi[2][23] , \xyi[2][22] ,
         \xyi[2][21] , \xyi[2][20] , \xyi[2][19] , \xyi[2][18] , \xyi[2][17] ,
         \xyi[2][16] , \xyi[2][15] , \xyi[2][14] , \xyi[2][13] , \xyi[2][12] ,
         \xyi[2][11] , \xyi[2][10] , \xyi[2][9] , \xyi[2][8] , \xyi[2][7] ,
         \xyi[2][6] , \xyi[2][5] , \xyi[2][4] , \xyi[2][3] , \xyi[2][2] ,
         \xyi[2][1] , \xyi[1][31] , \xyi[1][30] , \xyi[1][29] , \xyi[1][28] ,
         \xyi[1][27] , \xyi[1][26] , \xyi[1][25] , \xyi[1][24] , \xyi[1][23] ,
         \xyi[1][22] , \xyi[1][21] , \xyi[1][20] , \xyi[1][19] , \xyi[1][18] ,
         \xyi[1][17] , \xyi[1][16] , \xyi[1][15] , \xyi[1][14] , \xyi[1][13] ,
         \xyi[1][12] , \xyi[1][11] , \xyi[1][10] , \xyi[1][9] , \xyi[1][8] ,
         \xyi[1][7] , \xyi[1][6] , \xyi[1][5] , \xyi[1][4] , \xyi[1][3] ,
         \xyi[1][2] , \xyi[1][1] , \xyi[0][31] , \xyi[0][30] , \xyi[0][29] ,
         \xyi[0][28] , \xyi[0][27] , \xyi[0][26] , \xyi[0][25] , \xyi[0][24] ,
         \xyi[0][23] , \xyi[0][22] , \xyi[0][21] , \xyi[0][20] , \xyi[0][19] ,
         \xyi[0][18] , \xyi[0][17] , \xyi[0][16] , \xyi[0][15] , \xyi[0][14] ,
         \xyi[0][13] , \xyi[0][12] , \xyi[0][11] , \xyi[0][10] , \xyi[0][9] ,
         \xyi[0][8] , \xyi[0][7] , \xyi[0][6] , \xyi[0][5] , \xyi[0][4] ,
         \xyi[0][3] , \xyi[0][2] , \xyi[0][1] , \oi[3][31] , \oi[3][30] ,
         \oi[3][29] , \oi[3][28] , \oi[3][27] , \oi[3][26] , \oi[3][25] ,
         \oi[3][24] , \oi[3][23] , \oi[3][22] , \oi[3][21] , \oi[3][20] ,
         \oi[3][19] , \oi[3][18] , \oi[3][17] , \oi[3][16] , \oi[3][15] ,
         \oi[3][14] , \oi[3][13] , \oi[3][12] , \oi[3][11] , \oi[3][10] ,
         \oi[3][9] , \oi[3][8] , \oi[3][7] , \oi[3][6] , \oi[3][5] ,
         \oi[3][4] , \oi[3][3] , \oi[3][2] , \oi[3][1] , \oi[2][31] ,
         \oi[2][30] , \oi[2][29] , \oi[2][28] , \oi[2][27] , \oi[2][26] ,
         \oi[2][25] , \oi[2][24] , \oi[2][23] , \oi[2][22] , \oi[2][21] ,
         \oi[2][20] , \oi[2][19] , \oi[2][18] , \oi[2][17] , \oi[2][16] ,
         \oi[2][15] , \oi[2][14] , \oi[2][13] , \oi[2][12] , \oi[2][11] ,
         \oi[2][10] , \oi[2][9] , \oi[2][8] , \oi[2][7] , \oi[2][6] ,
         \oi[2][5] , \oi[2][4] , \oi[2][3] , \oi[2][2] , \oi[2][1] ,
         \oi[1][31] , \oi[1][30] , \oi[1][29] , \oi[1][28] , \oi[1][27] ,
         \oi[1][26] , \oi[1][25] , \oi[1][24] , \oi[1][23] , \oi[1][22] ,
         \oi[1][21] , \oi[1][20] , \oi[1][19] , \oi[1][18] , \oi[1][17] ,
         \oi[1][16] , \oi[1][15] , \oi[1][14] , \oi[1][13] , \oi[1][12] ,
         \oi[1][11] , \oi[1][10] , \oi[1][9] , \oi[1][8] , \oi[1][7] ,
         \oi[1][6] , \oi[1][5] , \oi[1][4] , \oi[1][3] , \oi[1][2] ,
         \oi[1][1] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5;
  assign o[0] = 1'b0;

  MULT_N32_0 \MMULT_ROW[0].MULT_  ( .A({x[31:1], 1'b0}), .B({1'b0, y[30:0]}), 
        .O({\xyi[0][31] , \xyi[0][30] , \xyi[0][29] , \xyi[0][28] , 
        \xyi[0][27] , \xyi[0][26] , \xyi[0][25] , \xyi[0][24] , \xyi[0][23] , 
        \xyi[0][22] , \xyi[0][21] , \xyi[0][20] , \xyi[0][19] , \xyi[0][18] , 
        \xyi[0][17] , \xyi[0][16] , \xyi[0][15] , \xyi[0][14] , \xyi[0][13] , 
        \xyi[0][12] , \xyi[0][11] , \xyi[0][10] , \xyi[0][9] , \xyi[0][8] , 
        \xyi[0][7] , \xyi[0][6] , \xyi[0][5] , \xyi[0][4] , \xyi[0][3] , 
        \xyi[0][2] , \xyi[0][1] , SYNOPSYS_UNCONNECTED__0}) );
  MULT_N32_2 \MMULT_ROW[1].MULT_  ( .A({x[63:33], 1'b0}), .B({1'b0, y[62:32]}), 
        .O({\xyi[1][31] , \xyi[1][30] , \xyi[1][29] , \xyi[1][28] , 
        \xyi[1][27] , \xyi[1][26] , \xyi[1][25] , \xyi[1][24] , \xyi[1][23] , 
        \xyi[1][22] , \xyi[1][21] , \xyi[1][20] , \xyi[1][19] , \xyi[1][18] , 
        \xyi[1][17] , \xyi[1][16] , \xyi[1][15] , \xyi[1][14] , \xyi[1][13] , 
        \xyi[1][12] , \xyi[1][11] , \xyi[1][10] , \xyi[1][9] , \xyi[1][8] , 
        \xyi[1][7] , \xyi[1][6] , \xyi[1][5] , \xyi[1][4] , \xyi[1][3] , 
        \xyi[1][2] , \xyi[1][1] , SYNOPSYS_UNCONNECTED__1}) );
  MULT_N32_1 \MMULT_ROW[2].MULT_  ( .A({x[95:65], 1'b0}), .B({1'b0, y[94:64]}), 
        .O({\xyi[2][31] , \xyi[2][30] , \xyi[2][29] , \xyi[2][28] , 
        \xyi[2][27] , \xyi[2][26] , \xyi[2][25] , \xyi[2][24] , \xyi[2][23] , 
        \xyi[2][22] , \xyi[2][21] , \xyi[2][20] , \xyi[2][19] , \xyi[2][18] , 
        \xyi[2][17] , \xyi[2][16] , \xyi[2][15] , \xyi[2][14] , \xyi[2][13] , 
        \xyi[2][12] , \xyi[2][11] , \xyi[2][10] , \xyi[2][9] , \xyi[2][8] , 
        \xyi[2][7] , \xyi[2][6] , \xyi[2][5] , \xyi[2][4] , \xyi[2][3] , 
        \xyi[2][2] , \xyi[2][1] , SYNOPSYS_UNCONNECTED__2}) );
  ADD_N32_0 \ADD_ROW[0].ADD_  ( .A({\xyi[0][31] , \xyi[0][30] , \xyi[0][29] , 
        \xyi[0][28] , \xyi[0][27] , \xyi[0][26] , \xyi[0][25] , \xyi[0][24] , 
        \xyi[0][23] , \xyi[0][22] , \xyi[0][21] , \xyi[0][20] , \xyi[0][19] , 
        \xyi[0][18] , \xyi[0][17] , \xyi[0][16] , \xyi[0][15] , \xyi[0][14] , 
        \xyi[0][13] , \xyi[0][12] , \xyi[0][11] , \xyi[0][10] , \xyi[0][9] , 
        \xyi[0][8] , \xyi[0][7] , \xyi[0][6] , \xyi[0][5] , \xyi[0][4] , 
        \xyi[0][3] , \xyi[0][2] , \xyi[0][1] , 1'b0}), .B({o[31:1], 1'b0}), 
        .CI(1'b0), .S({\oi[1][31] , \oi[1][30] , \oi[1][29] , \oi[1][28] , 
        \oi[1][27] , \oi[1][26] , \oi[1][25] , \oi[1][24] , \oi[1][23] , 
        \oi[1][22] , \oi[1][21] , \oi[1][20] , \oi[1][19] , \oi[1][18] , 
        \oi[1][17] , \oi[1][16] , \oi[1][15] , \oi[1][14] , \oi[1][13] , 
        \oi[1][12] , \oi[1][11] , \oi[1][10] , \oi[1][9] , \oi[1][8] , 
        \oi[1][7] , \oi[1][6] , \oi[1][5] , \oi[1][4] , \oi[1][3] , \oi[1][2] , 
        \oi[1][1] , SYNOPSYS_UNCONNECTED__3}) );
  ADD_N32_95 \ADD_ROW[1].ADD_  ( .A({\xyi[1][31] , \xyi[1][30] , \xyi[1][29] , 
        \xyi[1][28] , \xyi[1][27] , \xyi[1][26] , \xyi[1][25] , \xyi[1][24] , 
        \xyi[1][23] , \xyi[1][22] , \xyi[1][21] , \xyi[1][20] , \xyi[1][19] , 
        \xyi[1][18] , \xyi[1][17] , \xyi[1][16] , \xyi[1][15] , \xyi[1][14] , 
        \xyi[1][13] , \xyi[1][12] , \xyi[1][11] , \xyi[1][10] , \xyi[1][9] , 
        \xyi[1][8] , \xyi[1][7] , \xyi[1][6] , \xyi[1][5] , \xyi[1][4] , 
        \xyi[1][3] , \xyi[1][2] , \xyi[1][1] , 1'b0}), .B({\oi[1][31] , 
        \oi[1][30] , \oi[1][29] , \oi[1][28] , \oi[1][27] , \oi[1][26] , 
        \oi[1][25] , \oi[1][24] , \oi[1][23] , \oi[1][22] , \oi[1][21] , 
        \oi[1][20] , \oi[1][19] , \oi[1][18] , \oi[1][17] , \oi[1][16] , 
        \oi[1][15] , \oi[1][14] , \oi[1][13] , \oi[1][12] , \oi[1][11] , 
        \oi[1][10] , \oi[1][9] , \oi[1][8] , \oi[1][7] , \oi[1][6] , 
        \oi[1][5] , \oi[1][4] , \oi[1][3] , \oi[1][2] , \oi[1][1] , 1'b0}), 
        .CI(1'b0), .S({\oi[2][31] , \oi[2][30] , \oi[2][29] , \oi[2][28] , 
        \oi[2][27] , \oi[2][26] , \oi[2][25] , \oi[2][24] , \oi[2][23] , 
        \oi[2][22] , \oi[2][21] , \oi[2][20] , \oi[2][19] , \oi[2][18] , 
        \oi[2][17] , \oi[2][16] , \oi[2][15] , \oi[2][14] , \oi[2][13] , 
        \oi[2][12] , \oi[2][11] , \oi[2][10] , \oi[2][9] , \oi[2][8] , 
        \oi[2][7] , \oi[2][6] , \oi[2][5] , \oi[2][4] , \oi[2][3] , \oi[2][2] , 
        \oi[2][1] , SYNOPSYS_UNCONNECTED__4}) );
  ADD_N32_94 \ADD_ROW[2].ADD_  ( .A({\xyi[2][31] , \xyi[2][30] , \xyi[2][29] , 
        \xyi[2][28] , \xyi[2][27] , \xyi[2][26] , \xyi[2][25] , \xyi[2][24] , 
        \xyi[2][23] , \xyi[2][22] , \xyi[2][21] , \xyi[2][20] , \xyi[2][19] , 
        \xyi[2][18] , \xyi[2][17] , \xyi[2][16] , \xyi[2][15] , \xyi[2][14] , 
        \xyi[2][13] , \xyi[2][12] , \xyi[2][11] , \xyi[2][10] , \xyi[2][9] , 
        \xyi[2][8] , \xyi[2][7] , \xyi[2][6] , \xyi[2][5] , \xyi[2][4] , 
        \xyi[2][3] , \xyi[2][2] , \xyi[2][1] , 1'b0}), .B({\oi[2][31] , 
        \oi[2][30] , \oi[2][29] , \oi[2][28] , \oi[2][27] , \oi[2][26] , 
        \oi[2][25] , \oi[2][24] , \oi[2][23] , \oi[2][22] , \oi[2][21] , 
        \oi[2][20] , \oi[2][19] , \oi[2][18] , \oi[2][17] , \oi[2][16] , 
        \oi[2][15] , \oi[2][14] , \oi[2][13] , \oi[2][12] , \oi[2][11] , 
        \oi[2][10] , \oi[2][9] , \oi[2][8] , \oi[2][7] , \oi[2][6] , 
        \oi[2][5] , \oi[2][4] , \oi[2][3] , \oi[2][2] , \oi[2][1] , 1'b0}), 
        .CI(1'b0), .S({\oi[3][31] , \oi[3][30] , \oi[3][29] , \oi[3][28] , 
        \oi[3][27] , \oi[3][26] , \oi[3][25] , \oi[3][24] , \oi[3][23] , 
        \oi[3][22] , \oi[3][21] , \oi[3][20] , \oi[3][19] , \oi[3][18] , 
        \oi[3][17] , \oi[3][16] , \oi[3][15] , \oi[3][14] , \oi[3][13] , 
        \oi[3][12] , \oi[3][11] , \oi[3][10] , \oi[3][9] , \oi[3][8] , 
        \oi[3][7] , \oi[3][6] , \oi[3][5] , \oi[3][4] , \oi[3][3] , \oi[3][2] , 
        \oi[3][1] , SYNOPSYS_UNCONNECTED__5}) );
  DFF \o_reg[1]  ( .D(\oi[3][1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[1]) );
  DFF \o_reg[2]  ( .D(\oi[3][2] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[2]) );
  DFF \o_reg[3]  ( .D(\oi[3][3] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[3]) );
  DFF \o_reg[4]  ( .D(\oi[3][4] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[4]) );
  DFF \o_reg[5]  ( .D(\oi[3][5] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[5]) );
  DFF \o_reg[6]  ( .D(\oi[3][6] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[6]) );
  DFF \o_reg[7]  ( .D(\oi[3][7] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[7]) );
  DFF \o_reg[8]  ( .D(\oi[3][8] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[8]) );
  DFF \o_reg[9]  ( .D(\oi[3][9] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[9]) );
  DFF \o_reg[10]  ( .D(\oi[3][10] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[10])
         );
  DFF \o_reg[11]  ( .D(\oi[3][11] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[11])
         );
  DFF \o_reg[12]  ( .D(\oi[3][12] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[12])
         );
  DFF \o_reg[13]  ( .D(\oi[3][13] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[13])
         );
  DFF \o_reg[14]  ( .D(\oi[3][14] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[14])
         );
  DFF \o_reg[15]  ( .D(\oi[3][15] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[15])
         );
  DFF \o_reg[16]  ( .D(\oi[3][16] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[16])
         );
  DFF \o_reg[17]  ( .D(\oi[3][17] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[17])
         );
  DFF \o_reg[18]  ( .D(\oi[3][18] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[18])
         );
  DFF \o_reg[19]  ( .D(\oi[3][19] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[19])
         );
  DFF \o_reg[20]  ( .D(\oi[3][20] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[20])
         );
  DFF \o_reg[21]  ( .D(\oi[3][21] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[21])
         );
  DFF \o_reg[22]  ( .D(\oi[3][22] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[22])
         );
  DFF \o_reg[23]  ( .D(\oi[3][23] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[23])
         );
  DFF \o_reg[24]  ( .D(\oi[3][24] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[24])
         );
  DFF \o_reg[25]  ( .D(\oi[3][25] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[25])
         );
  DFF \o_reg[26]  ( .D(\oi[3][26] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[26])
         );
  DFF \o_reg[27]  ( .D(\oi[3][27] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[27])
         );
  DFF \o_reg[28]  ( .D(\oi[3][28] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[28])
         );
  DFF \o_reg[29]  ( .D(\oi[3][29] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[29])
         );
  DFF \o_reg[30]  ( .D(\oi[3][30] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[30])
         );
  DFF \o_reg[31]  ( .D(\oi[3][31] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[31])
         );
endmodule

