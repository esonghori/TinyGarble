
module SubBytes ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XNOR U2962 ( .A(n328), .B(n339), .Z(n341) );
  XNOR U2963 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2964 ( .A(n493), .B(n494), .Z(n646) );
  IV U2965 ( .A(x[1]), .Z(n1447) );
  XOR U2966 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2967 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2968 ( .A(n1446), .Z(n3) );
  AND U2969 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2970 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2971 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2972 ( .A(n2), .B(n1), .Z(n66) );
  IV U2973 ( .A(n66), .Z(n12) );
  XNOR U2974 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2975 ( .A(x[7]), .Z(n4) );
  XNOR U2976 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2977 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2978 ( .A(n4), .B(n3), .Z(n11) );
  IV U2979 ( .A(n11), .Z(n1083) );
  XOR U2980 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2981 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2982 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2983 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2984 ( .A(n5), .Z(n790) );
  NANDN U2985 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2986 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2987 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2988 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2989 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2990 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2991 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2992 ( .A(n10), .B(n9), .Z(n46) );
  IV U2993 ( .A(n46), .Z(n52) );
  AND U2994 ( .A(n12), .B(n11), .Z(n17) );
  XOR U2995 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U2996 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U2997 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U2998 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U2999 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3000 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3001 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3002 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3003 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3004 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3005 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3006 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3007 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3008 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3009 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3010 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3011 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3012 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3013 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3014 ( .A(n52), .B(n25), .Z(n36) );
  IV U3015 ( .A(n42), .Z(n43) );
  IV U3016 ( .A(n44), .Z(n50) );
  XOR U3017 ( .A(n26), .B(n800), .Z(n29) );
  AND U3018 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3019 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3020 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3021 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3022 ( .A(n33), .B(n32), .Z(n54) );
  IV U3023 ( .A(n54), .Z(n49) );
  XOR U3024 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3025 ( .A(n43), .B(n34), .Z(n35) );
  AND U3026 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3027 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3028 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3029 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3030 ( .A(n44), .B(n38), .Z(n39) );
  AND U3031 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3032 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3033 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3034 ( .A(n52), .B(n42), .Z(n48) );
  AND U3035 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3036 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3037 ( .A(n46), .B(n45), .Z(n47) );
  AND U3038 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3039 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3040 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3041 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3042 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3043 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3044 ( .A(n806), .B(n791), .Z(n793) );
  OR U3045 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3046 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3047 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3048 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3049 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3050 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3051 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3052 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3053 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3054 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3055 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3056 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3057 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3058 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3059 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3060 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3061 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3062 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3063 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3064 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3065 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3066 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3067 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3068 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3069 ( .A(n70), .Z(n142) );
  NANDN U3070 ( .A(n128), .B(n142), .Z(n80) );
  IV U3071 ( .A(n135), .Z(n91) );
  XNOR U3072 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3073 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3074 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3075 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3076 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3077 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3078 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3079 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3080 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3081 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3082 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3083 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3084 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3085 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3086 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3087 ( .A(n78), .B(n77), .Z(n115) );
  IV U3088 ( .A(n115), .Z(n108) );
  XNOR U3089 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3090 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3091 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3092 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3093 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3094 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3095 ( .A(n81), .B(n171), .Z(n84) );
  AND U3096 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3097 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3098 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3099 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3100 ( .A(n94), .B(n86), .Z(n118) );
  AND U3101 ( .A(n129), .B(n161), .Z(n89) );
  IV U3102 ( .A(x[97]), .Z(n136) );
  XNOR U3103 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3104 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3105 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3106 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3107 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3108 ( .A(n108), .B(n90), .Z(n99) );
  IV U3109 ( .A(n118), .Z(n102) );
  NAND U3110 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3111 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3112 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3113 ( .A(n97), .B(n96), .Z(n114) );
  IV U3114 ( .A(n107), .Z(n116) );
  XOR U3115 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3116 ( .A(n102), .B(n111), .Z(n98) );
  AND U3117 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3118 ( .A(n118), .B(n108), .Z(n104) );
  AND U3119 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3120 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3121 ( .A(n102), .B(n101), .Z(n103) );
  AND U3122 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3123 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3124 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3125 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3126 ( .A(n131), .B(n106), .Z(n173) );
  IV U3127 ( .A(n114), .Z(n120) );
  NAND U3128 ( .A(n120), .B(n107), .Z(n113) );
  AND U3129 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3130 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3131 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3132 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3133 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3134 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3135 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3136 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3137 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3138 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3139 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3140 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3141 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3142 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3143 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3144 ( .B(n163), .A(n126), .Z(n184) );
  IV U3145 ( .A(n127), .Z(n162) );
  OR U3146 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3147 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3148 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3149 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3150 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3151 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3152 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3153 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3154 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3155 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3156 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3157 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3158 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3159 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3160 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3161 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3162 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3163 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3164 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3165 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3166 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3167 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3168 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3169 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3170 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3171 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3172 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3173 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3174 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3175 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3176 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3177 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3178 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3179 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3180 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3181 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3182 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3183 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3184 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3185 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3186 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3187 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3188 ( .A(x[105]), .Z(n292) );
  XOR U3189 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3190 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3191 ( .A(n291), .Z(n188) );
  AND U3192 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3193 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3194 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3195 ( .A(n187), .B(n186), .Z(n251) );
  IV U3196 ( .A(n251), .Z(n197) );
  XNOR U3197 ( .A(n197), .B(n291), .Z(n250) );
  IV U3198 ( .A(x[111]), .Z(n189) );
  XNOR U3199 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3200 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3201 ( .A(n189), .B(n188), .Z(n196) );
  IV U3202 ( .A(n196), .Z(n280) );
  XOR U3203 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3204 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3205 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3206 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3207 ( .A(n190), .Z(n255) );
  NANDN U3208 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3209 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3210 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3211 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3212 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3213 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3214 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3215 ( .A(n195), .B(n194), .Z(n231) );
  IV U3216 ( .A(n231), .Z(n237) );
  AND U3217 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3218 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3219 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3220 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3221 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3222 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3223 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3224 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3225 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3226 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3227 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3228 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3229 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3230 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3231 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3232 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3233 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3234 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3235 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3236 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3237 ( .A(n237), .B(n210), .Z(n221) );
  IV U3238 ( .A(n227), .Z(n228) );
  IV U3239 ( .A(n229), .Z(n235) );
  XOR U3240 ( .A(n211), .B(n265), .Z(n214) );
  AND U3241 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3242 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3243 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3244 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3245 ( .A(n218), .B(n217), .Z(n239) );
  IV U3246 ( .A(n239), .Z(n234) );
  XOR U3247 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3248 ( .A(n228), .B(n219), .Z(n220) );
  AND U3249 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3250 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3251 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3252 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3253 ( .A(n229), .B(n223), .Z(n224) );
  AND U3254 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3255 ( .A(n299), .B(n281), .Z(n256) );
  OR U3256 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3257 ( .A(n237), .B(n227), .Z(n233) );
  AND U3258 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3259 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3260 ( .A(n231), .B(n230), .Z(n232) );
  AND U3261 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3262 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3263 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3264 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3265 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3266 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3267 ( .A(n271), .B(n256), .Z(n258) );
  OR U3268 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3269 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3270 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3271 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3272 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3273 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3274 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3275 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3276 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3277 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3278 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3279 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3280 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3281 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3282 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3283 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3284 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3285 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3286 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3287 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3288 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3289 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3290 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3291 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3292 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3293 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3294 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3295 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3296 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3297 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3298 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3299 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3300 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3301 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3302 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3303 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3304 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3305 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3306 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3307 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3308 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3309 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3310 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3311 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3312 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3313 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3314 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3315 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3316 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3317 ( .A(x[15]), .Z(n311) );
  IV U3318 ( .A(x[10]), .Z(n315) );
  XOR U3319 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3320 ( .A(n315), .B(n307), .Z(n352) );
  IV U3321 ( .A(n352), .Z(n309) );
  XOR U3322 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3323 ( .A(x[9]), .Z(n655) );
  XNOR U3324 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3325 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3326 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3327 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3328 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3329 ( .A(n314), .B(n497), .Z(n318) );
  IV U3330 ( .A(x[13]), .Z(n353) );
  XOR U3331 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3332 ( .A(n353), .B(n310), .Z(n325) );
  IV U3333 ( .A(n325), .Z(n656) );
  XOR U3334 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3335 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3336 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3337 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3338 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3339 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3340 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3341 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3342 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3343 ( .A(n333), .B(n312), .Z(n328) );
  IV U3344 ( .A(n313), .Z(n647) );
  IV U3345 ( .A(n314), .Z(n507) );
  XNOR U3346 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3347 ( .A(n507), .B(n321), .Z(n501) );
  IV U3348 ( .A(n316), .Z(n344) );
  NANDN U3349 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3350 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3351 ( .A(n648), .B(n497), .Z(n498) );
  OR U3352 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3353 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3354 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3355 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3356 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3357 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3358 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3359 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3360 ( .A(n647), .B(n324), .Z(n356) );
  IV U3361 ( .A(n356), .Z(n359) );
  NAND U3362 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3363 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3364 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3365 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3366 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3367 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3368 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3369 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3370 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3371 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3372 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3373 ( .A(n348), .B(n358), .Z(n336) );
  AND U3374 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3375 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3376 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3377 ( .A(n342), .B(n340), .Z(n354) );
  OR U3378 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3379 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3380 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3381 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3382 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3383 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3384 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3385 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3386 ( .A(n347), .B(n346), .Z(n361) );
  OR U3387 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3388 ( .A(n496), .B(n349), .Z(n504) );
  AND U3389 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3390 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3391 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3392 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3393 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3394 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3395 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3396 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3397 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3398 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3399 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3400 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3401 ( .A(n670), .B(n519), .Z(n654) );
  IV U3402 ( .A(n654), .Z(z[10]) );
  XNOR U3403 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3404 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3405 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3406 ( .A(x[113]), .Z(n475) );
  XOR U3407 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3408 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3409 ( .A(n474), .Z(n371) );
  AND U3410 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3411 ( .A(x[115]), .B(n475), .Z(n374) );
  XNOR U3412 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3413 ( .A(n370), .B(n369), .Z(n434) );
  IV U3414 ( .A(n434), .Z(n380) );
  XNOR U3415 ( .A(n380), .B(n474), .Z(n433) );
  IV U3416 ( .A(x[119]), .Z(n372) );
  XNOR U3417 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3418 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3419 ( .A(n372), .B(n371), .Z(n379) );
  IV U3420 ( .A(n379), .Z(n463) );
  XOR U3421 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3422 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3423 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3424 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3425 ( .A(n373), .Z(n438) );
  NANDN U3426 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3427 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3428 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3429 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3430 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3431 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3432 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3433 ( .A(n378), .B(n377), .Z(n414) );
  IV U3434 ( .A(n414), .Z(n420) );
  AND U3435 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3436 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3437 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3438 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3439 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3440 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3441 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3442 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3443 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3444 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3445 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3446 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3447 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3448 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3449 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3450 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3451 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3452 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3453 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3454 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3455 ( .A(n420), .B(n393), .Z(n404) );
  IV U3456 ( .A(n410), .Z(n411) );
  IV U3457 ( .A(n412), .Z(n418) );
  XOR U3458 ( .A(n394), .B(n448), .Z(n397) );
  AND U3459 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3460 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3461 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3462 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3463 ( .A(n401), .B(n400), .Z(n422) );
  IV U3464 ( .A(n422), .Z(n417) );
  XOR U3465 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3466 ( .A(n411), .B(n402), .Z(n403) );
  AND U3467 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3468 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3469 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3470 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3471 ( .A(n412), .B(n406), .Z(n407) );
  AND U3472 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3473 ( .A(n482), .B(n464), .Z(n439) );
  OR U3474 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3475 ( .A(n420), .B(n410), .Z(n416) );
  AND U3476 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3477 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3478 ( .A(n414), .B(n413), .Z(n415) );
  AND U3479 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3480 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3481 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3482 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3483 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3484 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3485 ( .A(n454), .B(n439), .Z(n441) );
  OR U3486 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3487 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3488 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3489 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3490 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3491 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3492 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3493 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3494 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3495 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3496 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3497 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3498 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3499 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3500 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3501 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3502 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3503 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3504 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3505 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3506 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3507 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3508 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3509 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3510 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3511 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3512 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3513 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3514 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3515 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3516 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3517 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3518 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3519 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3520 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3521 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3522 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3523 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3524 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3525 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3526 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3527 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3528 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3529 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3530 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3531 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3532 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3533 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3534 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3535 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3536 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3537 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3538 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3539 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3540 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3541 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3542 ( .A(n506), .B(n672), .Z(n509) );
  OR U3543 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3544 ( .A(n650), .B(n499), .Z(n671) );
  OR U3545 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3546 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3547 ( .A(n511), .B(n503), .Z(n678) );
  AND U3548 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3549 ( .A(n507), .B(n506), .Z(n675) );
  OR U3550 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3551 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3552 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3553 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3554 ( .A(n515), .B(n514), .Z(n660) );
  OR U3555 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3556 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3557 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3558 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3559 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3560 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3561 ( .A(x[121]), .Z(n628) );
  XOR U3562 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3563 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3564 ( .A(n627), .Z(n524) );
  AND U3565 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3566 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3567 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3568 ( .A(n523), .B(n522), .Z(n587) );
  IV U3569 ( .A(n587), .Z(n533) );
  XNOR U3570 ( .A(n533), .B(n627), .Z(n586) );
  IV U3571 ( .A(x[127]), .Z(n525) );
  XNOR U3572 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3573 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3574 ( .A(n525), .B(n524), .Z(n532) );
  IV U3575 ( .A(n532), .Z(n616) );
  XOR U3576 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3577 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3578 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3579 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3580 ( .A(n526), .Z(n591) );
  NANDN U3581 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3582 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3583 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3584 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3585 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3586 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3587 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3588 ( .A(n531), .B(n530), .Z(n567) );
  IV U3589 ( .A(n567), .Z(n573) );
  AND U3590 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3591 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3592 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3593 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3594 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3595 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3596 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3597 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3598 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3599 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3600 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3601 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3602 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3603 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3604 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3605 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3606 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3607 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3608 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3609 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3610 ( .A(n573), .B(n546), .Z(n557) );
  IV U3611 ( .A(n563), .Z(n564) );
  IV U3612 ( .A(n565), .Z(n571) );
  XOR U3613 ( .A(n547), .B(n601), .Z(n550) );
  AND U3614 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3615 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3616 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3617 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3618 ( .A(n554), .B(n553), .Z(n575) );
  IV U3619 ( .A(n575), .Z(n570) );
  XOR U3620 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3621 ( .A(n564), .B(n555), .Z(n556) );
  AND U3622 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3623 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3624 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3625 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3626 ( .A(n565), .B(n559), .Z(n560) );
  AND U3627 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3628 ( .A(n635), .B(n617), .Z(n592) );
  OR U3629 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3630 ( .A(n573), .B(n563), .Z(n569) );
  AND U3631 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3632 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3633 ( .A(n567), .B(n566), .Z(n568) );
  AND U3634 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3635 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3636 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3637 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3638 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3639 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3640 ( .A(n607), .B(n592), .Z(n594) );
  OR U3641 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3642 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3643 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3644 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3645 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3646 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3647 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3648 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3649 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3650 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3651 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3652 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3653 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3654 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3655 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3656 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3657 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3658 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3659 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3660 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3661 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3662 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3663 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3664 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3665 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3666 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3667 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3668 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3669 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3670 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3671 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3672 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3673 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3674 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3675 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3676 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3677 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3678 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3679 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3680 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3681 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3682 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3683 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3684 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3685 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3686 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3687 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3688 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3689 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3690 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3691 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3692 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3693 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3694 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3695 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3696 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3697 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3698 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3699 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3700 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3701 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3702 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3703 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3704 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3705 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3706 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3707 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3708 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3709 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3710 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3711 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3712 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3713 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3714 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3715 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3716 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3717 ( .A(x[17]), .Z(n815) );
  XOR U3718 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XOR U3719 ( .A(x[21]), .B(n685), .Z(n814) );
  IV U3720 ( .A(n814), .Z(n686) );
  AND U3721 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3722 ( .A(x[19]), .B(n815), .Z(n689) );
  XNOR U3723 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3724 ( .A(n685), .B(n684), .Z(n749) );
  IV U3725 ( .A(n749), .Z(n695) );
  XNOR U3726 ( .A(n695), .B(n814), .Z(n748) );
  IV U3727 ( .A(x[23]), .Z(n687) );
  XNOR U3728 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3729 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3730 ( .A(n687), .B(n686), .Z(n694) );
  IV U3731 ( .A(n694), .Z(n778) );
  XOR U3732 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3733 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3734 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3735 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3736 ( .A(n688), .Z(n753) );
  NANDN U3737 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3738 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3739 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3740 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3741 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3742 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3743 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3744 ( .A(n693), .B(n692), .Z(n729) );
  IV U3745 ( .A(n729), .Z(n735) );
  AND U3746 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3747 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3748 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3749 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3750 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3751 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3752 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3753 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3754 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3755 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3756 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3757 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3758 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3759 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3760 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3761 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3762 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3763 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3764 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3765 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3766 ( .A(n735), .B(n708), .Z(n719) );
  IV U3767 ( .A(n725), .Z(n726) );
  IV U3768 ( .A(n727), .Z(n733) );
  XOR U3769 ( .A(n709), .B(n763), .Z(n712) );
  AND U3770 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3771 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3772 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3773 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3774 ( .A(n716), .B(n715), .Z(n737) );
  IV U3775 ( .A(n737), .Z(n732) );
  XOR U3776 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3777 ( .A(n726), .B(n717), .Z(n718) );
  AND U3778 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3779 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3780 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3781 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3782 ( .A(n727), .B(n721), .Z(n722) );
  AND U3783 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3784 ( .A(n822), .B(n779), .Z(n754) );
  OR U3785 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3786 ( .A(n735), .B(n725), .Z(n731) );
  AND U3787 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3788 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3789 ( .A(n729), .B(n728), .Z(n730) );
  AND U3790 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3791 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3792 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3793 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3794 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3795 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3796 ( .A(n769), .B(n754), .Z(n756) );
  OR U3797 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3798 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3799 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3800 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3801 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3802 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3803 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3804 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3805 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3806 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3807 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3808 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3809 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3810 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3811 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3812 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3813 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3814 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3815 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3816 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3817 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3818 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3819 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3820 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3821 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3822 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3823 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3824 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3825 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3826 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3827 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3828 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3829 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3830 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3831 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3832 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3833 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3834 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3835 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3836 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3837 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3838 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3839 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3840 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3841 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3842 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3843 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3844 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3845 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3846 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3847 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3848 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3849 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3850 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3851 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3852 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3853 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3854 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3855 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3856 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3857 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3858 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3859 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3860 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3861 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3862 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3863 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3864 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3865 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3866 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3867 ( .A(x[25]), .Z(n939) );
  XOR U3868 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U3869 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3870 ( .A(n938), .Z(n835) );
  AND U3871 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3872 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3873 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3874 ( .A(n834), .B(n833), .Z(n898) );
  IV U3875 ( .A(n898), .Z(n844) );
  XNOR U3876 ( .A(n844), .B(n938), .Z(n897) );
  IV U3877 ( .A(x[31]), .Z(n836) );
  XNOR U3878 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3879 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3880 ( .A(n836), .B(n835), .Z(n843) );
  IV U3881 ( .A(n843), .Z(n927) );
  XOR U3882 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3883 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3884 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3885 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3886 ( .A(n837), .Z(n902) );
  NANDN U3887 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3888 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3889 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3890 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3891 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3892 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3893 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3894 ( .A(n842), .B(n841), .Z(n878) );
  IV U3895 ( .A(n878), .Z(n884) );
  AND U3896 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3897 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3898 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3899 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3900 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3901 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3902 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3903 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3904 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3905 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3906 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3907 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3908 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3909 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3910 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3911 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3912 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3913 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3914 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3915 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3916 ( .A(n884), .B(n857), .Z(n868) );
  IV U3917 ( .A(n874), .Z(n875) );
  IV U3918 ( .A(n876), .Z(n882) );
  XOR U3919 ( .A(n858), .B(n912), .Z(n861) );
  AND U3920 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3921 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3922 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3923 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3924 ( .A(n865), .B(n864), .Z(n886) );
  IV U3925 ( .A(n886), .Z(n881) );
  XOR U3926 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3927 ( .A(n875), .B(n866), .Z(n867) );
  AND U3928 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3929 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3930 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3931 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3932 ( .A(n876), .B(n870), .Z(n871) );
  AND U3933 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3934 ( .A(n946), .B(n928), .Z(n903) );
  OR U3935 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3936 ( .A(n884), .B(n874), .Z(n880) );
  AND U3937 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3938 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3939 ( .A(n878), .B(n877), .Z(n879) );
  AND U3940 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3941 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3942 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3943 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3944 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3945 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3946 ( .A(n918), .B(n903), .Z(n905) );
  OR U3947 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3948 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3949 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3950 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3951 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3952 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3953 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3954 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3955 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3956 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3957 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3958 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3959 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3960 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3961 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3962 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3963 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3964 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3965 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3966 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3967 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3968 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3969 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3970 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3971 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3972 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3973 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3974 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3975 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3976 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3977 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3978 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3979 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3980 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3981 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3982 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3983 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3984 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3985 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3986 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3987 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3988 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3989 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3990 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3991 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3992 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3993 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3994 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3995 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3996 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3997 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U3998 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U3999 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4000 ( .A(x[33]), .Z(n1065) );
  XOR U4001 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4002 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4003 ( .A(n1064), .Z(n961) );
  AND U4004 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4005 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4006 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4007 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4008 ( .A(n1024), .Z(n970) );
  XNOR U4009 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4010 ( .A(x[39]), .Z(n962) );
  XNOR U4011 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4012 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4013 ( .A(n962), .B(n961), .Z(n969) );
  IV U4014 ( .A(n969), .Z(n1053) );
  XOR U4015 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4016 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4017 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4018 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4019 ( .A(n963), .Z(n1028) );
  NANDN U4020 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4021 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4022 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4023 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4024 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4025 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4026 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4027 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4028 ( .A(n1004), .Z(n1010) );
  AND U4029 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4030 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4031 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4032 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4033 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4034 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4035 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4036 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4037 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4038 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4039 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4040 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4041 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4042 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4043 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4044 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4045 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4046 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4047 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4048 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4049 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4050 ( .A(n1000), .Z(n1001) );
  IV U4051 ( .A(n1002), .Z(n1008) );
  XOR U4052 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4053 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4054 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4055 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4056 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4057 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4058 ( .A(n1012), .Z(n1007) );
  XOR U4059 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4060 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4061 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4062 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4063 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4064 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4065 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4066 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4067 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4068 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4069 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4070 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4071 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4072 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4073 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4074 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4075 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4076 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4077 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4078 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4079 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4080 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4081 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4082 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4083 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4084 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4085 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4086 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4087 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4088 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4089 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4090 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4091 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4092 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4093 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4094 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4095 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4096 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4097 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4098 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4099 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4100 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4101 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4102 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4103 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4104 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4105 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4106 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4107 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4108 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4109 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4110 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4111 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4112 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4113 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4114 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4115 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4116 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4117 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4118 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4119 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4120 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4121 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4122 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4123 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4124 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4125 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4126 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4127 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4128 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4129 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4130 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4131 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4132 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4133 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4134 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4135 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4136 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4137 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4138 ( .A(x[41]), .Z(n1199) );
  XOR U4139 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4140 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4141 ( .A(n1198), .Z(n1095) );
  AND U4142 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4143 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4144 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4145 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4146 ( .A(n1158), .Z(n1104) );
  XNOR U4147 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4148 ( .A(x[47]), .Z(n1096) );
  XNOR U4149 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4150 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4151 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4152 ( .A(n1103), .Z(n1187) );
  XOR U4153 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4154 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4155 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4156 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4157 ( .A(n1097), .Z(n1162) );
  NANDN U4158 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4159 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4160 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4161 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4162 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4163 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4164 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4165 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4166 ( .A(n1138), .Z(n1144) );
  AND U4167 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4168 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4169 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4170 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4171 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4172 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4173 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4174 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4175 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4176 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4177 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4178 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4179 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4180 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4181 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4182 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4183 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4184 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4185 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4186 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4187 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4188 ( .A(n1134), .Z(n1135) );
  IV U4189 ( .A(n1136), .Z(n1142) );
  XOR U4190 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4191 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4192 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4193 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4194 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4195 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4196 ( .A(n1146), .Z(n1141) );
  XOR U4197 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4198 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4199 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4200 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4201 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4202 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4203 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4204 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4205 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4206 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4207 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4208 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4209 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4210 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4211 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4212 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4213 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4214 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4215 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4216 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4217 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4218 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4219 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4220 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4221 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4222 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4223 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4224 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4225 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4226 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4227 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4228 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4229 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4230 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4231 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4232 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4233 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4234 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4235 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4236 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4237 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4238 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4239 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4240 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4241 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4242 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4243 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4244 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4245 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4246 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4247 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4248 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4249 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4250 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4251 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4252 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4253 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4254 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4255 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4256 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4257 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4258 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4259 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4260 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4261 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4262 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4263 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4264 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4265 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4266 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4267 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4268 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4269 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4270 ( .A(x[49]), .Z(n1324) );
  XOR U4271 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4272 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4273 ( .A(n1323), .Z(n1219) );
  AND U4274 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4275 ( .A(x[51]), .B(n1324), .Z(n1222) );
  XNOR U4276 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4277 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4278 ( .A(n1282), .Z(n1228) );
  XNOR U4279 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4280 ( .A(x[55]), .Z(n1220) );
  XNOR U4281 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4282 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4283 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4284 ( .A(n1227), .Z(n1312) );
  XOR U4285 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4286 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4287 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4288 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4289 ( .A(n1221), .Z(n1286) );
  NANDN U4290 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4291 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4292 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4293 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4294 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4295 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4296 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4297 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4298 ( .A(n1262), .Z(n1268) );
  AND U4299 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4300 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4301 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4302 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4303 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4304 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4305 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4306 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4307 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4308 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4309 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4310 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4311 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4312 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4313 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4314 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4315 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4316 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4317 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4318 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4319 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4320 ( .A(n1258), .Z(n1259) );
  IV U4321 ( .A(n1260), .Z(n1266) );
  XOR U4322 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4323 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4324 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4325 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4326 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4327 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4328 ( .A(n1270), .Z(n1265) );
  XOR U4329 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4330 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4331 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4332 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4333 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4334 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4335 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4336 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4337 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4338 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4339 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4340 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4341 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4342 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4343 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4344 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4345 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4346 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4347 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4348 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4349 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4350 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4351 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4352 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4353 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4354 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4355 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4356 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4357 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4358 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4359 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4360 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4361 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4362 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4363 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4364 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4365 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4366 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4367 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4368 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4369 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4370 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4371 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4372 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4373 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4374 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4375 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4376 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4377 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4378 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4379 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4380 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4381 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4382 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4383 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4384 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4385 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4386 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4387 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4388 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4389 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4390 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4391 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4392 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4393 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4394 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4395 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4396 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4397 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4398 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4399 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4400 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4401 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4402 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4403 ( .A(x[57]), .Z(n1462) );
  XOR U4404 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4405 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4406 ( .A(n1461), .Z(n1344) );
  AND U4407 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4408 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4409 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4410 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4411 ( .A(n1407), .Z(n1353) );
  XNOR U4412 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4413 ( .A(x[63]), .Z(n1345) );
  XNOR U4414 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4415 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4416 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4417 ( .A(n1352), .Z(n1436) );
  XOR U4418 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4419 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4420 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4421 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4422 ( .A(n1346), .Z(n1411) );
  NANDN U4423 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4424 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4425 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4426 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4427 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4428 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4429 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4430 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4431 ( .A(n1387), .Z(n1393) );
  AND U4432 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4433 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4434 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4435 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4436 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4437 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4438 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4439 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4440 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4441 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4442 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4443 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4444 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4445 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4446 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4447 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4448 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4449 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4450 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4451 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4452 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4453 ( .A(n1383), .Z(n1384) );
  IV U4454 ( .A(n1385), .Z(n1391) );
  XOR U4455 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4456 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4457 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4458 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4459 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4460 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4461 ( .A(n1395), .Z(n1390) );
  XOR U4462 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4463 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4464 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4465 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4466 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4467 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4468 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4469 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4470 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4471 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4472 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4473 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4474 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4475 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4476 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4477 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4478 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4479 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4480 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4481 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4482 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4483 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4484 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4485 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4486 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4487 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4488 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4489 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4490 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4491 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4492 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4493 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4494 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4495 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4496 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4497 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4498 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4499 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4500 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4501 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4502 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4503 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4504 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4505 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4506 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4507 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4508 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4509 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4510 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4511 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4512 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4513 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4514 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4515 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4516 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4517 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4518 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4519 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4520 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4521 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4522 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4523 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4524 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4525 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4526 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4527 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4528 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4529 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4530 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4531 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4532 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4533 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4534 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4535 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4536 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4537 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4538 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4539 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4540 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4541 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4542 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4543 ( .A(x[65]), .Z(n1586) );
  XOR U4544 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4545 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4546 ( .A(n1585), .Z(n1482) );
  AND U4547 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4548 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4549 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4550 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4551 ( .A(n1545), .Z(n1491) );
  XNOR U4552 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4553 ( .A(x[71]), .Z(n1483) );
  XNOR U4554 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4555 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4556 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4557 ( .A(n1490), .Z(n1574) );
  XOR U4558 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4559 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4560 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4561 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4562 ( .A(n1484), .Z(n1549) );
  NANDN U4563 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4564 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4565 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4566 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4567 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4568 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4569 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4570 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4571 ( .A(n1525), .Z(n1531) );
  AND U4572 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4573 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4574 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4575 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4576 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4577 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4578 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4579 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4580 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4581 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4582 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4583 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4584 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4585 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4586 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4587 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4588 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4589 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4590 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4591 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4592 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4593 ( .A(n1521), .Z(n1522) );
  IV U4594 ( .A(n1523), .Z(n1529) );
  XOR U4595 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4596 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4597 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4598 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4599 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4600 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4601 ( .A(n1533), .Z(n1528) );
  XOR U4602 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4603 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4604 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4605 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4606 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4607 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4608 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4609 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4610 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4611 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4612 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4613 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4614 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4615 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4616 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4617 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4618 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4619 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4620 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4621 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4622 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4623 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4624 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4625 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4626 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4627 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4628 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4629 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4630 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4631 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4632 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4633 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4634 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4635 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4636 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4637 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4638 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4639 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4640 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4641 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4642 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4643 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4644 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4645 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4646 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4647 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4648 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4649 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4650 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4651 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4652 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4653 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4654 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4655 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4656 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4657 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4658 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4659 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4660 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4661 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4662 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4663 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4664 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4665 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4666 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4667 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4668 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4669 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4670 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4671 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4672 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4673 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4674 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4675 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4676 ( .A(x[73]), .Z(n1712) );
  XOR U4677 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4678 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4679 ( .A(n1711), .Z(n1608) );
  AND U4680 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4681 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4682 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4683 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4684 ( .A(n1671), .Z(n1617) );
  XNOR U4685 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4686 ( .A(x[79]), .Z(n1609) );
  XNOR U4687 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4688 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4689 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4690 ( .A(n1616), .Z(n1700) );
  XOR U4691 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4692 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4693 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4694 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4695 ( .A(n1610), .Z(n1675) );
  NANDN U4696 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4697 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4698 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4699 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4700 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4701 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4702 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4703 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4704 ( .A(n1651), .Z(n1657) );
  AND U4705 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4706 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4707 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4708 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4709 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4710 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4711 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4712 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4713 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4714 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4715 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4716 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4717 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4718 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4719 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4720 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4721 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4722 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4723 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4724 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4725 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4726 ( .A(n1647), .Z(n1648) );
  IV U4727 ( .A(n1649), .Z(n1655) );
  XOR U4728 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4729 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4730 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4731 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4732 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4733 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4734 ( .A(n1659), .Z(n1654) );
  XOR U4735 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4736 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4737 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4738 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4739 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4740 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4741 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4742 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4743 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4744 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4745 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4746 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4747 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4748 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4749 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4750 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4751 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4752 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4753 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4754 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4755 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4756 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4757 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4758 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4759 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4760 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4761 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4762 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4763 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4764 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4765 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4766 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4767 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4768 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4769 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4770 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4771 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4772 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4773 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4774 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4775 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4776 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4777 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4778 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4779 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4780 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4781 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4782 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4783 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4784 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4785 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4786 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4787 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4788 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4789 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4790 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4791 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4792 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4793 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4794 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4795 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4796 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4797 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4798 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4799 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4800 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4801 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4802 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4803 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4804 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4805 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4806 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4807 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4808 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4809 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4810 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4811 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4812 ( .A(n1838), .Z(n1735) );
  IV U4813 ( .A(x[81]), .Z(n1837) );
  NAND U4814 ( .A(n1735), .B(n1837), .Z(n1742) );
  XOR U4815 ( .A(x[83]), .B(x[81]), .Z(n1738) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module aes_seq_CC10 ( clk, rst, msg, key, out );
  input [127:0] msg;
  input [127:0] key;
  output [127:0] out;
  input clk, rst;
  wire   init, \w0[0][127] , \w0[0][126] , \w0[0][125] , \w0[0][124] ,
         \w0[0][123] , \w0[0][122] , \w0[0][121] , \w0[0][120] , \w0[0][119] ,
         \w0[0][118] , \w0[0][117] , \w0[0][116] , \w0[0][115] , \w0[0][114] ,
         \w0[0][113] , \w0[0][112] , \w0[0][111] , \w0[0][110] , \w0[0][109] ,
         \w0[0][108] , \w0[0][107] , \w0[0][106] , \w0[0][105] , \w0[0][104] ,
         \w0[0][103] , \w0[0][102] , \w0[0][101] , \w0[0][100] , \w0[0][99] ,
         \w0[0][98] , \w0[0][97] , \w0[0][96] , \w0[0][95] , \w0[0][94] ,
         \w0[0][93] , \w0[0][92] , \w0[0][91] , \w0[0][90] , \w0[0][89] ,
         \w0[0][88] , \w0[0][87] , \w0[0][86] , \w0[0][85] , \w0[0][84] ,
         \w0[0][83] , \w0[0][82] , \w0[0][81] , \w0[0][80] , \w0[0][79] ,
         \w0[0][78] , \w0[0][77] , \w0[0][76] , \w0[0][75] , \w0[0][74] ,
         \w0[0][73] , \w0[0][72] , \w0[0][71] , \w0[0][70] , \w0[0][69] ,
         \w0[0][68] , \w0[0][67] , \w0[0][66] , \w0[0][65] , \w0[0][64] ,
         \w0[0][63] , \w0[0][62] , \w0[0][61] , \w0[0][60] , \w0[0][59] ,
         \w0[0][58] , \w0[0][57] , \w0[0][56] , \w0[0][55] , \w0[0][54] ,
         \w0[0][53] , \w0[0][52] , \w0[0][51] , \w0[0][50] , \w0[0][49] ,
         \w0[0][48] , \w0[0][47] , \w0[0][46] , \w0[0][45] , \w0[0][44] ,
         \w0[0][43] , \w0[0][42] , \w0[0][41] , \w0[0][40] , \w0[0][39] ,
         \w0[0][38] , \w0[0][37] , \w0[0][36] , \w0[0][35] , \w0[0][34] ,
         \w0[0][33] , \w0[0][32] , \w0[0][31] , \w0[0][30] , \w0[0][29] ,
         \w0[0][28] , \w0[0][27] , \w0[0][26] , \w0[0][25] , \w0[0][24] ,
         \w0[0][23] , \w0[0][22] , \w0[0][21] , \w0[0][20] , \w0[0][19] ,
         \w0[0][18] , \w0[0][17] , \w0[0][16] , \w0[0][15] , \w0[0][14] ,
         \w0[0][13] , \w0[0][12] , \w0[0][11] , \w0[0][10] , \w0[0][9] ,
         \w0[0][8] , \w0[0][7] , \w0[0][6] , \w0[0][5] , \w0[0][4] ,
         \w0[0][3] , \w0[0][2] , \w0[0][1] , \w0[0][0] , \w1[0][127] ,
         \w1[0][126] , \w1[0][125] , \w1[0][124] , \w1[0][123] , \w1[0][122] ,
         \w1[0][121] , \w1[0][120] , \w1[0][119] , \w1[0][118] , \w1[0][117] ,
         \w1[0][116] , \w1[0][115] , \w1[0][114] , \w1[0][113] , \w1[0][112] ,
         \w1[0][111] , \w1[0][110] , \w1[0][109] , \w1[0][108] , \w1[0][107] ,
         \w1[0][106] , \w1[0][105] , \w1[0][104] , \w1[0][103] , \w1[0][102] ,
         \w1[0][101] , \w1[0][100] , \w1[0][99] , \w1[0][98] , \w1[0][97] ,
         \w1[0][96] , \w1[0][95] , \w1[0][94] , \w1[0][93] , \w1[0][92] ,
         \w1[0][91] , \w1[0][90] , \w1[0][89] , \w1[0][88] , \w1[0][87] ,
         \w1[0][86] , \w1[0][85] , \w1[0][84] , \w1[0][83] , \w1[0][82] ,
         \w1[0][81] , \w1[0][80] , \w1[0][79] , \w1[0][78] , \w1[0][77] ,
         \w1[0][76] , \w1[0][75] , \w1[0][74] , \w1[0][73] , \w1[0][72] ,
         \w1[0][71] , \w1[0][70] , \w1[0][69] , \w1[0][68] , \w1[0][67] ,
         \w1[0][66] , \w1[0][65] , \w1[0][64] , \w1[0][63] , \w1[0][62] ,
         \w1[0][61] , \w1[0][60] , \w1[0][59] , \w1[0][58] , \w1[0][57] ,
         \w1[0][56] , \w1[0][55] , \w1[0][54] , \w1[0][53] , \w1[0][52] ,
         \w1[0][51] , \w1[0][50] , \w1[0][49] , \w1[0][48] , \w1[0][47] ,
         \w1[0][46] , \w1[0][45] , \w1[0][44] , \w1[0][43] , \w1[0][42] ,
         \w1[0][41] , \w1[0][40] , \w1[0][39] , \w1[0][38] , \w1[0][37] ,
         \w1[0][36] , \w1[0][35] , \w1[0][34] , \w1[0][33] , \w1[0][32] ,
         \w1[0][31] , \w1[0][30] , \w1[0][29] , \w1[0][28] , \w1[0][27] ,
         \w1[0][26] , \w1[0][25] , \w1[0][24] , \w1[0][23] , \w1[0][22] ,
         \w1[0][21] , \w1[0][20] , \w1[0][19] , \w1[0][18] , \w1[0][17] ,
         \w1[0][16] , \w1[0][15] , \w1[0][14] , \w1[0][13] , \w1[0][12] ,
         \w1[0][11] , \w1[0][10] , \w1[0][9] , \w1[0][8] , \w1[0][7] ,
         \w1[0][6] , \w1[0][5] , \w1[0][4] , \w1[0][3] , \w1[0][2] ,
         \w1[0][1] , \w1[0][0] , \w3[0][127] , \w3[0][126] , \w3[0][125] ,
         \w3[0][124] , \w3[0][123] , \w3[0][122] , \w3[0][121] , \w3[0][120] ,
         \w3[0][119] , \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] ,
         \w3[0][114] , \w3[0][113] , \w3[0][112] , \w3[0][111] , \w3[0][110] ,
         \w3[0][109] , \w3[0][108] , \w3[0][107] , \w3[0][106] , \w3[0][105] ,
         \w3[0][104] , \w3[0][103] , \w3[0][102] , \w3[0][101] , \w3[0][100] ,
         \w3[0][99] , \w3[0][98] , \w3[0][97] , \w3[0][96] , \w3[0][95] ,
         \w3[0][94] , \w3[0][93] , \w3[0][92] , \w3[0][91] , \w3[0][90] ,
         \w3[0][89] , \w3[0][88] , \w3[0][87] , \w3[0][86] , \w3[0][85] ,
         \w3[0][84] , \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] ,
         \w3[0][79] , \w3[0][78] , \w3[0][77] , \w3[0][76] , \w3[0][75] ,
         \w3[0][74] , \w3[0][73] , \w3[0][72] , \w3[0][71] , \w3[0][70] ,
         \w3[0][69] , \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] ,
         \w3[0][64] , \w3[0][63] , \w3[0][62] , \w3[0][61] , \w3[0][60] ,
         \w3[0][59] , \w3[0][58] , \w3[0][57] , \w3[0][56] , \w3[0][55] ,
         \w3[0][54] , \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] ,
         \w3[0][49] , \w3[0][48] , \w3[0][47] , \w3[0][46] , \w3[0][45] ,
         \w3[0][44] , \w3[0][43] , \w3[0][42] , \w3[0][41] , \w3[0][40] ,
         \w3[0][39] , \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] ,
         \w3[0][34] , \w3[0][33] , \w3[0][32] , \w3[0][31] , \w3[0][30] ,
         \w3[0][29] , \w3[0][28] , \w3[0][27] , \w3[0][26] , \w3[0][25] ,
         \w3[0][24] , \w3[0][23] , \w3[0][22] , \w3[0][21] , \w3[0][20] ,
         \w3[0][19] , \w3[0][18] , \w3[0][17] , \w3[0][16] , \w3[0][15] ,
         \w3[0][14] , \w3[0][13] , \w3[0][12] , \w3[0][11] , \w3[0][10] ,
         \w3[0][9] , \w3[0][8] , \w3[0][7] , \w3[0][6] , \w3[0][5] ,
         \w3[0][4] , \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514;
  wire   [127:0] state;

  SubBytes \SUBBYTES[0].a  ( .x({\w1[0][127] , \w1[0][126] , \w1[0][125] , 
        \w1[0][124] , \w1[0][123] , \w1[0][122] , \w1[0][121] , \w1[0][120] , 
        \w1[0][119] , \w1[0][118] , \w1[0][117] , \w1[0][116] , \w1[0][115] , 
        \w1[0][114] , \w1[0][113] , \w1[0][112] , \w1[0][111] , \w1[0][110] , 
        \w1[0][109] , \w1[0][108] , \w1[0][107] , \w1[0][106] , \w1[0][105] , 
        \w1[0][104] , \w1[0][103] , \w1[0][102] , \w1[0][101] , \w1[0][100] , 
        \w1[0][99] , \w1[0][98] , \w1[0][97] , \w1[0][96] , \w1[0][95] , 
        \w1[0][94] , \w1[0][93] , \w1[0][92] , \w1[0][91] , \w1[0][90] , 
        \w1[0][89] , \w1[0][88] , \w1[0][87] , \w1[0][86] , \w1[0][85] , 
        \w1[0][84] , \w1[0][83] , \w1[0][82] , \w1[0][81] , \w1[0][80] , 
        \w1[0][79] , \w1[0][78] , \w1[0][77] , \w1[0][76] , \w1[0][75] , 
        \w1[0][74] , \w1[0][73] , \w1[0][72] , \w1[0][71] , \w1[0][70] , 
        \w1[0][69] , \w1[0][68] , \w1[0][67] , \w1[0][66] , \w1[0][65] , 
        \w1[0][64] , \w1[0][63] , \w1[0][62] , \w1[0][61] , \w1[0][60] , 
        \w1[0][59] , \w1[0][58] , \w1[0][57] , \w1[0][56] , \w1[0][55] , 
        \w1[0][54] , \w1[0][53] , \w1[0][52] , \w1[0][51] , \w1[0][50] , 
        \w1[0][49] , \w1[0][48] , \w1[0][47] , \w1[0][46] , \w1[0][45] , 
        \w1[0][44] , \w1[0][43] , \w1[0][42] , \w1[0][41] , \w1[0][40] , 
        \w1[0][39] , \w1[0][38] , \w1[0][37] , \w1[0][36] , \w1[0][35] , 
        \w1[0][34] , \w1[0][33] , \w1[0][32] , \w1[0][31] , \w1[0][30] , 
        \w1[0][29] , \w1[0][28] , \w1[0][27] , \w1[0][26] , \w1[0][25] , 
        \w1[0][24] , \w1[0][23] , \w1[0][22] , \w1[0][21] , \w1[0][20] , 
        \w1[0][19] , \w1[0][18] , \w1[0][17] , \w1[0][16] , \w1[0][15] , 
        \w1[0][14] , \w1[0][13] , \w1[0][12] , \w1[0][11] , \w1[0][10] , 
        \w1[0][9] , \w1[0][8] , \w1[0][7] , \w1[0][6] , \w1[0][5] , \w1[0][4] , 
        \w1[0][3] , \w1[0][2] , \w1[0][1] , \w1[0][0] }), .z({\w3[0][127] , 
        \w3[0][126] , \w3[0][125] , \w3[0][124] , \w3[0][123] , \w3[0][122] , 
        \w3[0][121] , \w3[0][120] , \w3[0][23] , \w3[0][22] , \w3[0][21] , 
        \w3[0][20] , \w3[0][19] , \w3[0][18] , \w3[0][17] , \w3[0][16] , 
        \w3[0][47] , \w3[0][46] , \w3[0][45] , \w3[0][44] , \w3[0][43] , 
        \w3[0][42] , \w3[0][41] , \w3[0][40] , \w3[0][71] , \w3[0][70] , 
        \w3[0][69] , \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] , 
        \w3[0][64] , \w3[0][95] , \w3[0][94] , \w3[0][93] , \w3[0][92] , 
        \w3[0][91] , \w3[0][90] , \w3[0][89] , \w3[0][88] , \w3[0][119] , 
        \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] , \w3[0][114] , 
        \w3[0][113] , \w3[0][112] , \w3[0][15] , \w3[0][14] , \w3[0][13] , 
        \w3[0][12] , \w3[0][11] , \w3[0][10] , \w3[0][9] , \w3[0][8] , 
        \w3[0][39] , \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] , 
        \w3[0][34] , \w3[0][33] , \w3[0][32] , \w3[0][63] , \w3[0][62] , 
        \w3[0][61] , \w3[0][60] , \w3[0][59] , \w3[0][58] , \w3[0][57] , 
        \w3[0][56] , \w3[0][87] , \w3[0][86] , \w3[0][85] , \w3[0][84] , 
        \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] , \w3[0][111] , 
        \w3[0][110] , \w3[0][109] , \w3[0][108] , \w3[0][107] , \w3[0][106] , 
        \w3[0][105] , \w3[0][104] , \w3[0][7] , \w3[0][6] , \w3[0][5] , 
        \w3[0][4] , \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , 
        \w3[0][31] , \w3[0][30] , \w3[0][29] , \w3[0][28] , \w3[0][27] , 
        \w3[0][26] , \w3[0][25] , \w3[0][24] , \w3[0][55] , \w3[0][54] , 
        \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] , \w3[0][49] , 
        \w3[0][48] , \w3[0][79] , \w3[0][78] , \w3[0][77] , \w3[0][76] , 
        \w3[0][75] , \w3[0][74] , \w3[0][73] , \w3[0][72] , \w3[0][103] , 
        \w3[0][102] , \w3[0][101] , \w3[0][100] , \w3[0][99] , \w3[0][98] , 
        \w3[0][97] , \w3[0][96] }) );
  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \state_reg[127]  ( .D(\w0[0][127] ), .CLK(clk), .RST(rst), .Q(state[127]) );
  DFF \state_reg[126]  ( .D(\w0[0][126] ), .CLK(clk), .RST(rst), .Q(state[126]) );
  DFF \state_reg[125]  ( .D(\w0[0][125] ), .CLK(clk), .RST(rst), .Q(state[125]) );
  DFF \state_reg[124]  ( .D(\w0[0][124] ), .CLK(clk), .RST(rst), .Q(state[124]) );
  DFF \state_reg[123]  ( .D(\w0[0][123] ), .CLK(clk), .RST(rst), .Q(state[123]) );
  DFF \state_reg[122]  ( .D(\w0[0][122] ), .CLK(clk), .RST(rst), .Q(state[122]) );
  DFF \state_reg[121]  ( .D(\w0[0][121] ), .CLK(clk), .RST(rst), .Q(state[121]) );
  DFF \state_reg[120]  ( .D(\w0[0][120] ), .CLK(clk), .RST(rst), .Q(state[120]) );
  DFF \state_reg[119]  ( .D(\w0[0][119] ), .CLK(clk), .RST(rst), .Q(state[119]) );
  DFF \state_reg[118]  ( .D(\w0[0][118] ), .CLK(clk), .RST(rst), .Q(state[118]) );
  DFF \state_reg[117]  ( .D(\w0[0][117] ), .CLK(clk), .RST(rst), .Q(state[117]) );
  DFF \state_reg[116]  ( .D(\w0[0][116] ), .CLK(clk), .RST(rst), .Q(state[116]) );
  DFF \state_reg[115]  ( .D(\w0[0][115] ), .CLK(clk), .RST(rst), .Q(state[115]) );
  DFF \state_reg[114]  ( .D(\w0[0][114] ), .CLK(clk), .RST(rst), .Q(state[114]) );
  DFF \state_reg[113]  ( .D(\w0[0][113] ), .CLK(clk), .RST(rst), .Q(state[113]) );
  DFF \state_reg[112]  ( .D(\w0[0][112] ), .CLK(clk), .RST(rst), .Q(state[112]) );
  DFF \state_reg[111]  ( .D(\w0[0][111] ), .CLK(clk), .RST(rst), .Q(state[111]) );
  DFF \state_reg[110]  ( .D(\w0[0][110] ), .CLK(clk), .RST(rst), .Q(state[110]) );
  DFF \state_reg[109]  ( .D(\w0[0][109] ), .CLK(clk), .RST(rst), .Q(state[109]) );
  DFF \state_reg[108]  ( .D(\w0[0][108] ), .CLK(clk), .RST(rst), .Q(state[108]) );
  DFF \state_reg[107]  ( .D(\w0[0][107] ), .CLK(clk), .RST(rst), .Q(state[107]) );
  DFF \state_reg[106]  ( .D(\w0[0][106] ), .CLK(clk), .RST(rst), .Q(state[106]) );
  DFF \state_reg[105]  ( .D(\w0[0][105] ), .CLK(clk), .RST(rst), .Q(state[105]) );
  DFF \state_reg[104]  ( .D(\w0[0][104] ), .CLK(clk), .RST(rst), .Q(state[104]) );
  DFF \state_reg[103]  ( .D(\w0[0][103] ), .CLK(clk), .RST(rst), .Q(state[103]) );
  DFF \state_reg[102]  ( .D(\w0[0][102] ), .CLK(clk), .RST(rst), .Q(state[102]) );
  DFF \state_reg[101]  ( .D(\w0[0][101] ), .CLK(clk), .RST(rst), .Q(state[101]) );
  DFF \state_reg[100]  ( .D(\w0[0][100] ), .CLK(clk), .RST(rst), .Q(state[100]) );
  DFF \state_reg[99]  ( .D(\w0[0][99] ), .CLK(clk), .RST(rst), .Q(state[99])
         );
  DFF \state_reg[98]  ( .D(\w0[0][98] ), .CLK(clk), .RST(rst), .Q(state[98])
         );
  DFF \state_reg[97]  ( .D(\w0[0][97] ), .CLK(clk), .RST(rst), .Q(state[97])
         );
  DFF \state_reg[96]  ( .D(\w0[0][96] ), .CLK(clk), .RST(rst), .Q(state[96])
         );
  DFF \state_reg[95]  ( .D(\w0[0][95] ), .CLK(clk), .RST(rst), .Q(state[95])
         );
  DFF \state_reg[94]  ( .D(\w0[0][94] ), .CLK(clk), .RST(rst), .Q(state[94])
         );
  DFF \state_reg[93]  ( .D(\w0[0][93] ), .CLK(clk), .RST(rst), .Q(state[93])
         );
  DFF \state_reg[92]  ( .D(\w0[0][92] ), .CLK(clk), .RST(rst), .Q(state[92])
         );
  DFF \state_reg[91]  ( .D(\w0[0][91] ), .CLK(clk), .RST(rst), .Q(state[91])
         );
  DFF \state_reg[90]  ( .D(\w0[0][90] ), .CLK(clk), .RST(rst), .Q(state[90])
         );
  DFF \state_reg[89]  ( .D(\w0[0][89] ), .CLK(clk), .RST(rst), .Q(state[89])
         );
  DFF \state_reg[88]  ( .D(\w0[0][88] ), .CLK(clk), .RST(rst), .Q(state[88])
         );
  DFF \state_reg[87]  ( .D(\w0[0][87] ), .CLK(clk), .RST(rst), .Q(state[87])
         );
  DFF \state_reg[86]  ( .D(\w0[0][86] ), .CLK(clk), .RST(rst), .Q(state[86])
         );
  DFF \state_reg[85]  ( .D(\w0[0][85] ), .CLK(clk), .RST(rst), .Q(state[85])
         );
  DFF \state_reg[84]  ( .D(\w0[0][84] ), .CLK(clk), .RST(rst), .Q(state[84])
         );
  DFF \state_reg[83]  ( .D(\w0[0][83] ), .CLK(clk), .RST(rst), .Q(state[83])
         );
  DFF \state_reg[82]  ( .D(\w0[0][82] ), .CLK(clk), .RST(rst), .Q(state[82])
         );
  DFF \state_reg[81]  ( .D(\w0[0][81] ), .CLK(clk), .RST(rst), .Q(state[81])
         );
  DFF \state_reg[80]  ( .D(\w0[0][80] ), .CLK(clk), .RST(rst), .Q(state[80])
         );
  DFF \state_reg[79]  ( .D(\w0[0][79] ), .CLK(clk), .RST(rst), .Q(state[79])
         );
  DFF \state_reg[78]  ( .D(\w0[0][78] ), .CLK(clk), .RST(rst), .Q(state[78])
         );
  DFF \state_reg[77]  ( .D(\w0[0][77] ), .CLK(clk), .RST(rst), .Q(state[77])
         );
  DFF \state_reg[76]  ( .D(\w0[0][76] ), .CLK(clk), .RST(rst), .Q(state[76])
         );
  DFF \state_reg[75]  ( .D(\w0[0][75] ), .CLK(clk), .RST(rst), .Q(state[75])
         );
  DFF \state_reg[74]  ( .D(\w0[0][74] ), .CLK(clk), .RST(rst), .Q(state[74])
         );
  DFF \state_reg[73]  ( .D(\w0[0][73] ), .CLK(clk), .RST(rst), .Q(state[73])
         );
  DFF \state_reg[72]  ( .D(\w0[0][72] ), .CLK(clk), .RST(rst), .Q(state[72])
         );
  DFF \state_reg[71]  ( .D(\w0[0][71] ), .CLK(clk), .RST(rst), .Q(state[71])
         );
  DFF \state_reg[70]  ( .D(\w0[0][70] ), .CLK(clk), .RST(rst), .Q(state[70])
         );
  DFF \state_reg[69]  ( .D(\w0[0][69] ), .CLK(clk), .RST(rst), .Q(state[69])
         );
  DFF \state_reg[68]  ( .D(\w0[0][68] ), .CLK(clk), .RST(rst), .Q(state[68])
         );
  DFF \state_reg[67]  ( .D(\w0[0][67] ), .CLK(clk), .RST(rst), .Q(state[67])
         );
  DFF \state_reg[66]  ( .D(\w0[0][66] ), .CLK(clk), .RST(rst), .Q(state[66])
         );
  DFF \state_reg[65]  ( .D(\w0[0][65] ), .CLK(clk), .RST(rst), .Q(state[65])
         );
  DFF \state_reg[64]  ( .D(\w0[0][64] ), .CLK(clk), .RST(rst), .Q(state[64])
         );
  DFF \state_reg[63]  ( .D(\w0[0][63] ), .CLK(clk), .RST(rst), .Q(state[63])
         );
  DFF \state_reg[62]  ( .D(\w0[0][62] ), .CLK(clk), .RST(rst), .Q(state[62])
         );
  DFF \state_reg[61]  ( .D(\w0[0][61] ), .CLK(clk), .RST(rst), .Q(state[61])
         );
  DFF \state_reg[60]  ( .D(\w0[0][60] ), .CLK(clk), .RST(rst), .Q(state[60])
         );
  DFF \state_reg[59]  ( .D(\w0[0][59] ), .CLK(clk), .RST(rst), .Q(state[59])
         );
  DFF \state_reg[58]  ( .D(\w0[0][58] ), .CLK(clk), .RST(rst), .Q(state[58])
         );
  DFF \state_reg[57]  ( .D(\w0[0][57] ), .CLK(clk), .RST(rst), .Q(state[57])
         );
  DFF \state_reg[56]  ( .D(\w0[0][56] ), .CLK(clk), .RST(rst), .Q(state[56])
         );
  DFF \state_reg[55]  ( .D(\w0[0][55] ), .CLK(clk), .RST(rst), .Q(state[55])
         );
  DFF \state_reg[54]  ( .D(\w0[0][54] ), .CLK(clk), .RST(rst), .Q(state[54])
         );
  DFF \state_reg[53]  ( .D(\w0[0][53] ), .CLK(clk), .RST(rst), .Q(state[53])
         );
  DFF \state_reg[52]  ( .D(\w0[0][52] ), .CLK(clk), .RST(rst), .Q(state[52])
         );
  DFF \state_reg[51]  ( .D(\w0[0][51] ), .CLK(clk), .RST(rst), .Q(state[51])
         );
  DFF \state_reg[50]  ( .D(\w0[0][50] ), .CLK(clk), .RST(rst), .Q(state[50])
         );
  DFF \state_reg[49]  ( .D(\w0[0][49] ), .CLK(clk), .RST(rst), .Q(state[49])
         );
  DFF \state_reg[48]  ( .D(\w0[0][48] ), .CLK(clk), .RST(rst), .Q(state[48])
         );
  DFF \state_reg[47]  ( .D(\w0[0][47] ), .CLK(clk), .RST(rst), .Q(state[47])
         );
  DFF \state_reg[46]  ( .D(\w0[0][46] ), .CLK(clk), .RST(rst), .Q(state[46])
         );
  DFF \state_reg[45]  ( .D(\w0[0][45] ), .CLK(clk), .RST(rst), .Q(state[45])
         );
  DFF \state_reg[44]  ( .D(\w0[0][44] ), .CLK(clk), .RST(rst), .Q(state[44])
         );
  DFF \state_reg[43]  ( .D(\w0[0][43] ), .CLK(clk), .RST(rst), .Q(state[43])
         );
  DFF \state_reg[42]  ( .D(\w0[0][42] ), .CLK(clk), .RST(rst), .Q(state[42])
         );
  DFF \state_reg[41]  ( .D(\w0[0][41] ), .CLK(clk), .RST(rst), .Q(state[41])
         );
  DFF \state_reg[40]  ( .D(\w0[0][40] ), .CLK(clk), .RST(rst), .Q(state[40])
         );
  DFF \state_reg[39]  ( .D(\w0[0][39] ), .CLK(clk), .RST(rst), .Q(state[39])
         );
  DFF \state_reg[38]  ( .D(\w0[0][38] ), .CLK(clk), .RST(rst), .Q(state[38])
         );
  DFF \state_reg[37]  ( .D(\w0[0][37] ), .CLK(clk), .RST(rst), .Q(state[37])
         );
  DFF \state_reg[36]  ( .D(\w0[0][36] ), .CLK(clk), .RST(rst), .Q(state[36])
         );
  DFF \state_reg[35]  ( .D(\w0[0][35] ), .CLK(clk), .RST(rst), .Q(state[35])
         );
  DFF \state_reg[34]  ( .D(\w0[0][34] ), .CLK(clk), .RST(rst), .Q(state[34])
         );
  DFF \state_reg[33]  ( .D(\w0[0][33] ), .CLK(clk), .RST(rst), .Q(state[33])
         );
  DFF \state_reg[32]  ( .D(\w0[0][32] ), .CLK(clk), .RST(rst), .Q(state[32])
         );
  DFF \state_reg[31]  ( .D(\w0[0][31] ), .CLK(clk), .RST(rst), .Q(state[31])
         );
  DFF \state_reg[30]  ( .D(\w0[0][30] ), .CLK(clk), .RST(rst), .Q(state[30])
         );
  DFF \state_reg[29]  ( .D(\w0[0][29] ), .CLK(clk), .RST(rst), .Q(state[29])
         );
  DFF \state_reg[28]  ( .D(\w0[0][28] ), .CLK(clk), .RST(rst), .Q(state[28])
         );
  DFF \state_reg[27]  ( .D(\w0[0][27] ), .CLK(clk), .RST(rst), .Q(state[27])
         );
  DFF \state_reg[26]  ( .D(\w0[0][26] ), .CLK(clk), .RST(rst), .Q(state[26])
         );
  DFF \state_reg[25]  ( .D(\w0[0][25] ), .CLK(clk), .RST(rst), .Q(state[25])
         );
  DFF \state_reg[24]  ( .D(\w0[0][24] ), .CLK(clk), .RST(rst), .Q(state[24])
         );
  DFF \state_reg[23]  ( .D(\w0[0][23] ), .CLK(clk), .RST(rst), .Q(state[23])
         );
  DFF \state_reg[22]  ( .D(\w0[0][22] ), .CLK(clk), .RST(rst), .Q(state[22])
         );
  DFF \state_reg[21]  ( .D(\w0[0][21] ), .CLK(clk), .RST(rst), .Q(state[21])
         );
  DFF \state_reg[20]  ( .D(\w0[0][20] ), .CLK(clk), .RST(rst), .Q(state[20])
         );
  DFF \state_reg[19]  ( .D(\w0[0][19] ), .CLK(clk), .RST(rst), .Q(state[19])
         );
  DFF \state_reg[18]  ( .D(\w0[0][18] ), .CLK(clk), .RST(rst), .Q(state[18])
         );
  DFF \state_reg[17]  ( .D(\w0[0][17] ), .CLK(clk), .RST(rst), .Q(state[17])
         );
  DFF \state_reg[16]  ( .D(\w0[0][16] ), .CLK(clk), .RST(rst), .Q(state[16])
         );
  DFF \state_reg[15]  ( .D(\w0[0][15] ), .CLK(clk), .RST(rst), .Q(state[15])
         );
  DFF \state_reg[14]  ( .D(\w0[0][14] ), .CLK(clk), .RST(rst), .Q(state[14])
         );
  DFF \state_reg[13]  ( .D(\w0[0][13] ), .CLK(clk), .RST(rst), .Q(state[13])
         );
  DFF \state_reg[12]  ( .D(\w0[0][12] ), .CLK(clk), .RST(rst), .Q(state[12])
         );
  DFF \state_reg[11]  ( .D(\w0[0][11] ), .CLK(clk), .RST(rst), .Q(state[11])
         );
  DFF \state_reg[10]  ( .D(\w0[0][10] ), .CLK(clk), .RST(rst), .Q(state[10])
         );
  DFF \state_reg[9]  ( .D(\w0[0][9] ), .CLK(clk), .RST(rst), .Q(state[9]) );
  DFF \state_reg[8]  ( .D(\w0[0][8] ), .CLK(clk), .RST(rst), .Q(state[8]) );
  DFF \state_reg[7]  ( .D(\w0[0][7] ), .CLK(clk), .RST(rst), .Q(state[7]) );
  DFF \state_reg[6]  ( .D(\w0[0][6] ), .CLK(clk), .RST(rst), .Q(state[6]) );
  DFF \state_reg[5]  ( .D(\w0[0][5] ), .CLK(clk), .RST(rst), .Q(state[5]) );
  DFF \state_reg[4]  ( .D(\w0[0][4] ), .CLK(clk), .RST(rst), .Q(state[4]) );
  DFF \state_reg[3]  ( .D(\w0[0][3] ), .CLK(clk), .RST(rst), .Q(state[3]) );
  DFF \state_reg[2]  ( .D(\w0[0][2] ), .CLK(clk), .RST(rst), .Q(state[2]) );
  DFF \state_reg[1]  ( .D(\w0[0][1] ), .CLK(clk), .RST(rst), .Q(state[1]) );
  DFF \state_reg[0]  ( .D(\w0[0][0] ), .CLK(clk), .RST(rst), .Q(state[0]) );
  IV U644 ( .A(init), .Z(n258) );
  XOR U645 ( .A(key[0]), .B(\w3[0][0] ), .Z(out[0]) );
  XOR U646 ( .A(key[100]), .B(\w3[0][100] ), .Z(out[100]) );
  XOR U647 ( .A(key[101]), .B(\w3[0][101] ), .Z(out[101]) );
  XOR U648 ( .A(key[102]), .B(\w3[0][102] ), .Z(out[102]) );
  XOR U649 ( .A(key[103]), .B(\w3[0][103] ), .Z(out[103]) );
  XOR U650 ( .A(key[104]), .B(\w3[0][104] ), .Z(out[104]) );
  XOR U651 ( .A(key[105]), .B(\w3[0][105] ), .Z(out[105]) );
  XOR U652 ( .A(key[106]), .B(\w3[0][106] ), .Z(out[106]) );
  XOR U653 ( .A(key[107]), .B(\w3[0][107] ), .Z(out[107]) );
  XOR U654 ( .A(key[108]), .B(\w3[0][108] ), .Z(out[108]) );
  XOR U655 ( .A(key[109]), .B(\w3[0][109] ), .Z(out[109]) );
  XOR U656 ( .A(key[10]), .B(\w3[0][10] ), .Z(out[10]) );
  XOR U657 ( .A(key[110]), .B(\w3[0][110] ), .Z(out[110]) );
  XOR U658 ( .A(key[111]), .B(\w3[0][111] ), .Z(out[111]) );
  XOR U659 ( .A(key[112]), .B(\w3[0][112] ), .Z(out[112]) );
  XOR U660 ( .A(key[113]), .B(\w3[0][113] ), .Z(out[113]) );
  XOR U661 ( .A(key[114]), .B(\w3[0][114] ), .Z(out[114]) );
  XOR U662 ( .A(key[115]), .B(\w3[0][115] ), .Z(out[115]) );
  XOR U663 ( .A(key[116]), .B(\w3[0][116] ), .Z(out[116]) );
  XOR U664 ( .A(key[117]), .B(\w3[0][117] ), .Z(out[117]) );
  XOR U665 ( .A(key[118]), .B(\w3[0][118] ), .Z(out[118]) );
  XOR U666 ( .A(key[119]), .B(\w3[0][119] ), .Z(out[119]) );
  XOR U667 ( .A(key[11]), .B(\w3[0][11] ), .Z(out[11]) );
  XOR U668 ( .A(key[120]), .B(\w3[0][120] ), .Z(out[120]) );
  XOR U669 ( .A(key[121]), .B(\w3[0][121] ), .Z(out[121]) );
  XOR U670 ( .A(key[122]), .B(\w3[0][122] ), .Z(out[122]) );
  XOR U671 ( .A(key[123]), .B(\w3[0][123] ), .Z(out[123]) );
  XOR U672 ( .A(key[124]), .B(\w3[0][124] ), .Z(out[124]) );
  XOR U673 ( .A(key[125]), .B(\w3[0][125] ), .Z(out[125]) );
  XOR U674 ( .A(key[126]), .B(\w3[0][126] ), .Z(out[126]) );
  XOR U675 ( .A(key[127]), .B(\w3[0][127] ), .Z(out[127]) );
  XOR U676 ( .A(key[12]), .B(\w3[0][12] ), .Z(out[12]) );
  XOR U677 ( .A(key[13]), .B(\w3[0][13] ), .Z(out[13]) );
  XOR U678 ( .A(key[14]), .B(\w3[0][14] ), .Z(out[14]) );
  XOR U679 ( .A(key[15]), .B(\w3[0][15] ), .Z(out[15]) );
  XOR U680 ( .A(key[16]), .B(\w3[0][16] ), .Z(out[16]) );
  XOR U681 ( .A(key[17]), .B(\w3[0][17] ), .Z(out[17]) );
  XOR U682 ( .A(key[18]), .B(\w3[0][18] ), .Z(out[18]) );
  XOR U683 ( .A(key[19]), .B(\w3[0][19] ), .Z(out[19]) );
  XOR U684 ( .A(key[1]), .B(\w3[0][1] ), .Z(out[1]) );
  XOR U685 ( .A(key[20]), .B(\w3[0][20] ), .Z(out[20]) );
  XOR U686 ( .A(key[21]), .B(\w3[0][21] ), .Z(out[21]) );
  XOR U687 ( .A(key[22]), .B(\w3[0][22] ), .Z(out[22]) );
  XOR U688 ( .A(key[23]), .B(\w3[0][23] ), .Z(out[23]) );
  XOR U689 ( .A(key[24]), .B(\w3[0][24] ), .Z(out[24]) );
  XOR U690 ( .A(key[25]), .B(\w3[0][25] ), .Z(out[25]) );
  XOR U691 ( .A(key[26]), .B(\w3[0][26] ), .Z(out[26]) );
  XOR U692 ( .A(key[27]), .B(\w3[0][27] ), .Z(out[27]) );
  XOR U693 ( .A(key[28]), .B(\w3[0][28] ), .Z(out[28]) );
  XOR U694 ( .A(key[29]), .B(\w3[0][29] ), .Z(out[29]) );
  XOR U695 ( .A(key[2]), .B(\w3[0][2] ), .Z(out[2]) );
  XOR U696 ( .A(key[30]), .B(\w3[0][30] ), .Z(out[30]) );
  XOR U697 ( .A(key[31]), .B(\w3[0][31] ), .Z(out[31]) );
  XOR U698 ( .A(key[32]), .B(\w3[0][32] ), .Z(out[32]) );
  XOR U699 ( .A(key[33]), .B(\w3[0][33] ), .Z(out[33]) );
  XOR U700 ( .A(key[34]), .B(\w3[0][34] ), .Z(out[34]) );
  XOR U701 ( .A(key[35]), .B(\w3[0][35] ), .Z(out[35]) );
  XOR U702 ( .A(key[36]), .B(\w3[0][36] ), .Z(out[36]) );
  XOR U703 ( .A(key[37]), .B(\w3[0][37] ), .Z(out[37]) );
  XOR U704 ( .A(key[38]), .B(\w3[0][38] ), .Z(out[38]) );
  XOR U705 ( .A(key[39]), .B(\w3[0][39] ), .Z(out[39]) );
  XOR U706 ( .A(key[3]), .B(\w3[0][3] ), .Z(out[3]) );
  XOR U707 ( .A(key[40]), .B(\w3[0][40] ), .Z(out[40]) );
  XOR U708 ( .A(key[41]), .B(\w3[0][41] ), .Z(out[41]) );
  XOR U709 ( .A(key[42]), .B(\w3[0][42] ), .Z(out[42]) );
  XOR U710 ( .A(key[43]), .B(\w3[0][43] ), .Z(out[43]) );
  XOR U711 ( .A(key[44]), .B(\w3[0][44] ), .Z(out[44]) );
  XOR U712 ( .A(key[45]), .B(\w3[0][45] ), .Z(out[45]) );
  XOR U713 ( .A(key[46]), .B(\w3[0][46] ), .Z(out[46]) );
  XOR U714 ( .A(key[47]), .B(\w3[0][47] ), .Z(out[47]) );
  XOR U715 ( .A(key[48]), .B(\w3[0][48] ), .Z(out[48]) );
  XOR U716 ( .A(key[49]), .B(\w3[0][49] ), .Z(out[49]) );
  XOR U717 ( .A(key[4]), .B(\w3[0][4] ), .Z(out[4]) );
  XOR U718 ( .A(key[50]), .B(\w3[0][50] ), .Z(out[50]) );
  XOR U719 ( .A(key[51]), .B(\w3[0][51] ), .Z(out[51]) );
  XOR U720 ( .A(key[52]), .B(\w3[0][52] ), .Z(out[52]) );
  XOR U721 ( .A(key[53]), .B(\w3[0][53] ), .Z(out[53]) );
  XOR U722 ( .A(key[54]), .B(\w3[0][54] ), .Z(out[54]) );
  XOR U723 ( .A(key[55]), .B(\w3[0][55] ), .Z(out[55]) );
  XOR U724 ( .A(key[56]), .B(\w3[0][56] ), .Z(out[56]) );
  XOR U725 ( .A(key[57]), .B(\w3[0][57] ), .Z(out[57]) );
  XOR U726 ( .A(key[58]), .B(\w3[0][58] ), .Z(out[58]) );
  XOR U727 ( .A(key[59]), .B(\w3[0][59] ), .Z(out[59]) );
  XOR U728 ( .A(key[5]), .B(\w3[0][5] ), .Z(out[5]) );
  XOR U729 ( .A(key[60]), .B(\w3[0][60] ), .Z(out[60]) );
  XOR U730 ( .A(key[61]), .B(\w3[0][61] ), .Z(out[61]) );
  XOR U731 ( .A(key[62]), .B(\w3[0][62] ), .Z(out[62]) );
  XOR U732 ( .A(key[63]), .B(\w3[0][63] ), .Z(out[63]) );
  XOR U733 ( .A(key[64]), .B(\w3[0][64] ), .Z(out[64]) );
  XOR U734 ( .A(key[65]), .B(\w3[0][65] ), .Z(out[65]) );
  XOR U735 ( .A(key[66]), .B(\w3[0][66] ), .Z(out[66]) );
  XOR U736 ( .A(key[67]), .B(\w3[0][67] ), .Z(out[67]) );
  XOR U737 ( .A(key[68]), .B(\w3[0][68] ), .Z(out[68]) );
  XOR U738 ( .A(key[69]), .B(\w3[0][69] ), .Z(out[69]) );
  XOR U739 ( .A(key[6]), .B(\w3[0][6] ), .Z(out[6]) );
  XOR U740 ( .A(key[70]), .B(\w3[0][70] ), .Z(out[70]) );
  XOR U741 ( .A(key[71]), .B(\w3[0][71] ), .Z(out[71]) );
  XOR U742 ( .A(key[72]), .B(\w3[0][72] ), .Z(out[72]) );
  XOR U743 ( .A(key[73]), .B(\w3[0][73] ), .Z(out[73]) );
  XOR U744 ( .A(key[74]), .B(\w3[0][74] ), .Z(out[74]) );
  XOR U745 ( .A(key[75]), .B(\w3[0][75] ), .Z(out[75]) );
  XOR U746 ( .A(key[76]), .B(\w3[0][76] ), .Z(out[76]) );
  XOR U747 ( .A(key[77]), .B(\w3[0][77] ), .Z(out[77]) );
  XOR U748 ( .A(key[78]), .B(\w3[0][78] ), .Z(out[78]) );
  XOR U749 ( .A(key[79]), .B(\w3[0][79] ), .Z(out[79]) );
  XOR U750 ( .A(key[7]), .B(\w3[0][7] ), .Z(out[7]) );
  XOR U751 ( .A(key[80]), .B(\w3[0][80] ), .Z(out[80]) );
  XOR U752 ( .A(key[81]), .B(\w3[0][81] ), .Z(out[81]) );
  XOR U753 ( .A(key[82]), .B(\w3[0][82] ), .Z(out[82]) );
  XOR U754 ( .A(key[83]), .B(\w3[0][83] ), .Z(out[83]) );
  XOR U755 ( .A(key[84]), .B(\w3[0][84] ), .Z(out[84]) );
  XOR U756 ( .A(key[85]), .B(\w3[0][85] ), .Z(out[85]) );
  XOR U757 ( .A(key[86]), .B(\w3[0][86] ), .Z(out[86]) );
  XOR U758 ( .A(key[87]), .B(\w3[0][87] ), .Z(out[87]) );
  XOR U759 ( .A(key[88]), .B(\w3[0][88] ), .Z(out[88]) );
  XOR U760 ( .A(key[89]), .B(\w3[0][89] ), .Z(out[89]) );
  XOR U761 ( .A(key[8]), .B(\w3[0][8] ), .Z(out[8]) );
  XOR U762 ( .A(key[90]), .B(\w3[0][90] ), .Z(out[90]) );
  XOR U763 ( .A(key[91]), .B(\w3[0][91] ), .Z(out[91]) );
  XOR U764 ( .A(key[92]), .B(\w3[0][92] ), .Z(out[92]) );
  XOR U765 ( .A(key[93]), .B(\w3[0][93] ), .Z(out[93]) );
  XOR U766 ( .A(key[94]), .B(\w3[0][94] ), .Z(out[94]) );
  XOR U767 ( .A(key[95]), .B(\w3[0][95] ), .Z(out[95]) );
  XOR U768 ( .A(key[96]), .B(\w3[0][96] ), .Z(out[96]) );
  XOR U769 ( .A(key[97]), .B(\w3[0][97] ), .Z(out[97]) );
  XOR U770 ( .A(key[98]), .B(\w3[0][98] ), .Z(out[98]) );
  XOR U771 ( .A(key[99]), .B(\w3[0][99] ), .Z(out[99]) );
  XOR U772 ( .A(key[9]), .B(\w3[0][9] ), .Z(out[9]) );
  NAND U773 ( .A(init), .B(state[0]), .Z(n260) );
  NAND U774 ( .A(n258), .B(msg[0]), .Z(n259) );
  NAND U775 ( .A(n260), .B(n259), .Z(\w0[0][0] ) );
  NAND U776 ( .A(init), .B(state[100]), .Z(n262) );
  NAND U777 ( .A(n258), .B(msg[100]), .Z(n261) );
  NAND U778 ( .A(n262), .B(n261), .Z(\w0[0][100] ) );
  NAND U779 ( .A(init), .B(state[101]), .Z(n264) );
  NAND U780 ( .A(n258), .B(msg[101]), .Z(n263) );
  NAND U781 ( .A(n264), .B(n263), .Z(\w0[0][101] ) );
  NAND U782 ( .A(init), .B(state[102]), .Z(n266) );
  NAND U783 ( .A(n258), .B(msg[102]), .Z(n265) );
  NAND U784 ( .A(n266), .B(n265), .Z(\w0[0][102] ) );
  NAND U785 ( .A(init), .B(state[103]), .Z(n268) );
  NAND U786 ( .A(n258), .B(msg[103]), .Z(n267) );
  NAND U787 ( .A(n268), .B(n267), .Z(\w0[0][103] ) );
  NAND U788 ( .A(init), .B(state[104]), .Z(n270) );
  NAND U789 ( .A(n258), .B(msg[104]), .Z(n269) );
  NAND U790 ( .A(n270), .B(n269), .Z(\w0[0][104] ) );
  NAND U791 ( .A(init), .B(state[105]), .Z(n272) );
  NAND U792 ( .A(n258), .B(msg[105]), .Z(n271) );
  NAND U793 ( .A(n272), .B(n271), .Z(\w0[0][105] ) );
  NAND U794 ( .A(init), .B(state[106]), .Z(n274) );
  NAND U795 ( .A(n258), .B(msg[106]), .Z(n273) );
  NAND U796 ( .A(n274), .B(n273), .Z(\w0[0][106] ) );
  NAND U797 ( .A(init), .B(state[107]), .Z(n276) );
  NAND U798 ( .A(n258), .B(msg[107]), .Z(n275) );
  NAND U799 ( .A(n276), .B(n275), .Z(\w0[0][107] ) );
  NAND U800 ( .A(init), .B(state[108]), .Z(n278) );
  NAND U801 ( .A(n258), .B(msg[108]), .Z(n277) );
  NAND U802 ( .A(n278), .B(n277), .Z(\w0[0][108] ) );
  NAND U803 ( .A(init), .B(state[109]), .Z(n280) );
  NAND U804 ( .A(n258), .B(msg[109]), .Z(n279) );
  NAND U805 ( .A(n280), .B(n279), .Z(\w0[0][109] ) );
  NAND U806 ( .A(init), .B(state[10]), .Z(n282) );
  NAND U807 ( .A(n258), .B(msg[10]), .Z(n281) );
  NAND U808 ( .A(n282), .B(n281), .Z(\w0[0][10] ) );
  NAND U809 ( .A(init), .B(state[110]), .Z(n284) );
  NAND U810 ( .A(n258), .B(msg[110]), .Z(n283) );
  NAND U811 ( .A(n284), .B(n283), .Z(\w0[0][110] ) );
  NAND U812 ( .A(init), .B(state[111]), .Z(n286) );
  NAND U813 ( .A(n258), .B(msg[111]), .Z(n285) );
  NAND U814 ( .A(n286), .B(n285), .Z(\w0[0][111] ) );
  NAND U815 ( .A(init), .B(state[112]), .Z(n288) );
  NAND U816 ( .A(n258), .B(msg[112]), .Z(n287) );
  NAND U817 ( .A(n288), .B(n287), .Z(\w0[0][112] ) );
  NAND U818 ( .A(init), .B(state[113]), .Z(n290) );
  NAND U819 ( .A(n258), .B(msg[113]), .Z(n289) );
  NAND U820 ( .A(n290), .B(n289), .Z(\w0[0][113] ) );
  NAND U821 ( .A(init), .B(state[114]), .Z(n292) );
  NAND U822 ( .A(n258), .B(msg[114]), .Z(n291) );
  NAND U823 ( .A(n292), .B(n291), .Z(\w0[0][114] ) );
  NAND U824 ( .A(init), .B(state[115]), .Z(n294) );
  NAND U825 ( .A(n258), .B(msg[115]), .Z(n293) );
  NAND U826 ( .A(n294), .B(n293), .Z(\w0[0][115] ) );
  NAND U827 ( .A(init), .B(state[116]), .Z(n296) );
  NAND U828 ( .A(n258), .B(msg[116]), .Z(n295) );
  NAND U829 ( .A(n296), .B(n295), .Z(\w0[0][116] ) );
  NAND U830 ( .A(init), .B(state[117]), .Z(n298) );
  NAND U831 ( .A(n258), .B(msg[117]), .Z(n297) );
  NAND U832 ( .A(n298), .B(n297), .Z(\w0[0][117] ) );
  NAND U833 ( .A(init), .B(state[118]), .Z(n300) );
  NAND U834 ( .A(n258), .B(msg[118]), .Z(n299) );
  NAND U835 ( .A(n300), .B(n299), .Z(\w0[0][118] ) );
  NAND U836 ( .A(init), .B(state[119]), .Z(n302) );
  NAND U837 ( .A(n258), .B(msg[119]), .Z(n301) );
  NAND U838 ( .A(n302), .B(n301), .Z(\w0[0][119] ) );
  NAND U839 ( .A(init), .B(state[11]), .Z(n304) );
  NAND U840 ( .A(n258), .B(msg[11]), .Z(n303) );
  NAND U841 ( .A(n304), .B(n303), .Z(\w0[0][11] ) );
  NAND U842 ( .A(init), .B(state[120]), .Z(n306) );
  NAND U843 ( .A(n258), .B(msg[120]), .Z(n305) );
  NAND U844 ( .A(n306), .B(n305), .Z(\w0[0][120] ) );
  NAND U845 ( .A(init), .B(state[121]), .Z(n308) );
  NAND U846 ( .A(n258), .B(msg[121]), .Z(n307) );
  NAND U847 ( .A(n308), .B(n307), .Z(\w0[0][121] ) );
  NAND U848 ( .A(init), .B(state[122]), .Z(n310) );
  NAND U849 ( .A(n258), .B(msg[122]), .Z(n309) );
  NAND U850 ( .A(n310), .B(n309), .Z(\w0[0][122] ) );
  NAND U851 ( .A(init), .B(state[123]), .Z(n312) );
  NAND U852 ( .A(n258), .B(msg[123]), .Z(n311) );
  NAND U853 ( .A(n312), .B(n311), .Z(\w0[0][123] ) );
  NAND U854 ( .A(init), .B(state[124]), .Z(n314) );
  NAND U855 ( .A(n258), .B(msg[124]), .Z(n313) );
  NAND U856 ( .A(n314), .B(n313), .Z(\w0[0][124] ) );
  NAND U857 ( .A(init), .B(state[125]), .Z(n316) );
  NAND U858 ( .A(n258), .B(msg[125]), .Z(n315) );
  NAND U859 ( .A(n316), .B(n315), .Z(\w0[0][125] ) );
  NAND U860 ( .A(init), .B(state[126]), .Z(n318) );
  NAND U861 ( .A(n258), .B(msg[126]), .Z(n317) );
  NAND U862 ( .A(n318), .B(n317), .Z(\w0[0][126] ) );
  NAND U863 ( .A(init), .B(state[127]), .Z(n320) );
  NAND U864 ( .A(n258), .B(msg[127]), .Z(n319) );
  NAND U865 ( .A(n320), .B(n319), .Z(\w0[0][127] ) );
  NAND U866 ( .A(init), .B(state[12]), .Z(n322) );
  NAND U867 ( .A(n258), .B(msg[12]), .Z(n321) );
  NAND U868 ( .A(n322), .B(n321), .Z(\w0[0][12] ) );
  NAND U869 ( .A(init), .B(state[13]), .Z(n324) );
  NAND U870 ( .A(n258), .B(msg[13]), .Z(n323) );
  NAND U871 ( .A(n324), .B(n323), .Z(\w0[0][13] ) );
  NAND U872 ( .A(init), .B(state[14]), .Z(n326) );
  NAND U873 ( .A(n258), .B(msg[14]), .Z(n325) );
  NAND U874 ( .A(n326), .B(n325), .Z(\w0[0][14] ) );
  NAND U875 ( .A(init), .B(state[15]), .Z(n328) );
  NAND U876 ( .A(n258), .B(msg[15]), .Z(n327) );
  NAND U877 ( .A(n328), .B(n327), .Z(\w0[0][15] ) );
  NAND U878 ( .A(init), .B(state[16]), .Z(n330) );
  NAND U879 ( .A(n258), .B(msg[16]), .Z(n329) );
  NAND U880 ( .A(n330), .B(n329), .Z(\w0[0][16] ) );
  NAND U881 ( .A(init), .B(state[17]), .Z(n332) );
  NAND U882 ( .A(n258), .B(msg[17]), .Z(n331) );
  NAND U883 ( .A(n332), .B(n331), .Z(\w0[0][17] ) );
  NAND U884 ( .A(init), .B(state[18]), .Z(n334) );
  NAND U885 ( .A(n258), .B(msg[18]), .Z(n333) );
  NAND U886 ( .A(n334), .B(n333), .Z(\w0[0][18] ) );
  NAND U887 ( .A(init), .B(state[19]), .Z(n336) );
  NAND U888 ( .A(n258), .B(msg[19]), .Z(n335) );
  NAND U889 ( .A(n336), .B(n335), .Z(\w0[0][19] ) );
  NAND U890 ( .A(init), .B(state[1]), .Z(n338) );
  NAND U891 ( .A(n258), .B(msg[1]), .Z(n337) );
  NAND U892 ( .A(n338), .B(n337), .Z(\w0[0][1] ) );
  NAND U893 ( .A(init), .B(state[20]), .Z(n340) );
  NAND U894 ( .A(n258), .B(msg[20]), .Z(n339) );
  NAND U895 ( .A(n340), .B(n339), .Z(\w0[0][20] ) );
  NAND U896 ( .A(init), .B(state[21]), .Z(n342) );
  NAND U897 ( .A(n258), .B(msg[21]), .Z(n341) );
  NAND U898 ( .A(n342), .B(n341), .Z(\w0[0][21] ) );
  NAND U899 ( .A(init), .B(state[22]), .Z(n344) );
  NAND U900 ( .A(n258), .B(msg[22]), .Z(n343) );
  NAND U901 ( .A(n344), .B(n343), .Z(\w0[0][22] ) );
  NAND U902 ( .A(init), .B(state[23]), .Z(n346) );
  NAND U903 ( .A(n258), .B(msg[23]), .Z(n345) );
  NAND U904 ( .A(n346), .B(n345), .Z(\w0[0][23] ) );
  NAND U905 ( .A(init), .B(state[24]), .Z(n348) );
  NAND U906 ( .A(n258), .B(msg[24]), .Z(n347) );
  NAND U907 ( .A(n348), .B(n347), .Z(\w0[0][24] ) );
  NAND U908 ( .A(init), .B(state[25]), .Z(n350) );
  NAND U909 ( .A(n258), .B(msg[25]), .Z(n349) );
  NAND U910 ( .A(n350), .B(n349), .Z(\w0[0][25] ) );
  NAND U911 ( .A(init), .B(state[26]), .Z(n352) );
  NAND U912 ( .A(n258), .B(msg[26]), .Z(n351) );
  NAND U913 ( .A(n352), .B(n351), .Z(\w0[0][26] ) );
  NAND U914 ( .A(init), .B(state[27]), .Z(n354) );
  NAND U915 ( .A(n258), .B(msg[27]), .Z(n353) );
  NAND U916 ( .A(n354), .B(n353), .Z(\w0[0][27] ) );
  NAND U917 ( .A(init), .B(state[28]), .Z(n356) );
  NAND U918 ( .A(n258), .B(msg[28]), .Z(n355) );
  NAND U919 ( .A(n356), .B(n355), .Z(\w0[0][28] ) );
  NAND U920 ( .A(init), .B(state[29]), .Z(n358) );
  NAND U921 ( .A(n258), .B(msg[29]), .Z(n357) );
  NAND U922 ( .A(n358), .B(n357), .Z(\w0[0][29] ) );
  NAND U923 ( .A(init), .B(state[2]), .Z(n360) );
  NAND U924 ( .A(n258), .B(msg[2]), .Z(n359) );
  NAND U925 ( .A(n360), .B(n359), .Z(\w0[0][2] ) );
  NAND U926 ( .A(init), .B(state[30]), .Z(n362) );
  NAND U927 ( .A(n258), .B(msg[30]), .Z(n361) );
  NAND U928 ( .A(n362), .B(n361), .Z(\w0[0][30] ) );
  NAND U929 ( .A(init), .B(state[31]), .Z(n364) );
  NAND U930 ( .A(n258), .B(msg[31]), .Z(n363) );
  NAND U931 ( .A(n364), .B(n363), .Z(\w0[0][31] ) );
  NAND U932 ( .A(init), .B(state[32]), .Z(n366) );
  NAND U933 ( .A(n258), .B(msg[32]), .Z(n365) );
  NAND U934 ( .A(n366), .B(n365), .Z(\w0[0][32] ) );
  NAND U935 ( .A(init), .B(state[33]), .Z(n368) );
  NAND U936 ( .A(n258), .B(msg[33]), .Z(n367) );
  NAND U937 ( .A(n368), .B(n367), .Z(\w0[0][33] ) );
  NAND U938 ( .A(init), .B(state[34]), .Z(n370) );
  NAND U939 ( .A(n258), .B(msg[34]), .Z(n369) );
  NAND U940 ( .A(n370), .B(n369), .Z(\w0[0][34] ) );
  NAND U941 ( .A(init), .B(state[35]), .Z(n372) );
  NAND U942 ( .A(n258), .B(msg[35]), .Z(n371) );
  NAND U943 ( .A(n372), .B(n371), .Z(\w0[0][35] ) );
  NAND U944 ( .A(init), .B(state[36]), .Z(n374) );
  NAND U945 ( .A(n258), .B(msg[36]), .Z(n373) );
  NAND U946 ( .A(n374), .B(n373), .Z(\w0[0][36] ) );
  NAND U947 ( .A(init), .B(state[37]), .Z(n376) );
  NAND U948 ( .A(n258), .B(msg[37]), .Z(n375) );
  NAND U949 ( .A(n376), .B(n375), .Z(\w0[0][37] ) );
  NAND U950 ( .A(init), .B(state[38]), .Z(n378) );
  NAND U951 ( .A(n258), .B(msg[38]), .Z(n377) );
  NAND U952 ( .A(n378), .B(n377), .Z(\w0[0][38] ) );
  NAND U953 ( .A(init), .B(state[39]), .Z(n380) );
  NAND U954 ( .A(n258), .B(msg[39]), .Z(n379) );
  NAND U955 ( .A(n380), .B(n379), .Z(\w0[0][39] ) );
  NAND U956 ( .A(init), .B(state[3]), .Z(n382) );
  NAND U957 ( .A(n258), .B(msg[3]), .Z(n381) );
  NAND U958 ( .A(n382), .B(n381), .Z(\w0[0][3] ) );
  NAND U959 ( .A(init), .B(state[40]), .Z(n384) );
  NAND U960 ( .A(n258), .B(msg[40]), .Z(n383) );
  NAND U961 ( .A(n384), .B(n383), .Z(\w0[0][40] ) );
  NAND U962 ( .A(init), .B(state[41]), .Z(n386) );
  NAND U963 ( .A(n258), .B(msg[41]), .Z(n385) );
  NAND U964 ( .A(n386), .B(n385), .Z(\w0[0][41] ) );
  NAND U965 ( .A(init), .B(state[42]), .Z(n388) );
  NAND U966 ( .A(n258), .B(msg[42]), .Z(n387) );
  NAND U967 ( .A(n388), .B(n387), .Z(\w0[0][42] ) );
  NAND U968 ( .A(init), .B(state[43]), .Z(n390) );
  NAND U969 ( .A(n258), .B(msg[43]), .Z(n389) );
  NAND U970 ( .A(n390), .B(n389), .Z(\w0[0][43] ) );
  NAND U971 ( .A(init), .B(state[44]), .Z(n392) );
  NAND U972 ( .A(n258), .B(msg[44]), .Z(n391) );
  NAND U973 ( .A(n392), .B(n391), .Z(\w0[0][44] ) );
  NAND U974 ( .A(init), .B(state[45]), .Z(n394) );
  NAND U975 ( .A(n258), .B(msg[45]), .Z(n393) );
  NAND U976 ( .A(n394), .B(n393), .Z(\w0[0][45] ) );
  NAND U977 ( .A(init), .B(state[46]), .Z(n396) );
  NAND U978 ( .A(n258), .B(msg[46]), .Z(n395) );
  NAND U979 ( .A(n396), .B(n395), .Z(\w0[0][46] ) );
  NAND U980 ( .A(init), .B(state[47]), .Z(n398) );
  NAND U981 ( .A(n258), .B(msg[47]), .Z(n397) );
  NAND U982 ( .A(n398), .B(n397), .Z(\w0[0][47] ) );
  NAND U983 ( .A(init), .B(state[48]), .Z(n400) );
  NAND U984 ( .A(n258), .B(msg[48]), .Z(n399) );
  NAND U985 ( .A(n400), .B(n399), .Z(\w0[0][48] ) );
  NAND U986 ( .A(init), .B(state[49]), .Z(n402) );
  NAND U987 ( .A(n258), .B(msg[49]), .Z(n401) );
  NAND U988 ( .A(n402), .B(n401), .Z(\w0[0][49] ) );
  NAND U989 ( .A(init), .B(state[4]), .Z(n404) );
  NAND U990 ( .A(n258), .B(msg[4]), .Z(n403) );
  NAND U991 ( .A(n404), .B(n403), .Z(\w0[0][4] ) );
  NAND U992 ( .A(init), .B(state[50]), .Z(n406) );
  NAND U993 ( .A(n258), .B(msg[50]), .Z(n405) );
  NAND U994 ( .A(n406), .B(n405), .Z(\w0[0][50] ) );
  NAND U995 ( .A(init), .B(state[51]), .Z(n408) );
  NAND U996 ( .A(n258), .B(msg[51]), .Z(n407) );
  NAND U997 ( .A(n408), .B(n407), .Z(\w0[0][51] ) );
  NAND U998 ( .A(init), .B(state[52]), .Z(n410) );
  NAND U999 ( .A(n258), .B(msg[52]), .Z(n409) );
  NAND U1000 ( .A(n410), .B(n409), .Z(\w0[0][52] ) );
  NAND U1001 ( .A(init), .B(state[53]), .Z(n412) );
  NAND U1002 ( .A(n258), .B(msg[53]), .Z(n411) );
  NAND U1003 ( .A(n412), .B(n411), .Z(\w0[0][53] ) );
  NAND U1004 ( .A(init), .B(state[54]), .Z(n414) );
  NAND U1005 ( .A(n258), .B(msg[54]), .Z(n413) );
  NAND U1006 ( .A(n414), .B(n413), .Z(\w0[0][54] ) );
  NAND U1007 ( .A(init), .B(state[55]), .Z(n416) );
  NAND U1008 ( .A(n258), .B(msg[55]), .Z(n415) );
  NAND U1009 ( .A(n416), .B(n415), .Z(\w0[0][55] ) );
  NAND U1010 ( .A(init), .B(state[56]), .Z(n418) );
  NAND U1011 ( .A(n258), .B(msg[56]), .Z(n417) );
  NAND U1012 ( .A(n418), .B(n417), .Z(\w0[0][56] ) );
  NAND U1013 ( .A(init), .B(state[57]), .Z(n420) );
  NAND U1014 ( .A(n258), .B(msg[57]), .Z(n419) );
  NAND U1015 ( .A(n420), .B(n419), .Z(\w0[0][57] ) );
  NAND U1016 ( .A(init), .B(state[58]), .Z(n422) );
  NAND U1017 ( .A(n258), .B(msg[58]), .Z(n421) );
  NAND U1018 ( .A(n422), .B(n421), .Z(\w0[0][58] ) );
  NAND U1019 ( .A(init), .B(state[59]), .Z(n424) );
  NAND U1020 ( .A(n258), .B(msg[59]), .Z(n423) );
  NAND U1021 ( .A(n424), .B(n423), .Z(\w0[0][59] ) );
  NAND U1022 ( .A(init), .B(state[5]), .Z(n426) );
  NAND U1023 ( .A(n258), .B(msg[5]), .Z(n425) );
  NAND U1024 ( .A(n426), .B(n425), .Z(\w0[0][5] ) );
  NAND U1025 ( .A(init), .B(state[60]), .Z(n428) );
  NAND U1026 ( .A(n258), .B(msg[60]), .Z(n427) );
  NAND U1027 ( .A(n428), .B(n427), .Z(\w0[0][60] ) );
  NAND U1028 ( .A(init), .B(state[61]), .Z(n430) );
  NAND U1029 ( .A(n258), .B(msg[61]), .Z(n429) );
  NAND U1030 ( .A(n430), .B(n429), .Z(\w0[0][61] ) );
  NAND U1031 ( .A(init), .B(state[62]), .Z(n432) );
  NAND U1032 ( .A(n258), .B(msg[62]), .Z(n431) );
  NAND U1033 ( .A(n432), .B(n431), .Z(\w0[0][62] ) );
  NAND U1034 ( .A(init), .B(state[63]), .Z(n434) );
  NAND U1035 ( .A(n258), .B(msg[63]), .Z(n433) );
  NAND U1036 ( .A(n434), .B(n433), .Z(\w0[0][63] ) );
  NAND U1037 ( .A(init), .B(state[64]), .Z(n436) );
  NAND U1038 ( .A(n258), .B(msg[64]), .Z(n435) );
  NAND U1039 ( .A(n436), .B(n435), .Z(\w0[0][64] ) );
  NAND U1040 ( .A(init), .B(state[65]), .Z(n438) );
  NAND U1041 ( .A(n258), .B(msg[65]), .Z(n437) );
  NAND U1042 ( .A(n438), .B(n437), .Z(\w0[0][65] ) );
  NAND U1043 ( .A(init), .B(state[66]), .Z(n440) );
  NAND U1044 ( .A(n258), .B(msg[66]), .Z(n439) );
  NAND U1045 ( .A(n440), .B(n439), .Z(\w0[0][66] ) );
  NAND U1046 ( .A(init), .B(state[67]), .Z(n442) );
  NAND U1047 ( .A(n258), .B(msg[67]), .Z(n441) );
  NAND U1048 ( .A(n442), .B(n441), .Z(\w0[0][67] ) );
  NAND U1049 ( .A(init), .B(state[68]), .Z(n444) );
  NAND U1050 ( .A(n258), .B(msg[68]), .Z(n443) );
  NAND U1051 ( .A(n444), .B(n443), .Z(\w0[0][68] ) );
  NAND U1052 ( .A(init), .B(state[69]), .Z(n446) );
  NAND U1053 ( .A(n258), .B(msg[69]), .Z(n445) );
  NAND U1054 ( .A(n446), .B(n445), .Z(\w0[0][69] ) );
  NAND U1055 ( .A(init), .B(state[6]), .Z(n448) );
  NAND U1056 ( .A(n258), .B(msg[6]), .Z(n447) );
  NAND U1057 ( .A(n448), .B(n447), .Z(\w0[0][6] ) );
  NAND U1058 ( .A(init), .B(state[70]), .Z(n450) );
  NAND U1059 ( .A(n258), .B(msg[70]), .Z(n449) );
  NAND U1060 ( .A(n450), .B(n449), .Z(\w0[0][70] ) );
  NAND U1061 ( .A(init), .B(state[71]), .Z(n452) );
  NAND U1062 ( .A(n258), .B(msg[71]), .Z(n451) );
  NAND U1063 ( .A(n452), .B(n451), .Z(\w0[0][71] ) );
  NAND U1064 ( .A(init), .B(state[72]), .Z(n454) );
  NAND U1065 ( .A(n258), .B(msg[72]), .Z(n453) );
  NAND U1066 ( .A(n454), .B(n453), .Z(\w0[0][72] ) );
  NAND U1067 ( .A(init), .B(state[73]), .Z(n456) );
  NAND U1068 ( .A(n258), .B(msg[73]), .Z(n455) );
  NAND U1069 ( .A(n456), .B(n455), .Z(\w0[0][73] ) );
  NAND U1070 ( .A(init), .B(state[74]), .Z(n458) );
  NAND U1071 ( .A(n258), .B(msg[74]), .Z(n457) );
  NAND U1072 ( .A(n458), .B(n457), .Z(\w0[0][74] ) );
  NAND U1073 ( .A(init), .B(state[75]), .Z(n460) );
  NAND U1074 ( .A(n258), .B(msg[75]), .Z(n459) );
  NAND U1075 ( .A(n460), .B(n459), .Z(\w0[0][75] ) );
  NAND U1076 ( .A(init), .B(state[76]), .Z(n462) );
  NAND U1077 ( .A(n258), .B(msg[76]), .Z(n461) );
  NAND U1078 ( .A(n462), .B(n461), .Z(\w0[0][76] ) );
  NAND U1079 ( .A(init), .B(state[77]), .Z(n464) );
  NAND U1080 ( .A(n258), .B(msg[77]), .Z(n463) );
  NAND U1081 ( .A(n464), .B(n463), .Z(\w0[0][77] ) );
  NAND U1082 ( .A(init), .B(state[78]), .Z(n466) );
  NAND U1083 ( .A(n258), .B(msg[78]), .Z(n465) );
  NAND U1084 ( .A(n466), .B(n465), .Z(\w0[0][78] ) );
  NAND U1085 ( .A(init), .B(state[79]), .Z(n468) );
  NAND U1086 ( .A(n258), .B(msg[79]), .Z(n467) );
  NAND U1087 ( .A(n468), .B(n467), .Z(\w0[0][79] ) );
  NAND U1088 ( .A(init), .B(state[7]), .Z(n470) );
  NAND U1089 ( .A(n258), .B(msg[7]), .Z(n469) );
  NAND U1090 ( .A(n470), .B(n469), .Z(\w0[0][7] ) );
  NAND U1091 ( .A(init), .B(state[80]), .Z(n472) );
  NAND U1092 ( .A(n258), .B(msg[80]), .Z(n471) );
  NAND U1093 ( .A(n472), .B(n471), .Z(\w0[0][80] ) );
  NAND U1094 ( .A(init), .B(state[81]), .Z(n474) );
  NAND U1095 ( .A(n258), .B(msg[81]), .Z(n473) );
  NAND U1096 ( .A(n474), .B(n473), .Z(\w0[0][81] ) );
  NAND U1097 ( .A(init), .B(state[82]), .Z(n476) );
  NAND U1098 ( .A(n258), .B(msg[82]), .Z(n475) );
  NAND U1099 ( .A(n476), .B(n475), .Z(\w0[0][82] ) );
  NAND U1100 ( .A(init), .B(state[83]), .Z(n478) );
  NAND U1101 ( .A(n258), .B(msg[83]), .Z(n477) );
  NAND U1102 ( .A(n478), .B(n477), .Z(\w0[0][83] ) );
  NAND U1103 ( .A(init), .B(state[84]), .Z(n480) );
  NAND U1104 ( .A(n258), .B(msg[84]), .Z(n479) );
  NAND U1105 ( .A(n480), .B(n479), .Z(\w0[0][84] ) );
  NAND U1106 ( .A(init), .B(state[85]), .Z(n482) );
  NAND U1107 ( .A(n258), .B(msg[85]), .Z(n481) );
  NAND U1108 ( .A(n482), .B(n481), .Z(\w0[0][85] ) );
  NAND U1109 ( .A(init), .B(state[86]), .Z(n484) );
  NAND U1110 ( .A(n258), .B(msg[86]), .Z(n483) );
  NAND U1111 ( .A(n484), .B(n483), .Z(\w0[0][86] ) );
  NAND U1112 ( .A(init), .B(state[87]), .Z(n486) );
  NAND U1113 ( .A(n258), .B(msg[87]), .Z(n485) );
  NAND U1114 ( .A(n486), .B(n485), .Z(\w0[0][87] ) );
  NAND U1115 ( .A(init), .B(state[88]), .Z(n488) );
  NAND U1116 ( .A(n258), .B(msg[88]), .Z(n487) );
  NAND U1117 ( .A(n488), .B(n487), .Z(\w0[0][88] ) );
  NAND U1118 ( .A(init), .B(state[89]), .Z(n490) );
  NAND U1119 ( .A(n258), .B(msg[89]), .Z(n489) );
  NAND U1120 ( .A(n490), .B(n489), .Z(\w0[0][89] ) );
  NAND U1121 ( .A(init), .B(state[8]), .Z(n492) );
  NAND U1122 ( .A(n258), .B(msg[8]), .Z(n491) );
  NAND U1123 ( .A(n492), .B(n491), .Z(\w0[0][8] ) );
  NAND U1124 ( .A(init), .B(state[90]), .Z(n494) );
  NAND U1125 ( .A(n258), .B(msg[90]), .Z(n493) );
  NAND U1126 ( .A(n494), .B(n493), .Z(\w0[0][90] ) );
  NAND U1127 ( .A(init), .B(state[91]), .Z(n496) );
  NAND U1128 ( .A(n258), .B(msg[91]), .Z(n495) );
  NAND U1129 ( .A(n496), .B(n495), .Z(\w0[0][91] ) );
  NAND U1130 ( .A(init), .B(state[92]), .Z(n498) );
  NAND U1131 ( .A(n258), .B(msg[92]), .Z(n497) );
  NAND U1132 ( .A(n498), .B(n497), .Z(\w0[0][92] ) );
  NAND U1133 ( .A(init), .B(state[93]), .Z(n500) );
  NAND U1134 ( .A(n258), .B(msg[93]), .Z(n499) );
  NAND U1135 ( .A(n500), .B(n499), .Z(\w0[0][93] ) );
  NAND U1136 ( .A(init), .B(state[94]), .Z(n502) );
  NAND U1137 ( .A(n258), .B(msg[94]), .Z(n501) );
  NAND U1138 ( .A(n502), .B(n501), .Z(\w0[0][94] ) );
  NAND U1139 ( .A(init), .B(state[95]), .Z(n504) );
  NAND U1140 ( .A(n258), .B(msg[95]), .Z(n503) );
  NAND U1141 ( .A(n504), .B(n503), .Z(\w0[0][95] ) );
  NAND U1142 ( .A(init), .B(state[96]), .Z(n506) );
  NAND U1143 ( .A(n258), .B(msg[96]), .Z(n505) );
  NAND U1144 ( .A(n506), .B(n505), .Z(\w0[0][96] ) );
  NAND U1145 ( .A(init), .B(state[97]), .Z(n508) );
  NAND U1146 ( .A(n258), .B(msg[97]), .Z(n507) );
  NAND U1147 ( .A(n508), .B(n507), .Z(\w0[0][97] ) );
  NAND U1148 ( .A(init), .B(state[98]), .Z(n510) );
  NAND U1149 ( .A(n258), .B(msg[98]), .Z(n509) );
  NAND U1150 ( .A(n510), .B(n509), .Z(\w0[0][98] ) );
  NAND U1151 ( .A(init), .B(state[99]), .Z(n512) );
  NAND U1152 ( .A(n258), .B(msg[99]), .Z(n511) );
  NAND U1153 ( .A(n512), .B(n511), .Z(\w0[0][99] ) );
  NAND U1154 ( .A(init), .B(state[9]), .Z(n514) );
  NAND U1155 ( .A(n258), .B(msg[9]), .Z(n513) );
  NAND U1156 ( .A(n514), .B(n513), .Z(\w0[0][9] ) );
  XOR U1157 ( .A(key[0]), .B(\w0[0][0] ), .Z(\w1[0][0] ) );
  XOR U1158 ( .A(key[100]), .B(\w0[0][100] ), .Z(\w1[0][100] ) );
  XOR U1159 ( .A(key[101]), .B(\w0[0][101] ), .Z(\w1[0][101] ) );
  XOR U1160 ( .A(key[102]), .B(\w0[0][102] ), .Z(\w1[0][102] ) );
  XOR U1161 ( .A(key[103]), .B(\w0[0][103] ), .Z(\w1[0][103] ) );
  XOR U1162 ( .A(key[104]), .B(\w0[0][104] ), .Z(\w1[0][104] ) );
  XOR U1163 ( .A(key[105]), .B(\w0[0][105] ), .Z(\w1[0][105] ) );
  XOR U1164 ( .A(key[106]), .B(\w0[0][106] ), .Z(\w1[0][106] ) );
  XOR U1165 ( .A(key[107]), .B(\w0[0][107] ), .Z(\w1[0][107] ) );
  XOR U1166 ( .A(key[108]), .B(\w0[0][108] ), .Z(\w1[0][108] ) );
  XOR U1167 ( .A(key[109]), .B(\w0[0][109] ), .Z(\w1[0][109] ) );
  XOR U1168 ( .A(key[10]), .B(\w0[0][10] ), .Z(\w1[0][10] ) );
  XOR U1169 ( .A(key[110]), .B(\w0[0][110] ), .Z(\w1[0][110] ) );
  XOR U1170 ( .A(key[111]), .B(\w0[0][111] ), .Z(\w1[0][111] ) );
  XOR U1171 ( .A(key[112]), .B(\w0[0][112] ), .Z(\w1[0][112] ) );
  XOR U1172 ( .A(key[113]), .B(\w0[0][113] ), .Z(\w1[0][113] ) );
  XOR U1173 ( .A(key[114]), .B(\w0[0][114] ), .Z(\w1[0][114] ) );
  XOR U1174 ( .A(key[115]), .B(\w0[0][115] ), .Z(\w1[0][115] ) );
  XOR U1175 ( .A(key[116]), .B(\w0[0][116] ), .Z(\w1[0][116] ) );
  XOR U1176 ( .A(key[117]), .B(\w0[0][117] ), .Z(\w1[0][117] ) );
  XOR U1177 ( .A(key[118]), .B(\w0[0][118] ), .Z(\w1[0][118] ) );
  XOR U1178 ( .A(key[119]), .B(\w0[0][119] ), .Z(\w1[0][119] ) );
  XOR U1179 ( .A(key[11]), .B(\w0[0][11] ), .Z(\w1[0][11] ) );
  XOR U1180 ( .A(key[120]), .B(\w0[0][120] ), .Z(\w1[0][120] ) );
  XOR U1181 ( .A(key[121]), .B(\w0[0][121] ), .Z(\w1[0][121] ) );
  XOR U1182 ( .A(key[122]), .B(\w0[0][122] ), .Z(\w1[0][122] ) );
  XOR U1183 ( .A(key[123]), .B(\w0[0][123] ), .Z(\w1[0][123] ) );
  XOR U1184 ( .A(key[124]), .B(\w0[0][124] ), .Z(\w1[0][124] ) );
  XOR U1185 ( .A(key[125]), .B(\w0[0][125] ), .Z(\w1[0][125] ) );
  XOR U1186 ( .A(key[126]), .B(\w0[0][126] ), .Z(\w1[0][126] ) );
  XOR U1187 ( .A(key[127]), .B(\w0[0][127] ), .Z(\w1[0][127] ) );
  XOR U1188 ( .A(key[12]), .B(\w0[0][12] ), .Z(\w1[0][12] ) );
  XOR U1189 ( .A(key[13]), .B(\w0[0][13] ), .Z(\w1[0][13] ) );
  XOR U1190 ( .A(key[14]), .B(\w0[0][14] ), .Z(\w1[0][14] ) );
  XOR U1191 ( .A(key[15]), .B(\w0[0][15] ), .Z(\w1[0][15] ) );
  XOR U1192 ( .A(key[16]), .B(\w0[0][16] ), .Z(\w1[0][16] ) );
  XOR U1193 ( .A(key[17]), .B(\w0[0][17] ), .Z(\w1[0][17] ) );
  XOR U1194 ( .A(key[18]), .B(\w0[0][18] ), .Z(\w1[0][18] ) );
  XOR U1195 ( .A(key[19]), .B(\w0[0][19] ), .Z(\w1[0][19] ) );
  XOR U1196 ( .A(key[1]), .B(\w0[0][1] ), .Z(\w1[0][1] ) );
  XOR U1197 ( .A(key[20]), .B(\w0[0][20] ), .Z(\w1[0][20] ) );
  XOR U1198 ( .A(key[21]), .B(\w0[0][21] ), .Z(\w1[0][21] ) );
  XOR U1199 ( .A(key[22]), .B(\w0[0][22] ), .Z(\w1[0][22] ) );
  XOR U1200 ( .A(key[23]), .B(\w0[0][23] ), .Z(\w1[0][23] ) );
  XOR U1201 ( .A(key[24]), .B(\w0[0][24] ), .Z(\w1[0][24] ) );
  XOR U1202 ( .A(key[25]), .B(\w0[0][25] ), .Z(\w1[0][25] ) );
  XOR U1203 ( .A(key[26]), .B(\w0[0][26] ), .Z(\w1[0][26] ) );
  XOR U1204 ( .A(key[27]), .B(\w0[0][27] ), .Z(\w1[0][27] ) );
  XOR U1205 ( .A(key[28]), .B(\w0[0][28] ), .Z(\w1[0][28] ) );
  XOR U1206 ( .A(key[29]), .B(\w0[0][29] ), .Z(\w1[0][29] ) );
  XOR U1207 ( .A(key[2]), .B(\w0[0][2] ), .Z(\w1[0][2] ) );
  XOR U1208 ( .A(key[30]), .B(\w0[0][30] ), .Z(\w1[0][30] ) );
  XOR U1209 ( .A(key[31]), .B(\w0[0][31] ), .Z(\w1[0][31] ) );
  XOR U1210 ( .A(key[32]), .B(\w0[0][32] ), .Z(\w1[0][32] ) );
  XOR U1211 ( .A(key[33]), .B(\w0[0][33] ), .Z(\w1[0][33] ) );
  XOR U1212 ( .A(key[34]), .B(\w0[0][34] ), .Z(\w1[0][34] ) );
  XOR U1213 ( .A(key[35]), .B(\w0[0][35] ), .Z(\w1[0][35] ) );
  XOR U1214 ( .A(key[36]), .B(\w0[0][36] ), .Z(\w1[0][36] ) );
  XOR U1215 ( .A(key[37]), .B(\w0[0][37] ), .Z(\w1[0][37] ) );
  XOR U1216 ( .A(key[38]), .B(\w0[0][38] ), .Z(\w1[0][38] ) );
  XOR U1217 ( .A(key[39]), .B(\w0[0][39] ), .Z(\w1[0][39] ) );
  XOR U1218 ( .A(key[3]), .B(\w0[0][3] ), .Z(\w1[0][3] ) );
  XOR U1219 ( .A(key[40]), .B(\w0[0][40] ), .Z(\w1[0][40] ) );
  XOR U1220 ( .A(key[41]), .B(\w0[0][41] ), .Z(\w1[0][41] ) );
  XOR U1221 ( .A(key[42]), .B(\w0[0][42] ), .Z(\w1[0][42] ) );
  XOR U1222 ( .A(key[43]), .B(\w0[0][43] ), .Z(\w1[0][43] ) );
  XOR U1223 ( .A(key[44]), .B(\w0[0][44] ), .Z(\w1[0][44] ) );
  XOR U1224 ( .A(key[45]), .B(\w0[0][45] ), .Z(\w1[0][45] ) );
  XOR U1225 ( .A(key[46]), .B(\w0[0][46] ), .Z(\w1[0][46] ) );
  XOR U1226 ( .A(key[47]), .B(\w0[0][47] ), .Z(\w1[0][47] ) );
  XOR U1227 ( .A(key[48]), .B(\w0[0][48] ), .Z(\w1[0][48] ) );
  XOR U1228 ( .A(key[49]), .B(\w0[0][49] ), .Z(\w1[0][49] ) );
  XOR U1229 ( .A(key[4]), .B(\w0[0][4] ), .Z(\w1[0][4] ) );
  XOR U1230 ( .A(key[50]), .B(\w0[0][50] ), .Z(\w1[0][50] ) );
  XOR U1231 ( .A(key[51]), .B(\w0[0][51] ), .Z(\w1[0][51] ) );
  XOR U1232 ( .A(key[52]), .B(\w0[0][52] ), .Z(\w1[0][52] ) );
  XOR U1233 ( .A(key[53]), .B(\w0[0][53] ), .Z(\w1[0][53] ) );
  XOR U1234 ( .A(key[54]), .B(\w0[0][54] ), .Z(\w1[0][54] ) );
  XOR U1235 ( .A(key[55]), .B(\w0[0][55] ), .Z(\w1[0][55] ) );
  XOR U1236 ( .A(key[56]), .B(\w0[0][56] ), .Z(\w1[0][56] ) );
  XOR U1237 ( .A(key[57]), .B(\w0[0][57] ), .Z(\w1[0][57] ) );
  XOR U1238 ( .A(key[58]), .B(\w0[0][58] ), .Z(\w1[0][58] ) );
  XOR U1239 ( .A(key[59]), .B(\w0[0][59] ), .Z(\w1[0][59] ) );
  XOR U1240 ( .A(key[5]), .B(\w0[0][5] ), .Z(\w1[0][5] ) );
  XOR U1241 ( .A(key[60]), .B(\w0[0][60] ), .Z(\w1[0][60] ) );
  XOR U1242 ( .A(key[61]), .B(\w0[0][61] ), .Z(\w1[0][61] ) );
  XOR U1243 ( .A(key[62]), .B(\w0[0][62] ), .Z(\w1[0][62] ) );
  XOR U1244 ( .A(key[63]), .B(\w0[0][63] ), .Z(\w1[0][63] ) );
  XOR U1245 ( .A(key[64]), .B(\w0[0][64] ), .Z(\w1[0][64] ) );
  XOR U1246 ( .A(key[65]), .B(\w0[0][65] ), .Z(\w1[0][65] ) );
  XOR U1247 ( .A(key[66]), .B(\w0[0][66] ), .Z(\w1[0][66] ) );
  XOR U1248 ( .A(key[67]), .B(\w0[0][67] ), .Z(\w1[0][67] ) );
  XOR U1249 ( .A(key[68]), .B(\w0[0][68] ), .Z(\w1[0][68] ) );
  XOR U1250 ( .A(key[69]), .B(\w0[0][69] ), .Z(\w1[0][69] ) );
  XOR U1251 ( .A(key[6]), .B(\w0[0][6] ), .Z(\w1[0][6] ) );
  XOR U1252 ( .A(key[70]), .B(\w0[0][70] ), .Z(\w1[0][70] ) );
  XOR U1253 ( .A(key[71]), .B(\w0[0][71] ), .Z(\w1[0][71] ) );
  XOR U1254 ( .A(key[72]), .B(\w0[0][72] ), .Z(\w1[0][72] ) );
  XOR U1255 ( .A(key[73]), .B(\w0[0][73] ), .Z(\w1[0][73] ) );
  XOR U1256 ( .A(key[74]), .B(\w0[0][74] ), .Z(\w1[0][74] ) );
  XOR U1257 ( .A(key[75]), .B(\w0[0][75] ), .Z(\w1[0][75] ) );
  XOR U1258 ( .A(key[76]), .B(\w0[0][76] ), .Z(\w1[0][76] ) );
  XOR U1259 ( .A(key[77]), .B(\w0[0][77] ), .Z(\w1[0][77] ) );
  XOR U1260 ( .A(key[78]), .B(\w0[0][78] ), .Z(\w1[0][78] ) );
  XOR U1261 ( .A(key[79]), .B(\w0[0][79] ), .Z(\w1[0][79] ) );
  XOR U1262 ( .A(key[7]), .B(\w0[0][7] ), .Z(\w1[0][7] ) );
  XOR U1263 ( .A(key[80]), .B(\w0[0][80] ), .Z(\w1[0][80] ) );
  XOR U1264 ( .A(key[81]), .B(\w0[0][81] ), .Z(\w1[0][81] ) );
  XOR U1265 ( .A(key[82]), .B(\w0[0][82] ), .Z(\w1[0][82] ) );
  XOR U1266 ( .A(key[83]), .B(\w0[0][83] ), .Z(\w1[0][83] ) );
  XOR U1267 ( .A(key[84]), .B(\w0[0][84] ), .Z(\w1[0][84] ) );
  XOR U1268 ( .A(key[85]), .B(\w0[0][85] ), .Z(\w1[0][85] ) );
  XOR U1269 ( .A(key[86]), .B(\w0[0][86] ), .Z(\w1[0][86] ) );
  XOR U1270 ( .A(key[87]), .B(\w0[0][87] ), .Z(\w1[0][87] ) );
  XOR U1271 ( .A(key[88]), .B(\w0[0][88] ), .Z(\w1[0][88] ) );
  XOR U1272 ( .A(key[89]), .B(\w0[0][89] ), .Z(\w1[0][89] ) );
  XOR U1273 ( .A(key[8]), .B(\w0[0][8] ), .Z(\w1[0][8] ) );
  XOR U1274 ( .A(key[90]), .B(\w0[0][90] ), .Z(\w1[0][90] ) );
  XOR U1275 ( .A(key[91]), .B(\w0[0][91] ), .Z(\w1[0][91] ) );
  XOR U1276 ( .A(key[92]), .B(\w0[0][92] ), .Z(\w1[0][92] ) );
  XOR U1277 ( .A(key[93]), .B(\w0[0][93] ), .Z(\w1[0][93] ) );
  XOR U1278 ( .A(key[94]), .B(\w0[0][94] ), .Z(\w1[0][94] ) );
  XOR U1279 ( .A(key[95]), .B(\w0[0][95] ), .Z(\w1[0][95] ) );
  XOR U1280 ( .A(key[96]), .B(\w0[0][96] ), .Z(\w1[0][96] ) );
  XOR U1281 ( .A(key[97]), .B(\w0[0][97] ), .Z(\w1[0][97] ) );
  XOR U1282 ( .A(key[98]), .B(\w0[0][98] ), .Z(\w1[0][98] ) );
  XOR U1283 ( .A(key[99]), .B(\w0[0][99] ), .Z(\w1[0][99] ) );
  XOR U1284 ( .A(key[9]), .B(\w0[0][9] ), .Z(\w1[0][9] ) );
endmodule

