
module compare_N16384_CC64 ( clk, rst, x, y, g, e );
  input [255:0] x;
  input [255:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  XOR U10 ( .A(x[1]), .B(n1090), .Z(n8) );
  NANDN U11 ( .A(y[1]), .B(n8), .Z(n9) );
  ANDN U12 ( .B(n9), .A(n1091), .Z(n10) );
  NAND U13 ( .A(n1090), .B(x[1]), .Z(n11) );
  AND U14 ( .A(n10), .B(n11), .Z(n12) );
  NANDN U15 ( .A(y[3]), .B(x[3]), .Z(n13) );
  NANDN U16 ( .A(n12), .B(n1092), .Z(n14) );
  NAND U17 ( .A(n13), .B(n14), .Z(n15) );
  OR U18 ( .A(n1093), .B(n15), .Z(n16) );
  ANDN U19 ( .B(n16), .A(n1089), .Z(n17) );
  NOR U20 ( .A(n1094), .B(n17), .Z(n18) );
  NANDN U21 ( .A(y[5]), .B(x[5]), .Z(n19) );
  NAND U22 ( .A(n18), .B(n19), .Z(n1095) );
  OR U23 ( .A(n1109), .B(n1110), .Z(n20) );
  AND U24 ( .A(n1111), .B(n20), .Z(n21) );
  NOR U25 ( .A(n1112), .B(n21), .Z(n22) );
  NANDN U26 ( .A(y[25]), .B(x[25]), .Z(n23) );
  NAND U27 ( .A(n22), .B(n23), .Z(n24) );
  NANDN U28 ( .A(n1081), .B(n24), .Z(n25) );
  NANDN U29 ( .A(y[27]), .B(x[27]), .Z(n26) );
  NAND U30 ( .A(n25), .B(n26), .Z(n27) );
  OR U31 ( .A(n1113), .B(n27), .Z(n28) );
  ANDN U32 ( .B(n28), .A(n1080), .Z(n29) );
  NOR U33 ( .A(n1114), .B(n29), .Z(n30) );
  NANDN U34 ( .A(y[29]), .B(x[29]), .Z(n31) );
  AND U35 ( .A(n30), .B(n31), .Z(n32) );
  OR U36 ( .A(n1079), .B(n32), .Z(n33) );
  NANDN U37 ( .A(y[31]), .B(x[31]), .Z(n34) );
  AND U38 ( .A(n33), .B(n34), .Z(n35) );
  NANDN U39 ( .A(n1115), .B(n35), .Z(n1116) );
  OR U40 ( .A(n1130), .B(n1131), .Z(n36) );
  ANDN U41 ( .B(n36), .A(n1072), .Z(n37) );
  NOR U42 ( .A(n1132), .B(n37), .Z(n38) );
  NANDN U43 ( .A(y[51]), .B(x[51]), .Z(n39) );
  NAND U44 ( .A(n38), .B(n39), .Z(n40) );
  NANDN U45 ( .A(n1071), .B(n40), .Z(n41) );
  NANDN U46 ( .A(y[53]), .B(x[53]), .Z(n42) );
  NAND U47 ( .A(n41), .B(n42), .Z(n43) );
  OR U48 ( .A(n1133), .B(n43), .Z(n44) );
  ANDN U49 ( .B(n44), .A(n1070), .Z(n45) );
  NOR U50 ( .A(n1134), .B(n45), .Z(n46) );
  NANDN U51 ( .A(y[55]), .B(x[55]), .Z(n47) );
  AND U52 ( .A(n46), .B(n47), .Z(n48) );
  NANDN U53 ( .A(n48), .B(n1135), .Z(n49) );
  NANDN U54 ( .A(y[57]), .B(x[57]), .Z(n50) );
  AND U55 ( .A(n49), .B(n50), .Z(n51) );
  NANDN U56 ( .A(n1136), .B(n51), .Z(n1137) );
  OR U57 ( .A(n1151), .B(n1152), .Z(n52) );
  ANDN U58 ( .B(n52), .A(n1062), .Z(n53) );
  NOR U59 ( .A(n1153), .B(n53), .Z(n54) );
  NANDN U60 ( .A(y[77]), .B(x[77]), .Z(n55) );
  NAND U61 ( .A(n54), .B(n55), .Z(n56) );
  NANDN U62 ( .A(n1061), .B(n56), .Z(n57) );
  NANDN U63 ( .A(y[79]), .B(x[79]), .Z(n58) );
  NAND U64 ( .A(n57), .B(n58), .Z(n59) );
  OR U65 ( .A(n1154), .B(n59), .Z(n60) );
  AND U66 ( .A(n1155), .B(n60), .Z(n61) );
  NOR U67 ( .A(n1156), .B(n61), .Z(n62) );
  NANDN U68 ( .A(y[81]), .B(x[81]), .Z(n63) );
  AND U69 ( .A(n62), .B(n63), .Z(n64) );
  OR U70 ( .A(n1060), .B(n64), .Z(n65) );
  NANDN U71 ( .A(y[83]), .B(x[83]), .Z(n66) );
  AND U72 ( .A(n65), .B(n66), .Z(n67) );
  NANDN U73 ( .A(n1157), .B(n67), .Z(n1158) );
  OR U74 ( .A(n1172), .B(n1173), .Z(n68) );
  ANDN U75 ( .B(n68), .A(n1052), .Z(n69) );
  NOR U76 ( .A(n1174), .B(n69), .Z(n70) );
  NANDN U77 ( .A(y[103]), .B(x[103]), .Z(n71) );
  AND U78 ( .A(n70), .B(n71), .Z(n72) );
  NANDN U79 ( .A(y[105]), .B(x[105]), .Z(n73) );
  NANDN U80 ( .A(n72), .B(n1175), .Z(n74) );
  NAND U81 ( .A(n73), .B(n74), .Z(n75) );
  OR U82 ( .A(n1176), .B(n75), .Z(n76) );
  ANDN U83 ( .B(n76), .A(n1051), .Z(n77) );
  NOR U84 ( .A(n1177), .B(n77), .Z(n78) );
  NANDN U85 ( .A(y[107]), .B(x[107]), .Z(n79) );
  AND U86 ( .A(n78), .B(n79), .Z(n80) );
  OR U87 ( .A(n1050), .B(n80), .Z(n81) );
  NANDN U88 ( .A(y[109]), .B(x[109]), .Z(n82) );
  AND U89 ( .A(n81), .B(n82), .Z(n83) );
  NANDN U90 ( .A(n1178), .B(n83), .Z(n1179) );
  OR U91 ( .A(n1193), .B(n1194), .Z(n84) );
  NAND U92 ( .A(n1195), .B(n84), .Z(n85) );
  ANDN U93 ( .B(n85), .A(n1196), .Z(n86) );
  NANDN U94 ( .A(y[129]), .B(x[129]), .Z(n87) );
  NAND U95 ( .A(n86), .B(n87), .Z(n88) );
  NANDN U96 ( .A(n1042), .B(n88), .Z(n89) );
  ANDN U97 ( .B(n89), .A(n1197), .Z(n90) );
  NANDN U98 ( .A(y[131]), .B(x[131]), .Z(n91) );
  AND U99 ( .A(n90), .B(n91), .Z(n92) );
  OR U100 ( .A(n1041), .B(n92), .Z(n93) );
  ANDN U101 ( .B(n93), .A(n1198), .Z(n94) );
  NANDN U102 ( .A(y[133]), .B(x[133]), .Z(n95) );
  NAND U103 ( .A(n94), .B(n95), .Z(n96) );
  ANDN U104 ( .B(n96), .A(n1040), .Z(n97) );
  NOR U105 ( .A(n1199), .B(n97), .Z(n98) );
  NANDN U106 ( .A(y[135]), .B(x[135]), .Z(n99) );
  NAND U107 ( .A(n98), .B(n99), .Z(n1200) );
  OR U108 ( .A(n1214), .B(n1215), .Z(n100) );
  NANDN U109 ( .A(n1033), .B(n100), .Z(n101) );
  ANDN U110 ( .B(n101), .A(n1216), .Z(n102) );
  NANDN U111 ( .A(y[155]), .B(x[155]), .Z(n103) );
  NAND U112 ( .A(n102), .B(n103), .Z(n104) );
  NANDN U113 ( .A(n1032), .B(n104), .Z(n105) );
  ANDN U114 ( .B(n105), .A(n1217), .Z(n106) );
  NANDN U115 ( .A(y[157]), .B(x[157]), .Z(n107) );
  AND U116 ( .A(n106), .B(n107), .Z(n108) );
  OR U117 ( .A(n1031), .B(n108), .Z(n109) );
  ANDN U118 ( .B(n109), .A(n1218), .Z(n110) );
  NANDN U119 ( .A(y[159]), .B(x[159]), .Z(n111) );
  NAND U120 ( .A(n110), .B(n111), .Z(n112) );
  AND U121 ( .A(n1219), .B(n112), .Z(n113) );
  NOR U122 ( .A(n1220), .B(n113), .Z(n114) );
  NANDN U123 ( .A(y[161]), .B(x[161]), .Z(n115) );
  NAND U124 ( .A(n114), .B(n115), .Z(n1221) );
  OR U125 ( .A(n1235), .B(n1236), .Z(n116) );
  NANDN U126 ( .A(n1023), .B(n116), .Z(n117) );
  ANDN U127 ( .B(n117), .A(n1237), .Z(n118) );
  NANDN U128 ( .A(y[181]), .B(x[181]), .Z(n119) );
  NAND U129 ( .A(n118), .B(n119), .Z(n120) );
  NANDN U130 ( .A(n1022), .B(n120), .Z(n121) );
  ANDN U131 ( .B(n121), .A(n1238), .Z(n122) );
  NANDN U132 ( .A(y[183]), .B(x[183]), .Z(n123) );
  AND U133 ( .A(n122), .B(n123), .Z(n124) );
  NANDN U134 ( .A(n124), .B(n1239), .Z(n125) );
  ANDN U135 ( .B(n125), .A(n1240), .Z(n126) );
  NANDN U136 ( .A(y[185]), .B(x[185]), .Z(n127) );
  NAND U137 ( .A(n126), .B(n127), .Z(n128) );
  ANDN U138 ( .B(n128), .A(n1021), .Z(n129) );
  NOR U139 ( .A(n1241), .B(n129), .Z(n130) );
  NANDN U140 ( .A(y[187]), .B(x[187]), .Z(n131) );
  NAND U141 ( .A(n130), .B(n131), .Z(n1242) );
  OR U142 ( .A(n1256), .B(n1257), .Z(n132) );
  NANDN U143 ( .A(n1013), .B(n132), .Z(n133) );
  ANDN U144 ( .B(n133), .A(n1258), .Z(n134) );
  NANDN U145 ( .A(y[207]), .B(x[207]), .Z(n135) );
  NAND U146 ( .A(n134), .B(n135), .Z(n136) );
  NAND U147 ( .A(n1259), .B(n136), .Z(n137) );
  ANDN U148 ( .B(n137), .A(n1260), .Z(n138) );
  NANDN U149 ( .A(y[209]), .B(x[209]), .Z(n139) );
  AND U150 ( .A(n138), .B(n139), .Z(n140) );
  OR U151 ( .A(n1012), .B(n140), .Z(n141) );
  ANDN U152 ( .B(n141), .A(n1261), .Z(n142) );
  NANDN U153 ( .A(y[211]), .B(x[211]), .Z(n143) );
  NAND U154 ( .A(n142), .B(n143), .Z(n144) );
  ANDN U155 ( .B(n144), .A(n1011), .Z(n145) );
  NOR U156 ( .A(n1262), .B(n145), .Z(n146) );
  NANDN U157 ( .A(y[213]), .B(x[213]), .Z(n147) );
  NAND U158 ( .A(n146), .B(n147), .Z(n1263) );
  OR U159 ( .A(n1277), .B(n1278), .Z(n148) );
  NAND U160 ( .A(n1279), .B(n148), .Z(n149) );
  ANDN U161 ( .B(n149), .A(n1280), .Z(n150) );
  NANDN U162 ( .A(y[233]), .B(x[233]), .Z(n151) );
  NAND U163 ( .A(n150), .B(n151), .Z(n152) );
  NANDN U164 ( .A(n1003), .B(n152), .Z(n153) );
  ANDN U165 ( .B(n153), .A(n1281), .Z(n154) );
  NANDN U166 ( .A(y[235]), .B(x[235]), .Z(n155) );
  AND U167 ( .A(n154), .B(n155), .Z(n156) );
  OR U168 ( .A(n1002), .B(n156), .Z(n157) );
  ANDN U169 ( .B(n157), .A(n1282), .Z(n158) );
  NANDN U170 ( .A(y[237]), .B(x[237]), .Z(n159) );
  NAND U171 ( .A(n158), .B(n159), .Z(n160) );
  ANDN U172 ( .B(n160), .A(n1001), .Z(n161) );
  NOR U173 ( .A(n1283), .B(n161), .Z(n162) );
  NANDN U174 ( .A(y[239]), .B(x[239]), .Z(n163) );
  NAND U175 ( .A(n162), .B(n163), .Z(n1284) );
  NAND U176 ( .A(n1096), .B(n1095), .Z(n164) );
  NANDN U177 ( .A(y[7]), .B(x[7]), .Z(n165) );
  NAND U178 ( .A(n164), .B(n165), .Z(n166) );
  OR U179 ( .A(n1097), .B(n166), .Z(n167) );
  AND U180 ( .A(n1098), .B(n167), .Z(n168) );
  NOR U181 ( .A(n1099), .B(n168), .Z(n169) );
  NANDN U182 ( .A(y[9]), .B(x[9]), .Z(n170) );
  NAND U183 ( .A(n169), .B(n170), .Z(n171) );
  NANDN U184 ( .A(n1087), .B(n171), .Z(n172) );
  NANDN U185 ( .A(y[11]), .B(x[11]), .Z(n173) );
  NAND U186 ( .A(n172), .B(n173), .Z(n174) );
  OR U187 ( .A(n1100), .B(n174), .Z(n175) );
  ANDN U188 ( .B(n175), .A(n1086), .Z(n176) );
  NOR U189 ( .A(n1101), .B(n176), .Z(n177) );
  NANDN U190 ( .A(y[13]), .B(x[13]), .Z(n178) );
  NAND U191 ( .A(n177), .B(n178), .Z(n179) );
  NANDN U192 ( .A(n1085), .B(n179), .Z(n1102) );
  NAND U193 ( .A(n1117), .B(n1116), .Z(n180) );
  NANDN U194 ( .A(y[33]), .B(x[33]), .Z(n181) );
  NAND U195 ( .A(n180), .B(n181), .Z(n182) );
  OR U196 ( .A(n1118), .B(n182), .Z(n183) );
  ANDN U197 ( .B(n183), .A(n1078), .Z(n184) );
  NOR U198 ( .A(n1119), .B(n184), .Z(n185) );
  NANDN U199 ( .A(y[35]), .B(x[35]), .Z(n186) );
  NAND U200 ( .A(n185), .B(n186), .Z(n187) );
  NANDN U201 ( .A(n1077), .B(n187), .Z(n188) );
  NANDN U202 ( .A(y[37]), .B(x[37]), .Z(n189) );
  NAND U203 ( .A(n188), .B(n189), .Z(n190) );
  OR U204 ( .A(n1120), .B(n190), .Z(n191) );
  ANDN U205 ( .B(n191), .A(n1076), .Z(n192) );
  NOR U206 ( .A(n1121), .B(n192), .Z(n193) );
  NANDN U207 ( .A(y[39]), .B(x[39]), .Z(n194) );
  NAND U208 ( .A(n193), .B(n194), .Z(n195) );
  NAND U209 ( .A(n1122), .B(n195), .Z(n1123) );
  NAND U210 ( .A(n1138), .B(n1137), .Z(n196) );
  NANDN U211 ( .A(y[59]), .B(x[59]), .Z(n197) );
  NAND U212 ( .A(n196), .B(n197), .Z(n198) );
  OR U213 ( .A(n1139), .B(n198), .Z(n199) );
  ANDN U214 ( .B(n199), .A(n1068), .Z(n200) );
  NOR U215 ( .A(n1140), .B(n200), .Z(n201) );
  NANDN U216 ( .A(y[61]), .B(x[61]), .Z(n202) );
  NAND U217 ( .A(n201), .B(n202), .Z(n203) );
  NANDN U218 ( .A(n1067), .B(n203), .Z(n204) );
  NANDN U219 ( .A(y[63]), .B(x[63]), .Z(n205) );
  NAND U220 ( .A(n204), .B(n205), .Z(n206) );
  OR U221 ( .A(n1141), .B(n206), .Z(n207) );
  AND U222 ( .A(n1142), .B(n207), .Z(n208) );
  NOR U223 ( .A(n1143), .B(n208), .Z(n209) );
  NANDN U224 ( .A(y[65]), .B(x[65]), .Z(n210) );
  NAND U225 ( .A(n209), .B(n210), .Z(n211) );
  NANDN U226 ( .A(n1066), .B(n211), .Z(n1144) );
  NAND U227 ( .A(n1159), .B(n1158), .Z(n212) );
  NANDN U228 ( .A(y[85]), .B(x[85]), .Z(n213) );
  NAND U229 ( .A(n212), .B(n213), .Z(n214) );
  OR U230 ( .A(n1160), .B(n214), .Z(n215) );
  ANDN U231 ( .B(n215), .A(n1058), .Z(n216) );
  NOR U232 ( .A(n1161), .B(n216), .Z(n217) );
  NANDN U233 ( .A(y[87]), .B(x[87]), .Z(n218) );
  AND U234 ( .A(n217), .B(n218), .Z(n219) );
  NANDN U235 ( .A(y[89]), .B(x[89]), .Z(n220) );
  NANDN U236 ( .A(n219), .B(n1162), .Z(n221) );
  NAND U237 ( .A(n220), .B(n221), .Z(n222) );
  OR U238 ( .A(n1163), .B(n222), .Z(n223) );
  ANDN U239 ( .B(n223), .A(n1057), .Z(n224) );
  NOR U240 ( .A(n1164), .B(n224), .Z(n225) );
  NANDN U241 ( .A(y[91]), .B(x[91]), .Z(n226) );
  NAND U242 ( .A(n225), .B(n226), .Z(n227) );
  NANDN U243 ( .A(n1056), .B(n227), .Z(n1165) );
  NAND U244 ( .A(n1180), .B(n1179), .Z(n228) );
  NANDN U245 ( .A(y[111]), .B(x[111]), .Z(n229) );
  NAND U246 ( .A(n228), .B(n229), .Z(n230) );
  OR U247 ( .A(n1181), .B(n230), .Z(n231) );
  AND U248 ( .A(n1182), .B(n231), .Z(n232) );
  NOR U249 ( .A(n1183), .B(n232), .Z(n233) );
  NANDN U250 ( .A(y[113]), .B(x[113]), .Z(n234) );
  NAND U251 ( .A(n233), .B(n234), .Z(n235) );
  NANDN U252 ( .A(n1048), .B(n235), .Z(n236) );
  NANDN U253 ( .A(y[115]), .B(x[115]), .Z(n237) );
  NAND U254 ( .A(n236), .B(n237), .Z(n238) );
  OR U255 ( .A(n1184), .B(n238), .Z(n239) );
  ANDN U256 ( .B(n239), .A(n1047), .Z(n240) );
  NOR U257 ( .A(n1185), .B(n240), .Z(n241) );
  NANDN U258 ( .A(y[117]), .B(x[117]), .Z(n242) );
  NAND U259 ( .A(n241), .B(n242), .Z(n243) );
  NANDN U260 ( .A(n1046), .B(n243), .Z(n1186) );
  NAND U261 ( .A(n1201), .B(n1200), .Z(n244) );
  ANDN U262 ( .B(n244), .A(n1202), .Z(n245) );
  NANDN U263 ( .A(y[137]), .B(x[137]), .Z(n246) );
  NAND U264 ( .A(n245), .B(n246), .Z(n247) );
  NANDN U265 ( .A(n1039), .B(n247), .Z(n248) );
  ANDN U266 ( .B(n248), .A(n1203), .Z(n249) );
  NANDN U267 ( .A(y[139]), .B(x[139]), .Z(n250) );
  AND U268 ( .A(n249), .B(n250), .Z(n251) );
  OR U269 ( .A(n1038), .B(n251), .Z(n252) );
  ANDN U270 ( .B(n252), .A(n1204), .Z(n253) );
  NANDN U271 ( .A(y[141]), .B(x[141]), .Z(n254) );
  NAND U272 ( .A(n253), .B(n254), .Z(n255) );
  ANDN U273 ( .B(n255), .A(n1037), .Z(n256) );
  NOR U274 ( .A(n1205), .B(n256), .Z(n257) );
  NANDN U275 ( .A(y[143]), .B(x[143]), .Z(n258) );
  NAND U276 ( .A(n257), .B(n258), .Z(n259) );
  NAND U277 ( .A(n1206), .B(n259), .Z(n1207) );
  NAND U278 ( .A(n1221), .B(n1222), .Z(n260) );
  ANDN U279 ( .B(n260), .A(n1223), .Z(n261) );
  NANDN U280 ( .A(y[163]), .B(x[163]), .Z(n262) );
  NAND U281 ( .A(n261), .B(n262), .Z(n263) );
  NANDN U282 ( .A(n1029), .B(n263), .Z(n264) );
  ANDN U283 ( .B(n264), .A(n1224), .Z(n265) );
  NANDN U284 ( .A(y[165]), .B(x[165]), .Z(n266) );
  AND U285 ( .A(n265), .B(n266), .Z(n267) );
  OR U286 ( .A(n1028), .B(n267), .Z(n268) );
  ANDN U287 ( .B(n268), .A(n1225), .Z(n269) );
  NANDN U288 ( .A(y[167]), .B(x[167]), .Z(n270) );
  NAND U289 ( .A(n269), .B(n270), .Z(n271) );
  AND U290 ( .A(n1226), .B(n271), .Z(n272) );
  NOR U291 ( .A(n1227), .B(n272), .Z(n273) );
  NANDN U292 ( .A(y[169]), .B(x[169]), .Z(n274) );
  NAND U293 ( .A(n273), .B(n274), .Z(n275) );
  NANDN U294 ( .A(n1027), .B(n275), .Z(n1228) );
  NAND U295 ( .A(n1242), .B(n1243), .Z(n276) );
  ANDN U296 ( .B(n276), .A(n1244), .Z(n277) );
  NANDN U297 ( .A(y[189]), .B(x[189]), .Z(n278) );
  NAND U298 ( .A(n277), .B(n278), .Z(n279) );
  NANDN U299 ( .A(n1019), .B(n279), .Z(n280) );
  ANDN U300 ( .B(n280), .A(n1245), .Z(n281) );
  NANDN U301 ( .A(y[191]), .B(x[191]), .Z(n282) );
  AND U302 ( .A(n281), .B(n282), .Z(n283) );
  NANDN U303 ( .A(n283), .B(n1246), .Z(n284) );
  ANDN U304 ( .B(n284), .A(n1247), .Z(n285) );
  NANDN U305 ( .A(y[193]), .B(x[193]), .Z(n286) );
  NAND U306 ( .A(n285), .B(n286), .Z(n287) );
  ANDN U307 ( .B(n287), .A(n1018), .Z(n288) );
  NOR U308 ( .A(n1248), .B(n288), .Z(n289) );
  NANDN U309 ( .A(y[195]), .B(x[195]), .Z(n290) );
  NAND U310 ( .A(n289), .B(n290), .Z(n291) );
  NANDN U311 ( .A(n1017), .B(n291), .Z(n1249) );
  NAND U312 ( .A(n1263), .B(n1264), .Z(n292) );
  ANDN U313 ( .B(n292), .A(n1265), .Z(n293) );
  NANDN U314 ( .A(y[215]), .B(x[215]), .Z(n294) );
  NAND U315 ( .A(n293), .B(n294), .Z(n295) );
  NAND U316 ( .A(n1266), .B(n295), .Z(n296) );
  ANDN U317 ( .B(n296), .A(n1267), .Z(n297) );
  NANDN U318 ( .A(y[217]), .B(x[217]), .Z(n298) );
  AND U319 ( .A(n297), .B(n298), .Z(n299) );
  OR U320 ( .A(n1009), .B(n299), .Z(n300) );
  ANDN U321 ( .B(n300), .A(n1268), .Z(n301) );
  NANDN U322 ( .A(y[219]), .B(x[219]), .Z(n302) );
  NAND U323 ( .A(n301), .B(n302), .Z(n303) );
  ANDN U324 ( .B(n303), .A(n1008), .Z(n304) );
  NOR U325 ( .A(n1269), .B(n304), .Z(n305) );
  NANDN U326 ( .A(y[221]), .B(x[221]), .Z(n306) );
  NAND U327 ( .A(n305), .B(n306), .Z(n307) );
  NANDN U328 ( .A(n1007), .B(n307), .Z(n1270) );
  NAND U329 ( .A(n1285), .B(n1284), .Z(n308) );
  ANDN U330 ( .B(n308), .A(n1286), .Z(n309) );
  NANDN U331 ( .A(y[241]), .B(x[241]), .Z(n310) );
  NAND U332 ( .A(n309), .B(n310), .Z(n311) );
  NANDN U333 ( .A(n1000), .B(n311), .Z(n312) );
  ANDN U334 ( .B(n312), .A(n1287), .Z(n313) );
  NANDN U335 ( .A(y[243]), .B(x[243]), .Z(n314) );
  AND U336 ( .A(n313), .B(n314), .Z(n315) );
  OR U337 ( .A(n999), .B(n315), .Z(n316) );
  ANDN U338 ( .B(n316), .A(n1288), .Z(n317) );
  NANDN U339 ( .A(y[245]), .B(x[245]), .Z(n318) );
  NAND U340 ( .A(n317), .B(n318), .Z(n319) );
  ANDN U341 ( .B(n319), .A(n998), .Z(n320) );
  NOR U342 ( .A(n1289), .B(n320), .Z(n321) );
  NANDN U343 ( .A(y[247]), .B(x[247]), .Z(n322) );
  NAND U344 ( .A(n321), .B(n322), .Z(n323) );
  NAND U345 ( .A(n1290), .B(n323), .Z(n1291) );
  NOR U346 ( .A(n1104), .B(n1103), .Z(n324) );
  NAND U347 ( .A(n1102), .B(n324), .Z(n325) );
  AND U348 ( .A(n1105), .B(n325), .Z(n326) );
  NOR U349 ( .A(n1106), .B(n326), .Z(n327) );
  NANDN U350 ( .A(y[17]), .B(x[17]), .Z(n328) );
  NAND U351 ( .A(n327), .B(n328), .Z(n329) );
  NANDN U352 ( .A(n1084), .B(n329), .Z(n330) );
  NANDN U353 ( .A(y[19]), .B(x[19]), .Z(n331) );
  NAND U354 ( .A(n330), .B(n331), .Z(n332) );
  OR U355 ( .A(n1107), .B(n332), .Z(n333) );
  ANDN U356 ( .B(n333), .A(n1083), .Z(n334) );
  NOR U357 ( .A(n1108), .B(n334), .Z(n335) );
  NANDN U358 ( .A(y[21]), .B(x[21]), .Z(n336) );
  NAND U359 ( .A(n335), .B(n336), .Z(n337) );
  NANDN U360 ( .A(n1082), .B(n337), .Z(n338) );
  NANDN U361 ( .A(y[23]), .B(x[23]), .Z(n339) );
  NAND U362 ( .A(n338), .B(n339), .Z(n1110) );
  NOR U363 ( .A(n1125), .B(n1124), .Z(n340) );
  NAND U364 ( .A(n1123), .B(n340), .Z(n341) );
  ANDN U365 ( .B(n341), .A(n1075), .Z(n342) );
  NOR U366 ( .A(n1126), .B(n342), .Z(n343) );
  NANDN U367 ( .A(y[43]), .B(x[43]), .Z(n344) );
  NAND U368 ( .A(n343), .B(n344), .Z(n345) );
  NANDN U369 ( .A(n1074), .B(n345), .Z(n346) );
  NANDN U370 ( .A(y[45]), .B(x[45]), .Z(n347) );
  NAND U371 ( .A(n346), .B(n347), .Z(n348) );
  OR U372 ( .A(n1127), .B(n348), .Z(n349) );
  ANDN U373 ( .B(n349), .A(n1073), .Z(n350) );
  NOR U374 ( .A(n1128), .B(n350), .Z(n351) );
  NANDN U375 ( .A(y[47]), .B(x[47]), .Z(n352) );
  AND U376 ( .A(n351), .B(n352), .Z(n353) );
  NANDN U377 ( .A(y[49]), .B(x[49]), .Z(n354) );
  NANDN U378 ( .A(n353), .B(n1129), .Z(n355) );
  NAND U379 ( .A(n354), .B(n355), .Z(n1131) );
  NOR U380 ( .A(n1146), .B(n1145), .Z(n356) );
  NAND U381 ( .A(n1144), .B(n356), .Z(n357) );
  ANDN U382 ( .B(n357), .A(n1065), .Z(n358) );
  NOR U383 ( .A(n1147), .B(n358), .Z(n359) );
  NANDN U384 ( .A(y[69]), .B(x[69]), .Z(n360) );
  NAND U385 ( .A(n359), .B(n360), .Z(n361) );
  NANDN U386 ( .A(n1064), .B(n361), .Z(n362) );
  NANDN U387 ( .A(y[71]), .B(x[71]), .Z(n363) );
  NAND U388 ( .A(n362), .B(n363), .Z(n364) );
  OR U389 ( .A(n1148), .B(n364), .Z(n365) );
  AND U390 ( .A(n1149), .B(n365), .Z(n366) );
  NOR U391 ( .A(n1150), .B(n366), .Z(n367) );
  NANDN U392 ( .A(y[73]), .B(x[73]), .Z(n368) );
  NAND U393 ( .A(n367), .B(n368), .Z(n369) );
  NANDN U394 ( .A(n1063), .B(n369), .Z(n370) );
  NANDN U395 ( .A(y[75]), .B(x[75]), .Z(n371) );
  NAND U396 ( .A(n370), .B(n371), .Z(n1152) );
  NOR U397 ( .A(n1167), .B(n1166), .Z(n372) );
  NAND U398 ( .A(n1165), .B(n372), .Z(n373) );
  NANDN U399 ( .A(n1055), .B(n373), .Z(n374) );
  ANDN U400 ( .B(n374), .A(n1168), .Z(n375) );
  NANDN U401 ( .A(y[95]), .B(x[95]), .Z(n376) );
  AND U402 ( .A(n375), .B(n376), .Z(n377) );
  NANDN U403 ( .A(y[97]), .B(x[97]), .Z(n378) );
  NANDN U404 ( .A(n377), .B(n1169), .Z(n379) );
  NAND U405 ( .A(n378), .B(n379), .Z(n380) );
  OR U406 ( .A(n1170), .B(n380), .Z(n381) );
  ANDN U407 ( .B(n381), .A(n1054), .Z(n382) );
  NOR U408 ( .A(n1171), .B(n382), .Z(n383) );
  NANDN U409 ( .A(y[99]), .B(x[99]), .Z(n384) );
  NAND U410 ( .A(n383), .B(n384), .Z(n385) );
  NANDN U411 ( .A(n1053), .B(n385), .Z(n386) );
  NANDN U412 ( .A(y[101]), .B(x[101]), .Z(n387) );
  NAND U413 ( .A(n386), .B(n387), .Z(n1173) );
  NOR U414 ( .A(n1188), .B(n1187), .Z(n388) );
  NAND U415 ( .A(n1186), .B(n388), .Z(n389) );
  AND U416 ( .A(n1189), .B(n389), .Z(n390) );
  NOR U417 ( .A(n1190), .B(n390), .Z(n391) );
  NANDN U418 ( .A(y[121]), .B(x[121]), .Z(n392) );
  NAND U419 ( .A(n391), .B(n392), .Z(n393) );
  NANDN U420 ( .A(n1045), .B(n393), .Z(n394) );
  NANDN U421 ( .A(y[123]), .B(x[123]), .Z(n395) );
  NAND U422 ( .A(n394), .B(n395), .Z(n396) );
  OR U423 ( .A(n1191), .B(n396), .Z(n397) );
  ANDN U424 ( .B(n397), .A(n1044), .Z(n398) );
  NOR U425 ( .A(n1192), .B(n398), .Z(n399) );
  NANDN U426 ( .A(y[125]), .B(x[125]), .Z(n400) );
  NAND U427 ( .A(n399), .B(n400), .Z(n401) );
  NANDN U428 ( .A(n1043), .B(n401), .Z(n402) );
  NANDN U429 ( .A(y[127]), .B(x[127]), .Z(n403) );
  NAND U430 ( .A(n402), .B(n403), .Z(n1194) );
  ANDN U431 ( .B(n1207), .A(n1208), .Z(n404) );
  NANDN U432 ( .A(y[145]), .B(x[145]), .Z(n405) );
  AND U433 ( .A(n404), .B(n405), .Z(n406) );
  OR U434 ( .A(n1036), .B(n406), .Z(n407) );
  ANDN U435 ( .B(n407), .A(n1209), .Z(n408) );
  NANDN U436 ( .A(y[147]), .B(x[147]), .Z(n409) );
  NAND U437 ( .A(n408), .B(n409), .Z(n410) );
  NANDN U438 ( .A(n1035), .B(n410), .Z(n411) );
  ANDN U439 ( .B(n411), .A(n1210), .Z(n412) );
  NANDN U440 ( .A(y[149]), .B(x[149]), .Z(n413) );
  AND U441 ( .A(n412), .B(n413), .Z(n414) );
  OR U442 ( .A(n1034), .B(n414), .Z(n415) );
  ANDN U443 ( .B(n415), .A(n1211), .Z(n416) );
  NANDN U444 ( .A(y[151]), .B(x[151]), .Z(n417) );
  NAND U445 ( .A(n416), .B(n417), .Z(n418) );
  NAND U446 ( .A(n1212), .B(n418), .Z(n419) );
  NANDN U447 ( .A(n1213), .B(n419), .Z(n1215) );
  ANDN U448 ( .B(n1228), .A(n1229), .Z(n420) );
  NANDN U449 ( .A(y[171]), .B(x[171]), .Z(n421) );
  AND U450 ( .A(n420), .B(n421), .Z(n422) );
  OR U451 ( .A(n1026), .B(n422), .Z(n423) );
  ANDN U452 ( .B(n423), .A(n1230), .Z(n424) );
  NANDN U453 ( .A(y[173]), .B(x[173]), .Z(n425) );
  NAND U454 ( .A(n424), .B(n425), .Z(n426) );
  NANDN U455 ( .A(n1025), .B(n426), .Z(n427) );
  ANDN U456 ( .B(n427), .A(n1231), .Z(n428) );
  NANDN U457 ( .A(y[175]), .B(x[175]), .Z(n429) );
  AND U458 ( .A(n428), .B(n429), .Z(n430) );
  NANDN U459 ( .A(n430), .B(n1232), .Z(n431) );
  ANDN U460 ( .B(n431), .A(n1233), .Z(n432) );
  NANDN U461 ( .A(y[177]), .B(x[177]), .Z(n433) );
  NAND U462 ( .A(n432), .B(n433), .Z(n434) );
  NANDN U463 ( .A(n1024), .B(n434), .Z(n435) );
  NANDN U464 ( .A(n1234), .B(n435), .Z(n1236) );
  ANDN U465 ( .B(n1249), .A(n1250), .Z(n436) );
  NANDN U466 ( .A(y[197]), .B(x[197]), .Z(n437) );
  AND U467 ( .A(n436), .B(n437), .Z(n438) );
  OR U468 ( .A(n1016), .B(n438), .Z(n439) );
  ANDN U469 ( .B(n439), .A(n1251), .Z(n440) );
  NANDN U470 ( .A(y[199]), .B(x[199]), .Z(n441) );
  NAND U471 ( .A(n440), .B(n441), .Z(n442) );
  NAND U472 ( .A(n1252), .B(n442), .Z(n443) );
  ANDN U473 ( .B(n443), .A(n1253), .Z(n444) );
  NANDN U474 ( .A(y[201]), .B(x[201]), .Z(n445) );
  AND U475 ( .A(n444), .B(n445), .Z(n446) );
  OR U476 ( .A(n1015), .B(n446), .Z(n447) );
  ANDN U477 ( .B(n447), .A(n1254), .Z(n448) );
  NANDN U478 ( .A(y[203]), .B(x[203]), .Z(n449) );
  NAND U479 ( .A(n448), .B(n449), .Z(n450) );
  NANDN U480 ( .A(n1014), .B(n450), .Z(n451) );
  NANDN U481 ( .A(n1255), .B(n451), .Z(n1257) );
  ANDN U482 ( .B(n1270), .A(n1271), .Z(n452) );
  NANDN U483 ( .A(y[223]), .B(x[223]), .Z(n453) );
  AND U484 ( .A(n452), .B(n453), .Z(n454) );
  NANDN U485 ( .A(n454), .B(n1272), .Z(n455) );
  ANDN U486 ( .B(n455), .A(n1273), .Z(n456) );
  NANDN U487 ( .A(y[225]), .B(x[225]), .Z(n457) );
  NAND U488 ( .A(n456), .B(n457), .Z(n458) );
  NANDN U489 ( .A(n1006), .B(n458), .Z(n459) );
  ANDN U490 ( .B(n459), .A(n1274), .Z(n460) );
  NANDN U491 ( .A(y[227]), .B(x[227]), .Z(n461) );
  AND U492 ( .A(n460), .B(n461), .Z(n462) );
  OR U493 ( .A(n1005), .B(n462), .Z(n463) );
  ANDN U494 ( .B(n463), .A(n1275), .Z(n464) );
  NANDN U495 ( .A(y[229]), .B(x[229]), .Z(n465) );
  NAND U496 ( .A(n464), .B(n465), .Z(n466) );
  NANDN U497 ( .A(n1004), .B(n466), .Z(n467) );
  NANDN U498 ( .A(n1276), .B(n467), .Z(n1278) );
  AND U499 ( .A(e), .B(n1296), .Z(n468) );
  NOR U500 ( .A(n1293), .B(n1292), .Z(n469) );
  NAND U501 ( .A(n1291), .B(n469), .Z(n470) );
  ANDN U502 ( .B(n470), .A(n997), .Z(n471) );
  NOR U503 ( .A(n1294), .B(n471), .Z(n472) );
  NANDN U504 ( .A(y[251]), .B(x[251]), .Z(n473) );
  NAND U505 ( .A(n472), .B(n473), .Z(n474) );
  ANDN U506 ( .B(n474), .A(n996), .Z(n475) );
  NOR U507 ( .A(n1295), .B(n475), .Z(n476) );
  NANDN U508 ( .A(y[253]), .B(x[253]), .Z(n477) );
  NAND U509 ( .A(n476), .B(n477), .Z(n478) );
  NANDN U510 ( .A(n995), .B(n478), .Z(n479) );
  NANDN U511 ( .A(y[255]), .B(x[255]), .Z(n480) );
  NAND U512 ( .A(n479), .B(n480), .Z(n481) );
  NAND U513 ( .A(n481), .B(n468), .Z(n482) );
  NANDN U514 ( .A(n468), .B(g), .Z(n483) );
  NAND U515 ( .A(n482), .B(n483), .Z(n4) );
  IV U516 ( .A(ebreg), .Z(e) );
  XNOR U517 ( .A(y[85]), .B(x[85]), .Z(n485) );
  NANDN U518 ( .A(x[84]), .B(y[84]), .Z(n484) );
  NAND U519 ( .A(n485), .B(n484), .Z(n1059) );
  XNOR U520 ( .A(y[81]), .B(x[81]), .Z(n487) );
  NANDN U521 ( .A(x[80]), .B(y[80]), .Z(n486) );
  AND U522 ( .A(n487), .B(n486), .Z(n1155) );
  XNOR U523 ( .A(y[83]), .B(x[83]), .Z(n489) );
  NANDN U524 ( .A(x[82]), .B(y[82]), .Z(n488) );
  NAND U525 ( .A(n489), .B(n488), .Z(n1060) );
  ANDN U526 ( .B(n1155), .A(n1060), .Z(n492) );
  XNOR U527 ( .A(y[87]), .B(x[87]), .Z(n491) );
  NANDN U528 ( .A(x[86]), .B(y[86]), .Z(n490) );
  NAND U529 ( .A(n491), .B(n490), .Z(n1058) );
  ANDN U530 ( .B(n492), .A(n1058), .Z(n493) );
  NANDN U531 ( .A(n1059), .B(n493), .Z(n529) );
  XNOR U532 ( .A(y[69]), .B(x[69]), .Z(n495) );
  NANDN U533 ( .A(x[68]), .B(y[68]), .Z(n494) );
  NAND U534 ( .A(n495), .B(n494), .Z(n1065) );
  XNOR U535 ( .A(y[65]), .B(x[65]), .Z(n497) );
  NANDN U536 ( .A(x[64]), .B(y[64]), .Z(n496) );
  AND U537 ( .A(n497), .B(n496), .Z(n1142) );
  XNOR U538 ( .A(y[67]), .B(x[67]), .Z(n499) );
  NANDN U539 ( .A(x[66]), .B(y[66]), .Z(n498) );
  NAND U540 ( .A(n499), .B(n498), .Z(n1066) );
  ANDN U541 ( .B(n1142), .A(n1066), .Z(n502) );
  XNOR U542 ( .A(y[71]), .B(x[71]), .Z(n501) );
  NANDN U543 ( .A(x[70]), .B(y[70]), .Z(n500) );
  NAND U544 ( .A(n501), .B(n500), .Z(n1064) );
  ANDN U545 ( .B(n502), .A(n1064), .Z(n503) );
  NANDN U546 ( .A(n1065), .B(n503), .Z(n515) );
  XNOR U547 ( .A(y[77]), .B(x[77]), .Z(n505) );
  NANDN U548 ( .A(x[76]), .B(y[76]), .Z(n504) );
  NAND U549 ( .A(n505), .B(n504), .Z(n1062) );
  XNOR U550 ( .A(y[73]), .B(x[73]), .Z(n507) );
  NANDN U551 ( .A(x[72]), .B(y[72]), .Z(n506) );
  AND U552 ( .A(n507), .B(n506), .Z(n1149) );
  XNOR U553 ( .A(y[75]), .B(x[75]), .Z(n509) );
  NANDN U554 ( .A(x[74]), .B(y[74]), .Z(n508) );
  NAND U555 ( .A(n509), .B(n508), .Z(n1063) );
  ANDN U556 ( .B(n1149), .A(n1063), .Z(n512) );
  XNOR U557 ( .A(y[79]), .B(x[79]), .Z(n511) );
  NANDN U558 ( .A(x[78]), .B(y[78]), .Z(n510) );
  NAND U559 ( .A(n511), .B(n510), .Z(n1061) );
  ANDN U560 ( .B(n512), .A(n1061), .Z(n513) );
  NANDN U561 ( .A(n1062), .B(n513), .Z(n514) );
  NOR U562 ( .A(n515), .B(n514), .Z(n527) );
  XNOR U563 ( .A(y[93]), .B(x[93]), .Z(n517) );
  NANDN U564 ( .A(x[92]), .B(y[92]), .Z(n516) );
  NAND U565 ( .A(n517), .B(n516), .Z(n1056) );
  XNOR U566 ( .A(y[89]), .B(x[89]), .Z(n519) );
  NANDN U567 ( .A(x[88]), .B(y[88]), .Z(n518) );
  AND U568 ( .A(n519), .B(n518), .Z(n1162) );
  XNOR U569 ( .A(y[91]), .B(x[91]), .Z(n521) );
  NANDN U570 ( .A(x[90]), .B(y[90]), .Z(n520) );
  NAND U571 ( .A(n521), .B(n520), .Z(n1057) );
  ANDN U572 ( .B(n1162), .A(n1057), .Z(n524) );
  XNOR U573 ( .A(y[95]), .B(x[95]), .Z(n523) );
  NANDN U574 ( .A(x[94]), .B(y[94]), .Z(n522) );
  NAND U575 ( .A(n523), .B(n522), .Z(n1055) );
  ANDN U576 ( .B(n524), .A(n1055), .Z(n525) );
  NANDN U577 ( .A(n1056), .B(n525), .Z(n526) );
  ANDN U578 ( .B(n527), .A(n526), .Z(n528) );
  NANDN U579 ( .A(n529), .B(n528), .Z(n674) );
  XNOR U580 ( .A(y[21]), .B(x[21]), .Z(n531) );
  NANDN U581 ( .A(x[20]), .B(y[20]), .Z(n530) );
  NAND U582 ( .A(n531), .B(n530), .Z(n1083) );
  XNOR U583 ( .A(y[17]), .B(x[17]), .Z(n533) );
  NANDN U584 ( .A(x[16]), .B(y[16]), .Z(n532) );
  AND U585 ( .A(n533), .B(n532), .Z(n1105) );
  XNOR U586 ( .A(y[19]), .B(x[19]), .Z(n535) );
  NANDN U587 ( .A(x[18]), .B(y[18]), .Z(n534) );
  NAND U588 ( .A(n535), .B(n534), .Z(n1084) );
  ANDN U589 ( .B(n1105), .A(n1084), .Z(n538) );
  XNOR U590 ( .A(y[23]), .B(x[23]), .Z(n537) );
  NANDN U591 ( .A(x[22]), .B(y[22]), .Z(n536) );
  NAND U592 ( .A(n537), .B(n536), .Z(n1082) );
  ANDN U593 ( .B(n538), .A(n1082), .Z(n539) );
  NANDN U594 ( .A(n1083), .B(n539), .Z(n576) );
  XNOR U595 ( .A(y[7]), .B(x[7]), .Z(n541) );
  NANDN U596 ( .A(x[6]), .B(y[6]), .Z(n540) );
  NAND U597 ( .A(n541), .B(n540), .Z(n1088) );
  XNOR U598 ( .A(y[3]), .B(x[3]), .Z(n543) );
  NANDN U599 ( .A(x[2]), .B(y[2]), .Z(n542) );
  AND U600 ( .A(n543), .B(n542), .Z(n1092) );
  XNOR U601 ( .A(y[5]), .B(x[5]), .Z(n545) );
  NANDN U602 ( .A(x[4]), .B(y[4]), .Z(n544) );
  NAND U603 ( .A(n545), .B(n544), .Z(n1089) );
  ANDN U604 ( .B(n1092), .A(n1089), .Z(n549) );
  XNOR U605 ( .A(y[1]), .B(x[1]), .Z(n547) );
  NANDN U606 ( .A(x[0]), .B(y[0]), .Z(n546) );
  NAND U607 ( .A(n547), .B(n546), .Z(n548) );
  ANDN U608 ( .B(n549), .A(n548), .Z(n550) );
  NANDN U609 ( .A(n1088), .B(n550), .Z(n562) );
  XNOR U610 ( .A(y[13]), .B(x[13]), .Z(n552) );
  NANDN U611 ( .A(x[12]), .B(y[12]), .Z(n551) );
  NAND U612 ( .A(n552), .B(n551), .Z(n1086) );
  XNOR U613 ( .A(y[9]), .B(x[9]), .Z(n554) );
  NANDN U614 ( .A(x[8]), .B(y[8]), .Z(n553) );
  AND U615 ( .A(n554), .B(n553), .Z(n1098) );
  XNOR U616 ( .A(y[11]), .B(x[11]), .Z(n556) );
  NANDN U617 ( .A(x[10]), .B(y[10]), .Z(n555) );
  NAND U618 ( .A(n556), .B(n555), .Z(n1087) );
  ANDN U619 ( .B(n1098), .A(n1087), .Z(n559) );
  XNOR U620 ( .A(y[15]), .B(x[15]), .Z(n558) );
  NANDN U621 ( .A(x[14]), .B(y[14]), .Z(n557) );
  NAND U622 ( .A(n558), .B(n557), .Z(n1085) );
  ANDN U623 ( .B(n559), .A(n1085), .Z(n560) );
  NANDN U624 ( .A(n1086), .B(n560), .Z(n561) );
  NOR U625 ( .A(n562), .B(n561), .Z(n574) );
  XNOR U626 ( .A(y[29]), .B(x[29]), .Z(n564) );
  NANDN U627 ( .A(x[28]), .B(y[28]), .Z(n563) );
  NAND U628 ( .A(n564), .B(n563), .Z(n1080) );
  XNOR U629 ( .A(y[25]), .B(x[25]), .Z(n566) );
  NANDN U630 ( .A(x[24]), .B(y[24]), .Z(n565) );
  AND U631 ( .A(n566), .B(n565), .Z(n1111) );
  XNOR U632 ( .A(y[27]), .B(x[27]), .Z(n568) );
  NANDN U633 ( .A(x[26]), .B(y[26]), .Z(n567) );
  NAND U634 ( .A(n568), .B(n567), .Z(n1081) );
  ANDN U635 ( .B(n1111), .A(n1081), .Z(n571) );
  XNOR U636 ( .A(y[31]), .B(x[31]), .Z(n570) );
  NANDN U637 ( .A(x[30]), .B(y[30]), .Z(n569) );
  NAND U638 ( .A(n570), .B(n569), .Z(n1079) );
  ANDN U639 ( .B(n571), .A(n1079), .Z(n572) );
  NANDN U640 ( .A(n1080), .B(n572), .Z(n573) );
  ANDN U641 ( .B(n574), .A(n573), .Z(n575) );
  NANDN U642 ( .A(n576), .B(n575), .Z(n624) );
  XNOR U643 ( .A(y[53]), .B(x[53]), .Z(n578) );
  NANDN U644 ( .A(x[52]), .B(y[52]), .Z(n577) );
  NAND U645 ( .A(n578), .B(n577), .Z(n1071) );
  XNOR U646 ( .A(y[49]), .B(x[49]), .Z(n580) );
  NANDN U647 ( .A(x[48]), .B(y[48]), .Z(n579) );
  AND U648 ( .A(n580), .B(n579), .Z(n1129) );
  XNOR U649 ( .A(y[51]), .B(x[51]), .Z(n582) );
  NANDN U650 ( .A(x[50]), .B(y[50]), .Z(n581) );
  NAND U651 ( .A(n582), .B(n581), .Z(n1072) );
  ANDN U652 ( .B(n1129), .A(n1072), .Z(n585) );
  XNOR U653 ( .A(y[55]), .B(x[55]), .Z(n584) );
  NANDN U654 ( .A(x[54]), .B(y[54]), .Z(n583) );
  NAND U655 ( .A(n584), .B(n583), .Z(n1070) );
  ANDN U656 ( .B(n585), .A(n1070), .Z(n586) );
  NANDN U657 ( .A(n1071), .B(n586), .Z(n622) );
  XNOR U658 ( .A(y[37]), .B(x[37]), .Z(n588) );
  NANDN U659 ( .A(x[36]), .B(y[36]), .Z(n587) );
  NAND U660 ( .A(n588), .B(n587), .Z(n1077) );
  XNOR U661 ( .A(y[33]), .B(x[33]), .Z(n590) );
  NANDN U662 ( .A(x[32]), .B(y[32]), .Z(n589) );
  AND U663 ( .A(n590), .B(n589), .Z(n1117) );
  XNOR U664 ( .A(y[35]), .B(x[35]), .Z(n592) );
  NANDN U665 ( .A(x[34]), .B(y[34]), .Z(n591) );
  NAND U666 ( .A(n592), .B(n591), .Z(n1078) );
  ANDN U667 ( .B(n1117), .A(n1078), .Z(n595) );
  XNOR U668 ( .A(y[39]), .B(x[39]), .Z(n594) );
  NANDN U669 ( .A(x[38]), .B(y[38]), .Z(n593) );
  NAND U670 ( .A(n594), .B(n593), .Z(n1076) );
  ANDN U671 ( .B(n595), .A(n1076), .Z(n596) );
  NANDN U672 ( .A(n1077), .B(n596), .Z(n608) );
  XNOR U673 ( .A(y[45]), .B(x[45]), .Z(n598) );
  NANDN U674 ( .A(x[44]), .B(y[44]), .Z(n597) );
  NAND U675 ( .A(n598), .B(n597), .Z(n1074) );
  XNOR U676 ( .A(y[41]), .B(x[41]), .Z(n600) );
  NANDN U677 ( .A(x[40]), .B(y[40]), .Z(n599) );
  AND U678 ( .A(n600), .B(n599), .Z(n1122) );
  XNOR U679 ( .A(y[43]), .B(x[43]), .Z(n602) );
  NANDN U680 ( .A(x[42]), .B(y[42]), .Z(n601) );
  NAND U681 ( .A(n602), .B(n601), .Z(n1075) );
  ANDN U682 ( .B(n1122), .A(n1075), .Z(n605) );
  XNOR U683 ( .A(y[47]), .B(x[47]), .Z(n604) );
  NANDN U684 ( .A(x[46]), .B(y[46]), .Z(n603) );
  NAND U685 ( .A(n604), .B(n603), .Z(n1073) );
  ANDN U686 ( .B(n605), .A(n1073), .Z(n606) );
  NANDN U687 ( .A(n1074), .B(n606), .Z(n607) );
  NOR U688 ( .A(n608), .B(n607), .Z(n620) );
  XNOR U689 ( .A(y[61]), .B(x[61]), .Z(n610) );
  NANDN U690 ( .A(x[60]), .B(y[60]), .Z(n609) );
  NAND U691 ( .A(n610), .B(n609), .Z(n1068) );
  XNOR U692 ( .A(y[57]), .B(x[57]), .Z(n612) );
  NANDN U693 ( .A(x[56]), .B(y[56]), .Z(n611) );
  AND U694 ( .A(n612), .B(n611), .Z(n1135) );
  XNOR U695 ( .A(y[59]), .B(x[59]), .Z(n614) );
  NANDN U696 ( .A(x[58]), .B(y[58]), .Z(n613) );
  NAND U697 ( .A(n614), .B(n613), .Z(n1069) );
  ANDN U698 ( .B(n1135), .A(n1069), .Z(n617) );
  XNOR U699 ( .A(y[63]), .B(x[63]), .Z(n616) );
  NANDN U700 ( .A(x[62]), .B(y[62]), .Z(n615) );
  NAND U701 ( .A(n616), .B(n615), .Z(n1067) );
  ANDN U702 ( .B(n617), .A(n1067), .Z(n618) );
  NANDN U703 ( .A(n1068), .B(n618), .Z(n619) );
  ANDN U704 ( .B(n620), .A(n619), .Z(n621) );
  NANDN U705 ( .A(n622), .B(n621), .Z(n623) );
  NOR U706 ( .A(n624), .B(n623), .Z(n672) );
  XNOR U707 ( .A(y[117]), .B(x[117]), .Z(n626) );
  NANDN U708 ( .A(x[116]), .B(y[116]), .Z(n625) );
  NAND U709 ( .A(n626), .B(n625), .Z(n1047) );
  XNOR U710 ( .A(y[113]), .B(x[113]), .Z(n628) );
  NANDN U711 ( .A(x[112]), .B(y[112]), .Z(n627) );
  AND U712 ( .A(n628), .B(n627), .Z(n1182) );
  XNOR U713 ( .A(y[115]), .B(x[115]), .Z(n630) );
  NANDN U714 ( .A(x[114]), .B(y[114]), .Z(n629) );
  NAND U715 ( .A(n630), .B(n629), .Z(n1048) );
  ANDN U716 ( .B(n1182), .A(n1048), .Z(n633) );
  XNOR U717 ( .A(y[119]), .B(x[119]), .Z(n632) );
  NANDN U718 ( .A(x[118]), .B(y[118]), .Z(n631) );
  NAND U719 ( .A(n632), .B(n631), .Z(n1046) );
  ANDN U720 ( .B(n633), .A(n1046), .Z(n634) );
  NANDN U721 ( .A(n1047), .B(n634), .Z(n670) );
  XNOR U722 ( .A(y[101]), .B(x[101]), .Z(n636) );
  NANDN U723 ( .A(x[100]), .B(y[100]), .Z(n635) );
  NAND U724 ( .A(n636), .B(n635), .Z(n1053) );
  XNOR U725 ( .A(y[97]), .B(x[97]), .Z(n638) );
  NANDN U726 ( .A(x[96]), .B(y[96]), .Z(n637) );
  AND U727 ( .A(n638), .B(n637), .Z(n1169) );
  XNOR U728 ( .A(y[99]), .B(x[99]), .Z(n640) );
  NANDN U729 ( .A(x[98]), .B(y[98]), .Z(n639) );
  NAND U730 ( .A(n640), .B(n639), .Z(n1054) );
  ANDN U731 ( .B(n1169), .A(n1054), .Z(n643) );
  XNOR U732 ( .A(y[103]), .B(x[103]), .Z(n642) );
  NANDN U733 ( .A(x[102]), .B(y[102]), .Z(n641) );
  NAND U734 ( .A(n642), .B(n641), .Z(n1052) );
  ANDN U735 ( .B(n643), .A(n1052), .Z(n644) );
  NANDN U736 ( .A(n1053), .B(n644), .Z(n656) );
  XNOR U737 ( .A(y[109]), .B(x[109]), .Z(n646) );
  NANDN U738 ( .A(x[108]), .B(y[108]), .Z(n645) );
  NAND U739 ( .A(n646), .B(n645), .Z(n1050) );
  XNOR U740 ( .A(y[105]), .B(x[105]), .Z(n648) );
  NANDN U741 ( .A(x[104]), .B(y[104]), .Z(n647) );
  AND U742 ( .A(n648), .B(n647), .Z(n1175) );
  XNOR U743 ( .A(y[107]), .B(x[107]), .Z(n650) );
  NANDN U744 ( .A(x[106]), .B(y[106]), .Z(n649) );
  NAND U745 ( .A(n650), .B(n649), .Z(n1051) );
  ANDN U746 ( .B(n1175), .A(n1051), .Z(n653) );
  XNOR U747 ( .A(y[111]), .B(x[111]), .Z(n652) );
  NANDN U748 ( .A(x[110]), .B(y[110]), .Z(n651) );
  NAND U749 ( .A(n652), .B(n651), .Z(n1049) );
  ANDN U750 ( .B(n653), .A(n1049), .Z(n654) );
  NANDN U751 ( .A(n1050), .B(n654), .Z(n655) );
  NOR U752 ( .A(n656), .B(n655), .Z(n668) );
  XNOR U753 ( .A(y[125]), .B(x[125]), .Z(n658) );
  NANDN U754 ( .A(x[124]), .B(y[124]), .Z(n657) );
  NAND U755 ( .A(n658), .B(n657), .Z(n1044) );
  XNOR U756 ( .A(y[121]), .B(x[121]), .Z(n660) );
  NANDN U757 ( .A(x[120]), .B(y[120]), .Z(n659) );
  AND U758 ( .A(n660), .B(n659), .Z(n1189) );
  XNOR U759 ( .A(y[123]), .B(x[123]), .Z(n662) );
  NANDN U760 ( .A(x[122]), .B(y[122]), .Z(n661) );
  NAND U761 ( .A(n662), .B(n661), .Z(n1045) );
  ANDN U762 ( .B(n1189), .A(n1045), .Z(n665) );
  XNOR U763 ( .A(y[127]), .B(x[127]), .Z(n664) );
  NANDN U764 ( .A(x[126]), .B(y[126]), .Z(n663) );
  NAND U765 ( .A(n664), .B(n663), .Z(n1043) );
  ANDN U766 ( .B(n665), .A(n1043), .Z(n666) );
  NANDN U767 ( .A(n1044), .B(n666), .Z(n667) );
  ANDN U768 ( .B(n668), .A(n667), .Z(n669) );
  NANDN U769 ( .A(n670), .B(n669), .Z(n671) );
  ANDN U770 ( .B(n672), .A(n671), .Z(n673) );
  NANDN U771 ( .A(n674), .B(n673), .Z(n994) );
  XNOR U772 ( .A(x[189]), .B(y[189]), .Z(n676) );
  NANDN U773 ( .A(x[188]), .B(y[188]), .Z(n675) );
  NAND U774 ( .A(n676), .B(n675), .Z(n1020) );
  XNOR U775 ( .A(x[185]), .B(y[185]), .Z(n678) );
  NANDN U776 ( .A(x[184]), .B(y[184]), .Z(n677) );
  AND U777 ( .A(n678), .B(n677), .Z(n1239) );
  XNOR U778 ( .A(x[187]), .B(y[187]), .Z(n680) );
  NANDN U779 ( .A(x[186]), .B(y[186]), .Z(n679) );
  NAND U780 ( .A(n680), .B(n679), .Z(n1021) );
  ANDN U781 ( .B(n1239), .A(n1021), .Z(n683) );
  XNOR U782 ( .A(x[191]), .B(y[191]), .Z(n682) );
  NANDN U783 ( .A(x[190]), .B(y[190]), .Z(n681) );
  NAND U784 ( .A(n682), .B(n681), .Z(n1019) );
  ANDN U785 ( .B(n683), .A(n1019), .Z(n684) );
  NANDN U786 ( .A(n1020), .B(n684), .Z(n720) );
  XNOR U787 ( .A(x[173]), .B(y[173]), .Z(n686) );
  NANDN U788 ( .A(x[172]), .B(y[172]), .Z(n685) );
  NAND U789 ( .A(n686), .B(n685), .Z(n1026) );
  XNOR U790 ( .A(x[169]), .B(y[169]), .Z(n688) );
  NANDN U791 ( .A(x[168]), .B(y[168]), .Z(n687) );
  AND U792 ( .A(n688), .B(n687), .Z(n1226) );
  XNOR U793 ( .A(x[171]), .B(y[171]), .Z(n690) );
  NANDN U794 ( .A(x[170]), .B(y[170]), .Z(n689) );
  NAND U795 ( .A(n690), .B(n689), .Z(n1027) );
  ANDN U796 ( .B(n1226), .A(n1027), .Z(n693) );
  XNOR U797 ( .A(x[175]), .B(y[175]), .Z(n692) );
  NANDN U798 ( .A(x[174]), .B(y[174]), .Z(n691) );
  NAND U799 ( .A(n692), .B(n691), .Z(n1025) );
  ANDN U800 ( .B(n693), .A(n1025), .Z(n694) );
  NANDN U801 ( .A(n1026), .B(n694), .Z(n706) );
  XNOR U802 ( .A(x[165]), .B(y[165]), .Z(n696) );
  NANDN U803 ( .A(x[164]), .B(y[164]), .Z(n695) );
  NAND U804 ( .A(n696), .B(n695), .Z(n1029) );
  XNOR U805 ( .A(x[161]), .B(y[161]), .Z(n698) );
  NANDN U806 ( .A(x[160]), .B(y[160]), .Z(n697) );
  AND U807 ( .A(n698), .B(n697), .Z(n1219) );
  XNOR U808 ( .A(x[163]), .B(y[163]), .Z(n700) );
  NANDN U809 ( .A(x[162]), .B(y[162]), .Z(n699) );
  NAND U810 ( .A(n700), .B(n699), .Z(n1030) );
  ANDN U811 ( .B(n1219), .A(n1030), .Z(n703) );
  XNOR U812 ( .A(x[167]), .B(y[167]), .Z(n702) );
  NANDN U813 ( .A(x[166]), .B(y[166]), .Z(n701) );
  NAND U814 ( .A(n702), .B(n701), .Z(n1028) );
  ANDN U815 ( .B(n703), .A(n1028), .Z(n704) );
  NANDN U816 ( .A(n1029), .B(n704), .Z(n705) );
  NOR U817 ( .A(n706), .B(n705), .Z(n718) );
  XNOR U818 ( .A(x[181]), .B(y[181]), .Z(n708) );
  NANDN U819 ( .A(x[180]), .B(y[180]), .Z(n707) );
  NAND U820 ( .A(n708), .B(n707), .Z(n1023) );
  XNOR U821 ( .A(x[177]), .B(y[177]), .Z(n710) );
  NANDN U822 ( .A(x[176]), .B(y[176]), .Z(n709) );
  AND U823 ( .A(n710), .B(n709), .Z(n1232) );
  XNOR U824 ( .A(x[179]), .B(y[179]), .Z(n712) );
  NANDN U825 ( .A(x[178]), .B(y[178]), .Z(n711) );
  NAND U826 ( .A(n712), .B(n711), .Z(n1024) );
  ANDN U827 ( .B(n1232), .A(n1024), .Z(n715) );
  XNOR U828 ( .A(x[183]), .B(y[183]), .Z(n714) );
  NANDN U829 ( .A(x[182]), .B(y[182]), .Z(n713) );
  NAND U830 ( .A(n714), .B(n713), .Z(n1022) );
  ANDN U831 ( .B(n715), .A(n1022), .Z(n716) );
  NANDN U832 ( .A(n1023), .B(n716), .Z(n717) );
  ANDN U833 ( .B(n718), .A(n717), .Z(n719) );
  NANDN U834 ( .A(n720), .B(n719), .Z(n768) );
  XNOR U835 ( .A(x[157]), .B(y[157]), .Z(n722) );
  NANDN U836 ( .A(x[156]), .B(y[156]), .Z(n721) );
  NAND U837 ( .A(n722), .B(n721), .Z(n1032) );
  XNOR U838 ( .A(x[153]), .B(y[153]), .Z(n724) );
  NANDN U839 ( .A(x[152]), .B(y[152]), .Z(n723) );
  AND U840 ( .A(n724), .B(n723), .Z(n1212) );
  XNOR U841 ( .A(x[155]), .B(y[155]), .Z(n726) );
  NANDN U842 ( .A(x[154]), .B(y[154]), .Z(n725) );
  NAND U843 ( .A(n726), .B(n725), .Z(n1033) );
  ANDN U844 ( .B(n1212), .A(n1033), .Z(n729) );
  XNOR U845 ( .A(x[159]), .B(y[159]), .Z(n728) );
  NANDN U846 ( .A(x[158]), .B(y[158]), .Z(n727) );
  NAND U847 ( .A(n728), .B(n727), .Z(n1031) );
  ANDN U848 ( .B(n729), .A(n1031), .Z(n730) );
  NANDN U849 ( .A(n1032), .B(n730), .Z(n766) );
  XNOR U850 ( .A(x[141]), .B(y[141]), .Z(n732) );
  NANDN U851 ( .A(x[140]), .B(y[140]), .Z(n731) );
  NAND U852 ( .A(n732), .B(n731), .Z(n1038) );
  XNOR U853 ( .A(x[137]), .B(y[137]), .Z(n734) );
  NANDN U854 ( .A(x[136]), .B(y[136]), .Z(n733) );
  AND U855 ( .A(n734), .B(n733), .Z(n1201) );
  XNOR U856 ( .A(x[139]), .B(y[139]), .Z(n736) );
  NANDN U857 ( .A(x[138]), .B(y[138]), .Z(n735) );
  NAND U858 ( .A(n736), .B(n735), .Z(n1039) );
  ANDN U859 ( .B(n1201), .A(n1039), .Z(n739) );
  XNOR U860 ( .A(x[143]), .B(y[143]), .Z(n738) );
  NANDN U861 ( .A(x[142]), .B(y[142]), .Z(n737) );
  NAND U862 ( .A(n738), .B(n737), .Z(n1037) );
  ANDN U863 ( .B(n739), .A(n1037), .Z(n740) );
  NANDN U864 ( .A(n1038), .B(n740), .Z(n752) );
  XNOR U865 ( .A(x[133]), .B(y[133]), .Z(n742) );
  NANDN U866 ( .A(x[132]), .B(y[132]), .Z(n741) );
  NAND U867 ( .A(n742), .B(n741), .Z(n1041) );
  XNOR U868 ( .A(x[129]), .B(y[129]), .Z(n744) );
  NANDN U869 ( .A(x[128]), .B(y[128]), .Z(n743) );
  AND U870 ( .A(n744), .B(n743), .Z(n1195) );
  XNOR U871 ( .A(x[131]), .B(y[131]), .Z(n746) );
  NANDN U872 ( .A(x[130]), .B(y[130]), .Z(n745) );
  NAND U873 ( .A(n746), .B(n745), .Z(n1042) );
  ANDN U874 ( .B(n1195), .A(n1042), .Z(n749) );
  XNOR U875 ( .A(x[135]), .B(y[135]), .Z(n748) );
  NANDN U876 ( .A(x[134]), .B(y[134]), .Z(n747) );
  NAND U877 ( .A(n748), .B(n747), .Z(n1040) );
  ANDN U878 ( .B(n749), .A(n1040), .Z(n750) );
  NANDN U879 ( .A(n1041), .B(n750), .Z(n751) );
  NOR U880 ( .A(n752), .B(n751), .Z(n764) );
  XNOR U881 ( .A(x[149]), .B(y[149]), .Z(n754) );
  NANDN U882 ( .A(x[148]), .B(y[148]), .Z(n753) );
  NAND U883 ( .A(n754), .B(n753), .Z(n1035) );
  XNOR U884 ( .A(x[145]), .B(y[145]), .Z(n756) );
  NANDN U885 ( .A(x[144]), .B(y[144]), .Z(n755) );
  AND U886 ( .A(n756), .B(n755), .Z(n1206) );
  XNOR U887 ( .A(x[147]), .B(y[147]), .Z(n758) );
  NANDN U888 ( .A(x[146]), .B(y[146]), .Z(n757) );
  NAND U889 ( .A(n758), .B(n757), .Z(n1036) );
  ANDN U890 ( .B(n1206), .A(n1036), .Z(n761) );
  XNOR U891 ( .A(x[151]), .B(y[151]), .Z(n760) );
  NANDN U892 ( .A(x[150]), .B(y[150]), .Z(n759) );
  NAND U893 ( .A(n760), .B(n759), .Z(n1034) );
  ANDN U894 ( .B(n761), .A(n1034), .Z(n762) );
  NANDN U895 ( .A(n1035), .B(n762), .Z(n763) );
  ANDN U896 ( .B(n764), .A(n763), .Z(n765) );
  NANDN U897 ( .A(n766), .B(n765), .Z(n767) );
  NOR U898 ( .A(n768), .B(n767), .Z(n992) );
  ANDN U899 ( .B(x[252]), .A(y[252]), .Z(n1294) );
  ANDN U900 ( .B(x[248]), .A(y[248]), .Z(n1289) );
  ANDN U901 ( .B(x[250]), .A(y[250]), .Z(n1292) );
  NOR U902 ( .A(n1289), .B(n1292), .Z(n769) );
  ANDN U903 ( .B(x[254]), .A(y[254]), .Z(n1295) );
  ANDN U904 ( .B(n769), .A(n1295), .Z(n770) );
  NANDN U905 ( .A(n1294), .B(n770), .Z(n782) );
  ANDN U906 ( .B(x[236]), .A(y[236]), .Z(n1281) );
  ANDN U907 ( .B(x[232]), .A(y[232]), .Z(n1276) );
  ANDN U908 ( .B(x[234]), .A(y[234]), .Z(n1280) );
  NOR U909 ( .A(n1276), .B(n1280), .Z(n771) );
  ANDN U910 ( .B(x[238]), .A(y[238]), .Z(n1282) );
  ANDN U911 ( .B(n771), .A(n1282), .Z(n772) );
  NANDN U912 ( .A(n1281), .B(n772), .Z(n776) );
  ANDN U913 ( .B(x[228]), .A(y[228]), .Z(n1274) );
  ANDN U914 ( .B(x[224]), .A(y[224]), .Z(n1271) );
  ANDN U915 ( .B(x[226]), .A(y[226]), .Z(n1273) );
  NOR U916 ( .A(n1271), .B(n1273), .Z(n773) );
  ANDN U917 ( .B(x[230]), .A(y[230]), .Z(n1275) );
  ANDN U918 ( .B(n773), .A(n1275), .Z(n774) );
  NANDN U919 ( .A(n1274), .B(n774), .Z(n775) );
  NOR U920 ( .A(n776), .B(n775), .Z(n780) );
  ANDN U921 ( .B(x[244]), .A(y[244]), .Z(n1287) );
  ANDN U922 ( .B(x[240]), .A(y[240]), .Z(n1283) );
  ANDN U923 ( .B(x[242]), .A(y[242]), .Z(n1286) );
  NOR U924 ( .A(n1283), .B(n1286), .Z(n777) );
  ANDN U925 ( .B(x[246]), .A(y[246]), .Z(n1288) );
  ANDN U926 ( .B(n777), .A(n1288), .Z(n778) );
  NANDN U927 ( .A(n1287), .B(n778), .Z(n779) );
  ANDN U928 ( .B(n780), .A(n779), .Z(n781) );
  NANDN U929 ( .A(n782), .B(n781), .Z(n830) );
  ANDN U930 ( .B(x[188]), .A(y[188]), .Z(n1241) );
  ANDN U931 ( .B(x[184]), .A(y[184]), .Z(n1238) );
  ANDN U932 ( .B(x[186]), .A(y[186]), .Z(n1240) );
  NOR U933 ( .A(n1238), .B(n1240), .Z(n783) );
  ANDN U934 ( .B(x[190]), .A(y[190]), .Z(n1244) );
  ANDN U935 ( .B(n783), .A(n1244), .Z(n784) );
  NANDN U936 ( .A(n1241), .B(n784), .Z(n796) );
  ANDN U937 ( .B(x[172]), .A(y[172]), .Z(n1229) );
  ANDN U938 ( .B(x[168]), .A(y[168]), .Z(n1225) );
  ANDN U939 ( .B(x[170]), .A(y[170]), .Z(n1227) );
  NOR U940 ( .A(n1225), .B(n1227), .Z(n785) );
  ANDN U941 ( .B(x[174]), .A(y[174]), .Z(n1230) );
  ANDN U942 ( .B(n785), .A(n1230), .Z(n786) );
  NANDN U943 ( .A(n1229), .B(n786), .Z(n790) );
  ANDN U944 ( .B(x[164]), .A(y[164]), .Z(n1223) );
  ANDN U945 ( .B(x[160]), .A(y[160]), .Z(n1218) );
  ANDN U946 ( .B(x[162]), .A(y[162]), .Z(n1220) );
  NOR U947 ( .A(n1218), .B(n1220), .Z(n787) );
  ANDN U948 ( .B(x[166]), .A(y[166]), .Z(n1224) );
  ANDN U949 ( .B(n787), .A(n1224), .Z(n788) );
  NANDN U950 ( .A(n1223), .B(n788), .Z(n789) );
  NOR U951 ( .A(n790), .B(n789), .Z(n794) );
  ANDN U952 ( .B(x[180]), .A(y[180]), .Z(n1234) );
  ANDN U953 ( .B(x[176]), .A(y[176]), .Z(n1231) );
  ANDN U954 ( .B(x[178]), .A(y[178]), .Z(n1233) );
  NOR U955 ( .A(n1231), .B(n1233), .Z(n791) );
  ANDN U956 ( .B(x[182]), .A(y[182]), .Z(n1237) );
  ANDN U957 ( .B(n791), .A(n1237), .Z(n792) );
  NANDN U958 ( .A(n1234), .B(n792), .Z(n793) );
  ANDN U959 ( .B(n794), .A(n793), .Z(n795) );
  NANDN U960 ( .A(n796), .B(n795), .Z(n812) );
  ANDN U961 ( .B(x[156]), .A(y[156]), .Z(n1216) );
  ANDN U962 ( .B(x[152]), .A(y[152]), .Z(n1211) );
  ANDN U963 ( .B(x[154]), .A(y[154]), .Z(n1213) );
  NOR U964 ( .A(n1211), .B(n1213), .Z(n797) );
  ANDN U965 ( .B(x[158]), .A(y[158]), .Z(n1217) );
  ANDN U966 ( .B(n797), .A(n1217), .Z(n798) );
  NANDN U967 ( .A(n1216), .B(n798), .Z(n810) );
  ANDN U968 ( .B(x[140]), .A(y[140]), .Z(n1203) );
  ANDN U969 ( .B(x[136]), .A(y[136]), .Z(n1199) );
  ANDN U970 ( .B(x[138]), .A(y[138]), .Z(n1202) );
  NOR U971 ( .A(n1199), .B(n1202), .Z(n799) );
  ANDN U972 ( .B(x[142]), .A(y[142]), .Z(n1204) );
  ANDN U973 ( .B(n799), .A(n1204), .Z(n800) );
  NANDN U974 ( .A(n1203), .B(n800), .Z(n804) );
  ANDN U975 ( .B(x[132]), .A(y[132]), .Z(n1197) );
  ANDN U976 ( .B(x[128]), .A(y[128]), .Z(n1193) );
  ANDN U977 ( .B(x[130]), .A(y[130]), .Z(n1196) );
  NOR U978 ( .A(n1193), .B(n1196), .Z(n801) );
  ANDN U979 ( .B(x[134]), .A(y[134]), .Z(n1198) );
  ANDN U980 ( .B(n801), .A(n1198), .Z(n802) );
  NANDN U981 ( .A(n1197), .B(n802), .Z(n803) );
  NOR U982 ( .A(n804), .B(n803), .Z(n808) );
  ANDN U983 ( .B(x[148]), .A(y[148]), .Z(n1209) );
  ANDN U984 ( .B(x[144]), .A(y[144]), .Z(n1205) );
  ANDN U985 ( .B(x[146]), .A(y[146]), .Z(n1208) );
  NOR U986 ( .A(n1205), .B(n1208), .Z(n805) );
  ANDN U987 ( .B(x[150]), .A(y[150]), .Z(n1210) );
  ANDN U988 ( .B(n805), .A(n1210), .Z(n806) );
  NANDN U989 ( .A(n1209), .B(n806), .Z(n807) );
  ANDN U990 ( .B(n808), .A(n807), .Z(n809) );
  NANDN U991 ( .A(n810), .B(n809), .Z(n811) );
  NOR U992 ( .A(n812), .B(n811), .Z(n828) );
  ANDN U993 ( .B(x[220]), .A(y[220]), .Z(n1268) );
  ANDN U994 ( .B(x[216]), .A(y[216]), .Z(n1265) );
  ANDN U995 ( .B(x[218]), .A(y[218]), .Z(n1267) );
  NOR U996 ( .A(n1265), .B(n1267), .Z(n813) );
  ANDN U997 ( .B(x[222]), .A(y[222]), .Z(n1269) );
  ANDN U998 ( .B(n813), .A(n1269), .Z(n814) );
  NANDN U999 ( .A(n1268), .B(n814), .Z(n826) );
  ANDN U1000 ( .B(x[204]), .A(y[204]), .Z(n1254) );
  ANDN U1001 ( .B(x[200]), .A(y[200]), .Z(n1251) );
  ANDN U1002 ( .B(x[202]), .A(y[202]), .Z(n1253) );
  NOR U1003 ( .A(n1251), .B(n1253), .Z(n815) );
  ANDN U1004 ( .B(x[206]), .A(y[206]), .Z(n1255) );
  ANDN U1005 ( .B(n815), .A(n1255), .Z(n816) );
  NANDN U1006 ( .A(n1254), .B(n816), .Z(n820) );
  ANDN U1007 ( .B(x[196]), .A(y[196]), .Z(n1248) );
  ANDN U1008 ( .B(x[192]), .A(y[192]), .Z(n1245) );
  ANDN U1009 ( .B(x[194]), .A(y[194]), .Z(n1247) );
  NOR U1010 ( .A(n1245), .B(n1247), .Z(n817) );
  ANDN U1011 ( .B(x[198]), .A(y[198]), .Z(n1250) );
  ANDN U1012 ( .B(n817), .A(n1250), .Z(n818) );
  NANDN U1013 ( .A(n1248), .B(n818), .Z(n819) );
  NOR U1014 ( .A(n820), .B(n819), .Z(n824) );
  ANDN U1015 ( .B(x[212]), .A(y[212]), .Z(n1261) );
  ANDN U1016 ( .B(x[208]), .A(y[208]), .Z(n1258) );
  ANDN U1017 ( .B(x[210]), .A(y[210]), .Z(n1260) );
  NOR U1018 ( .A(n1258), .B(n1260), .Z(n821) );
  ANDN U1019 ( .B(x[214]), .A(y[214]), .Z(n1262) );
  ANDN U1020 ( .B(n821), .A(n1262), .Z(n822) );
  NANDN U1021 ( .A(n1261), .B(n822), .Z(n823) );
  ANDN U1022 ( .B(n824), .A(n823), .Z(n825) );
  NANDN U1023 ( .A(n826), .B(n825), .Z(n827) );
  ANDN U1024 ( .B(n828), .A(n827), .Z(n829) );
  NANDN U1025 ( .A(n830), .B(n829), .Z(n990) );
  XNOR U1026 ( .A(x[253]), .B(y[253]), .Z(n832) );
  NANDN U1027 ( .A(x[252]), .B(y[252]), .Z(n831) );
  NAND U1028 ( .A(n832), .B(n831), .Z(n996) );
  XNOR U1029 ( .A(x[249]), .B(y[249]), .Z(n834) );
  NANDN U1030 ( .A(x[248]), .B(y[248]), .Z(n833) );
  AND U1031 ( .A(n834), .B(n833), .Z(n1290) );
  XNOR U1032 ( .A(x[251]), .B(y[251]), .Z(n836) );
  NANDN U1033 ( .A(x[250]), .B(y[250]), .Z(n835) );
  NAND U1034 ( .A(n836), .B(n835), .Z(n997) );
  ANDN U1035 ( .B(n1290), .A(n997), .Z(n839) );
  XNOR U1036 ( .A(x[255]), .B(y[255]), .Z(n838) );
  NANDN U1037 ( .A(x[254]), .B(y[254]), .Z(n837) );
  NAND U1038 ( .A(n838), .B(n837), .Z(n995) );
  ANDN U1039 ( .B(n839), .A(n995), .Z(n840) );
  NANDN U1040 ( .A(n996), .B(n840), .Z(n876) );
  XNOR U1041 ( .A(x[237]), .B(y[237]), .Z(n842) );
  NANDN U1042 ( .A(x[236]), .B(y[236]), .Z(n841) );
  NAND U1043 ( .A(n842), .B(n841), .Z(n1002) );
  XNOR U1044 ( .A(x[233]), .B(y[233]), .Z(n844) );
  NANDN U1045 ( .A(x[232]), .B(y[232]), .Z(n843) );
  AND U1046 ( .A(n844), .B(n843), .Z(n1279) );
  XNOR U1047 ( .A(x[235]), .B(y[235]), .Z(n846) );
  NANDN U1048 ( .A(x[234]), .B(y[234]), .Z(n845) );
  NAND U1049 ( .A(n846), .B(n845), .Z(n1003) );
  ANDN U1050 ( .B(n1279), .A(n1003), .Z(n849) );
  XNOR U1051 ( .A(x[239]), .B(y[239]), .Z(n848) );
  NANDN U1052 ( .A(x[238]), .B(y[238]), .Z(n847) );
  NAND U1053 ( .A(n848), .B(n847), .Z(n1001) );
  ANDN U1054 ( .B(n849), .A(n1001), .Z(n850) );
  NANDN U1055 ( .A(n1002), .B(n850), .Z(n862) );
  XNOR U1056 ( .A(x[229]), .B(y[229]), .Z(n852) );
  NANDN U1057 ( .A(x[228]), .B(y[228]), .Z(n851) );
  NAND U1058 ( .A(n852), .B(n851), .Z(n1005) );
  XNOR U1059 ( .A(x[225]), .B(y[225]), .Z(n854) );
  NANDN U1060 ( .A(x[224]), .B(y[224]), .Z(n853) );
  AND U1061 ( .A(n854), .B(n853), .Z(n1272) );
  XNOR U1062 ( .A(x[227]), .B(y[227]), .Z(n856) );
  NANDN U1063 ( .A(x[226]), .B(y[226]), .Z(n855) );
  NAND U1064 ( .A(n856), .B(n855), .Z(n1006) );
  ANDN U1065 ( .B(n1272), .A(n1006), .Z(n859) );
  XNOR U1066 ( .A(x[231]), .B(y[231]), .Z(n858) );
  NANDN U1067 ( .A(x[230]), .B(y[230]), .Z(n857) );
  NAND U1068 ( .A(n858), .B(n857), .Z(n1004) );
  ANDN U1069 ( .B(n859), .A(n1004), .Z(n860) );
  NANDN U1070 ( .A(n1005), .B(n860), .Z(n861) );
  NOR U1071 ( .A(n862), .B(n861), .Z(n874) );
  XNOR U1072 ( .A(x[245]), .B(y[245]), .Z(n864) );
  NANDN U1073 ( .A(x[244]), .B(y[244]), .Z(n863) );
  NAND U1074 ( .A(n864), .B(n863), .Z(n999) );
  XNOR U1075 ( .A(x[241]), .B(y[241]), .Z(n866) );
  NANDN U1076 ( .A(x[240]), .B(y[240]), .Z(n865) );
  AND U1077 ( .A(n866), .B(n865), .Z(n1285) );
  XNOR U1078 ( .A(x[243]), .B(y[243]), .Z(n868) );
  NANDN U1079 ( .A(x[242]), .B(y[242]), .Z(n867) );
  NAND U1080 ( .A(n868), .B(n867), .Z(n1000) );
  ANDN U1081 ( .B(n1285), .A(n1000), .Z(n871) );
  XNOR U1082 ( .A(x[247]), .B(y[247]), .Z(n870) );
  NANDN U1083 ( .A(x[246]), .B(y[246]), .Z(n869) );
  NAND U1084 ( .A(n870), .B(n869), .Z(n998) );
  ANDN U1085 ( .B(n871), .A(n998), .Z(n872) );
  NANDN U1086 ( .A(n999), .B(n872), .Z(n873) );
  ANDN U1087 ( .B(n874), .A(n873), .Z(n875) );
  NANDN U1088 ( .A(n876), .B(n875), .Z(n924) );
  XNOR U1089 ( .A(x[221]), .B(y[221]), .Z(n878) );
  NANDN U1090 ( .A(x[220]), .B(y[220]), .Z(n877) );
  NAND U1091 ( .A(n878), .B(n877), .Z(n1008) );
  XNOR U1092 ( .A(x[217]), .B(y[217]), .Z(n880) );
  NANDN U1093 ( .A(x[216]), .B(y[216]), .Z(n879) );
  AND U1094 ( .A(n880), .B(n879), .Z(n1266) );
  XNOR U1095 ( .A(x[219]), .B(y[219]), .Z(n882) );
  NANDN U1096 ( .A(x[218]), .B(y[218]), .Z(n881) );
  NAND U1097 ( .A(n882), .B(n881), .Z(n1009) );
  ANDN U1098 ( .B(n1266), .A(n1009), .Z(n885) );
  XNOR U1099 ( .A(x[223]), .B(y[223]), .Z(n884) );
  NANDN U1100 ( .A(x[222]), .B(y[222]), .Z(n883) );
  NAND U1101 ( .A(n884), .B(n883), .Z(n1007) );
  ANDN U1102 ( .B(n885), .A(n1007), .Z(n886) );
  NANDN U1103 ( .A(n1008), .B(n886), .Z(n922) );
  XNOR U1104 ( .A(x[205]), .B(y[205]), .Z(n888) );
  NANDN U1105 ( .A(x[204]), .B(y[204]), .Z(n887) );
  NAND U1106 ( .A(n888), .B(n887), .Z(n1014) );
  XNOR U1107 ( .A(x[201]), .B(y[201]), .Z(n890) );
  NANDN U1108 ( .A(x[200]), .B(y[200]), .Z(n889) );
  AND U1109 ( .A(n890), .B(n889), .Z(n1252) );
  XNOR U1110 ( .A(x[203]), .B(y[203]), .Z(n892) );
  NANDN U1111 ( .A(x[202]), .B(y[202]), .Z(n891) );
  NAND U1112 ( .A(n892), .B(n891), .Z(n1015) );
  ANDN U1113 ( .B(n1252), .A(n1015), .Z(n895) );
  XNOR U1114 ( .A(x[207]), .B(y[207]), .Z(n894) );
  NANDN U1115 ( .A(x[206]), .B(y[206]), .Z(n893) );
  NAND U1116 ( .A(n894), .B(n893), .Z(n1013) );
  ANDN U1117 ( .B(n895), .A(n1013), .Z(n896) );
  NANDN U1118 ( .A(n1014), .B(n896), .Z(n908) );
  XNOR U1119 ( .A(x[197]), .B(y[197]), .Z(n898) );
  NANDN U1120 ( .A(x[196]), .B(y[196]), .Z(n897) );
  NAND U1121 ( .A(n898), .B(n897), .Z(n1017) );
  XNOR U1122 ( .A(x[193]), .B(y[193]), .Z(n900) );
  NANDN U1123 ( .A(x[192]), .B(y[192]), .Z(n899) );
  AND U1124 ( .A(n900), .B(n899), .Z(n1246) );
  XNOR U1125 ( .A(x[195]), .B(y[195]), .Z(n902) );
  NANDN U1126 ( .A(x[194]), .B(y[194]), .Z(n901) );
  NAND U1127 ( .A(n902), .B(n901), .Z(n1018) );
  ANDN U1128 ( .B(n1246), .A(n1018), .Z(n905) );
  XNOR U1129 ( .A(x[199]), .B(y[199]), .Z(n904) );
  NANDN U1130 ( .A(x[198]), .B(y[198]), .Z(n903) );
  NAND U1131 ( .A(n904), .B(n903), .Z(n1016) );
  ANDN U1132 ( .B(n905), .A(n1016), .Z(n906) );
  NANDN U1133 ( .A(n1017), .B(n906), .Z(n907) );
  NOR U1134 ( .A(n908), .B(n907), .Z(n920) );
  XNOR U1135 ( .A(x[213]), .B(y[213]), .Z(n910) );
  NANDN U1136 ( .A(x[212]), .B(y[212]), .Z(n909) );
  NAND U1137 ( .A(n910), .B(n909), .Z(n1011) );
  XNOR U1138 ( .A(x[209]), .B(y[209]), .Z(n912) );
  NANDN U1139 ( .A(x[208]), .B(y[208]), .Z(n911) );
  AND U1140 ( .A(n912), .B(n911), .Z(n1259) );
  XNOR U1141 ( .A(x[211]), .B(y[211]), .Z(n914) );
  NANDN U1142 ( .A(x[210]), .B(y[210]), .Z(n913) );
  NAND U1143 ( .A(n914), .B(n913), .Z(n1012) );
  ANDN U1144 ( .B(n1259), .A(n1012), .Z(n917) );
  XNOR U1145 ( .A(x[215]), .B(y[215]), .Z(n916) );
  NANDN U1146 ( .A(x[214]), .B(y[214]), .Z(n915) );
  NAND U1147 ( .A(n916), .B(n915), .Z(n1010) );
  ANDN U1148 ( .B(n917), .A(n1010), .Z(n918) );
  NANDN U1149 ( .A(n1011), .B(n918), .Z(n919) );
  ANDN U1150 ( .B(n920), .A(n919), .Z(n921) );
  NANDN U1151 ( .A(n922), .B(n921), .Z(n923) );
  NOR U1152 ( .A(n924), .B(n923), .Z(n988) );
  ANDN U1153 ( .B(x[124]), .A(y[124]), .Z(n1191) );
  ANDN U1154 ( .B(x[120]), .A(y[120]), .Z(n1188) );
  ANDN U1155 ( .B(x[122]), .A(y[122]), .Z(n1190) );
  NOR U1156 ( .A(n1188), .B(n1190), .Z(n925) );
  ANDN U1157 ( .B(x[126]), .A(y[126]), .Z(n1192) );
  ANDN U1158 ( .B(n925), .A(n1192), .Z(n926) );
  NANDN U1159 ( .A(n1191), .B(n926), .Z(n938) );
  ANDN U1160 ( .B(x[108]), .A(y[108]), .Z(n1177) );
  ANDN U1161 ( .B(x[104]), .A(y[104]), .Z(n1174) );
  ANDN U1162 ( .B(x[106]), .A(y[106]), .Z(n1176) );
  NOR U1163 ( .A(n1174), .B(n1176), .Z(n927) );
  ANDN U1164 ( .B(x[110]), .A(y[110]), .Z(n1178) );
  ANDN U1165 ( .B(n927), .A(n1178), .Z(n928) );
  NANDN U1166 ( .A(n1177), .B(n928), .Z(n932) );
  ANDN U1167 ( .B(x[100]), .A(y[100]), .Z(n1171) );
  ANDN U1168 ( .B(x[96]), .A(y[96]), .Z(n1168) );
  ANDN U1169 ( .B(x[98]), .A(y[98]), .Z(n1170) );
  NOR U1170 ( .A(n1168), .B(n1170), .Z(n929) );
  ANDN U1171 ( .B(x[102]), .A(y[102]), .Z(n1172) );
  ANDN U1172 ( .B(n929), .A(n1172), .Z(n930) );
  NANDN U1173 ( .A(n1171), .B(n930), .Z(n931) );
  NOR U1174 ( .A(n932), .B(n931), .Z(n936) );
  ANDN U1175 ( .B(x[116]), .A(y[116]), .Z(n1184) );
  ANDN U1176 ( .B(x[112]), .A(y[112]), .Z(n1181) );
  ANDN U1177 ( .B(x[114]), .A(y[114]), .Z(n1183) );
  NOR U1178 ( .A(n1181), .B(n1183), .Z(n933) );
  ANDN U1179 ( .B(x[118]), .A(y[118]), .Z(n1185) );
  ANDN U1180 ( .B(n933), .A(n1185), .Z(n934) );
  NANDN U1181 ( .A(n1184), .B(n934), .Z(n935) );
  ANDN U1182 ( .B(n936), .A(n935), .Z(n937) );
  NANDN U1183 ( .A(n938), .B(n937), .Z(n986) );
  ANDN U1184 ( .B(x[60]), .A(y[60]), .Z(n1139) );
  ANDN U1185 ( .B(x[56]), .A(y[56]), .Z(n1134) );
  ANDN U1186 ( .B(x[58]), .A(y[58]), .Z(n1136) );
  NOR U1187 ( .A(n1134), .B(n1136), .Z(n939) );
  ANDN U1188 ( .B(x[62]), .A(y[62]), .Z(n1140) );
  ANDN U1189 ( .B(n939), .A(n1140), .Z(n940) );
  NANDN U1190 ( .A(n1139), .B(n940), .Z(n952) );
  ANDN U1191 ( .B(x[44]), .A(y[44]), .Z(n1126) );
  ANDN U1192 ( .B(x[40]), .A(y[40]), .Z(n1121) );
  ANDN U1193 ( .B(x[42]), .A(y[42]), .Z(n1125) );
  NOR U1194 ( .A(n1121), .B(n1125), .Z(n941) );
  ANDN U1195 ( .B(x[46]), .A(y[46]), .Z(n1127) );
  ANDN U1196 ( .B(n941), .A(n1127), .Z(n942) );
  NANDN U1197 ( .A(n1126), .B(n942), .Z(n946) );
  ANDN U1198 ( .B(x[36]), .A(y[36]), .Z(n1119) );
  ANDN U1199 ( .B(x[32]), .A(y[32]), .Z(n1115) );
  ANDN U1200 ( .B(x[34]), .A(y[34]), .Z(n1118) );
  NOR U1201 ( .A(n1115), .B(n1118), .Z(n943) );
  ANDN U1202 ( .B(x[38]), .A(y[38]), .Z(n1120) );
  ANDN U1203 ( .B(n943), .A(n1120), .Z(n944) );
  NANDN U1204 ( .A(n1119), .B(n944), .Z(n945) );
  NOR U1205 ( .A(n946), .B(n945), .Z(n950) );
  ANDN U1206 ( .B(x[52]), .A(y[52]), .Z(n1132) );
  ANDN U1207 ( .B(x[48]), .A(y[48]), .Z(n1128) );
  ANDN U1208 ( .B(x[50]), .A(y[50]), .Z(n1130) );
  NOR U1209 ( .A(n1128), .B(n1130), .Z(n947) );
  ANDN U1210 ( .B(x[54]), .A(y[54]), .Z(n1133) );
  ANDN U1211 ( .B(n947), .A(n1133), .Z(n948) );
  NANDN U1212 ( .A(n1132), .B(n948), .Z(n949) );
  ANDN U1213 ( .B(n950), .A(n949), .Z(n951) );
  NANDN U1214 ( .A(n952), .B(n951), .Z(n968) );
  ANDN U1215 ( .B(x[28]), .A(y[28]), .Z(n1113) );
  ANDN U1216 ( .B(x[24]), .A(y[24]), .Z(n1109) );
  ANDN U1217 ( .B(x[26]), .A(y[26]), .Z(n1112) );
  NOR U1218 ( .A(n1109), .B(n1112), .Z(n953) );
  ANDN U1219 ( .B(x[30]), .A(y[30]), .Z(n1114) );
  ANDN U1220 ( .B(n953), .A(n1114), .Z(n954) );
  NANDN U1221 ( .A(n1113), .B(n954), .Z(n966) );
  ANDN U1222 ( .B(x[12]), .A(y[12]), .Z(n1100) );
  ANDN U1223 ( .B(x[8]), .A(y[8]), .Z(n1097) );
  ANDN U1224 ( .B(x[10]), .A(y[10]), .Z(n1099) );
  NOR U1225 ( .A(n1097), .B(n1099), .Z(n955) );
  ANDN U1226 ( .B(x[14]), .A(y[14]), .Z(n1101) );
  ANDN U1227 ( .B(n955), .A(n1101), .Z(n956) );
  NANDN U1228 ( .A(n1100), .B(n956), .Z(n960) );
  ANDN U1229 ( .B(x[2]), .A(y[2]), .Z(n1091) );
  ANDN U1230 ( .B(x[4]), .A(y[4]), .Z(n1093) );
  ANDN U1231 ( .B(x[0]), .A(y[0]), .Z(n1090) );
  NOR U1232 ( .A(n1093), .B(n1090), .Z(n957) );
  ANDN U1233 ( .B(x[6]), .A(y[6]), .Z(n1094) );
  ANDN U1234 ( .B(n957), .A(n1094), .Z(n958) );
  NANDN U1235 ( .A(n1091), .B(n958), .Z(n959) );
  NOR U1236 ( .A(n960), .B(n959), .Z(n964) );
  ANDN U1237 ( .B(x[20]), .A(y[20]), .Z(n1107) );
  ANDN U1238 ( .B(x[16]), .A(y[16]), .Z(n1104) );
  ANDN U1239 ( .B(x[18]), .A(y[18]), .Z(n1106) );
  NOR U1240 ( .A(n1104), .B(n1106), .Z(n961) );
  ANDN U1241 ( .B(x[22]), .A(y[22]), .Z(n1108) );
  ANDN U1242 ( .B(n961), .A(n1108), .Z(n962) );
  NANDN U1243 ( .A(n1107), .B(n962), .Z(n963) );
  ANDN U1244 ( .B(n964), .A(n963), .Z(n965) );
  NANDN U1245 ( .A(n966), .B(n965), .Z(n967) );
  NOR U1246 ( .A(n968), .B(n967), .Z(n984) );
  ANDN U1247 ( .B(x[92]), .A(y[92]), .Z(n1164) );
  ANDN U1248 ( .B(x[88]), .A(y[88]), .Z(n1161) );
  ANDN U1249 ( .B(x[90]), .A(y[90]), .Z(n1163) );
  NOR U1250 ( .A(n1161), .B(n1163), .Z(n969) );
  ANDN U1251 ( .B(x[94]), .A(y[94]), .Z(n1167) );
  ANDN U1252 ( .B(n969), .A(n1167), .Z(n970) );
  NANDN U1253 ( .A(n1164), .B(n970), .Z(n982) );
  ANDN U1254 ( .B(x[76]), .A(y[76]), .Z(n1151) );
  ANDN U1255 ( .B(x[72]), .A(y[72]), .Z(n1148) );
  ANDN U1256 ( .B(x[74]), .A(y[74]), .Z(n1150) );
  NOR U1257 ( .A(n1148), .B(n1150), .Z(n971) );
  ANDN U1258 ( .B(x[78]), .A(y[78]), .Z(n1153) );
  ANDN U1259 ( .B(n971), .A(n1153), .Z(n972) );
  NANDN U1260 ( .A(n1151), .B(n972), .Z(n976) );
  ANDN U1261 ( .B(x[68]), .A(y[68]), .Z(n1146) );
  ANDN U1262 ( .B(x[64]), .A(y[64]), .Z(n1141) );
  ANDN U1263 ( .B(x[66]), .A(y[66]), .Z(n1143) );
  NOR U1264 ( .A(n1141), .B(n1143), .Z(n973) );
  ANDN U1265 ( .B(x[70]), .A(y[70]), .Z(n1147) );
  ANDN U1266 ( .B(n973), .A(n1147), .Z(n974) );
  NANDN U1267 ( .A(n1146), .B(n974), .Z(n975) );
  NOR U1268 ( .A(n976), .B(n975), .Z(n980) );
  ANDN U1269 ( .B(x[84]), .A(y[84]), .Z(n1157) );
  ANDN U1270 ( .B(x[80]), .A(y[80]), .Z(n1154) );
  ANDN U1271 ( .B(x[82]), .A(y[82]), .Z(n1156) );
  NOR U1272 ( .A(n1154), .B(n1156), .Z(n977) );
  ANDN U1273 ( .B(x[86]), .A(y[86]), .Z(n1160) );
  ANDN U1274 ( .B(n977), .A(n1160), .Z(n978) );
  NANDN U1275 ( .A(n1157), .B(n978), .Z(n979) );
  ANDN U1276 ( .B(n980), .A(n979), .Z(n981) );
  NANDN U1277 ( .A(n982), .B(n981), .Z(n983) );
  ANDN U1278 ( .B(n984), .A(n983), .Z(n985) );
  NANDN U1279 ( .A(n986), .B(n985), .Z(n987) );
  ANDN U1280 ( .B(n988), .A(n987), .Z(n989) );
  NANDN U1281 ( .A(n990), .B(n989), .Z(n991) );
  ANDN U1282 ( .B(n992), .A(n991), .Z(n993) );
  NANDN U1283 ( .A(n994), .B(n993), .Z(n1296) );
  NANDN U1284 ( .A(n1296), .B(e), .Z(n5) );
  IV U1285 ( .A(n1010), .Z(n1264) );
  IV U1286 ( .A(n1020), .Z(n1243) );
  IV U1287 ( .A(n1030), .Z(n1222) );
  ANDN U1288 ( .B(x[119]), .A(y[119]), .Z(n1187) );
  IV U1289 ( .A(n1049), .Z(n1180) );
  ANDN U1290 ( .B(x[93]), .A(y[93]), .Z(n1166) );
  IV U1291 ( .A(n1059), .Z(n1159) );
  ANDN U1292 ( .B(x[67]), .A(y[67]), .Z(n1145) );
  IV U1293 ( .A(n1069), .Z(n1138) );
  ANDN U1294 ( .B(x[41]), .A(y[41]), .Z(n1124) );
  ANDN U1295 ( .B(x[15]), .A(y[15]), .Z(n1103) );
  IV U1296 ( .A(n1088), .Z(n1096) );
  ANDN U1297 ( .B(x[153]), .A(y[153]), .Z(n1214) );
  ANDN U1298 ( .B(x[179]), .A(y[179]), .Z(n1235) );
  ANDN U1299 ( .B(x[205]), .A(y[205]), .Z(n1256) );
  ANDN U1300 ( .B(x[231]), .A(y[231]), .Z(n1277) );
  ANDN U1301 ( .B(x[249]), .A(y[249]), .Z(n1293) );
endmodule

