
module sum_N1024_CC4 ( clk, rst, a, b, c );
  input [255:0] a;
  input [255:0] b;
  output [255:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR U3 ( .A(a[3]), .B(n1013), .Z(n71) );
  XOR U4 ( .A(a[6]), .B(n1004), .Z(n38) );
  XOR U5 ( .A(a[9]), .B(n995), .Z(n5) );
  XOR U6 ( .A(a[12]), .B(n986), .Z(n605) );
  XOR U7 ( .A(a[15]), .B(n977), .Z(n482) );
  XOR U8 ( .A(a[18]), .B(n968), .Z(n359) );
  XOR U9 ( .A(a[21]), .B(n959), .Z(n235) );
  XOR U10 ( .A(a[24]), .B(n950), .Z(n112) );
  XOR U11 ( .A(a[27]), .B(n941), .Z(n85) );
  XOR U12 ( .A(a[30]), .B(n932), .Z(n81) );
  XOR U13 ( .A(a[33]), .B(n923), .Z(n78) );
  XOR U14 ( .A(a[36]), .B(n914), .Z(n75) );
  XOR U15 ( .A(a[39]), .B(n905), .Z(n72) );
  XOR U16 ( .A(a[42]), .B(n896), .Z(n68) );
  XOR U17 ( .A(a[45]), .B(n887), .Z(n65) );
  XOR U18 ( .A(a[48]), .B(n878), .Z(n62) );
  XOR U19 ( .A(a[51]), .B(n869), .Z(n58) );
  XOR U20 ( .A(a[54]), .B(n860), .Z(n55) );
  XOR U21 ( .A(a[57]), .B(n851), .Z(n52) );
  XOR U22 ( .A(a[60]), .B(n842), .Z(n48) );
  XOR U23 ( .A(a[63]), .B(n833), .Z(n45) );
  XOR U24 ( .A(a[66]), .B(n824), .Z(n42) );
  XOR U25 ( .A(a[69]), .B(n815), .Z(n39) );
  XOR U26 ( .A(a[72]), .B(n806), .Z(n35) );
  XOR U27 ( .A(a[75]), .B(n797), .Z(n32) );
  XOR U28 ( .A(a[78]), .B(n788), .Z(n29) );
  XOR U29 ( .A(a[81]), .B(n779), .Z(n25) );
  XOR U30 ( .A(a[84]), .B(n770), .Z(n22) );
  XOR U31 ( .A(a[87]), .B(n761), .Z(n19) );
  XOR U32 ( .A(a[90]), .B(n752), .Z(n15) );
  XOR U33 ( .A(a[93]), .B(n743), .Z(n12) );
  XOR U34 ( .A(a[96]), .B(n734), .Z(n9) );
  XOR U35 ( .A(a[99]), .B(n725), .Z(n6) );
  XOR U36 ( .A(a[102]), .B(n713), .Z(n715) );
  XOR U37 ( .A(a[105]), .B(n701), .Z(n703) );
  XOR U38 ( .A(a[108]), .B(n689), .Z(n691) );
  XOR U39 ( .A(a[111]), .B(n676), .Z(n678) );
  XOR U40 ( .A(a[114]), .B(n664), .Z(n666) );
  XOR U41 ( .A(a[117]), .B(n652), .Z(n654) );
  XOR U42 ( .A(a[120]), .B(n639), .Z(n641) );
  XOR U43 ( .A(a[123]), .B(n627), .Z(n629) );
  XOR U44 ( .A(a[126]), .B(n615), .Z(n617) );
  XOR U45 ( .A(a[129]), .B(n602), .Z(n604) );
  XOR U46 ( .A(a[132]), .B(n590), .Z(n592) );
  XOR U47 ( .A(a[135]), .B(n578), .Z(n580) );
  XOR U48 ( .A(a[138]), .B(n566), .Z(n568) );
  XOR U49 ( .A(a[141]), .B(n553), .Z(n555) );
  XOR U50 ( .A(a[144]), .B(n541), .Z(n543) );
  XOR U51 ( .A(a[147]), .B(n529), .Z(n531) );
  XOR U52 ( .A(a[150]), .B(n516), .Z(n518) );
  XOR U53 ( .A(a[153]), .B(n504), .Z(n506) );
  XOR U54 ( .A(a[156]), .B(n492), .Z(n494) );
  XOR U55 ( .A(a[159]), .B(n479), .Z(n481) );
  XOR U56 ( .A(a[162]), .B(n467), .Z(n469) );
  XOR U57 ( .A(a[165]), .B(n455), .Z(n457) );
  XOR U58 ( .A(a[168]), .B(n443), .Z(n445) );
  XOR U59 ( .A(a[171]), .B(n430), .Z(n432) );
  XOR U60 ( .A(a[174]), .B(n418), .Z(n420) );
  XOR U61 ( .A(a[177]), .B(n406), .Z(n408) );
  XOR U62 ( .A(a[180]), .B(n393), .Z(n395) );
  XOR U63 ( .A(a[183]), .B(n381), .Z(n383) );
  XOR U64 ( .A(a[186]), .B(n369), .Z(n371) );
  XOR U65 ( .A(a[189]), .B(n356), .Z(n358) );
  XOR U66 ( .A(a[192]), .B(n344), .Z(n346) );
  XOR U67 ( .A(a[195]), .B(n332), .Z(n334) );
  XOR U68 ( .A(a[198]), .B(n320), .Z(n322) );
  XOR U69 ( .A(a[201]), .B(n306), .Z(n308) );
  XOR U70 ( .A(a[204]), .B(n294), .Z(n296) );
  XOR U71 ( .A(a[207]), .B(n282), .Z(n284) );
  XOR U72 ( .A(a[210]), .B(n269), .Z(n271) );
  XOR U73 ( .A(a[213]), .B(n257), .Z(n259) );
  XOR U74 ( .A(a[216]), .B(n245), .Z(n247) );
  XOR U75 ( .A(a[219]), .B(n232), .Z(n234) );
  XOR U76 ( .A(a[222]), .B(n220), .Z(n222) );
  XOR U77 ( .A(a[225]), .B(n208), .Z(n210) );
  XOR U78 ( .A(a[228]), .B(n196), .Z(n198) );
  XOR U79 ( .A(a[231]), .B(n183), .Z(n185) );
  XOR U80 ( .A(a[234]), .B(n171), .Z(n173) );
  XOR U81 ( .A(a[237]), .B(n159), .Z(n161) );
  XOR U82 ( .A(a[240]), .B(n146), .Z(n148) );
  XOR U83 ( .A(a[243]), .B(n134), .Z(n136) );
  XOR U84 ( .A(a[246]), .B(n122), .Z(n124) );
  XOR U85 ( .A(a[249]), .B(n109), .Z(n111) );
  XOR U86 ( .A(a[252]), .B(n97), .Z(n99) );
  XOR U87 ( .A(a[1]), .B(n1019), .Z(n317) );
  XOR U88 ( .A(a[4]), .B(n1010), .Z(n60) );
  XOR U89 ( .A(a[7]), .B(n1001), .Z(n27) );
  XOR U90 ( .A(a[10]), .B(n992), .Z(n687) );
  XOR U91 ( .A(a[13]), .B(n983), .Z(n564) );
  XOR U92 ( .A(a[16]), .B(n974), .Z(n441) );
  XOR U93 ( .A(a[19]), .B(n965), .Z(n318) );
  XOR U94 ( .A(a[22]), .B(n956), .Z(n194) );
  XOR U95 ( .A(a[25]), .B(n947), .Z(n87) );
  XOR U96 ( .A(a[28]), .B(n938), .Z(n84) );
  XOR U97 ( .A(a[31]), .B(n929), .Z(n80) );
  XOR U98 ( .A(a[34]), .B(n920), .Z(n77) );
  XOR U99 ( .A(a[37]), .B(n911), .Z(n74) );
  XOR U100 ( .A(a[40]), .B(n902), .Z(n70) );
  XOR U101 ( .A(a[43]), .B(n893), .Z(n67) );
  XOR U102 ( .A(a[46]), .B(n884), .Z(n64) );
  XOR U103 ( .A(a[49]), .B(n875), .Z(n61) );
  XOR U104 ( .A(a[52]), .B(n866), .Z(n57) );
  XOR U105 ( .A(a[55]), .B(n857), .Z(n54) );
  XOR U106 ( .A(a[58]), .B(n848), .Z(n51) );
  XOR U107 ( .A(a[61]), .B(n839), .Z(n47) );
  XOR U108 ( .A(a[64]), .B(n830), .Z(n44) );
  XOR U109 ( .A(a[67]), .B(n821), .Z(n41) );
  XOR U110 ( .A(a[70]), .B(n812), .Z(n37) );
  XOR U111 ( .A(a[73]), .B(n803), .Z(n34) );
  XOR U112 ( .A(a[76]), .B(n794), .Z(n31) );
  XOR U113 ( .A(a[79]), .B(n785), .Z(n28) );
  XOR U114 ( .A(a[82]), .B(n776), .Z(n24) );
  XOR U115 ( .A(a[85]), .B(n767), .Z(n21) );
  XOR U116 ( .A(a[88]), .B(n758), .Z(n18) );
  XOR U117 ( .A(a[91]), .B(n749), .Z(n14) );
  XOR U118 ( .A(a[94]), .B(n740), .Z(n11) );
  XOR U119 ( .A(a[97]), .B(n731), .Z(n8) );
  XOR U120 ( .A(a[100]), .B(n721), .Z(n723) );
  XOR U121 ( .A(a[103]), .B(n709), .Z(n711) );
  XOR U122 ( .A(a[106]), .B(n697), .Z(n699) );
  XOR U123 ( .A(a[109]), .B(n684), .Z(n686) );
  XOR U124 ( .A(a[112]), .B(n672), .Z(n674) );
  XOR U125 ( .A(a[115]), .B(n660), .Z(n662) );
  XOR U126 ( .A(a[118]), .B(n648), .Z(n650) );
  XOR U127 ( .A(a[121]), .B(n635), .Z(n637) );
  XOR U128 ( .A(a[124]), .B(n623), .Z(n625) );
  XOR U129 ( .A(a[127]), .B(n611), .Z(n613) );
  XOR U130 ( .A(a[130]), .B(n598), .Z(n600) );
  XOR U131 ( .A(a[133]), .B(n586), .Z(n588) );
  XOR U132 ( .A(a[136]), .B(n574), .Z(n576) );
  XOR U133 ( .A(a[139]), .B(n561), .Z(n563) );
  XOR U134 ( .A(a[142]), .B(n549), .Z(n551) );
  XOR U135 ( .A(a[145]), .B(n537), .Z(n539) );
  XOR U136 ( .A(a[148]), .B(n525), .Z(n527) );
  XOR U137 ( .A(a[151]), .B(n512), .Z(n514) );
  XOR U138 ( .A(a[154]), .B(n500), .Z(n502) );
  XOR U139 ( .A(a[157]), .B(n488), .Z(n490) );
  XOR U140 ( .A(a[160]), .B(n475), .Z(n477) );
  XOR U141 ( .A(a[163]), .B(n463), .Z(n465) );
  XOR U142 ( .A(a[166]), .B(n451), .Z(n453) );
  XOR U143 ( .A(a[169]), .B(n438), .Z(n440) );
  XOR U144 ( .A(a[172]), .B(n426), .Z(n428) );
  XOR U145 ( .A(a[175]), .B(n414), .Z(n416) );
  XOR U146 ( .A(a[178]), .B(n402), .Z(n404) );
  XOR U147 ( .A(a[181]), .B(n389), .Z(n391) );
  XOR U148 ( .A(a[184]), .B(n377), .Z(n379) );
  XOR U149 ( .A(a[187]), .B(n365), .Z(n367) );
  XOR U150 ( .A(a[190]), .B(n352), .Z(n354) );
  XOR U151 ( .A(a[193]), .B(n340), .Z(n342) );
  XOR U152 ( .A(a[196]), .B(n328), .Z(n330) );
  XOR U153 ( .A(a[199]), .B(n314), .Z(n316) );
  XOR U154 ( .A(a[202]), .B(n302), .Z(n304) );
  XOR U155 ( .A(a[205]), .B(n290), .Z(n292) );
  XOR U156 ( .A(a[208]), .B(n278), .Z(n280) );
  XOR U157 ( .A(a[211]), .B(n265), .Z(n267) );
  XOR U158 ( .A(a[214]), .B(n253), .Z(n255) );
  XOR U159 ( .A(a[217]), .B(n241), .Z(n243) );
  XOR U160 ( .A(a[220]), .B(n228), .Z(n230) );
  XOR U161 ( .A(a[223]), .B(n216), .Z(n218) );
  XOR U162 ( .A(a[226]), .B(n204), .Z(n206) );
  XOR U163 ( .A(a[229]), .B(n191), .Z(n193) );
  XOR U164 ( .A(a[232]), .B(n179), .Z(n181) );
  XOR U165 ( .A(a[235]), .B(n167), .Z(n169) );
  XOR U166 ( .A(a[238]), .B(n155), .Z(n157) );
  XOR U167 ( .A(a[241]), .B(n142), .Z(n144) );
  XOR U168 ( .A(a[244]), .B(n130), .Z(n132) );
  XOR U169 ( .A(a[247]), .B(n118), .Z(n120) );
  XOR U170 ( .A(a[250]), .B(n105), .Z(n107) );
  XOR U171 ( .A(a[253]), .B(n93), .Z(n95) );
  XOR U172 ( .A(a[2]), .B(n1016), .Z(n82) );
  XOR U173 ( .A(a[5]), .B(n1007), .Z(n49) );
  XOR U174 ( .A(a[8]), .B(n998), .Z(n16) );
  XOR U175 ( .A(a[11]), .B(n989), .Z(n646) );
  XOR U176 ( .A(a[14]), .B(n980), .Z(n523) );
  XOR U177 ( .A(a[17]), .B(n971), .Z(n400) );
  XOR U178 ( .A(a[20]), .B(n962), .Z(n276) );
  XOR U179 ( .A(a[23]), .B(n953), .Z(n153) );
  XOR U180 ( .A(a[26]), .B(n944), .Z(n86) );
  XOR U181 ( .A(a[29]), .B(n935), .Z(n83) );
  XOR U182 ( .A(a[32]), .B(n926), .Z(n79) );
  XOR U183 ( .A(a[35]), .B(n917), .Z(n76) );
  XOR U184 ( .A(a[38]), .B(n908), .Z(n73) );
  XOR U185 ( .A(a[41]), .B(n899), .Z(n69) );
  XOR U186 ( .A(a[44]), .B(n890), .Z(n66) );
  XOR U187 ( .A(a[47]), .B(n881), .Z(n63) );
  XOR U188 ( .A(a[50]), .B(n872), .Z(n59) );
  XOR U189 ( .A(a[53]), .B(n863), .Z(n56) );
  XOR U190 ( .A(a[56]), .B(n854), .Z(n53) );
  XOR U191 ( .A(a[59]), .B(n845), .Z(n50) );
  XOR U192 ( .A(a[62]), .B(n836), .Z(n46) );
  XOR U193 ( .A(a[65]), .B(n827), .Z(n43) );
  XOR U194 ( .A(a[68]), .B(n818), .Z(n40) );
  XOR U195 ( .A(a[71]), .B(n809), .Z(n36) );
  XOR U196 ( .A(a[74]), .B(n800), .Z(n33) );
  XOR U197 ( .A(a[77]), .B(n791), .Z(n30) );
  XOR U198 ( .A(a[80]), .B(n782), .Z(n26) );
  XOR U199 ( .A(a[83]), .B(n773), .Z(n23) );
  XOR U200 ( .A(a[86]), .B(n764), .Z(n20) );
  XOR U201 ( .A(a[89]), .B(n755), .Z(n17) );
  XOR U202 ( .A(a[92]), .B(n746), .Z(n13) );
  XOR U203 ( .A(a[95]), .B(n737), .Z(n10) );
  XOR U204 ( .A(a[98]), .B(n728), .Z(n7) );
  XOR U205 ( .A(a[101]), .B(n717), .Z(n719) );
  XOR U206 ( .A(a[104]), .B(n705), .Z(n707) );
  XOR U207 ( .A(a[107]), .B(n693), .Z(n695) );
  XOR U208 ( .A(a[110]), .B(n680), .Z(n682) );
  XOR U209 ( .A(a[113]), .B(n668), .Z(n670) );
  XOR U210 ( .A(a[116]), .B(n656), .Z(n658) );
  XOR U211 ( .A(a[119]), .B(n643), .Z(n645) );
  XOR U212 ( .A(a[122]), .B(n631), .Z(n633) );
  XOR U213 ( .A(a[125]), .B(n619), .Z(n621) );
  XOR U214 ( .A(a[128]), .B(n607), .Z(n609) );
  XOR U215 ( .A(a[131]), .B(n594), .Z(n596) );
  XOR U216 ( .A(a[134]), .B(n582), .Z(n584) );
  XOR U217 ( .A(a[137]), .B(n570), .Z(n572) );
  XOR U218 ( .A(a[140]), .B(n557), .Z(n559) );
  XOR U219 ( .A(a[143]), .B(n545), .Z(n547) );
  XOR U220 ( .A(a[146]), .B(n533), .Z(n535) );
  XOR U221 ( .A(a[149]), .B(n520), .Z(n522) );
  XOR U222 ( .A(a[152]), .B(n508), .Z(n510) );
  XOR U223 ( .A(a[155]), .B(n496), .Z(n498) );
  XOR U224 ( .A(a[158]), .B(n484), .Z(n486) );
  XOR U225 ( .A(a[161]), .B(n471), .Z(n473) );
  XOR U226 ( .A(a[164]), .B(n459), .Z(n461) );
  XOR U227 ( .A(a[167]), .B(n447), .Z(n449) );
  XOR U228 ( .A(a[170]), .B(n434), .Z(n436) );
  XOR U229 ( .A(a[173]), .B(n422), .Z(n424) );
  XOR U230 ( .A(a[176]), .B(n410), .Z(n412) );
  XOR U231 ( .A(a[179]), .B(n397), .Z(n399) );
  XOR U232 ( .A(a[182]), .B(n385), .Z(n387) );
  XOR U233 ( .A(a[185]), .B(n373), .Z(n375) );
  XOR U234 ( .A(a[188]), .B(n361), .Z(n363) );
  XOR U235 ( .A(a[191]), .B(n348), .Z(n350) );
  XOR U236 ( .A(a[194]), .B(n336), .Z(n338) );
  XOR U237 ( .A(a[197]), .B(n324), .Z(n326) );
  XOR U238 ( .A(a[200]), .B(n310), .Z(n312) );
  XOR U239 ( .A(a[203]), .B(n298), .Z(n300) );
  XOR U240 ( .A(a[206]), .B(n286), .Z(n288) );
  XOR U241 ( .A(a[209]), .B(n273), .Z(n275) );
  XOR U242 ( .A(a[212]), .B(n261), .Z(n263) );
  XOR U243 ( .A(a[215]), .B(n249), .Z(n251) );
  XOR U244 ( .A(a[218]), .B(n237), .Z(n239) );
  XOR U245 ( .A(a[221]), .B(n224), .Z(n226) );
  XOR U246 ( .A(a[224]), .B(n212), .Z(n214) );
  XOR U247 ( .A(a[227]), .B(n200), .Z(n202) );
  XOR U248 ( .A(a[230]), .B(n187), .Z(n189) );
  XOR U249 ( .A(a[233]), .B(n175), .Z(n177) );
  XOR U250 ( .A(a[236]), .B(n163), .Z(n165) );
  XOR U251 ( .A(a[239]), .B(n150), .Z(n152) );
  XOR U252 ( .A(a[242]), .B(n138), .Z(n140) );
  XOR U253 ( .A(a[245]), .B(n126), .Z(n128) );
  XOR U254 ( .A(a[248]), .B(n114), .Z(n116) );
  XOR U255 ( .A(a[251]), .B(n101), .Z(n103) );
  XOR U256 ( .A(a[254]), .B(n89), .Z(n91) );
  XOR U257 ( .A(n1), .B(n2), .Z(carry_on_d) );
  ANDN U258 ( .B(n3), .A(n4), .Z(n1) );
  XOR U259 ( .A(b[255]), .B(n2), .Z(n3) );
  XNOR U260 ( .A(b[9]), .B(n5), .Z(c[9]) );
  XNOR U261 ( .A(b[99]), .B(n6), .Z(c[99]) );
  XNOR U262 ( .A(b[98]), .B(n7), .Z(c[98]) );
  XNOR U263 ( .A(b[97]), .B(n8), .Z(c[97]) );
  XNOR U264 ( .A(b[96]), .B(n9), .Z(c[96]) );
  XNOR U265 ( .A(b[95]), .B(n10), .Z(c[95]) );
  XNOR U266 ( .A(b[94]), .B(n11), .Z(c[94]) );
  XNOR U267 ( .A(b[93]), .B(n12), .Z(c[93]) );
  XNOR U268 ( .A(b[92]), .B(n13), .Z(c[92]) );
  XNOR U269 ( .A(b[91]), .B(n14), .Z(c[91]) );
  XNOR U270 ( .A(b[90]), .B(n15), .Z(c[90]) );
  XNOR U271 ( .A(b[8]), .B(n16), .Z(c[8]) );
  XNOR U272 ( .A(b[89]), .B(n17), .Z(c[89]) );
  XNOR U273 ( .A(b[88]), .B(n18), .Z(c[88]) );
  XNOR U274 ( .A(b[87]), .B(n19), .Z(c[87]) );
  XNOR U275 ( .A(b[86]), .B(n20), .Z(c[86]) );
  XNOR U276 ( .A(b[85]), .B(n21), .Z(c[85]) );
  XNOR U277 ( .A(b[84]), .B(n22), .Z(c[84]) );
  XNOR U278 ( .A(b[83]), .B(n23), .Z(c[83]) );
  XNOR U279 ( .A(b[82]), .B(n24), .Z(c[82]) );
  XNOR U280 ( .A(b[81]), .B(n25), .Z(c[81]) );
  XNOR U281 ( .A(b[80]), .B(n26), .Z(c[80]) );
  XNOR U282 ( .A(b[7]), .B(n27), .Z(c[7]) );
  XNOR U283 ( .A(b[79]), .B(n28), .Z(c[79]) );
  XNOR U284 ( .A(b[78]), .B(n29), .Z(c[78]) );
  XNOR U285 ( .A(b[77]), .B(n30), .Z(c[77]) );
  XNOR U286 ( .A(b[76]), .B(n31), .Z(c[76]) );
  XNOR U287 ( .A(b[75]), .B(n32), .Z(c[75]) );
  XNOR U288 ( .A(b[74]), .B(n33), .Z(c[74]) );
  XNOR U289 ( .A(b[73]), .B(n34), .Z(c[73]) );
  XNOR U290 ( .A(b[72]), .B(n35), .Z(c[72]) );
  XNOR U291 ( .A(b[71]), .B(n36), .Z(c[71]) );
  XNOR U292 ( .A(b[70]), .B(n37), .Z(c[70]) );
  XNOR U293 ( .A(b[6]), .B(n38), .Z(c[6]) );
  XNOR U294 ( .A(b[69]), .B(n39), .Z(c[69]) );
  XNOR U295 ( .A(b[68]), .B(n40), .Z(c[68]) );
  XNOR U296 ( .A(b[67]), .B(n41), .Z(c[67]) );
  XNOR U297 ( .A(b[66]), .B(n42), .Z(c[66]) );
  XNOR U298 ( .A(b[65]), .B(n43), .Z(c[65]) );
  XNOR U299 ( .A(b[64]), .B(n44), .Z(c[64]) );
  XNOR U300 ( .A(b[63]), .B(n45), .Z(c[63]) );
  XNOR U301 ( .A(b[62]), .B(n46), .Z(c[62]) );
  XNOR U302 ( .A(b[61]), .B(n47), .Z(c[61]) );
  XNOR U303 ( .A(b[60]), .B(n48), .Z(c[60]) );
  XNOR U304 ( .A(b[5]), .B(n49), .Z(c[5]) );
  XNOR U305 ( .A(b[59]), .B(n50), .Z(c[59]) );
  XNOR U306 ( .A(b[58]), .B(n51), .Z(c[58]) );
  XNOR U307 ( .A(b[57]), .B(n52), .Z(c[57]) );
  XNOR U308 ( .A(b[56]), .B(n53), .Z(c[56]) );
  XNOR U309 ( .A(b[55]), .B(n54), .Z(c[55]) );
  XNOR U310 ( .A(b[54]), .B(n55), .Z(c[54]) );
  XNOR U311 ( .A(b[53]), .B(n56), .Z(c[53]) );
  XNOR U312 ( .A(b[52]), .B(n57), .Z(c[52]) );
  XNOR U313 ( .A(b[51]), .B(n58), .Z(c[51]) );
  XNOR U314 ( .A(b[50]), .B(n59), .Z(c[50]) );
  XNOR U315 ( .A(b[4]), .B(n60), .Z(c[4]) );
  XNOR U316 ( .A(b[49]), .B(n61), .Z(c[49]) );
  XNOR U317 ( .A(b[48]), .B(n62), .Z(c[48]) );
  XNOR U318 ( .A(b[47]), .B(n63), .Z(c[47]) );
  XNOR U319 ( .A(b[46]), .B(n64), .Z(c[46]) );
  XNOR U320 ( .A(b[45]), .B(n65), .Z(c[45]) );
  XNOR U321 ( .A(b[44]), .B(n66), .Z(c[44]) );
  XNOR U322 ( .A(b[43]), .B(n67), .Z(c[43]) );
  XNOR U323 ( .A(b[42]), .B(n68), .Z(c[42]) );
  XNOR U324 ( .A(b[41]), .B(n69), .Z(c[41]) );
  XNOR U325 ( .A(b[40]), .B(n70), .Z(c[40]) );
  XNOR U326 ( .A(b[3]), .B(n71), .Z(c[3]) );
  XNOR U327 ( .A(b[39]), .B(n72), .Z(c[39]) );
  XNOR U328 ( .A(b[38]), .B(n73), .Z(c[38]) );
  XNOR U329 ( .A(b[37]), .B(n74), .Z(c[37]) );
  XNOR U330 ( .A(b[36]), .B(n75), .Z(c[36]) );
  XNOR U331 ( .A(b[35]), .B(n76), .Z(c[35]) );
  XNOR U332 ( .A(b[34]), .B(n77), .Z(c[34]) );
  XNOR U333 ( .A(b[33]), .B(n78), .Z(c[33]) );
  XNOR U334 ( .A(b[32]), .B(n79), .Z(c[32]) );
  XNOR U335 ( .A(b[31]), .B(n80), .Z(c[31]) );
  XNOR U336 ( .A(b[30]), .B(n81), .Z(c[30]) );
  XNOR U337 ( .A(b[2]), .B(n82), .Z(c[2]) );
  XNOR U338 ( .A(b[29]), .B(n83), .Z(c[29]) );
  XNOR U339 ( .A(b[28]), .B(n84), .Z(c[28]) );
  XNOR U340 ( .A(b[27]), .B(n85), .Z(c[27]) );
  XNOR U341 ( .A(b[26]), .B(n86), .Z(c[26]) );
  XNOR U342 ( .A(b[25]), .B(n87), .Z(c[25]) );
  XNOR U343 ( .A(b[255]), .B(n4), .Z(c[255]) );
  XNOR U344 ( .A(a[255]), .B(n2), .Z(n4) );
  XNOR U345 ( .A(n88), .B(n89), .Z(n2) );
  ANDN U346 ( .B(n90), .A(n91), .Z(n88) );
  XNOR U347 ( .A(b[254]), .B(n89), .Z(n90) );
  XNOR U348 ( .A(b[254]), .B(n91), .Z(c[254]) );
  XOR U349 ( .A(n92), .B(n93), .Z(n89) );
  ANDN U350 ( .B(n94), .A(n95), .Z(n92) );
  XNOR U351 ( .A(b[253]), .B(n93), .Z(n94) );
  XNOR U352 ( .A(b[253]), .B(n95), .Z(c[253]) );
  XOR U353 ( .A(n96), .B(n97), .Z(n93) );
  ANDN U354 ( .B(n98), .A(n99), .Z(n96) );
  XNOR U355 ( .A(b[252]), .B(n97), .Z(n98) );
  XNOR U356 ( .A(b[252]), .B(n99), .Z(c[252]) );
  XOR U357 ( .A(n100), .B(n101), .Z(n97) );
  ANDN U358 ( .B(n102), .A(n103), .Z(n100) );
  XNOR U359 ( .A(b[251]), .B(n101), .Z(n102) );
  XNOR U360 ( .A(b[251]), .B(n103), .Z(c[251]) );
  XOR U361 ( .A(n104), .B(n105), .Z(n101) );
  ANDN U362 ( .B(n106), .A(n107), .Z(n104) );
  XNOR U363 ( .A(b[250]), .B(n105), .Z(n106) );
  XNOR U364 ( .A(b[250]), .B(n107), .Z(c[250]) );
  XOR U365 ( .A(n108), .B(n109), .Z(n105) );
  ANDN U366 ( .B(n110), .A(n111), .Z(n108) );
  XNOR U367 ( .A(b[249]), .B(n109), .Z(n110) );
  XNOR U368 ( .A(b[24]), .B(n112), .Z(c[24]) );
  XNOR U369 ( .A(b[249]), .B(n111), .Z(c[249]) );
  XOR U370 ( .A(n113), .B(n114), .Z(n109) );
  ANDN U371 ( .B(n115), .A(n116), .Z(n113) );
  XNOR U372 ( .A(b[248]), .B(n114), .Z(n115) );
  XNOR U373 ( .A(b[248]), .B(n116), .Z(c[248]) );
  XOR U374 ( .A(n117), .B(n118), .Z(n114) );
  ANDN U375 ( .B(n119), .A(n120), .Z(n117) );
  XNOR U376 ( .A(b[247]), .B(n118), .Z(n119) );
  XNOR U377 ( .A(b[247]), .B(n120), .Z(c[247]) );
  XOR U378 ( .A(n121), .B(n122), .Z(n118) );
  ANDN U379 ( .B(n123), .A(n124), .Z(n121) );
  XNOR U380 ( .A(b[246]), .B(n122), .Z(n123) );
  XNOR U381 ( .A(b[246]), .B(n124), .Z(c[246]) );
  XOR U382 ( .A(n125), .B(n126), .Z(n122) );
  ANDN U383 ( .B(n127), .A(n128), .Z(n125) );
  XNOR U384 ( .A(b[245]), .B(n126), .Z(n127) );
  XNOR U385 ( .A(b[245]), .B(n128), .Z(c[245]) );
  XOR U386 ( .A(n129), .B(n130), .Z(n126) );
  ANDN U387 ( .B(n131), .A(n132), .Z(n129) );
  XNOR U388 ( .A(b[244]), .B(n130), .Z(n131) );
  XNOR U389 ( .A(b[244]), .B(n132), .Z(c[244]) );
  XOR U390 ( .A(n133), .B(n134), .Z(n130) );
  ANDN U391 ( .B(n135), .A(n136), .Z(n133) );
  XNOR U392 ( .A(b[243]), .B(n134), .Z(n135) );
  XNOR U393 ( .A(b[243]), .B(n136), .Z(c[243]) );
  XOR U394 ( .A(n137), .B(n138), .Z(n134) );
  ANDN U395 ( .B(n139), .A(n140), .Z(n137) );
  XNOR U396 ( .A(b[242]), .B(n138), .Z(n139) );
  XNOR U397 ( .A(b[242]), .B(n140), .Z(c[242]) );
  XOR U398 ( .A(n141), .B(n142), .Z(n138) );
  ANDN U399 ( .B(n143), .A(n144), .Z(n141) );
  XNOR U400 ( .A(b[241]), .B(n142), .Z(n143) );
  XNOR U401 ( .A(b[241]), .B(n144), .Z(c[241]) );
  XOR U402 ( .A(n145), .B(n146), .Z(n142) );
  ANDN U403 ( .B(n147), .A(n148), .Z(n145) );
  XNOR U404 ( .A(b[240]), .B(n146), .Z(n147) );
  XNOR U405 ( .A(b[240]), .B(n148), .Z(c[240]) );
  XOR U406 ( .A(n149), .B(n150), .Z(n146) );
  ANDN U407 ( .B(n151), .A(n152), .Z(n149) );
  XNOR U408 ( .A(b[239]), .B(n150), .Z(n151) );
  XNOR U409 ( .A(b[23]), .B(n153), .Z(c[23]) );
  XNOR U410 ( .A(b[239]), .B(n152), .Z(c[239]) );
  XOR U411 ( .A(n154), .B(n155), .Z(n150) );
  ANDN U412 ( .B(n156), .A(n157), .Z(n154) );
  XNOR U413 ( .A(b[238]), .B(n155), .Z(n156) );
  XNOR U414 ( .A(b[238]), .B(n157), .Z(c[238]) );
  XOR U415 ( .A(n158), .B(n159), .Z(n155) );
  ANDN U416 ( .B(n160), .A(n161), .Z(n158) );
  XNOR U417 ( .A(b[237]), .B(n159), .Z(n160) );
  XNOR U418 ( .A(b[237]), .B(n161), .Z(c[237]) );
  XOR U419 ( .A(n162), .B(n163), .Z(n159) );
  ANDN U420 ( .B(n164), .A(n165), .Z(n162) );
  XNOR U421 ( .A(b[236]), .B(n163), .Z(n164) );
  XNOR U422 ( .A(b[236]), .B(n165), .Z(c[236]) );
  XOR U423 ( .A(n166), .B(n167), .Z(n163) );
  ANDN U424 ( .B(n168), .A(n169), .Z(n166) );
  XNOR U425 ( .A(b[235]), .B(n167), .Z(n168) );
  XNOR U426 ( .A(b[235]), .B(n169), .Z(c[235]) );
  XOR U427 ( .A(n170), .B(n171), .Z(n167) );
  ANDN U428 ( .B(n172), .A(n173), .Z(n170) );
  XNOR U429 ( .A(b[234]), .B(n171), .Z(n172) );
  XNOR U430 ( .A(b[234]), .B(n173), .Z(c[234]) );
  XOR U431 ( .A(n174), .B(n175), .Z(n171) );
  ANDN U432 ( .B(n176), .A(n177), .Z(n174) );
  XNOR U433 ( .A(b[233]), .B(n175), .Z(n176) );
  XNOR U434 ( .A(b[233]), .B(n177), .Z(c[233]) );
  XOR U435 ( .A(n178), .B(n179), .Z(n175) );
  ANDN U436 ( .B(n180), .A(n181), .Z(n178) );
  XNOR U437 ( .A(b[232]), .B(n179), .Z(n180) );
  XNOR U438 ( .A(b[232]), .B(n181), .Z(c[232]) );
  XOR U439 ( .A(n182), .B(n183), .Z(n179) );
  ANDN U440 ( .B(n184), .A(n185), .Z(n182) );
  XNOR U441 ( .A(b[231]), .B(n183), .Z(n184) );
  XNOR U442 ( .A(b[231]), .B(n185), .Z(c[231]) );
  XOR U443 ( .A(n186), .B(n187), .Z(n183) );
  ANDN U444 ( .B(n188), .A(n189), .Z(n186) );
  XNOR U445 ( .A(b[230]), .B(n187), .Z(n188) );
  XNOR U446 ( .A(b[230]), .B(n189), .Z(c[230]) );
  XOR U447 ( .A(n190), .B(n191), .Z(n187) );
  ANDN U448 ( .B(n192), .A(n193), .Z(n190) );
  XNOR U449 ( .A(b[229]), .B(n191), .Z(n192) );
  XNOR U450 ( .A(b[22]), .B(n194), .Z(c[22]) );
  XNOR U451 ( .A(b[229]), .B(n193), .Z(c[229]) );
  XOR U452 ( .A(n195), .B(n196), .Z(n191) );
  ANDN U453 ( .B(n197), .A(n198), .Z(n195) );
  XNOR U454 ( .A(b[228]), .B(n196), .Z(n197) );
  XNOR U455 ( .A(b[228]), .B(n198), .Z(c[228]) );
  XOR U456 ( .A(n199), .B(n200), .Z(n196) );
  ANDN U457 ( .B(n201), .A(n202), .Z(n199) );
  XNOR U458 ( .A(b[227]), .B(n200), .Z(n201) );
  XNOR U459 ( .A(b[227]), .B(n202), .Z(c[227]) );
  XOR U460 ( .A(n203), .B(n204), .Z(n200) );
  ANDN U461 ( .B(n205), .A(n206), .Z(n203) );
  XNOR U462 ( .A(b[226]), .B(n204), .Z(n205) );
  XNOR U463 ( .A(b[226]), .B(n206), .Z(c[226]) );
  XOR U464 ( .A(n207), .B(n208), .Z(n204) );
  ANDN U465 ( .B(n209), .A(n210), .Z(n207) );
  XNOR U466 ( .A(b[225]), .B(n208), .Z(n209) );
  XNOR U467 ( .A(b[225]), .B(n210), .Z(c[225]) );
  XOR U468 ( .A(n211), .B(n212), .Z(n208) );
  ANDN U469 ( .B(n213), .A(n214), .Z(n211) );
  XNOR U470 ( .A(b[224]), .B(n212), .Z(n213) );
  XNOR U471 ( .A(b[224]), .B(n214), .Z(c[224]) );
  XOR U472 ( .A(n215), .B(n216), .Z(n212) );
  ANDN U473 ( .B(n217), .A(n218), .Z(n215) );
  XNOR U474 ( .A(b[223]), .B(n216), .Z(n217) );
  XNOR U475 ( .A(b[223]), .B(n218), .Z(c[223]) );
  XOR U476 ( .A(n219), .B(n220), .Z(n216) );
  ANDN U477 ( .B(n221), .A(n222), .Z(n219) );
  XNOR U478 ( .A(b[222]), .B(n220), .Z(n221) );
  XNOR U479 ( .A(b[222]), .B(n222), .Z(c[222]) );
  XOR U480 ( .A(n223), .B(n224), .Z(n220) );
  ANDN U481 ( .B(n225), .A(n226), .Z(n223) );
  XNOR U482 ( .A(b[221]), .B(n224), .Z(n225) );
  XNOR U483 ( .A(b[221]), .B(n226), .Z(c[221]) );
  XOR U484 ( .A(n227), .B(n228), .Z(n224) );
  ANDN U485 ( .B(n229), .A(n230), .Z(n227) );
  XNOR U486 ( .A(b[220]), .B(n228), .Z(n229) );
  XNOR U487 ( .A(b[220]), .B(n230), .Z(c[220]) );
  XOR U488 ( .A(n231), .B(n232), .Z(n228) );
  ANDN U489 ( .B(n233), .A(n234), .Z(n231) );
  XNOR U490 ( .A(b[219]), .B(n232), .Z(n233) );
  XNOR U491 ( .A(b[21]), .B(n235), .Z(c[21]) );
  XNOR U492 ( .A(b[219]), .B(n234), .Z(c[219]) );
  XOR U493 ( .A(n236), .B(n237), .Z(n232) );
  ANDN U494 ( .B(n238), .A(n239), .Z(n236) );
  XNOR U495 ( .A(b[218]), .B(n237), .Z(n238) );
  XNOR U496 ( .A(b[218]), .B(n239), .Z(c[218]) );
  XOR U497 ( .A(n240), .B(n241), .Z(n237) );
  ANDN U498 ( .B(n242), .A(n243), .Z(n240) );
  XNOR U499 ( .A(b[217]), .B(n241), .Z(n242) );
  XNOR U500 ( .A(b[217]), .B(n243), .Z(c[217]) );
  XOR U501 ( .A(n244), .B(n245), .Z(n241) );
  ANDN U502 ( .B(n246), .A(n247), .Z(n244) );
  XNOR U503 ( .A(b[216]), .B(n245), .Z(n246) );
  XNOR U504 ( .A(b[216]), .B(n247), .Z(c[216]) );
  XOR U505 ( .A(n248), .B(n249), .Z(n245) );
  ANDN U506 ( .B(n250), .A(n251), .Z(n248) );
  XNOR U507 ( .A(b[215]), .B(n249), .Z(n250) );
  XNOR U508 ( .A(b[215]), .B(n251), .Z(c[215]) );
  XOR U509 ( .A(n252), .B(n253), .Z(n249) );
  ANDN U510 ( .B(n254), .A(n255), .Z(n252) );
  XNOR U511 ( .A(b[214]), .B(n253), .Z(n254) );
  XNOR U512 ( .A(b[214]), .B(n255), .Z(c[214]) );
  XOR U513 ( .A(n256), .B(n257), .Z(n253) );
  ANDN U514 ( .B(n258), .A(n259), .Z(n256) );
  XNOR U515 ( .A(b[213]), .B(n257), .Z(n258) );
  XNOR U516 ( .A(b[213]), .B(n259), .Z(c[213]) );
  XOR U517 ( .A(n260), .B(n261), .Z(n257) );
  ANDN U518 ( .B(n262), .A(n263), .Z(n260) );
  XNOR U519 ( .A(b[212]), .B(n261), .Z(n262) );
  XNOR U520 ( .A(b[212]), .B(n263), .Z(c[212]) );
  XOR U521 ( .A(n264), .B(n265), .Z(n261) );
  ANDN U522 ( .B(n266), .A(n267), .Z(n264) );
  XNOR U523 ( .A(b[211]), .B(n265), .Z(n266) );
  XNOR U524 ( .A(b[211]), .B(n267), .Z(c[211]) );
  XOR U525 ( .A(n268), .B(n269), .Z(n265) );
  ANDN U526 ( .B(n270), .A(n271), .Z(n268) );
  XNOR U527 ( .A(b[210]), .B(n269), .Z(n270) );
  XNOR U528 ( .A(b[210]), .B(n271), .Z(c[210]) );
  XOR U529 ( .A(n272), .B(n273), .Z(n269) );
  ANDN U530 ( .B(n274), .A(n275), .Z(n272) );
  XNOR U531 ( .A(b[209]), .B(n273), .Z(n274) );
  XNOR U532 ( .A(b[20]), .B(n276), .Z(c[20]) );
  XNOR U533 ( .A(b[209]), .B(n275), .Z(c[209]) );
  XOR U534 ( .A(n277), .B(n278), .Z(n273) );
  ANDN U535 ( .B(n279), .A(n280), .Z(n277) );
  XNOR U536 ( .A(b[208]), .B(n278), .Z(n279) );
  XNOR U537 ( .A(b[208]), .B(n280), .Z(c[208]) );
  XOR U538 ( .A(n281), .B(n282), .Z(n278) );
  ANDN U539 ( .B(n283), .A(n284), .Z(n281) );
  XNOR U540 ( .A(b[207]), .B(n282), .Z(n283) );
  XNOR U541 ( .A(b[207]), .B(n284), .Z(c[207]) );
  XOR U542 ( .A(n285), .B(n286), .Z(n282) );
  ANDN U543 ( .B(n287), .A(n288), .Z(n285) );
  XNOR U544 ( .A(b[206]), .B(n286), .Z(n287) );
  XNOR U545 ( .A(b[206]), .B(n288), .Z(c[206]) );
  XOR U546 ( .A(n289), .B(n290), .Z(n286) );
  ANDN U547 ( .B(n291), .A(n292), .Z(n289) );
  XNOR U548 ( .A(b[205]), .B(n290), .Z(n291) );
  XNOR U549 ( .A(b[205]), .B(n292), .Z(c[205]) );
  XOR U550 ( .A(n293), .B(n294), .Z(n290) );
  ANDN U551 ( .B(n295), .A(n296), .Z(n293) );
  XNOR U552 ( .A(b[204]), .B(n294), .Z(n295) );
  XNOR U553 ( .A(b[204]), .B(n296), .Z(c[204]) );
  XOR U554 ( .A(n297), .B(n298), .Z(n294) );
  ANDN U555 ( .B(n299), .A(n300), .Z(n297) );
  XNOR U556 ( .A(b[203]), .B(n298), .Z(n299) );
  XNOR U557 ( .A(b[203]), .B(n300), .Z(c[203]) );
  XOR U558 ( .A(n301), .B(n302), .Z(n298) );
  ANDN U559 ( .B(n303), .A(n304), .Z(n301) );
  XNOR U560 ( .A(b[202]), .B(n302), .Z(n303) );
  XNOR U561 ( .A(b[202]), .B(n304), .Z(c[202]) );
  XOR U562 ( .A(n305), .B(n306), .Z(n302) );
  ANDN U563 ( .B(n307), .A(n308), .Z(n305) );
  XNOR U564 ( .A(b[201]), .B(n306), .Z(n307) );
  XNOR U565 ( .A(b[201]), .B(n308), .Z(c[201]) );
  XOR U566 ( .A(n309), .B(n310), .Z(n306) );
  ANDN U567 ( .B(n311), .A(n312), .Z(n309) );
  XNOR U568 ( .A(b[200]), .B(n310), .Z(n311) );
  XNOR U569 ( .A(b[200]), .B(n312), .Z(c[200]) );
  XOR U570 ( .A(n313), .B(n314), .Z(n310) );
  ANDN U571 ( .B(n315), .A(n316), .Z(n313) );
  XNOR U572 ( .A(b[199]), .B(n314), .Z(n315) );
  XNOR U573 ( .A(b[1]), .B(n317), .Z(c[1]) );
  XNOR U574 ( .A(b[19]), .B(n318), .Z(c[19]) );
  XNOR U575 ( .A(b[199]), .B(n316), .Z(c[199]) );
  XOR U576 ( .A(n319), .B(n320), .Z(n314) );
  ANDN U577 ( .B(n321), .A(n322), .Z(n319) );
  XNOR U578 ( .A(b[198]), .B(n320), .Z(n321) );
  XNOR U579 ( .A(b[198]), .B(n322), .Z(c[198]) );
  XOR U580 ( .A(n323), .B(n324), .Z(n320) );
  ANDN U581 ( .B(n325), .A(n326), .Z(n323) );
  XNOR U582 ( .A(b[197]), .B(n324), .Z(n325) );
  XNOR U583 ( .A(b[197]), .B(n326), .Z(c[197]) );
  XOR U584 ( .A(n327), .B(n328), .Z(n324) );
  ANDN U585 ( .B(n329), .A(n330), .Z(n327) );
  XNOR U586 ( .A(b[196]), .B(n328), .Z(n329) );
  XNOR U587 ( .A(b[196]), .B(n330), .Z(c[196]) );
  XOR U588 ( .A(n331), .B(n332), .Z(n328) );
  ANDN U589 ( .B(n333), .A(n334), .Z(n331) );
  XNOR U590 ( .A(b[195]), .B(n332), .Z(n333) );
  XNOR U591 ( .A(b[195]), .B(n334), .Z(c[195]) );
  XOR U592 ( .A(n335), .B(n336), .Z(n332) );
  ANDN U593 ( .B(n337), .A(n338), .Z(n335) );
  XNOR U594 ( .A(b[194]), .B(n336), .Z(n337) );
  XNOR U595 ( .A(b[194]), .B(n338), .Z(c[194]) );
  XOR U596 ( .A(n339), .B(n340), .Z(n336) );
  ANDN U597 ( .B(n341), .A(n342), .Z(n339) );
  XNOR U598 ( .A(b[193]), .B(n340), .Z(n341) );
  XNOR U599 ( .A(b[193]), .B(n342), .Z(c[193]) );
  XOR U600 ( .A(n343), .B(n344), .Z(n340) );
  ANDN U601 ( .B(n345), .A(n346), .Z(n343) );
  XNOR U602 ( .A(b[192]), .B(n344), .Z(n345) );
  XNOR U603 ( .A(b[192]), .B(n346), .Z(c[192]) );
  XOR U604 ( .A(n347), .B(n348), .Z(n344) );
  ANDN U605 ( .B(n349), .A(n350), .Z(n347) );
  XNOR U606 ( .A(b[191]), .B(n348), .Z(n349) );
  XNOR U607 ( .A(b[191]), .B(n350), .Z(c[191]) );
  XOR U608 ( .A(n351), .B(n352), .Z(n348) );
  ANDN U609 ( .B(n353), .A(n354), .Z(n351) );
  XNOR U610 ( .A(b[190]), .B(n352), .Z(n353) );
  XNOR U611 ( .A(b[190]), .B(n354), .Z(c[190]) );
  XOR U612 ( .A(n355), .B(n356), .Z(n352) );
  ANDN U613 ( .B(n357), .A(n358), .Z(n355) );
  XNOR U614 ( .A(b[189]), .B(n356), .Z(n357) );
  XNOR U615 ( .A(b[18]), .B(n359), .Z(c[18]) );
  XNOR U616 ( .A(b[189]), .B(n358), .Z(c[189]) );
  XOR U617 ( .A(n360), .B(n361), .Z(n356) );
  ANDN U618 ( .B(n362), .A(n363), .Z(n360) );
  XNOR U619 ( .A(b[188]), .B(n361), .Z(n362) );
  XNOR U620 ( .A(b[188]), .B(n363), .Z(c[188]) );
  XOR U621 ( .A(n364), .B(n365), .Z(n361) );
  ANDN U622 ( .B(n366), .A(n367), .Z(n364) );
  XNOR U623 ( .A(b[187]), .B(n365), .Z(n366) );
  XNOR U624 ( .A(b[187]), .B(n367), .Z(c[187]) );
  XOR U625 ( .A(n368), .B(n369), .Z(n365) );
  ANDN U626 ( .B(n370), .A(n371), .Z(n368) );
  XNOR U627 ( .A(b[186]), .B(n369), .Z(n370) );
  XNOR U628 ( .A(b[186]), .B(n371), .Z(c[186]) );
  XOR U629 ( .A(n372), .B(n373), .Z(n369) );
  ANDN U630 ( .B(n374), .A(n375), .Z(n372) );
  XNOR U631 ( .A(b[185]), .B(n373), .Z(n374) );
  XNOR U632 ( .A(b[185]), .B(n375), .Z(c[185]) );
  XOR U633 ( .A(n376), .B(n377), .Z(n373) );
  ANDN U634 ( .B(n378), .A(n379), .Z(n376) );
  XNOR U635 ( .A(b[184]), .B(n377), .Z(n378) );
  XNOR U636 ( .A(b[184]), .B(n379), .Z(c[184]) );
  XOR U637 ( .A(n380), .B(n381), .Z(n377) );
  ANDN U638 ( .B(n382), .A(n383), .Z(n380) );
  XNOR U639 ( .A(b[183]), .B(n381), .Z(n382) );
  XNOR U640 ( .A(b[183]), .B(n383), .Z(c[183]) );
  XOR U641 ( .A(n384), .B(n385), .Z(n381) );
  ANDN U642 ( .B(n386), .A(n387), .Z(n384) );
  XNOR U643 ( .A(b[182]), .B(n385), .Z(n386) );
  XNOR U644 ( .A(b[182]), .B(n387), .Z(c[182]) );
  XOR U645 ( .A(n388), .B(n389), .Z(n385) );
  ANDN U646 ( .B(n390), .A(n391), .Z(n388) );
  XNOR U647 ( .A(b[181]), .B(n389), .Z(n390) );
  XNOR U648 ( .A(b[181]), .B(n391), .Z(c[181]) );
  XOR U649 ( .A(n392), .B(n393), .Z(n389) );
  ANDN U650 ( .B(n394), .A(n395), .Z(n392) );
  XNOR U651 ( .A(b[180]), .B(n393), .Z(n394) );
  XNOR U652 ( .A(b[180]), .B(n395), .Z(c[180]) );
  XOR U653 ( .A(n396), .B(n397), .Z(n393) );
  ANDN U654 ( .B(n398), .A(n399), .Z(n396) );
  XNOR U655 ( .A(b[179]), .B(n397), .Z(n398) );
  XNOR U656 ( .A(b[17]), .B(n400), .Z(c[17]) );
  XNOR U657 ( .A(b[179]), .B(n399), .Z(c[179]) );
  XOR U658 ( .A(n401), .B(n402), .Z(n397) );
  ANDN U659 ( .B(n403), .A(n404), .Z(n401) );
  XNOR U660 ( .A(b[178]), .B(n402), .Z(n403) );
  XNOR U661 ( .A(b[178]), .B(n404), .Z(c[178]) );
  XOR U662 ( .A(n405), .B(n406), .Z(n402) );
  ANDN U663 ( .B(n407), .A(n408), .Z(n405) );
  XNOR U664 ( .A(b[177]), .B(n406), .Z(n407) );
  XNOR U665 ( .A(b[177]), .B(n408), .Z(c[177]) );
  XOR U666 ( .A(n409), .B(n410), .Z(n406) );
  ANDN U667 ( .B(n411), .A(n412), .Z(n409) );
  XNOR U668 ( .A(b[176]), .B(n410), .Z(n411) );
  XNOR U669 ( .A(b[176]), .B(n412), .Z(c[176]) );
  XOR U670 ( .A(n413), .B(n414), .Z(n410) );
  ANDN U671 ( .B(n415), .A(n416), .Z(n413) );
  XNOR U672 ( .A(b[175]), .B(n414), .Z(n415) );
  XNOR U673 ( .A(b[175]), .B(n416), .Z(c[175]) );
  XOR U674 ( .A(n417), .B(n418), .Z(n414) );
  ANDN U675 ( .B(n419), .A(n420), .Z(n417) );
  XNOR U676 ( .A(b[174]), .B(n418), .Z(n419) );
  XNOR U677 ( .A(b[174]), .B(n420), .Z(c[174]) );
  XOR U678 ( .A(n421), .B(n422), .Z(n418) );
  ANDN U679 ( .B(n423), .A(n424), .Z(n421) );
  XNOR U680 ( .A(b[173]), .B(n422), .Z(n423) );
  XNOR U681 ( .A(b[173]), .B(n424), .Z(c[173]) );
  XOR U682 ( .A(n425), .B(n426), .Z(n422) );
  ANDN U683 ( .B(n427), .A(n428), .Z(n425) );
  XNOR U684 ( .A(b[172]), .B(n426), .Z(n427) );
  XNOR U685 ( .A(b[172]), .B(n428), .Z(c[172]) );
  XOR U686 ( .A(n429), .B(n430), .Z(n426) );
  ANDN U687 ( .B(n431), .A(n432), .Z(n429) );
  XNOR U688 ( .A(b[171]), .B(n430), .Z(n431) );
  XNOR U689 ( .A(b[171]), .B(n432), .Z(c[171]) );
  XOR U690 ( .A(n433), .B(n434), .Z(n430) );
  ANDN U691 ( .B(n435), .A(n436), .Z(n433) );
  XNOR U692 ( .A(b[170]), .B(n434), .Z(n435) );
  XNOR U693 ( .A(b[170]), .B(n436), .Z(c[170]) );
  XOR U694 ( .A(n437), .B(n438), .Z(n434) );
  ANDN U695 ( .B(n439), .A(n440), .Z(n437) );
  XNOR U696 ( .A(b[169]), .B(n438), .Z(n439) );
  XNOR U697 ( .A(b[16]), .B(n441), .Z(c[16]) );
  XNOR U698 ( .A(b[169]), .B(n440), .Z(c[169]) );
  XOR U699 ( .A(n442), .B(n443), .Z(n438) );
  ANDN U700 ( .B(n444), .A(n445), .Z(n442) );
  XNOR U701 ( .A(b[168]), .B(n443), .Z(n444) );
  XNOR U702 ( .A(b[168]), .B(n445), .Z(c[168]) );
  XOR U703 ( .A(n446), .B(n447), .Z(n443) );
  ANDN U704 ( .B(n448), .A(n449), .Z(n446) );
  XNOR U705 ( .A(b[167]), .B(n447), .Z(n448) );
  XNOR U706 ( .A(b[167]), .B(n449), .Z(c[167]) );
  XOR U707 ( .A(n450), .B(n451), .Z(n447) );
  ANDN U708 ( .B(n452), .A(n453), .Z(n450) );
  XNOR U709 ( .A(b[166]), .B(n451), .Z(n452) );
  XNOR U710 ( .A(b[166]), .B(n453), .Z(c[166]) );
  XOR U711 ( .A(n454), .B(n455), .Z(n451) );
  ANDN U712 ( .B(n456), .A(n457), .Z(n454) );
  XNOR U713 ( .A(b[165]), .B(n455), .Z(n456) );
  XNOR U714 ( .A(b[165]), .B(n457), .Z(c[165]) );
  XOR U715 ( .A(n458), .B(n459), .Z(n455) );
  ANDN U716 ( .B(n460), .A(n461), .Z(n458) );
  XNOR U717 ( .A(b[164]), .B(n459), .Z(n460) );
  XNOR U718 ( .A(b[164]), .B(n461), .Z(c[164]) );
  XOR U719 ( .A(n462), .B(n463), .Z(n459) );
  ANDN U720 ( .B(n464), .A(n465), .Z(n462) );
  XNOR U721 ( .A(b[163]), .B(n463), .Z(n464) );
  XNOR U722 ( .A(b[163]), .B(n465), .Z(c[163]) );
  XOR U723 ( .A(n466), .B(n467), .Z(n463) );
  ANDN U724 ( .B(n468), .A(n469), .Z(n466) );
  XNOR U725 ( .A(b[162]), .B(n467), .Z(n468) );
  XNOR U726 ( .A(b[162]), .B(n469), .Z(c[162]) );
  XOR U727 ( .A(n470), .B(n471), .Z(n467) );
  ANDN U728 ( .B(n472), .A(n473), .Z(n470) );
  XNOR U729 ( .A(b[161]), .B(n471), .Z(n472) );
  XNOR U730 ( .A(b[161]), .B(n473), .Z(c[161]) );
  XOR U731 ( .A(n474), .B(n475), .Z(n471) );
  ANDN U732 ( .B(n476), .A(n477), .Z(n474) );
  XNOR U733 ( .A(b[160]), .B(n475), .Z(n476) );
  XNOR U734 ( .A(b[160]), .B(n477), .Z(c[160]) );
  XOR U735 ( .A(n478), .B(n479), .Z(n475) );
  ANDN U736 ( .B(n480), .A(n481), .Z(n478) );
  XNOR U737 ( .A(b[159]), .B(n479), .Z(n480) );
  XNOR U738 ( .A(b[15]), .B(n482), .Z(c[15]) );
  XNOR U739 ( .A(b[159]), .B(n481), .Z(c[159]) );
  XOR U740 ( .A(n483), .B(n484), .Z(n479) );
  ANDN U741 ( .B(n485), .A(n486), .Z(n483) );
  XNOR U742 ( .A(b[158]), .B(n484), .Z(n485) );
  XNOR U743 ( .A(b[158]), .B(n486), .Z(c[158]) );
  XOR U744 ( .A(n487), .B(n488), .Z(n484) );
  ANDN U745 ( .B(n489), .A(n490), .Z(n487) );
  XNOR U746 ( .A(b[157]), .B(n488), .Z(n489) );
  XNOR U747 ( .A(b[157]), .B(n490), .Z(c[157]) );
  XOR U748 ( .A(n491), .B(n492), .Z(n488) );
  ANDN U749 ( .B(n493), .A(n494), .Z(n491) );
  XNOR U750 ( .A(b[156]), .B(n492), .Z(n493) );
  XNOR U751 ( .A(b[156]), .B(n494), .Z(c[156]) );
  XOR U752 ( .A(n495), .B(n496), .Z(n492) );
  ANDN U753 ( .B(n497), .A(n498), .Z(n495) );
  XNOR U754 ( .A(b[155]), .B(n496), .Z(n497) );
  XNOR U755 ( .A(b[155]), .B(n498), .Z(c[155]) );
  XOR U756 ( .A(n499), .B(n500), .Z(n496) );
  ANDN U757 ( .B(n501), .A(n502), .Z(n499) );
  XNOR U758 ( .A(b[154]), .B(n500), .Z(n501) );
  XNOR U759 ( .A(b[154]), .B(n502), .Z(c[154]) );
  XOR U760 ( .A(n503), .B(n504), .Z(n500) );
  ANDN U761 ( .B(n505), .A(n506), .Z(n503) );
  XNOR U762 ( .A(b[153]), .B(n504), .Z(n505) );
  XNOR U763 ( .A(b[153]), .B(n506), .Z(c[153]) );
  XOR U764 ( .A(n507), .B(n508), .Z(n504) );
  ANDN U765 ( .B(n509), .A(n510), .Z(n507) );
  XNOR U766 ( .A(b[152]), .B(n508), .Z(n509) );
  XNOR U767 ( .A(b[152]), .B(n510), .Z(c[152]) );
  XOR U768 ( .A(n511), .B(n512), .Z(n508) );
  ANDN U769 ( .B(n513), .A(n514), .Z(n511) );
  XNOR U770 ( .A(b[151]), .B(n512), .Z(n513) );
  XNOR U771 ( .A(b[151]), .B(n514), .Z(c[151]) );
  XOR U772 ( .A(n515), .B(n516), .Z(n512) );
  ANDN U773 ( .B(n517), .A(n518), .Z(n515) );
  XNOR U774 ( .A(b[150]), .B(n516), .Z(n517) );
  XNOR U775 ( .A(b[150]), .B(n518), .Z(c[150]) );
  XOR U776 ( .A(n519), .B(n520), .Z(n516) );
  ANDN U777 ( .B(n521), .A(n522), .Z(n519) );
  XNOR U778 ( .A(b[149]), .B(n520), .Z(n521) );
  XNOR U779 ( .A(b[14]), .B(n523), .Z(c[14]) );
  XNOR U780 ( .A(b[149]), .B(n522), .Z(c[149]) );
  XOR U781 ( .A(n524), .B(n525), .Z(n520) );
  ANDN U782 ( .B(n526), .A(n527), .Z(n524) );
  XNOR U783 ( .A(b[148]), .B(n525), .Z(n526) );
  XNOR U784 ( .A(b[148]), .B(n527), .Z(c[148]) );
  XOR U785 ( .A(n528), .B(n529), .Z(n525) );
  ANDN U786 ( .B(n530), .A(n531), .Z(n528) );
  XNOR U787 ( .A(b[147]), .B(n529), .Z(n530) );
  XNOR U788 ( .A(b[147]), .B(n531), .Z(c[147]) );
  XOR U789 ( .A(n532), .B(n533), .Z(n529) );
  ANDN U790 ( .B(n534), .A(n535), .Z(n532) );
  XNOR U791 ( .A(b[146]), .B(n533), .Z(n534) );
  XNOR U792 ( .A(b[146]), .B(n535), .Z(c[146]) );
  XOR U793 ( .A(n536), .B(n537), .Z(n533) );
  ANDN U794 ( .B(n538), .A(n539), .Z(n536) );
  XNOR U795 ( .A(b[145]), .B(n537), .Z(n538) );
  XNOR U796 ( .A(b[145]), .B(n539), .Z(c[145]) );
  XOR U797 ( .A(n540), .B(n541), .Z(n537) );
  ANDN U798 ( .B(n542), .A(n543), .Z(n540) );
  XNOR U799 ( .A(b[144]), .B(n541), .Z(n542) );
  XNOR U800 ( .A(b[144]), .B(n543), .Z(c[144]) );
  XOR U801 ( .A(n544), .B(n545), .Z(n541) );
  ANDN U802 ( .B(n546), .A(n547), .Z(n544) );
  XNOR U803 ( .A(b[143]), .B(n545), .Z(n546) );
  XNOR U804 ( .A(b[143]), .B(n547), .Z(c[143]) );
  XOR U805 ( .A(n548), .B(n549), .Z(n545) );
  ANDN U806 ( .B(n550), .A(n551), .Z(n548) );
  XNOR U807 ( .A(b[142]), .B(n549), .Z(n550) );
  XNOR U808 ( .A(b[142]), .B(n551), .Z(c[142]) );
  XOR U809 ( .A(n552), .B(n553), .Z(n549) );
  ANDN U810 ( .B(n554), .A(n555), .Z(n552) );
  XNOR U811 ( .A(b[141]), .B(n553), .Z(n554) );
  XNOR U812 ( .A(b[141]), .B(n555), .Z(c[141]) );
  XOR U813 ( .A(n556), .B(n557), .Z(n553) );
  ANDN U814 ( .B(n558), .A(n559), .Z(n556) );
  XNOR U815 ( .A(b[140]), .B(n557), .Z(n558) );
  XNOR U816 ( .A(b[140]), .B(n559), .Z(c[140]) );
  XOR U817 ( .A(n560), .B(n561), .Z(n557) );
  ANDN U818 ( .B(n562), .A(n563), .Z(n560) );
  XNOR U819 ( .A(b[139]), .B(n561), .Z(n562) );
  XNOR U820 ( .A(b[13]), .B(n564), .Z(c[13]) );
  XNOR U821 ( .A(b[139]), .B(n563), .Z(c[139]) );
  XOR U822 ( .A(n565), .B(n566), .Z(n561) );
  ANDN U823 ( .B(n567), .A(n568), .Z(n565) );
  XNOR U824 ( .A(b[138]), .B(n566), .Z(n567) );
  XNOR U825 ( .A(b[138]), .B(n568), .Z(c[138]) );
  XOR U826 ( .A(n569), .B(n570), .Z(n566) );
  ANDN U827 ( .B(n571), .A(n572), .Z(n569) );
  XNOR U828 ( .A(b[137]), .B(n570), .Z(n571) );
  XNOR U829 ( .A(b[137]), .B(n572), .Z(c[137]) );
  XOR U830 ( .A(n573), .B(n574), .Z(n570) );
  ANDN U831 ( .B(n575), .A(n576), .Z(n573) );
  XNOR U832 ( .A(b[136]), .B(n574), .Z(n575) );
  XNOR U833 ( .A(b[136]), .B(n576), .Z(c[136]) );
  XOR U834 ( .A(n577), .B(n578), .Z(n574) );
  ANDN U835 ( .B(n579), .A(n580), .Z(n577) );
  XNOR U836 ( .A(b[135]), .B(n578), .Z(n579) );
  XNOR U837 ( .A(b[135]), .B(n580), .Z(c[135]) );
  XOR U838 ( .A(n581), .B(n582), .Z(n578) );
  ANDN U839 ( .B(n583), .A(n584), .Z(n581) );
  XNOR U840 ( .A(b[134]), .B(n582), .Z(n583) );
  XNOR U841 ( .A(b[134]), .B(n584), .Z(c[134]) );
  XOR U842 ( .A(n585), .B(n586), .Z(n582) );
  ANDN U843 ( .B(n587), .A(n588), .Z(n585) );
  XNOR U844 ( .A(b[133]), .B(n586), .Z(n587) );
  XNOR U845 ( .A(b[133]), .B(n588), .Z(c[133]) );
  XOR U846 ( .A(n589), .B(n590), .Z(n586) );
  ANDN U847 ( .B(n591), .A(n592), .Z(n589) );
  XNOR U848 ( .A(b[132]), .B(n590), .Z(n591) );
  XNOR U849 ( .A(b[132]), .B(n592), .Z(c[132]) );
  XOR U850 ( .A(n593), .B(n594), .Z(n590) );
  ANDN U851 ( .B(n595), .A(n596), .Z(n593) );
  XNOR U852 ( .A(b[131]), .B(n594), .Z(n595) );
  XNOR U853 ( .A(b[131]), .B(n596), .Z(c[131]) );
  XOR U854 ( .A(n597), .B(n598), .Z(n594) );
  ANDN U855 ( .B(n599), .A(n600), .Z(n597) );
  XNOR U856 ( .A(b[130]), .B(n598), .Z(n599) );
  XNOR U857 ( .A(b[130]), .B(n600), .Z(c[130]) );
  XOR U858 ( .A(n601), .B(n602), .Z(n598) );
  ANDN U859 ( .B(n603), .A(n604), .Z(n601) );
  XNOR U860 ( .A(b[129]), .B(n602), .Z(n603) );
  XNOR U861 ( .A(b[12]), .B(n605), .Z(c[12]) );
  XNOR U862 ( .A(b[129]), .B(n604), .Z(c[129]) );
  XOR U863 ( .A(n606), .B(n607), .Z(n602) );
  ANDN U864 ( .B(n608), .A(n609), .Z(n606) );
  XNOR U865 ( .A(b[128]), .B(n607), .Z(n608) );
  XNOR U866 ( .A(b[128]), .B(n609), .Z(c[128]) );
  XOR U867 ( .A(n610), .B(n611), .Z(n607) );
  ANDN U868 ( .B(n612), .A(n613), .Z(n610) );
  XNOR U869 ( .A(b[127]), .B(n611), .Z(n612) );
  XNOR U870 ( .A(b[127]), .B(n613), .Z(c[127]) );
  XOR U871 ( .A(n614), .B(n615), .Z(n611) );
  ANDN U872 ( .B(n616), .A(n617), .Z(n614) );
  XNOR U873 ( .A(b[126]), .B(n615), .Z(n616) );
  XNOR U874 ( .A(b[126]), .B(n617), .Z(c[126]) );
  XOR U875 ( .A(n618), .B(n619), .Z(n615) );
  ANDN U876 ( .B(n620), .A(n621), .Z(n618) );
  XNOR U877 ( .A(b[125]), .B(n619), .Z(n620) );
  XNOR U878 ( .A(b[125]), .B(n621), .Z(c[125]) );
  XOR U879 ( .A(n622), .B(n623), .Z(n619) );
  ANDN U880 ( .B(n624), .A(n625), .Z(n622) );
  XNOR U881 ( .A(b[124]), .B(n623), .Z(n624) );
  XNOR U882 ( .A(b[124]), .B(n625), .Z(c[124]) );
  XOR U883 ( .A(n626), .B(n627), .Z(n623) );
  ANDN U884 ( .B(n628), .A(n629), .Z(n626) );
  XNOR U885 ( .A(b[123]), .B(n627), .Z(n628) );
  XNOR U886 ( .A(b[123]), .B(n629), .Z(c[123]) );
  XOR U887 ( .A(n630), .B(n631), .Z(n627) );
  ANDN U888 ( .B(n632), .A(n633), .Z(n630) );
  XNOR U889 ( .A(b[122]), .B(n631), .Z(n632) );
  XNOR U890 ( .A(b[122]), .B(n633), .Z(c[122]) );
  XOR U891 ( .A(n634), .B(n635), .Z(n631) );
  ANDN U892 ( .B(n636), .A(n637), .Z(n634) );
  XNOR U893 ( .A(b[121]), .B(n635), .Z(n636) );
  XNOR U894 ( .A(b[121]), .B(n637), .Z(c[121]) );
  XOR U895 ( .A(n638), .B(n639), .Z(n635) );
  ANDN U896 ( .B(n640), .A(n641), .Z(n638) );
  XNOR U897 ( .A(b[120]), .B(n639), .Z(n640) );
  XNOR U898 ( .A(b[120]), .B(n641), .Z(c[120]) );
  XOR U899 ( .A(n642), .B(n643), .Z(n639) );
  ANDN U900 ( .B(n644), .A(n645), .Z(n642) );
  XNOR U901 ( .A(b[119]), .B(n643), .Z(n644) );
  XNOR U902 ( .A(b[11]), .B(n646), .Z(c[11]) );
  XNOR U903 ( .A(b[119]), .B(n645), .Z(c[119]) );
  XOR U904 ( .A(n647), .B(n648), .Z(n643) );
  ANDN U905 ( .B(n649), .A(n650), .Z(n647) );
  XNOR U906 ( .A(b[118]), .B(n648), .Z(n649) );
  XNOR U907 ( .A(b[118]), .B(n650), .Z(c[118]) );
  XOR U908 ( .A(n651), .B(n652), .Z(n648) );
  ANDN U909 ( .B(n653), .A(n654), .Z(n651) );
  XNOR U910 ( .A(b[117]), .B(n652), .Z(n653) );
  XNOR U911 ( .A(b[117]), .B(n654), .Z(c[117]) );
  XOR U912 ( .A(n655), .B(n656), .Z(n652) );
  ANDN U913 ( .B(n657), .A(n658), .Z(n655) );
  XNOR U914 ( .A(b[116]), .B(n656), .Z(n657) );
  XNOR U915 ( .A(b[116]), .B(n658), .Z(c[116]) );
  XOR U916 ( .A(n659), .B(n660), .Z(n656) );
  ANDN U917 ( .B(n661), .A(n662), .Z(n659) );
  XNOR U918 ( .A(b[115]), .B(n660), .Z(n661) );
  XNOR U919 ( .A(b[115]), .B(n662), .Z(c[115]) );
  XOR U920 ( .A(n663), .B(n664), .Z(n660) );
  ANDN U921 ( .B(n665), .A(n666), .Z(n663) );
  XNOR U922 ( .A(b[114]), .B(n664), .Z(n665) );
  XNOR U923 ( .A(b[114]), .B(n666), .Z(c[114]) );
  XOR U924 ( .A(n667), .B(n668), .Z(n664) );
  ANDN U925 ( .B(n669), .A(n670), .Z(n667) );
  XNOR U926 ( .A(b[113]), .B(n668), .Z(n669) );
  XNOR U927 ( .A(b[113]), .B(n670), .Z(c[113]) );
  XOR U928 ( .A(n671), .B(n672), .Z(n668) );
  ANDN U929 ( .B(n673), .A(n674), .Z(n671) );
  XNOR U930 ( .A(b[112]), .B(n672), .Z(n673) );
  XNOR U931 ( .A(b[112]), .B(n674), .Z(c[112]) );
  XOR U932 ( .A(n675), .B(n676), .Z(n672) );
  ANDN U933 ( .B(n677), .A(n678), .Z(n675) );
  XNOR U934 ( .A(b[111]), .B(n676), .Z(n677) );
  XNOR U935 ( .A(b[111]), .B(n678), .Z(c[111]) );
  XOR U936 ( .A(n679), .B(n680), .Z(n676) );
  ANDN U937 ( .B(n681), .A(n682), .Z(n679) );
  XNOR U938 ( .A(b[110]), .B(n680), .Z(n681) );
  XNOR U939 ( .A(b[110]), .B(n682), .Z(c[110]) );
  XOR U940 ( .A(n683), .B(n684), .Z(n680) );
  ANDN U941 ( .B(n685), .A(n686), .Z(n683) );
  XNOR U942 ( .A(b[109]), .B(n684), .Z(n685) );
  XNOR U943 ( .A(b[10]), .B(n687), .Z(c[10]) );
  XNOR U944 ( .A(b[109]), .B(n686), .Z(c[109]) );
  XOR U945 ( .A(n688), .B(n689), .Z(n684) );
  ANDN U946 ( .B(n690), .A(n691), .Z(n688) );
  XNOR U947 ( .A(b[108]), .B(n689), .Z(n690) );
  XNOR U948 ( .A(b[108]), .B(n691), .Z(c[108]) );
  XOR U949 ( .A(n692), .B(n693), .Z(n689) );
  ANDN U950 ( .B(n694), .A(n695), .Z(n692) );
  XNOR U951 ( .A(b[107]), .B(n693), .Z(n694) );
  XNOR U952 ( .A(b[107]), .B(n695), .Z(c[107]) );
  XOR U953 ( .A(n696), .B(n697), .Z(n693) );
  ANDN U954 ( .B(n698), .A(n699), .Z(n696) );
  XNOR U955 ( .A(b[106]), .B(n697), .Z(n698) );
  XNOR U956 ( .A(b[106]), .B(n699), .Z(c[106]) );
  XOR U957 ( .A(n700), .B(n701), .Z(n697) );
  ANDN U958 ( .B(n702), .A(n703), .Z(n700) );
  XNOR U959 ( .A(b[105]), .B(n701), .Z(n702) );
  XNOR U960 ( .A(b[105]), .B(n703), .Z(c[105]) );
  XOR U961 ( .A(n704), .B(n705), .Z(n701) );
  ANDN U962 ( .B(n706), .A(n707), .Z(n704) );
  XNOR U963 ( .A(b[104]), .B(n705), .Z(n706) );
  XNOR U964 ( .A(b[104]), .B(n707), .Z(c[104]) );
  XOR U965 ( .A(n708), .B(n709), .Z(n705) );
  ANDN U966 ( .B(n710), .A(n711), .Z(n708) );
  XNOR U967 ( .A(b[103]), .B(n709), .Z(n710) );
  XNOR U968 ( .A(b[103]), .B(n711), .Z(c[103]) );
  XOR U969 ( .A(n712), .B(n713), .Z(n709) );
  ANDN U970 ( .B(n714), .A(n715), .Z(n712) );
  XNOR U971 ( .A(b[102]), .B(n713), .Z(n714) );
  XNOR U972 ( .A(b[102]), .B(n715), .Z(c[102]) );
  XOR U973 ( .A(n716), .B(n717), .Z(n713) );
  ANDN U974 ( .B(n718), .A(n719), .Z(n716) );
  XNOR U975 ( .A(b[101]), .B(n717), .Z(n718) );
  XNOR U976 ( .A(b[101]), .B(n719), .Z(c[101]) );
  XOR U977 ( .A(n720), .B(n721), .Z(n717) );
  ANDN U978 ( .B(n722), .A(n723), .Z(n720) );
  XNOR U979 ( .A(b[100]), .B(n721), .Z(n722) );
  XNOR U980 ( .A(b[100]), .B(n723), .Z(c[100]) );
  XOR U981 ( .A(n724), .B(n725), .Z(n721) );
  ANDN U982 ( .B(n726), .A(n6), .Z(n724) );
  XNOR U983 ( .A(b[99]), .B(n725), .Z(n726) );
  XOR U984 ( .A(n727), .B(n728), .Z(n725) );
  ANDN U985 ( .B(n729), .A(n7), .Z(n727) );
  XNOR U986 ( .A(b[98]), .B(n728), .Z(n729) );
  XOR U987 ( .A(n730), .B(n731), .Z(n728) );
  ANDN U988 ( .B(n732), .A(n8), .Z(n730) );
  XNOR U989 ( .A(b[97]), .B(n731), .Z(n732) );
  XOR U990 ( .A(n733), .B(n734), .Z(n731) );
  ANDN U991 ( .B(n735), .A(n9), .Z(n733) );
  XNOR U992 ( .A(b[96]), .B(n734), .Z(n735) );
  XOR U993 ( .A(n736), .B(n737), .Z(n734) );
  ANDN U994 ( .B(n738), .A(n10), .Z(n736) );
  XNOR U995 ( .A(b[95]), .B(n737), .Z(n738) );
  XOR U996 ( .A(n739), .B(n740), .Z(n737) );
  ANDN U997 ( .B(n741), .A(n11), .Z(n739) );
  XNOR U998 ( .A(b[94]), .B(n740), .Z(n741) );
  XOR U999 ( .A(n742), .B(n743), .Z(n740) );
  ANDN U1000 ( .B(n744), .A(n12), .Z(n742) );
  XNOR U1001 ( .A(b[93]), .B(n743), .Z(n744) );
  XOR U1002 ( .A(n745), .B(n746), .Z(n743) );
  ANDN U1003 ( .B(n747), .A(n13), .Z(n745) );
  XNOR U1004 ( .A(b[92]), .B(n746), .Z(n747) );
  XOR U1005 ( .A(n748), .B(n749), .Z(n746) );
  ANDN U1006 ( .B(n750), .A(n14), .Z(n748) );
  XNOR U1007 ( .A(b[91]), .B(n749), .Z(n750) );
  XOR U1008 ( .A(n751), .B(n752), .Z(n749) );
  ANDN U1009 ( .B(n753), .A(n15), .Z(n751) );
  XNOR U1010 ( .A(b[90]), .B(n752), .Z(n753) );
  XOR U1011 ( .A(n754), .B(n755), .Z(n752) );
  ANDN U1012 ( .B(n756), .A(n17), .Z(n754) );
  XNOR U1013 ( .A(b[89]), .B(n755), .Z(n756) );
  XOR U1014 ( .A(n757), .B(n758), .Z(n755) );
  ANDN U1015 ( .B(n759), .A(n18), .Z(n757) );
  XNOR U1016 ( .A(b[88]), .B(n758), .Z(n759) );
  XOR U1017 ( .A(n760), .B(n761), .Z(n758) );
  ANDN U1018 ( .B(n762), .A(n19), .Z(n760) );
  XNOR U1019 ( .A(b[87]), .B(n761), .Z(n762) );
  XOR U1020 ( .A(n763), .B(n764), .Z(n761) );
  ANDN U1021 ( .B(n765), .A(n20), .Z(n763) );
  XNOR U1022 ( .A(b[86]), .B(n764), .Z(n765) );
  XOR U1023 ( .A(n766), .B(n767), .Z(n764) );
  ANDN U1024 ( .B(n768), .A(n21), .Z(n766) );
  XNOR U1025 ( .A(b[85]), .B(n767), .Z(n768) );
  XOR U1026 ( .A(n769), .B(n770), .Z(n767) );
  ANDN U1027 ( .B(n771), .A(n22), .Z(n769) );
  XNOR U1028 ( .A(b[84]), .B(n770), .Z(n771) );
  XOR U1029 ( .A(n772), .B(n773), .Z(n770) );
  ANDN U1030 ( .B(n774), .A(n23), .Z(n772) );
  XNOR U1031 ( .A(b[83]), .B(n773), .Z(n774) );
  XOR U1032 ( .A(n775), .B(n776), .Z(n773) );
  ANDN U1033 ( .B(n777), .A(n24), .Z(n775) );
  XNOR U1034 ( .A(b[82]), .B(n776), .Z(n777) );
  XOR U1035 ( .A(n778), .B(n779), .Z(n776) );
  ANDN U1036 ( .B(n780), .A(n25), .Z(n778) );
  XNOR U1037 ( .A(b[81]), .B(n779), .Z(n780) );
  XOR U1038 ( .A(n781), .B(n782), .Z(n779) );
  ANDN U1039 ( .B(n783), .A(n26), .Z(n781) );
  XNOR U1040 ( .A(b[80]), .B(n782), .Z(n783) );
  XOR U1041 ( .A(n784), .B(n785), .Z(n782) );
  ANDN U1042 ( .B(n786), .A(n28), .Z(n784) );
  XNOR U1043 ( .A(b[79]), .B(n785), .Z(n786) );
  XOR U1044 ( .A(n787), .B(n788), .Z(n785) );
  ANDN U1045 ( .B(n789), .A(n29), .Z(n787) );
  XNOR U1046 ( .A(b[78]), .B(n788), .Z(n789) );
  XOR U1047 ( .A(n790), .B(n791), .Z(n788) );
  ANDN U1048 ( .B(n792), .A(n30), .Z(n790) );
  XNOR U1049 ( .A(b[77]), .B(n791), .Z(n792) );
  XOR U1050 ( .A(n793), .B(n794), .Z(n791) );
  ANDN U1051 ( .B(n795), .A(n31), .Z(n793) );
  XNOR U1052 ( .A(b[76]), .B(n794), .Z(n795) );
  XOR U1053 ( .A(n796), .B(n797), .Z(n794) );
  ANDN U1054 ( .B(n798), .A(n32), .Z(n796) );
  XNOR U1055 ( .A(b[75]), .B(n797), .Z(n798) );
  XOR U1056 ( .A(n799), .B(n800), .Z(n797) );
  ANDN U1057 ( .B(n801), .A(n33), .Z(n799) );
  XNOR U1058 ( .A(b[74]), .B(n800), .Z(n801) );
  XOR U1059 ( .A(n802), .B(n803), .Z(n800) );
  ANDN U1060 ( .B(n804), .A(n34), .Z(n802) );
  XNOR U1061 ( .A(b[73]), .B(n803), .Z(n804) );
  XOR U1062 ( .A(n805), .B(n806), .Z(n803) );
  ANDN U1063 ( .B(n807), .A(n35), .Z(n805) );
  XNOR U1064 ( .A(b[72]), .B(n806), .Z(n807) );
  XOR U1065 ( .A(n808), .B(n809), .Z(n806) );
  ANDN U1066 ( .B(n810), .A(n36), .Z(n808) );
  XNOR U1067 ( .A(b[71]), .B(n809), .Z(n810) );
  XOR U1068 ( .A(n811), .B(n812), .Z(n809) );
  ANDN U1069 ( .B(n813), .A(n37), .Z(n811) );
  XNOR U1070 ( .A(b[70]), .B(n812), .Z(n813) );
  XOR U1071 ( .A(n814), .B(n815), .Z(n812) );
  ANDN U1072 ( .B(n816), .A(n39), .Z(n814) );
  XNOR U1073 ( .A(b[69]), .B(n815), .Z(n816) );
  XOR U1074 ( .A(n817), .B(n818), .Z(n815) );
  ANDN U1075 ( .B(n819), .A(n40), .Z(n817) );
  XNOR U1076 ( .A(b[68]), .B(n818), .Z(n819) );
  XOR U1077 ( .A(n820), .B(n821), .Z(n818) );
  ANDN U1078 ( .B(n822), .A(n41), .Z(n820) );
  XNOR U1079 ( .A(b[67]), .B(n821), .Z(n822) );
  XOR U1080 ( .A(n823), .B(n824), .Z(n821) );
  ANDN U1081 ( .B(n825), .A(n42), .Z(n823) );
  XNOR U1082 ( .A(b[66]), .B(n824), .Z(n825) );
  XOR U1083 ( .A(n826), .B(n827), .Z(n824) );
  ANDN U1084 ( .B(n828), .A(n43), .Z(n826) );
  XNOR U1085 ( .A(b[65]), .B(n827), .Z(n828) );
  XOR U1086 ( .A(n829), .B(n830), .Z(n827) );
  ANDN U1087 ( .B(n831), .A(n44), .Z(n829) );
  XNOR U1088 ( .A(b[64]), .B(n830), .Z(n831) );
  XOR U1089 ( .A(n832), .B(n833), .Z(n830) );
  ANDN U1090 ( .B(n834), .A(n45), .Z(n832) );
  XNOR U1091 ( .A(b[63]), .B(n833), .Z(n834) );
  XOR U1092 ( .A(n835), .B(n836), .Z(n833) );
  ANDN U1093 ( .B(n837), .A(n46), .Z(n835) );
  XNOR U1094 ( .A(b[62]), .B(n836), .Z(n837) );
  XOR U1095 ( .A(n838), .B(n839), .Z(n836) );
  ANDN U1096 ( .B(n840), .A(n47), .Z(n838) );
  XNOR U1097 ( .A(b[61]), .B(n839), .Z(n840) );
  XOR U1098 ( .A(n841), .B(n842), .Z(n839) );
  ANDN U1099 ( .B(n843), .A(n48), .Z(n841) );
  XNOR U1100 ( .A(b[60]), .B(n842), .Z(n843) );
  XOR U1101 ( .A(n844), .B(n845), .Z(n842) );
  ANDN U1102 ( .B(n846), .A(n50), .Z(n844) );
  XNOR U1103 ( .A(b[59]), .B(n845), .Z(n846) );
  XOR U1104 ( .A(n847), .B(n848), .Z(n845) );
  ANDN U1105 ( .B(n849), .A(n51), .Z(n847) );
  XNOR U1106 ( .A(b[58]), .B(n848), .Z(n849) );
  XOR U1107 ( .A(n850), .B(n851), .Z(n848) );
  ANDN U1108 ( .B(n852), .A(n52), .Z(n850) );
  XNOR U1109 ( .A(b[57]), .B(n851), .Z(n852) );
  XOR U1110 ( .A(n853), .B(n854), .Z(n851) );
  ANDN U1111 ( .B(n855), .A(n53), .Z(n853) );
  XNOR U1112 ( .A(b[56]), .B(n854), .Z(n855) );
  XOR U1113 ( .A(n856), .B(n857), .Z(n854) );
  ANDN U1114 ( .B(n858), .A(n54), .Z(n856) );
  XNOR U1115 ( .A(b[55]), .B(n857), .Z(n858) );
  XOR U1116 ( .A(n859), .B(n860), .Z(n857) );
  ANDN U1117 ( .B(n861), .A(n55), .Z(n859) );
  XNOR U1118 ( .A(b[54]), .B(n860), .Z(n861) );
  XOR U1119 ( .A(n862), .B(n863), .Z(n860) );
  ANDN U1120 ( .B(n864), .A(n56), .Z(n862) );
  XNOR U1121 ( .A(b[53]), .B(n863), .Z(n864) );
  XOR U1122 ( .A(n865), .B(n866), .Z(n863) );
  ANDN U1123 ( .B(n867), .A(n57), .Z(n865) );
  XNOR U1124 ( .A(b[52]), .B(n866), .Z(n867) );
  XOR U1125 ( .A(n868), .B(n869), .Z(n866) );
  ANDN U1126 ( .B(n870), .A(n58), .Z(n868) );
  XNOR U1127 ( .A(b[51]), .B(n869), .Z(n870) );
  XOR U1128 ( .A(n871), .B(n872), .Z(n869) );
  ANDN U1129 ( .B(n873), .A(n59), .Z(n871) );
  XNOR U1130 ( .A(b[50]), .B(n872), .Z(n873) );
  XOR U1131 ( .A(n874), .B(n875), .Z(n872) );
  ANDN U1132 ( .B(n876), .A(n61), .Z(n874) );
  XNOR U1133 ( .A(b[49]), .B(n875), .Z(n876) );
  XOR U1134 ( .A(n877), .B(n878), .Z(n875) );
  ANDN U1135 ( .B(n879), .A(n62), .Z(n877) );
  XNOR U1136 ( .A(b[48]), .B(n878), .Z(n879) );
  XOR U1137 ( .A(n880), .B(n881), .Z(n878) );
  ANDN U1138 ( .B(n882), .A(n63), .Z(n880) );
  XNOR U1139 ( .A(b[47]), .B(n881), .Z(n882) );
  XOR U1140 ( .A(n883), .B(n884), .Z(n881) );
  ANDN U1141 ( .B(n885), .A(n64), .Z(n883) );
  XNOR U1142 ( .A(b[46]), .B(n884), .Z(n885) );
  XOR U1143 ( .A(n886), .B(n887), .Z(n884) );
  ANDN U1144 ( .B(n888), .A(n65), .Z(n886) );
  XNOR U1145 ( .A(b[45]), .B(n887), .Z(n888) );
  XOR U1146 ( .A(n889), .B(n890), .Z(n887) );
  ANDN U1147 ( .B(n891), .A(n66), .Z(n889) );
  XNOR U1148 ( .A(b[44]), .B(n890), .Z(n891) );
  XOR U1149 ( .A(n892), .B(n893), .Z(n890) );
  ANDN U1150 ( .B(n894), .A(n67), .Z(n892) );
  XNOR U1151 ( .A(b[43]), .B(n893), .Z(n894) );
  XOR U1152 ( .A(n895), .B(n896), .Z(n893) );
  ANDN U1153 ( .B(n897), .A(n68), .Z(n895) );
  XNOR U1154 ( .A(b[42]), .B(n896), .Z(n897) );
  XOR U1155 ( .A(n898), .B(n899), .Z(n896) );
  ANDN U1156 ( .B(n900), .A(n69), .Z(n898) );
  XNOR U1157 ( .A(b[41]), .B(n899), .Z(n900) );
  XOR U1158 ( .A(n901), .B(n902), .Z(n899) );
  ANDN U1159 ( .B(n903), .A(n70), .Z(n901) );
  XNOR U1160 ( .A(b[40]), .B(n902), .Z(n903) );
  XOR U1161 ( .A(n904), .B(n905), .Z(n902) );
  ANDN U1162 ( .B(n906), .A(n72), .Z(n904) );
  XNOR U1163 ( .A(b[39]), .B(n905), .Z(n906) );
  XOR U1164 ( .A(n907), .B(n908), .Z(n905) );
  ANDN U1165 ( .B(n909), .A(n73), .Z(n907) );
  XNOR U1166 ( .A(b[38]), .B(n908), .Z(n909) );
  XOR U1167 ( .A(n910), .B(n911), .Z(n908) );
  ANDN U1168 ( .B(n912), .A(n74), .Z(n910) );
  XNOR U1169 ( .A(b[37]), .B(n911), .Z(n912) );
  XOR U1170 ( .A(n913), .B(n914), .Z(n911) );
  ANDN U1171 ( .B(n915), .A(n75), .Z(n913) );
  XNOR U1172 ( .A(b[36]), .B(n914), .Z(n915) );
  XOR U1173 ( .A(n916), .B(n917), .Z(n914) );
  ANDN U1174 ( .B(n918), .A(n76), .Z(n916) );
  XNOR U1175 ( .A(b[35]), .B(n917), .Z(n918) );
  XOR U1176 ( .A(n919), .B(n920), .Z(n917) );
  ANDN U1177 ( .B(n921), .A(n77), .Z(n919) );
  XNOR U1178 ( .A(b[34]), .B(n920), .Z(n921) );
  XOR U1179 ( .A(n922), .B(n923), .Z(n920) );
  ANDN U1180 ( .B(n924), .A(n78), .Z(n922) );
  XNOR U1181 ( .A(b[33]), .B(n923), .Z(n924) );
  XOR U1182 ( .A(n925), .B(n926), .Z(n923) );
  ANDN U1183 ( .B(n927), .A(n79), .Z(n925) );
  XNOR U1184 ( .A(b[32]), .B(n926), .Z(n927) );
  XOR U1185 ( .A(n928), .B(n929), .Z(n926) );
  ANDN U1186 ( .B(n930), .A(n80), .Z(n928) );
  XNOR U1187 ( .A(b[31]), .B(n929), .Z(n930) );
  XOR U1188 ( .A(n931), .B(n932), .Z(n929) );
  ANDN U1189 ( .B(n933), .A(n81), .Z(n931) );
  XNOR U1190 ( .A(b[30]), .B(n932), .Z(n933) );
  XOR U1191 ( .A(n934), .B(n935), .Z(n932) );
  ANDN U1192 ( .B(n936), .A(n83), .Z(n934) );
  XNOR U1193 ( .A(b[29]), .B(n935), .Z(n936) );
  XOR U1194 ( .A(n937), .B(n938), .Z(n935) );
  ANDN U1195 ( .B(n939), .A(n84), .Z(n937) );
  XNOR U1196 ( .A(b[28]), .B(n938), .Z(n939) );
  XOR U1197 ( .A(n940), .B(n941), .Z(n938) );
  ANDN U1198 ( .B(n942), .A(n85), .Z(n940) );
  XNOR U1199 ( .A(b[27]), .B(n941), .Z(n942) );
  XOR U1200 ( .A(n943), .B(n944), .Z(n941) );
  ANDN U1201 ( .B(n945), .A(n86), .Z(n943) );
  XNOR U1202 ( .A(b[26]), .B(n944), .Z(n945) );
  XOR U1203 ( .A(n946), .B(n947), .Z(n944) );
  ANDN U1204 ( .B(n948), .A(n87), .Z(n946) );
  XNOR U1205 ( .A(b[25]), .B(n947), .Z(n948) );
  XOR U1206 ( .A(n949), .B(n950), .Z(n947) );
  ANDN U1207 ( .B(n951), .A(n112), .Z(n949) );
  XNOR U1208 ( .A(b[24]), .B(n950), .Z(n951) );
  XOR U1209 ( .A(n952), .B(n953), .Z(n950) );
  ANDN U1210 ( .B(n954), .A(n153), .Z(n952) );
  XNOR U1211 ( .A(b[23]), .B(n953), .Z(n954) );
  XOR U1212 ( .A(n955), .B(n956), .Z(n953) );
  ANDN U1213 ( .B(n957), .A(n194), .Z(n955) );
  XNOR U1214 ( .A(b[22]), .B(n956), .Z(n957) );
  XOR U1215 ( .A(n958), .B(n959), .Z(n956) );
  ANDN U1216 ( .B(n960), .A(n235), .Z(n958) );
  XNOR U1217 ( .A(b[21]), .B(n959), .Z(n960) );
  XOR U1218 ( .A(n961), .B(n962), .Z(n959) );
  ANDN U1219 ( .B(n963), .A(n276), .Z(n961) );
  XNOR U1220 ( .A(b[20]), .B(n962), .Z(n963) );
  XOR U1221 ( .A(n964), .B(n965), .Z(n962) );
  ANDN U1222 ( .B(n966), .A(n318), .Z(n964) );
  XNOR U1223 ( .A(b[19]), .B(n965), .Z(n966) );
  XOR U1224 ( .A(n967), .B(n968), .Z(n965) );
  ANDN U1225 ( .B(n969), .A(n359), .Z(n967) );
  XNOR U1226 ( .A(b[18]), .B(n968), .Z(n969) );
  XOR U1227 ( .A(n970), .B(n971), .Z(n968) );
  ANDN U1228 ( .B(n972), .A(n400), .Z(n970) );
  XNOR U1229 ( .A(b[17]), .B(n971), .Z(n972) );
  XOR U1230 ( .A(n973), .B(n974), .Z(n971) );
  ANDN U1231 ( .B(n975), .A(n441), .Z(n973) );
  XNOR U1232 ( .A(b[16]), .B(n974), .Z(n975) );
  XOR U1233 ( .A(n976), .B(n977), .Z(n974) );
  ANDN U1234 ( .B(n978), .A(n482), .Z(n976) );
  XNOR U1235 ( .A(b[15]), .B(n977), .Z(n978) );
  XOR U1236 ( .A(n979), .B(n980), .Z(n977) );
  ANDN U1237 ( .B(n981), .A(n523), .Z(n979) );
  XNOR U1238 ( .A(b[14]), .B(n980), .Z(n981) );
  XOR U1239 ( .A(n982), .B(n983), .Z(n980) );
  ANDN U1240 ( .B(n984), .A(n564), .Z(n982) );
  XNOR U1241 ( .A(b[13]), .B(n983), .Z(n984) );
  XOR U1242 ( .A(n985), .B(n986), .Z(n983) );
  ANDN U1243 ( .B(n987), .A(n605), .Z(n985) );
  XNOR U1244 ( .A(b[12]), .B(n986), .Z(n987) );
  XOR U1245 ( .A(n988), .B(n989), .Z(n986) );
  ANDN U1246 ( .B(n990), .A(n646), .Z(n988) );
  XNOR U1247 ( .A(b[11]), .B(n989), .Z(n990) );
  XOR U1248 ( .A(n991), .B(n992), .Z(n989) );
  ANDN U1249 ( .B(n993), .A(n687), .Z(n991) );
  XNOR U1250 ( .A(b[10]), .B(n992), .Z(n993) );
  XOR U1251 ( .A(n994), .B(n995), .Z(n992) );
  ANDN U1252 ( .B(n996), .A(n5), .Z(n994) );
  XNOR U1253 ( .A(b[9]), .B(n995), .Z(n996) );
  XOR U1254 ( .A(n997), .B(n998), .Z(n995) );
  ANDN U1255 ( .B(n999), .A(n16), .Z(n997) );
  XNOR U1256 ( .A(b[8]), .B(n998), .Z(n999) );
  XOR U1257 ( .A(n1000), .B(n1001), .Z(n998) );
  ANDN U1258 ( .B(n1002), .A(n27), .Z(n1000) );
  XNOR U1259 ( .A(b[7]), .B(n1001), .Z(n1002) );
  XOR U1260 ( .A(n1003), .B(n1004), .Z(n1001) );
  ANDN U1261 ( .B(n1005), .A(n38), .Z(n1003) );
  XNOR U1262 ( .A(b[6]), .B(n1004), .Z(n1005) );
  XOR U1263 ( .A(n1006), .B(n1007), .Z(n1004) );
  ANDN U1264 ( .B(n1008), .A(n49), .Z(n1006) );
  XNOR U1265 ( .A(b[5]), .B(n1007), .Z(n1008) );
  XOR U1266 ( .A(n1009), .B(n1010), .Z(n1007) );
  ANDN U1267 ( .B(n1011), .A(n60), .Z(n1009) );
  XNOR U1268 ( .A(b[4]), .B(n1010), .Z(n1011) );
  XOR U1269 ( .A(n1012), .B(n1013), .Z(n1010) );
  ANDN U1270 ( .B(n1014), .A(n71), .Z(n1012) );
  XNOR U1271 ( .A(b[3]), .B(n1013), .Z(n1014) );
  XOR U1272 ( .A(n1015), .B(n1016), .Z(n1013) );
  ANDN U1273 ( .B(n1017), .A(n82), .Z(n1015) );
  XNOR U1274 ( .A(b[2]), .B(n1016), .Z(n1017) );
  XOR U1275 ( .A(n1018), .B(n1019), .Z(n1016) );
  ANDN U1276 ( .B(n1020), .A(n317), .Z(n1018) );
  XNOR U1277 ( .A(b[1]), .B(n1019), .Z(n1020) );
  XOR U1278 ( .A(carry_on), .B(n1021), .Z(n1019) );
  NANDN U1279 ( .A(n1022), .B(n1023), .Z(n1021) );
  XOR U1280 ( .A(carry_on), .B(b[0]), .Z(n1023) );
  XNOR U1281 ( .A(b[0]), .B(n1022), .Z(c[0]) );
  XNOR U1282 ( .A(a[0]), .B(carry_on), .Z(n1022) );
endmodule

