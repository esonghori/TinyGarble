
module mult_N256_CC32 ( clk, rst, a, b, c );
  input [255:0] a;
  input [7:0] b;
  output [511:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570;
  wire   [511:0] sreg;

  DFF \sreg_reg[503]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(sreg[503]) );
  DFF \sreg_reg[502]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(sreg[502]) );
  DFF \sreg_reg[501]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(sreg[501]) );
  DFF \sreg_reg[500]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(sreg[500]) );
  DFF \sreg_reg[499]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(sreg[499]) );
  DFF \sreg_reg[498]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(sreg[498]) );
  DFF \sreg_reg[497]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(sreg[497]) );
  DFF \sreg_reg[496]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(sreg[496]) );
  DFF \sreg_reg[495]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(sreg[495]) );
  DFF \sreg_reg[494]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(sreg[494]) );
  DFF \sreg_reg[493]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(sreg[493]) );
  DFF \sreg_reg[492]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(sreg[492]) );
  DFF \sreg_reg[491]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(sreg[491]) );
  DFF \sreg_reg[490]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(sreg[490]) );
  DFF \sreg_reg[489]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(sreg[489]) );
  DFF \sreg_reg[488]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(sreg[488]) );
  DFF \sreg_reg[487]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(sreg[487]) );
  DFF \sreg_reg[486]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(sreg[486]) );
  DFF \sreg_reg[485]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(sreg[485]) );
  DFF \sreg_reg[484]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(sreg[484]) );
  DFF \sreg_reg[483]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(sreg[483]) );
  DFF \sreg_reg[482]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(sreg[482]) );
  DFF \sreg_reg[481]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(sreg[481]) );
  DFF \sreg_reg[480]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(sreg[480]) );
  DFF \sreg_reg[479]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[478]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[477]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[476]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[475]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[474]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[473]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[472]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[471]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[470]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[469]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[468]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[467]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[466]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[465]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[464]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[463]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[462]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[461]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[460]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[459]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[458]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[457]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[456]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[455]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[454]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[453]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[452]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[451]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[450]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[449]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[448]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[447]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[446]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[445]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[444]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[443]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[442]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[441]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[440]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[439]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[438]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[437]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[436]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[435]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[434]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[433]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[432]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[431]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[430]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[429]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[428]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[427]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[426]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[425]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[424]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[423]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[422]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[421]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[420]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[419]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[418]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[417]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[416]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[415]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[414]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[413]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[412]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[411]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[410]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[409]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[408]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[407]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[406]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[405]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[404]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[403]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[402]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[401]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[400]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[399]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[398]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[397]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[396]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[395]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[394]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[393]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[392]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[391]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[390]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[389]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[388]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[387]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[386]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[385]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[384]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[383]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[382]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[381]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[380]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[379]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[378]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[377]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[376]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[375]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[374]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[373]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[372]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[371]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[370]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[369]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[368]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[367]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[366]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[365]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[364]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[363]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[362]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[361]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[360]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[359]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[358]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[357]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[356]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[355]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[354]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[353]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[352]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[351]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[350]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[349]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[348]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[347]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[346]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[345]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[344]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[343]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[342]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[341]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[340]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[339]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[338]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[337]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[336]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[335]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[334]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[333]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[332]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[331]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[330]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[329]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[328]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[327]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[326]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[325]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[324]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[323]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[322]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[321]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[320]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[319]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[318]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[317]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[316]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[315]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[314]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[313]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[312]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[311]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[310]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[309]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[308]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[307]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[306]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[305]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[304]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[303]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[302]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[301]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[300]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[299]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[298]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[297]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[296]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[295]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[294]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[293]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[292]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[291]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[290]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[289]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[288]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[287]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[286]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[285]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[284]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[283]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[282]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[281]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[280]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[279]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[278]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[277]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[276]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[275]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[274]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[273]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[272]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[271]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[270]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[269]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[268]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[267]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[266]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[265]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[264]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[263]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[262]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[261]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[260]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[259]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[258]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[257]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[256]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[255]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(sreg[255]) );
  DFF \sreg_reg[254]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[253]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[252]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[251]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[250]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[249]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[248]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[247]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[0]) );
  OR U11 ( .A(n79), .B(n80), .Z(n1) );
  NANDN U12 ( .A(n77), .B(n78), .Z(n2) );
  AND U13 ( .A(n1), .B(n2), .Z(n101) );
  XNOR U14 ( .A(n10304), .B(n10305), .Z(n10299) );
  XNOR U15 ( .A(n10344), .B(n10345), .Z(n10337) );
  XNOR U16 ( .A(n10414), .B(n10413), .Z(n10407) );
  XNOR U17 ( .A(n10476), .B(n10475), .Z(n10493) );
  XOR U18 ( .A(n62), .B(n60), .Z(n3) );
  NANDN U19 ( .A(n61), .B(n3), .Z(n4) );
  NAND U20 ( .A(n62), .B(n60), .Z(n5) );
  AND U21 ( .A(n4), .B(n5), .Z(n80) );
  XNOR U22 ( .A(n10337), .B(n10336), .Z(n10339) );
  XNOR U23 ( .A(n10299), .B(n10298), .Z(n10291) );
  XOR U24 ( .A(n10407), .B(n10406), .Z(n10409) );
  XNOR U25 ( .A(n10449), .B(n10448), .Z(n10441) );
  XOR U26 ( .A(n10493), .B(n10492), .Z(n10494) );
  XOR U27 ( .A(sreg[252]), .B(n75), .Z(n6) );
  NANDN U28 ( .A(n76), .B(n6), .Z(n7) );
  NAND U29 ( .A(sreg[252]), .B(n75), .Z(n8) );
  AND U30 ( .A(n7), .B(n8), .Z(n124) );
  NAND U31 ( .A(b[0]), .B(a[206]), .Z(n9) );
  XNOR U32 ( .A(b[1]), .B(n9), .Z(n10) );
  NANDN U33 ( .A(b[0]), .B(a[205]), .Z(n11) );
  AND U34 ( .A(n10), .B(n11), .Z(n8342) );
  NANDN U35 ( .A(b[0]), .B(a[255]), .Z(n12) );
  AND U36 ( .A(b[1]), .B(n12), .Z(n10386) );
  XOR U37 ( .A(n10291), .B(n10290), .Z(n10293) );
  XOR U38 ( .A(n10441), .B(n10440), .Z(n10443) );
  XNOR U39 ( .A(n10366), .B(n10365), .Z(n10368) );
  XNOR U40 ( .A(n10401), .B(n10400), .Z(n10403) );
  XNOR U41 ( .A(n10501), .B(n10500), .Z(n10503) );
  XNOR U42 ( .A(n10535), .B(n10534), .Z(n10537) );
  NAND U43 ( .A(n72), .B(n73), .Z(n13) );
  XOR U44 ( .A(n72), .B(n73), .Z(n14) );
  NAND U45 ( .A(n14), .B(sreg[251]), .Z(n15) );
  NAND U46 ( .A(n13), .B(n15), .Z(n75) );
  NAND U47 ( .A(n128), .B(n129), .Z(n16) );
  XOR U48 ( .A(n128), .B(n129), .Z(n17) );
  NAND U49 ( .A(n17), .B(sreg[254]), .Z(n18) );
  NAND U50 ( .A(n16), .B(n18), .Z(n164) );
  NAND U51 ( .A(n63), .B(n22), .Z(n19) );
  NAND U52 ( .A(n104), .B(n10424), .Z(n20) );
  NAND U53 ( .A(n139), .B(n10507), .Z(n21) );
  XNOR U54 ( .A(b[1]), .B(b[2]), .Z(n22) );
  IV U55 ( .A(n19), .Z(n23) );
  IV U56 ( .A(n22), .Z(n24) );
  IV U57 ( .A(n20), .Z(n25) );
  IV U58 ( .A(n21), .Z(n26) );
  AND U59 ( .A(b[0]), .B(a[0]), .Z(n28) );
  XOR U60 ( .A(n28), .B(sreg[248]), .Z(c[248]) );
  AND U61 ( .A(b[0]), .B(a[1]), .Z(n37) );
  NAND U62 ( .A(a[0]), .B(b[1]), .Z(n27) );
  XOR U63 ( .A(n37), .B(n27), .Z(n29) );
  XNOR U64 ( .A(sreg[249]), .B(n29), .Z(n31) );
  AND U65 ( .A(n28), .B(sreg[248]), .Z(n30) );
  XOR U66 ( .A(n31), .B(n30), .Z(c[249]) );
  NANDN U67 ( .A(n29), .B(sreg[249]), .Z(n33) );
  NAND U68 ( .A(n31), .B(n30), .Z(n32) );
  AND U69 ( .A(n33), .B(n32), .Z(n39) );
  XNOR U70 ( .A(n39), .B(sreg[250]), .Z(n41) );
  AND U71 ( .A(a[0]), .B(n24), .Z(n57) );
  NAND U72 ( .A(b[0]), .B(a[2]), .Z(n34) );
  XNOR U73 ( .A(b[1]), .B(n34), .Z(n36) );
  NANDN U74 ( .A(b[0]), .B(a[1]), .Z(n35) );
  NAND U75 ( .A(n36), .B(n35), .Z(n44) );
  XNOR U76 ( .A(n57), .B(n44), .Z(n45) );
  NOR U77 ( .A(n37), .B(a[0]), .Z(n38) );
  NAND U78 ( .A(b[1]), .B(n38), .Z(n46) );
  XNOR U79 ( .A(n45), .B(n46), .Z(n40) );
  XOR U80 ( .A(n41), .B(n40), .Z(c[250]) );
  NANDN U81 ( .A(n39), .B(sreg[250]), .Z(n43) );
  NAND U82 ( .A(n41), .B(n40), .Z(n42) );
  NAND U83 ( .A(n43), .B(n42), .Z(n73) );
  NANDN U84 ( .A(n44), .B(n57), .Z(n48) );
  NANDN U85 ( .A(n46), .B(n45), .Z(n47) );
  NAND U86 ( .A(n48), .B(n47), .Z(n62) );
  NAND U87 ( .A(b[0]), .B(a[3]), .Z(n49) );
  XNOR U88 ( .A(b[1]), .B(n49), .Z(n51) );
  NANDN U89 ( .A(b[0]), .B(a[2]), .Z(n50) );
  NAND U90 ( .A(n51), .B(n50), .Z(n70) );
  XOR U91 ( .A(b[3]), .B(b[2]), .Z(n63) );
  XOR U92 ( .A(b[3]), .B(a[0]), .Z(n52) );
  NAND U93 ( .A(n63), .B(n52), .Z(n53) );
  NANDN U94 ( .A(n53), .B(n22), .Z(n55) );
  XOR U95 ( .A(b[3]), .B(a[1]), .Z(n64) );
  NANDN U96 ( .A(n22), .B(n64), .Z(n54) );
  AND U97 ( .A(n55), .B(n54), .Z(n71) );
  XNOR U98 ( .A(n70), .B(n71), .Z(n61) );
  NAND U99 ( .A(b[1]), .B(b[2]), .Z(n56) );
  NAND U100 ( .A(b[3]), .B(n56), .Z(n10479) );
  NOR U101 ( .A(n10479), .B(n57), .Z(n60) );
  XOR U102 ( .A(n61), .B(n60), .Z(n58) );
  XNOR U103 ( .A(n62), .B(n58), .Z(n72) );
  XNOR U104 ( .A(sreg[251]), .B(n72), .Z(n59) );
  XNOR U105 ( .A(n73), .B(n59), .Z(c[251]) );
  NAND U106 ( .A(n23), .B(n64), .Z(n66) );
  XOR U107 ( .A(b[3]), .B(a[2]), .Z(n81) );
  NAND U108 ( .A(n24), .B(n81), .Z(n65) );
  AND U109 ( .A(n66), .B(n65), .Z(n95) );
  XNOR U110 ( .A(b[3]), .B(b[4]), .Z(n10424) );
  IV U111 ( .A(n10424), .Z(n10456) );
  AND U112 ( .A(a[0]), .B(n10456), .Z(n92) );
  NAND U113 ( .A(b[0]), .B(a[4]), .Z(n67) );
  XNOR U114 ( .A(b[1]), .B(n67), .Z(n69) );
  NANDN U115 ( .A(b[0]), .B(a[3]), .Z(n68) );
  NAND U116 ( .A(n69), .B(n68), .Z(n93) );
  XNOR U117 ( .A(n92), .B(n93), .Z(n94) );
  XNOR U118 ( .A(n95), .B(n94), .Z(n78) );
  OR U119 ( .A(n71), .B(n70), .Z(n77) );
  XOR U120 ( .A(n78), .B(n77), .Z(n79) );
  XNOR U121 ( .A(n80), .B(n79), .Z(n76) );
  XOR U122 ( .A(n75), .B(sreg[252]), .Z(n74) );
  XNOR U123 ( .A(n76), .B(n74), .Z(c[252]) );
  NAND U124 ( .A(n23), .B(n81), .Z(n83) );
  XOR U125 ( .A(b[3]), .B(a[3]), .Z(n110) );
  NAND U126 ( .A(n24), .B(n110), .Z(n82) );
  AND U127 ( .A(n83), .B(n82), .Z(n117) );
  NAND U128 ( .A(b[3]), .B(b[4]), .Z(n84) );
  NAND U129 ( .A(b[5]), .B(n84), .Z(n10524) );
  NOR U130 ( .A(n10524), .B(n92), .Z(n116) );
  XNOR U131 ( .A(n117), .B(n116), .Z(n119) );
  NAND U132 ( .A(b[0]), .B(a[5]), .Z(n85) );
  XNOR U133 ( .A(b[1]), .B(n85), .Z(n87) );
  NANDN U134 ( .A(b[0]), .B(a[4]), .Z(n86) );
  NAND U135 ( .A(n87), .B(n86), .Z(n108) );
  XOR U136 ( .A(b[5]), .B(b[4]), .Z(n104) );
  XOR U137 ( .A(b[5]), .B(a[0]), .Z(n88) );
  NAND U138 ( .A(n104), .B(n88), .Z(n89) );
  NANDN U139 ( .A(n89), .B(n10424), .Z(n91) );
  XOR U140 ( .A(b[5]), .B(a[1]), .Z(n105) );
  NANDN U141 ( .A(n10424), .B(n105), .Z(n90) );
  NAND U142 ( .A(n91), .B(n90), .Z(n109) );
  XNOR U143 ( .A(n108), .B(n109), .Z(n118) );
  XOR U144 ( .A(n119), .B(n118), .Z(n99) );
  NANDN U145 ( .A(n93), .B(n92), .Z(n97) );
  NANDN U146 ( .A(n95), .B(n94), .Z(n96) );
  AND U147 ( .A(n97), .B(n96), .Z(n98) );
  XNOR U148 ( .A(n99), .B(n98), .Z(n100) );
  XOR U149 ( .A(n101), .B(n100), .Z(n122) );
  XNOR U150 ( .A(n122), .B(sreg[253]), .Z(n123) );
  XNOR U151 ( .A(n124), .B(n123), .Z(c[253]) );
  NANDN U152 ( .A(n99), .B(n98), .Z(n103) );
  NAND U153 ( .A(n101), .B(n100), .Z(n102) );
  AND U154 ( .A(n103), .B(n102), .Z(n132) );
  NAND U155 ( .A(n25), .B(n105), .Z(n107) );
  XOR U156 ( .A(b[5]), .B(a[2]), .Z(n136) );
  NAND U157 ( .A(n10456), .B(n136), .Z(n106) );
  AND U158 ( .A(n107), .B(n106), .Z(n157) );
  ANDN U159 ( .B(n109), .A(n108), .Z(n156) );
  XNOR U160 ( .A(n157), .B(n156), .Z(n159) );
  NAND U161 ( .A(n23), .B(n110), .Z(n112) );
  XOR U162 ( .A(b[3]), .B(a[4]), .Z(n147) );
  NAND U163 ( .A(n24), .B(n147), .Z(n111) );
  AND U164 ( .A(n112), .B(n111), .Z(n153) );
  XNOR U165 ( .A(b[5]), .B(b[6]), .Z(n10507) );
  IV U166 ( .A(n10507), .Z(n10531) );
  AND U167 ( .A(a[0]), .B(n10531), .Z(n150) );
  NAND U168 ( .A(b[0]), .B(a[6]), .Z(n113) );
  XNOR U169 ( .A(b[1]), .B(n113), .Z(n115) );
  NANDN U170 ( .A(b[0]), .B(a[5]), .Z(n114) );
  NAND U171 ( .A(n115), .B(n114), .Z(n151) );
  XNOR U172 ( .A(n150), .B(n151), .Z(n152) );
  XNOR U173 ( .A(n153), .B(n152), .Z(n158) );
  XOR U174 ( .A(n159), .B(n158), .Z(n131) );
  NANDN U175 ( .A(n117), .B(n116), .Z(n121) );
  NAND U176 ( .A(n119), .B(n118), .Z(n120) );
  AND U177 ( .A(n121), .B(n120), .Z(n130) );
  XOR U178 ( .A(n131), .B(n130), .Z(n133) );
  XNOR U179 ( .A(n132), .B(n133), .Z(n129) );
  NANDN U180 ( .A(n122), .B(sreg[253]), .Z(n126) );
  NANDN U181 ( .A(n124), .B(n123), .Z(n125) );
  NAND U182 ( .A(n126), .B(n125), .Z(n128) );
  XNOR U183 ( .A(sreg[254]), .B(n128), .Z(n127) );
  XNOR U184 ( .A(n129), .B(n127), .Z(c[254]) );
  NANDN U185 ( .A(n131), .B(n130), .Z(n135) );
  OR U186 ( .A(n133), .B(n132), .Z(n134) );
  AND U187 ( .A(n135), .B(n134), .Z(n195) );
  NAND U188 ( .A(n25), .B(n136), .Z(n138) );
  XOR U189 ( .A(b[5]), .B(a[3]), .Z(n184) );
  NAND U190 ( .A(n10456), .B(n184), .Z(n137) );
  AND U191 ( .A(n138), .B(n137), .Z(n174) );
  XOR U192 ( .A(b[6]), .B(b[7]), .Z(n139) );
  XOR U193 ( .A(b[7]), .B(a[0]), .Z(n140) );
  NAND U194 ( .A(n26), .B(n140), .Z(n142) );
  XOR U195 ( .A(b[7]), .B(a[1]), .Z(n175) );
  NAND U196 ( .A(n10531), .B(n175), .Z(n141) );
  AND U197 ( .A(n142), .B(n141), .Z(n173) );
  XOR U198 ( .A(n174), .B(n173), .Z(n190) );
  ANDN U199 ( .B(b[7]), .A(n150), .Z(n143) );
  AND U200 ( .A(b[5]), .B(b[6]), .Z(n10558) );
  ANDN U201 ( .B(n143), .A(n10558), .Z(n188) );
  NAND U202 ( .A(b[0]), .B(a[7]), .Z(n144) );
  XNOR U203 ( .A(b[1]), .B(n144), .Z(n146) );
  NANDN U204 ( .A(b[0]), .B(a[6]), .Z(n145) );
  NAND U205 ( .A(n146), .B(n145), .Z(n187) );
  XNOR U206 ( .A(n188), .B(n187), .Z(n189) );
  XNOR U207 ( .A(n190), .B(n189), .Z(n167) );
  NANDN U208 ( .A(n19), .B(n147), .Z(n149) );
  XNOR U209 ( .A(b[3]), .B(a[5]), .Z(n178) );
  OR U210 ( .A(n178), .B(n22), .Z(n148) );
  NAND U211 ( .A(n149), .B(n148), .Z(n168) );
  XNOR U212 ( .A(n167), .B(n168), .Z(n169) );
  NANDN U213 ( .A(n151), .B(n150), .Z(n155) );
  NANDN U214 ( .A(n153), .B(n152), .Z(n154) );
  NAND U215 ( .A(n155), .B(n154), .Z(n170) );
  XNOR U216 ( .A(n169), .B(n170), .Z(n193) );
  NANDN U217 ( .A(n157), .B(n156), .Z(n161) );
  NAND U218 ( .A(n159), .B(n158), .Z(n160) );
  NAND U219 ( .A(n161), .B(n160), .Z(n194) );
  XOR U220 ( .A(n193), .B(n194), .Z(n196) );
  XOR U221 ( .A(n195), .B(n196), .Z(n162) );
  XNOR U222 ( .A(n162), .B(sreg[255]), .Z(n163) );
  XOR U223 ( .A(n164), .B(n163), .Z(c[255]) );
  NANDN U224 ( .A(n162), .B(sreg[255]), .Z(n166) );
  NAND U225 ( .A(n164), .B(n163), .Z(n165) );
  AND U226 ( .A(n166), .B(n165), .Z(n203) );
  IV U227 ( .A(n203), .Z(n200) );
  NANDN U228 ( .A(n168), .B(n167), .Z(n172) );
  NANDN U229 ( .A(n170), .B(n169), .Z(n171) );
  AND U230 ( .A(n172), .B(n171), .Z(n236) );
  NOR U231 ( .A(n174), .B(n173), .Z(n226) );
  NANDN U232 ( .A(n21), .B(n175), .Z(n177) );
  XNOR U233 ( .A(b[7]), .B(a[2]), .Z(n212) );
  OR U234 ( .A(n212), .B(n10507), .Z(n176) );
  AND U235 ( .A(n177), .B(n176), .Z(n224) );
  OR U236 ( .A(n178), .B(n19), .Z(n180) );
  XNOR U237 ( .A(b[3]), .B(a[6]), .Z(n215) );
  OR U238 ( .A(n215), .B(n22), .Z(n179) );
  NAND U239 ( .A(n180), .B(n179), .Z(n225) );
  XOR U240 ( .A(n224), .B(n225), .Z(n227) );
  XOR U241 ( .A(n226), .B(n227), .Z(n231) );
  NAND U242 ( .A(b[0]), .B(a[8]), .Z(n181) );
  XNOR U243 ( .A(b[1]), .B(n181), .Z(n183) );
  NANDN U244 ( .A(b[0]), .B(a[7]), .Z(n182) );
  NAND U245 ( .A(n183), .B(n182), .Z(n209) );
  NAND U246 ( .A(n25), .B(n184), .Z(n186) );
  XOR U247 ( .A(b[5]), .B(a[4]), .Z(n221) );
  NAND U248 ( .A(n10456), .B(n221), .Z(n185) );
  AND U249 ( .A(n186), .B(n185), .Z(n207) );
  AND U250 ( .A(b[7]), .B(a[0]), .Z(n206) );
  XNOR U251 ( .A(n207), .B(n206), .Z(n208) );
  XNOR U252 ( .A(n209), .B(n208), .Z(n230) );
  XNOR U253 ( .A(n231), .B(n230), .Z(n232) );
  NANDN U254 ( .A(n188), .B(n187), .Z(n192) );
  NANDN U255 ( .A(n190), .B(n189), .Z(n191) );
  NAND U256 ( .A(n192), .B(n191), .Z(n233) );
  XOR U257 ( .A(n232), .B(n233), .Z(n237) );
  XNOR U258 ( .A(n236), .B(n237), .Z(n238) );
  NANDN U259 ( .A(n194), .B(n193), .Z(n198) );
  OR U260 ( .A(n196), .B(n195), .Z(n197) );
  NAND U261 ( .A(n198), .B(n197), .Z(n239) );
  XNOR U262 ( .A(n238), .B(n239), .Z(n201) );
  XNOR U263 ( .A(sreg[256]), .B(n201), .Z(n199) );
  XNOR U264 ( .A(n200), .B(n199), .Z(c[256]) );
  AND U265 ( .A(sreg[256]), .B(n200), .Z(n202) );
  OR U266 ( .A(n202), .B(n201), .Z(n205) );
  ANDN U267 ( .B(n203), .A(sreg[256]), .Z(n204) );
  ANDN U268 ( .B(n205), .A(n204), .Z(n280) );
  NANDN U269 ( .A(n207), .B(n206), .Z(n211) );
  NANDN U270 ( .A(n209), .B(n208), .Z(n210) );
  AND U271 ( .A(n211), .B(n210), .Z(n273) );
  OR U272 ( .A(n212), .B(n21), .Z(n214) );
  XOR U273 ( .A(b[7]), .B(a[3]), .Z(n248) );
  NAND U274 ( .A(n10531), .B(n248), .Z(n213) );
  AND U275 ( .A(n214), .B(n213), .Z(n267) );
  OR U276 ( .A(n215), .B(n19), .Z(n217) );
  XOR U277 ( .A(b[3]), .B(a[7]), .Z(n251) );
  NAND U278 ( .A(n24), .B(n251), .Z(n216) );
  NAND U279 ( .A(n217), .B(n216), .Z(n266) );
  XNOR U280 ( .A(n267), .B(n266), .Z(n268) );
  NAND U281 ( .A(b[0]), .B(a[9]), .Z(n218) );
  XNOR U282 ( .A(b[1]), .B(n218), .Z(n220) );
  NANDN U283 ( .A(b[0]), .B(a[8]), .Z(n219) );
  NAND U284 ( .A(n220), .B(n219), .Z(n263) );
  NAND U285 ( .A(n25), .B(n221), .Z(n223) );
  XOR U286 ( .A(b[5]), .B(a[5]), .Z(n257) );
  NAND U287 ( .A(n10456), .B(n257), .Z(n222) );
  AND U288 ( .A(n223), .B(n222), .Z(n261) );
  AND U289 ( .A(b[7]), .B(a[1]), .Z(n260) );
  XNOR U290 ( .A(n261), .B(n260), .Z(n262) );
  XOR U291 ( .A(n263), .B(n262), .Z(n269) );
  XNOR U292 ( .A(n268), .B(n269), .Z(n272) );
  XNOR U293 ( .A(n273), .B(n272), .Z(n275) );
  NANDN U294 ( .A(n225), .B(n224), .Z(n229) );
  OR U295 ( .A(n227), .B(n226), .Z(n228) );
  AND U296 ( .A(n229), .B(n228), .Z(n274) );
  XOR U297 ( .A(n275), .B(n274), .Z(n243) );
  NANDN U298 ( .A(n231), .B(n230), .Z(n235) );
  NANDN U299 ( .A(n233), .B(n232), .Z(n234) );
  AND U300 ( .A(n235), .B(n234), .Z(n242) );
  XNOR U301 ( .A(n243), .B(n242), .Z(n245) );
  NANDN U302 ( .A(n237), .B(n236), .Z(n241) );
  NANDN U303 ( .A(n239), .B(n238), .Z(n240) );
  AND U304 ( .A(n241), .B(n240), .Z(n244) );
  XOR U305 ( .A(n245), .B(n244), .Z(n278) );
  XNOR U306 ( .A(n278), .B(sreg[257]), .Z(n279) );
  XOR U307 ( .A(n280), .B(n279), .Z(c[257]) );
  NANDN U308 ( .A(n243), .B(n242), .Z(n247) );
  NAND U309 ( .A(n245), .B(n244), .Z(n246) );
  AND U310 ( .A(n247), .B(n246), .Z(n290) );
  NAND U311 ( .A(n26), .B(n248), .Z(n250) );
  XOR U312 ( .A(b[7]), .B(a[4]), .Z(n300) );
  NAND U313 ( .A(n10531), .B(n300), .Z(n249) );
  AND U314 ( .A(n250), .B(n249), .Z(n319) );
  NAND U315 ( .A(n23), .B(n251), .Z(n253) );
  XOR U316 ( .A(b[3]), .B(a[8]), .Z(n303) );
  NAND U317 ( .A(n24), .B(n303), .Z(n252) );
  NAND U318 ( .A(n253), .B(n252), .Z(n318) );
  XNOR U319 ( .A(n319), .B(n318), .Z(n321) );
  NAND U320 ( .A(b[0]), .B(a[10]), .Z(n254) );
  XNOR U321 ( .A(b[1]), .B(n254), .Z(n256) );
  NANDN U322 ( .A(b[0]), .B(a[9]), .Z(n255) );
  NAND U323 ( .A(n256), .B(n255), .Z(n315) );
  NAND U324 ( .A(n25), .B(n257), .Z(n259) );
  XOR U325 ( .A(b[5]), .B(a[6]), .Z(n309) );
  NAND U326 ( .A(n10456), .B(n309), .Z(n258) );
  AND U327 ( .A(n259), .B(n258), .Z(n313) );
  AND U328 ( .A(b[7]), .B(a[2]), .Z(n312) );
  XNOR U329 ( .A(n313), .B(n312), .Z(n314) );
  XNOR U330 ( .A(n315), .B(n314), .Z(n320) );
  XOR U331 ( .A(n321), .B(n320), .Z(n295) );
  NANDN U332 ( .A(n261), .B(n260), .Z(n265) );
  NANDN U333 ( .A(n263), .B(n262), .Z(n264) );
  AND U334 ( .A(n265), .B(n264), .Z(n294) );
  XNOR U335 ( .A(n295), .B(n294), .Z(n296) );
  NANDN U336 ( .A(n267), .B(n266), .Z(n271) );
  NANDN U337 ( .A(n269), .B(n268), .Z(n270) );
  NAND U338 ( .A(n271), .B(n270), .Z(n297) );
  XNOR U339 ( .A(n296), .B(n297), .Z(n288) );
  NANDN U340 ( .A(n273), .B(n272), .Z(n277) );
  NAND U341 ( .A(n275), .B(n274), .Z(n276) );
  NAND U342 ( .A(n277), .B(n276), .Z(n289) );
  XOR U343 ( .A(n288), .B(n289), .Z(n291) );
  XOR U344 ( .A(n290), .B(n291), .Z(n283) );
  XNOR U345 ( .A(n283), .B(sreg[258]), .Z(n285) );
  NANDN U346 ( .A(n278), .B(sreg[257]), .Z(n282) );
  NAND U347 ( .A(n280), .B(n279), .Z(n281) );
  NAND U348 ( .A(n282), .B(n281), .Z(n284) );
  XOR U349 ( .A(n285), .B(n284), .Z(c[258]) );
  NANDN U350 ( .A(n283), .B(sreg[258]), .Z(n287) );
  NAND U351 ( .A(n285), .B(n284), .Z(n286) );
  AND U352 ( .A(n287), .B(n286), .Z(n362) );
  NANDN U353 ( .A(n289), .B(n288), .Z(n293) );
  OR U354 ( .A(n291), .B(n290), .Z(n292) );
  AND U355 ( .A(n293), .B(n292), .Z(n327) );
  NANDN U356 ( .A(n295), .B(n294), .Z(n299) );
  NANDN U357 ( .A(n297), .B(n296), .Z(n298) );
  AND U358 ( .A(n299), .B(n298), .Z(n325) );
  NAND U359 ( .A(n26), .B(n300), .Z(n302) );
  XOR U360 ( .A(b[7]), .B(a[5]), .Z(n336) );
  NAND U361 ( .A(n10531), .B(n336), .Z(n301) );
  AND U362 ( .A(n302), .B(n301), .Z(n355) );
  NAND U363 ( .A(n23), .B(n303), .Z(n305) );
  XOR U364 ( .A(b[3]), .B(a[9]), .Z(n339) );
  NAND U365 ( .A(n24), .B(n339), .Z(n304) );
  NAND U366 ( .A(n305), .B(n304), .Z(n354) );
  XNOR U367 ( .A(n355), .B(n354), .Z(n357) );
  NAND U368 ( .A(b[0]), .B(a[11]), .Z(n306) );
  XNOR U369 ( .A(b[1]), .B(n306), .Z(n308) );
  NANDN U370 ( .A(b[0]), .B(a[10]), .Z(n307) );
  NAND U371 ( .A(n308), .B(n307), .Z(n351) );
  NAND U372 ( .A(n25), .B(n309), .Z(n311) );
  XOR U373 ( .A(b[5]), .B(a[7]), .Z(n345) );
  NAND U374 ( .A(n10456), .B(n345), .Z(n310) );
  AND U375 ( .A(n311), .B(n310), .Z(n349) );
  AND U376 ( .A(b[7]), .B(a[3]), .Z(n348) );
  XNOR U377 ( .A(n349), .B(n348), .Z(n350) );
  XNOR U378 ( .A(n351), .B(n350), .Z(n356) );
  XOR U379 ( .A(n357), .B(n356), .Z(n331) );
  NANDN U380 ( .A(n313), .B(n312), .Z(n317) );
  NANDN U381 ( .A(n315), .B(n314), .Z(n316) );
  AND U382 ( .A(n317), .B(n316), .Z(n330) );
  XNOR U383 ( .A(n331), .B(n330), .Z(n332) );
  NANDN U384 ( .A(n319), .B(n318), .Z(n323) );
  NAND U385 ( .A(n321), .B(n320), .Z(n322) );
  NAND U386 ( .A(n323), .B(n322), .Z(n333) );
  XNOR U387 ( .A(n332), .B(n333), .Z(n324) );
  XNOR U388 ( .A(n325), .B(n324), .Z(n326) );
  XNOR U389 ( .A(n327), .B(n326), .Z(n360) );
  XNOR U390 ( .A(sreg[259]), .B(n360), .Z(n361) );
  XNOR U391 ( .A(n362), .B(n361), .Z(c[259]) );
  NANDN U392 ( .A(n325), .B(n324), .Z(n329) );
  NANDN U393 ( .A(n327), .B(n326), .Z(n328) );
  AND U394 ( .A(n329), .B(n328), .Z(n367) );
  NANDN U395 ( .A(n331), .B(n330), .Z(n335) );
  NANDN U396 ( .A(n333), .B(n332), .Z(n334) );
  AND U397 ( .A(n335), .B(n334), .Z(n366) );
  NAND U398 ( .A(n26), .B(n336), .Z(n338) );
  XOR U399 ( .A(b[7]), .B(a[6]), .Z(n377) );
  NAND U400 ( .A(n10531), .B(n377), .Z(n337) );
  AND U401 ( .A(n338), .B(n337), .Z(n396) );
  NAND U402 ( .A(n23), .B(n339), .Z(n341) );
  XOR U403 ( .A(b[3]), .B(a[10]), .Z(n380) );
  NAND U404 ( .A(n24), .B(n380), .Z(n340) );
  NAND U405 ( .A(n341), .B(n340), .Z(n395) );
  XNOR U406 ( .A(n396), .B(n395), .Z(n398) );
  NAND U407 ( .A(b[0]), .B(a[12]), .Z(n342) );
  XNOR U408 ( .A(b[1]), .B(n342), .Z(n344) );
  NANDN U409 ( .A(b[0]), .B(a[11]), .Z(n343) );
  NAND U410 ( .A(n344), .B(n343), .Z(n392) );
  NAND U411 ( .A(n25), .B(n345), .Z(n347) );
  XOR U412 ( .A(b[5]), .B(a[8]), .Z(n383) );
  NAND U413 ( .A(n10456), .B(n383), .Z(n346) );
  AND U414 ( .A(n347), .B(n346), .Z(n390) );
  AND U415 ( .A(b[7]), .B(a[4]), .Z(n389) );
  XNOR U416 ( .A(n390), .B(n389), .Z(n391) );
  XNOR U417 ( .A(n392), .B(n391), .Z(n397) );
  XOR U418 ( .A(n398), .B(n397), .Z(n372) );
  NANDN U419 ( .A(n349), .B(n348), .Z(n353) );
  NANDN U420 ( .A(n351), .B(n350), .Z(n352) );
  AND U421 ( .A(n353), .B(n352), .Z(n371) );
  XNOR U422 ( .A(n372), .B(n371), .Z(n373) );
  NANDN U423 ( .A(n355), .B(n354), .Z(n359) );
  NAND U424 ( .A(n357), .B(n356), .Z(n358) );
  NAND U425 ( .A(n359), .B(n358), .Z(n374) );
  XNOR U426 ( .A(n373), .B(n374), .Z(n365) );
  XOR U427 ( .A(n366), .B(n365), .Z(n368) );
  XOR U428 ( .A(n367), .B(n368), .Z(n401) );
  XNOR U429 ( .A(n401), .B(sreg[260]), .Z(n403) );
  NANDN U430 ( .A(sreg[259]), .B(n360), .Z(n364) );
  NAND U431 ( .A(n362), .B(n361), .Z(n363) );
  AND U432 ( .A(n364), .B(n363), .Z(n402) );
  XOR U433 ( .A(n403), .B(n402), .Z(c[260]) );
  NANDN U434 ( .A(n366), .B(n365), .Z(n370) );
  OR U435 ( .A(n368), .B(n367), .Z(n369) );
  AND U436 ( .A(n370), .B(n369), .Z(n413) );
  NANDN U437 ( .A(n372), .B(n371), .Z(n376) );
  NANDN U438 ( .A(n374), .B(n373), .Z(n375) );
  AND U439 ( .A(n376), .B(n375), .Z(n412) );
  NAND U440 ( .A(n26), .B(n377), .Z(n379) );
  XOR U441 ( .A(b[7]), .B(a[7]), .Z(n423) );
  NAND U442 ( .A(n10531), .B(n423), .Z(n378) );
  AND U443 ( .A(n379), .B(n378), .Z(n442) );
  NAND U444 ( .A(n23), .B(n380), .Z(n382) );
  XOR U445 ( .A(b[3]), .B(a[11]), .Z(n426) );
  NAND U446 ( .A(n24), .B(n426), .Z(n381) );
  NAND U447 ( .A(n382), .B(n381), .Z(n441) );
  XNOR U448 ( .A(n442), .B(n441), .Z(n444) );
  NAND U449 ( .A(n25), .B(n383), .Z(n385) );
  XOR U450 ( .A(b[5]), .B(a[9]), .Z(n432) );
  NAND U451 ( .A(n10456), .B(n432), .Z(n384) );
  AND U452 ( .A(n385), .B(n384), .Z(n436) );
  AND U453 ( .A(b[7]), .B(a[5]), .Z(n435) );
  XNOR U454 ( .A(n436), .B(n435), .Z(n437) );
  NAND U455 ( .A(b[0]), .B(a[13]), .Z(n386) );
  XNOR U456 ( .A(b[1]), .B(n386), .Z(n388) );
  NANDN U457 ( .A(b[0]), .B(a[12]), .Z(n387) );
  NAND U458 ( .A(n388), .B(n387), .Z(n438) );
  XNOR U459 ( .A(n437), .B(n438), .Z(n443) );
  XOR U460 ( .A(n444), .B(n443), .Z(n418) );
  NANDN U461 ( .A(n390), .B(n389), .Z(n394) );
  NANDN U462 ( .A(n392), .B(n391), .Z(n393) );
  AND U463 ( .A(n394), .B(n393), .Z(n417) );
  XNOR U464 ( .A(n418), .B(n417), .Z(n419) );
  NANDN U465 ( .A(n396), .B(n395), .Z(n400) );
  NAND U466 ( .A(n398), .B(n397), .Z(n399) );
  NAND U467 ( .A(n400), .B(n399), .Z(n420) );
  XNOR U468 ( .A(n419), .B(n420), .Z(n411) );
  XOR U469 ( .A(n412), .B(n411), .Z(n414) );
  XOR U470 ( .A(n413), .B(n414), .Z(n406) );
  XNOR U471 ( .A(n406), .B(sreg[261]), .Z(n408) );
  NANDN U472 ( .A(n401), .B(sreg[260]), .Z(n405) );
  NAND U473 ( .A(n403), .B(n402), .Z(n404) );
  NAND U474 ( .A(n405), .B(n404), .Z(n407) );
  XOR U475 ( .A(n408), .B(n407), .Z(c[261]) );
  NANDN U476 ( .A(n406), .B(sreg[261]), .Z(n410) );
  NAND U477 ( .A(n408), .B(n407), .Z(n409) );
  AND U478 ( .A(n410), .B(n409), .Z(n485) );
  NANDN U479 ( .A(n412), .B(n411), .Z(n416) );
  OR U480 ( .A(n414), .B(n413), .Z(n415) );
  AND U481 ( .A(n416), .B(n415), .Z(n450) );
  NANDN U482 ( .A(n418), .B(n417), .Z(n422) );
  NANDN U483 ( .A(n420), .B(n419), .Z(n421) );
  AND U484 ( .A(n422), .B(n421), .Z(n448) );
  NAND U485 ( .A(n26), .B(n423), .Z(n425) );
  XOR U486 ( .A(b[7]), .B(a[8]), .Z(n459) );
  NAND U487 ( .A(n10531), .B(n459), .Z(n424) );
  AND U488 ( .A(n425), .B(n424), .Z(n478) );
  NAND U489 ( .A(n23), .B(n426), .Z(n428) );
  XOR U490 ( .A(b[3]), .B(a[12]), .Z(n462) );
  NAND U491 ( .A(n24), .B(n462), .Z(n427) );
  NAND U492 ( .A(n428), .B(n427), .Z(n477) );
  XNOR U493 ( .A(n478), .B(n477), .Z(n480) );
  NAND U494 ( .A(b[0]), .B(a[14]), .Z(n429) );
  XNOR U495 ( .A(b[1]), .B(n429), .Z(n431) );
  NANDN U496 ( .A(b[0]), .B(a[13]), .Z(n430) );
  NAND U497 ( .A(n431), .B(n430), .Z(n474) );
  NAND U498 ( .A(n25), .B(n432), .Z(n434) );
  XOR U499 ( .A(b[5]), .B(a[10]), .Z(n468) );
  NAND U500 ( .A(n10456), .B(n468), .Z(n433) );
  AND U501 ( .A(n434), .B(n433), .Z(n472) );
  AND U502 ( .A(b[7]), .B(a[6]), .Z(n471) );
  XNOR U503 ( .A(n472), .B(n471), .Z(n473) );
  XNOR U504 ( .A(n474), .B(n473), .Z(n479) );
  XOR U505 ( .A(n480), .B(n479), .Z(n454) );
  NANDN U506 ( .A(n436), .B(n435), .Z(n440) );
  NANDN U507 ( .A(n438), .B(n437), .Z(n439) );
  AND U508 ( .A(n440), .B(n439), .Z(n453) );
  XNOR U509 ( .A(n454), .B(n453), .Z(n455) );
  NANDN U510 ( .A(n442), .B(n441), .Z(n446) );
  NAND U511 ( .A(n444), .B(n443), .Z(n445) );
  NAND U512 ( .A(n446), .B(n445), .Z(n456) );
  XNOR U513 ( .A(n455), .B(n456), .Z(n447) );
  XNOR U514 ( .A(n448), .B(n447), .Z(n449) );
  XNOR U515 ( .A(n450), .B(n449), .Z(n483) );
  XNOR U516 ( .A(sreg[262]), .B(n483), .Z(n484) );
  XNOR U517 ( .A(n485), .B(n484), .Z(c[262]) );
  NANDN U518 ( .A(n448), .B(n447), .Z(n452) );
  NANDN U519 ( .A(n450), .B(n449), .Z(n451) );
  AND U520 ( .A(n452), .B(n451), .Z(n496) );
  NANDN U521 ( .A(n454), .B(n453), .Z(n458) );
  NANDN U522 ( .A(n456), .B(n455), .Z(n457) );
  AND U523 ( .A(n458), .B(n457), .Z(n494) );
  NAND U524 ( .A(n26), .B(n459), .Z(n461) );
  XOR U525 ( .A(b[7]), .B(a[9]), .Z(n505) );
  NAND U526 ( .A(n10531), .B(n505), .Z(n460) );
  AND U527 ( .A(n461), .B(n460), .Z(n524) );
  NAND U528 ( .A(n23), .B(n462), .Z(n464) );
  XOR U529 ( .A(b[3]), .B(a[13]), .Z(n508) );
  NAND U530 ( .A(n24), .B(n508), .Z(n463) );
  NAND U531 ( .A(n464), .B(n463), .Z(n523) );
  XNOR U532 ( .A(n524), .B(n523), .Z(n526) );
  NAND U533 ( .A(b[0]), .B(a[15]), .Z(n465) );
  XNOR U534 ( .A(b[1]), .B(n465), .Z(n467) );
  NANDN U535 ( .A(b[0]), .B(a[14]), .Z(n466) );
  NAND U536 ( .A(n467), .B(n466), .Z(n520) );
  NAND U537 ( .A(n25), .B(n468), .Z(n470) );
  XOR U538 ( .A(b[5]), .B(a[11]), .Z(n511) );
  NAND U539 ( .A(n10456), .B(n511), .Z(n469) );
  AND U540 ( .A(n470), .B(n469), .Z(n518) );
  AND U541 ( .A(b[7]), .B(a[7]), .Z(n517) );
  XNOR U542 ( .A(n518), .B(n517), .Z(n519) );
  XNOR U543 ( .A(n520), .B(n519), .Z(n525) );
  XOR U544 ( .A(n526), .B(n525), .Z(n500) );
  NANDN U545 ( .A(n472), .B(n471), .Z(n476) );
  NANDN U546 ( .A(n474), .B(n473), .Z(n475) );
  AND U547 ( .A(n476), .B(n475), .Z(n499) );
  XNOR U548 ( .A(n500), .B(n499), .Z(n501) );
  NANDN U549 ( .A(n478), .B(n477), .Z(n482) );
  NAND U550 ( .A(n480), .B(n479), .Z(n481) );
  NAND U551 ( .A(n482), .B(n481), .Z(n502) );
  XNOR U552 ( .A(n501), .B(n502), .Z(n493) );
  XNOR U553 ( .A(n494), .B(n493), .Z(n495) );
  XNOR U554 ( .A(n496), .B(n495), .Z(n488) );
  XNOR U555 ( .A(sreg[263]), .B(n488), .Z(n490) );
  NANDN U556 ( .A(sreg[262]), .B(n483), .Z(n487) );
  NAND U557 ( .A(n485), .B(n484), .Z(n486) );
  NAND U558 ( .A(n487), .B(n486), .Z(n489) );
  XNOR U559 ( .A(n490), .B(n489), .Z(c[263]) );
  NANDN U560 ( .A(sreg[263]), .B(n488), .Z(n492) );
  NAND U561 ( .A(n490), .B(n489), .Z(n491) );
  AND U562 ( .A(n492), .B(n491), .Z(n531) );
  NANDN U563 ( .A(n494), .B(n493), .Z(n498) );
  NANDN U564 ( .A(n496), .B(n495), .Z(n497) );
  AND U565 ( .A(n498), .B(n497), .Z(n536) );
  NANDN U566 ( .A(n500), .B(n499), .Z(n504) );
  NANDN U567 ( .A(n502), .B(n501), .Z(n503) );
  AND U568 ( .A(n504), .B(n503), .Z(n535) );
  NAND U569 ( .A(n26), .B(n505), .Z(n507) );
  XOR U570 ( .A(b[7]), .B(a[10]), .Z(n546) );
  NAND U571 ( .A(n10531), .B(n546), .Z(n506) );
  AND U572 ( .A(n507), .B(n506), .Z(n565) );
  NAND U573 ( .A(n23), .B(n508), .Z(n510) );
  XOR U574 ( .A(b[3]), .B(a[14]), .Z(n549) );
  NAND U575 ( .A(n24), .B(n549), .Z(n509) );
  NAND U576 ( .A(n510), .B(n509), .Z(n564) );
  XNOR U577 ( .A(n565), .B(n564), .Z(n567) );
  NAND U578 ( .A(n25), .B(n511), .Z(n513) );
  XOR U579 ( .A(b[5]), .B(a[12]), .Z(n555) );
  NAND U580 ( .A(n10456), .B(n555), .Z(n512) );
  AND U581 ( .A(n513), .B(n512), .Z(n559) );
  AND U582 ( .A(b[7]), .B(a[8]), .Z(n558) );
  XNOR U583 ( .A(n559), .B(n558), .Z(n560) );
  NAND U584 ( .A(b[0]), .B(a[16]), .Z(n514) );
  XNOR U585 ( .A(b[1]), .B(n514), .Z(n516) );
  NANDN U586 ( .A(b[0]), .B(a[15]), .Z(n515) );
  NAND U587 ( .A(n516), .B(n515), .Z(n561) );
  XNOR U588 ( .A(n560), .B(n561), .Z(n566) );
  XOR U589 ( .A(n567), .B(n566), .Z(n541) );
  NANDN U590 ( .A(n518), .B(n517), .Z(n522) );
  NANDN U591 ( .A(n520), .B(n519), .Z(n521) );
  AND U592 ( .A(n522), .B(n521), .Z(n540) );
  XNOR U593 ( .A(n541), .B(n540), .Z(n542) );
  NANDN U594 ( .A(n524), .B(n523), .Z(n528) );
  NAND U595 ( .A(n526), .B(n525), .Z(n527) );
  NAND U596 ( .A(n528), .B(n527), .Z(n543) );
  XNOR U597 ( .A(n542), .B(n543), .Z(n534) );
  XOR U598 ( .A(n535), .B(n534), .Z(n537) );
  XOR U599 ( .A(n536), .B(n537), .Z(n529) );
  XNOR U600 ( .A(n529), .B(sreg[264]), .Z(n530) );
  XOR U601 ( .A(n531), .B(n530), .Z(c[264]) );
  NANDN U602 ( .A(n529), .B(sreg[264]), .Z(n533) );
  NAND U603 ( .A(n531), .B(n530), .Z(n532) );
  AND U604 ( .A(n533), .B(n532), .Z(n608) );
  NANDN U605 ( .A(n535), .B(n534), .Z(n539) );
  OR U606 ( .A(n537), .B(n536), .Z(n538) );
  AND U607 ( .A(n539), .B(n538), .Z(n573) );
  NANDN U608 ( .A(n541), .B(n540), .Z(n545) );
  NANDN U609 ( .A(n543), .B(n542), .Z(n544) );
  AND U610 ( .A(n545), .B(n544), .Z(n571) );
  NAND U611 ( .A(n26), .B(n546), .Z(n548) );
  XOR U612 ( .A(b[7]), .B(a[11]), .Z(n582) );
  NAND U613 ( .A(n10531), .B(n582), .Z(n547) );
  AND U614 ( .A(n548), .B(n547), .Z(n601) );
  NAND U615 ( .A(n23), .B(n549), .Z(n551) );
  XOR U616 ( .A(b[3]), .B(a[15]), .Z(n585) );
  NAND U617 ( .A(n24), .B(n585), .Z(n550) );
  NAND U618 ( .A(n551), .B(n550), .Z(n600) );
  XNOR U619 ( .A(n601), .B(n600), .Z(n603) );
  NAND U620 ( .A(b[0]), .B(a[17]), .Z(n552) );
  XNOR U621 ( .A(b[1]), .B(n552), .Z(n554) );
  NANDN U622 ( .A(b[0]), .B(a[16]), .Z(n553) );
  NAND U623 ( .A(n554), .B(n553), .Z(n597) );
  NAND U624 ( .A(n25), .B(n555), .Z(n557) );
  XOR U625 ( .A(b[5]), .B(a[13]), .Z(n591) );
  NAND U626 ( .A(n10456), .B(n591), .Z(n556) );
  AND U627 ( .A(n557), .B(n556), .Z(n595) );
  AND U628 ( .A(b[7]), .B(a[9]), .Z(n594) );
  XNOR U629 ( .A(n595), .B(n594), .Z(n596) );
  XNOR U630 ( .A(n597), .B(n596), .Z(n602) );
  XOR U631 ( .A(n603), .B(n602), .Z(n577) );
  NANDN U632 ( .A(n559), .B(n558), .Z(n563) );
  NANDN U633 ( .A(n561), .B(n560), .Z(n562) );
  AND U634 ( .A(n563), .B(n562), .Z(n576) );
  XNOR U635 ( .A(n577), .B(n576), .Z(n578) );
  NANDN U636 ( .A(n565), .B(n564), .Z(n569) );
  NAND U637 ( .A(n567), .B(n566), .Z(n568) );
  NAND U638 ( .A(n569), .B(n568), .Z(n579) );
  XNOR U639 ( .A(n578), .B(n579), .Z(n570) );
  XNOR U640 ( .A(n571), .B(n570), .Z(n572) );
  XNOR U641 ( .A(n573), .B(n572), .Z(n606) );
  XNOR U642 ( .A(sreg[265]), .B(n606), .Z(n607) );
  XNOR U643 ( .A(n608), .B(n607), .Z(c[265]) );
  NANDN U644 ( .A(n571), .B(n570), .Z(n575) );
  NANDN U645 ( .A(n573), .B(n572), .Z(n574) );
  AND U646 ( .A(n575), .B(n574), .Z(n619) );
  NANDN U647 ( .A(n577), .B(n576), .Z(n581) );
  NANDN U648 ( .A(n579), .B(n578), .Z(n580) );
  AND U649 ( .A(n581), .B(n580), .Z(n617) );
  NAND U650 ( .A(n26), .B(n582), .Z(n584) );
  XOR U651 ( .A(b[7]), .B(a[12]), .Z(n628) );
  NAND U652 ( .A(n10531), .B(n628), .Z(n583) );
  AND U653 ( .A(n584), .B(n583), .Z(n647) );
  NAND U654 ( .A(n23), .B(n585), .Z(n587) );
  XOR U655 ( .A(b[3]), .B(a[16]), .Z(n631) );
  NAND U656 ( .A(n24), .B(n631), .Z(n586) );
  NAND U657 ( .A(n587), .B(n586), .Z(n646) );
  XNOR U658 ( .A(n647), .B(n646), .Z(n649) );
  NAND U659 ( .A(b[0]), .B(a[18]), .Z(n588) );
  XNOR U660 ( .A(b[1]), .B(n588), .Z(n590) );
  NANDN U661 ( .A(b[0]), .B(a[17]), .Z(n589) );
  NAND U662 ( .A(n590), .B(n589), .Z(n643) );
  NAND U663 ( .A(n25), .B(n591), .Z(n593) );
  XOR U664 ( .A(b[5]), .B(a[14]), .Z(n637) );
  NAND U665 ( .A(n10456), .B(n637), .Z(n592) );
  AND U666 ( .A(n593), .B(n592), .Z(n641) );
  AND U667 ( .A(b[7]), .B(a[10]), .Z(n640) );
  XNOR U668 ( .A(n641), .B(n640), .Z(n642) );
  XNOR U669 ( .A(n643), .B(n642), .Z(n648) );
  XOR U670 ( .A(n649), .B(n648), .Z(n623) );
  NANDN U671 ( .A(n595), .B(n594), .Z(n599) );
  NANDN U672 ( .A(n597), .B(n596), .Z(n598) );
  AND U673 ( .A(n599), .B(n598), .Z(n622) );
  XNOR U674 ( .A(n623), .B(n622), .Z(n624) );
  NANDN U675 ( .A(n601), .B(n600), .Z(n605) );
  NAND U676 ( .A(n603), .B(n602), .Z(n604) );
  NAND U677 ( .A(n605), .B(n604), .Z(n625) );
  XNOR U678 ( .A(n624), .B(n625), .Z(n616) );
  XNOR U679 ( .A(n617), .B(n616), .Z(n618) );
  XNOR U680 ( .A(n619), .B(n618), .Z(n611) );
  XNOR U681 ( .A(sreg[266]), .B(n611), .Z(n613) );
  NANDN U682 ( .A(sreg[265]), .B(n606), .Z(n610) );
  NAND U683 ( .A(n608), .B(n607), .Z(n609) );
  NAND U684 ( .A(n610), .B(n609), .Z(n612) );
  XNOR U685 ( .A(n613), .B(n612), .Z(c[266]) );
  NANDN U686 ( .A(sreg[266]), .B(n611), .Z(n615) );
  NAND U687 ( .A(n613), .B(n612), .Z(n614) );
  AND U688 ( .A(n615), .B(n614), .Z(n654) );
  NANDN U689 ( .A(n617), .B(n616), .Z(n621) );
  NANDN U690 ( .A(n619), .B(n618), .Z(n620) );
  AND U691 ( .A(n621), .B(n620), .Z(n659) );
  NANDN U692 ( .A(n623), .B(n622), .Z(n627) );
  NANDN U693 ( .A(n625), .B(n624), .Z(n626) );
  AND U694 ( .A(n627), .B(n626), .Z(n658) );
  NAND U695 ( .A(n26), .B(n628), .Z(n630) );
  XOR U696 ( .A(b[7]), .B(a[13]), .Z(n669) );
  NAND U697 ( .A(n10531), .B(n669), .Z(n629) );
  AND U698 ( .A(n630), .B(n629), .Z(n688) );
  NAND U699 ( .A(n23), .B(n631), .Z(n633) );
  XOR U700 ( .A(b[3]), .B(a[17]), .Z(n672) );
  NAND U701 ( .A(n24), .B(n672), .Z(n632) );
  NAND U702 ( .A(n633), .B(n632), .Z(n687) );
  XNOR U703 ( .A(n688), .B(n687), .Z(n690) );
  NAND U704 ( .A(b[0]), .B(a[19]), .Z(n634) );
  XNOR U705 ( .A(b[1]), .B(n634), .Z(n636) );
  NANDN U706 ( .A(b[0]), .B(a[18]), .Z(n635) );
  NAND U707 ( .A(n636), .B(n635), .Z(n684) );
  NAND U708 ( .A(n25), .B(n637), .Z(n639) );
  XOR U709 ( .A(b[5]), .B(a[15]), .Z(n675) );
  NAND U710 ( .A(n10456), .B(n675), .Z(n638) );
  AND U711 ( .A(n639), .B(n638), .Z(n682) );
  AND U712 ( .A(b[7]), .B(a[11]), .Z(n681) );
  XNOR U713 ( .A(n682), .B(n681), .Z(n683) );
  XNOR U714 ( .A(n684), .B(n683), .Z(n689) );
  XOR U715 ( .A(n690), .B(n689), .Z(n664) );
  NANDN U716 ( .A(n641), .B(n640), .Z(n645) );
  NANDN U717 ( .A(n643), .B(n642), .Z(n644) );
  AND U718 ( .A(n645), .B(n644), .Z(n663) );
  XNOR U719 ( .A(n664), .B(n663), .Z(n665) );
  NANDN U720 ( .A(n647), .B(n646), .Z(n651) );
  NAND U721 ( .A(n649), .B(n648), .Z(n650) );
  NAND U722 ( .A(n651), .B(n650), .Z(n666) );
  XNOR U723 ( .A(n665), .B(n666), .Z(n657) );
  XOR U724 ( .A(n658), .B(n657), .Z(n660) );
  XOR U725 ( .A(n659), .B(n660), .Z(n652) );
  XNOR U726 ( .A(n652), .B(sreg[267]), .Z(n653) );
  XOR U727 ( .A(n654), .B(n653), .Z(c[267]) );
  NANDN U728 ( .A(n652), .B(sreg[267]), .Z(n656) );
  NAND U729 ( .A(n654), .B(n653), .Z(n655) );
  AND U730 ( .A(n656), .B(n655), .Z(n731) );
  NANDN U731 ( .A(n658), .B(n657), .Z(n662) );
  OR U732 ( .A(n660), .B(n659), .Z(n661) );
  AND U733 ( .A(n662), .B(n661), .Z(n696) );
  NANDN U734 ( .A(n664), .B(n663), .Z(n668) );
  NANDN U735 ( .A(n666), .B(n665), .Z(n667) );
  AND U736 ( .A(n668), .B(n667), .Z(n694) );
  NAND U737 ( .A(n26), .B(n669), .Z(n671) );
  XOR U738 ( .A(b[7]), .B(a[14]), .Z(n705) );
  NAND U739 ( .A(n10531), .B(n705), .Z(n670) );
  AND U740 ( .A(n671), .B(n670), .Z(n724) );
  NAND U741 ( .A(n23), .B(n672), .Z(n674) );
  XOR U742 ( .A(b[3]), .B(a[18]), .Z(n708) );
  NAND U743 ( .A(n24), .B(n708), .Z(n673) );
  NAND U744 ( .A(n674), .B(n673), .Z(n723) );
  XNOR U745 ( .A(n724), .B(n723), .Z(n726) );
  NAND U746 ( .A(n25), .B(n675), .Z(n677) );
  XOR U747 ( .A(b[5]), .B(a[16]), .Z(n714) );
  NAND U748 ( .A(n10456), .B(n714), .Z(n676) );
  AND U749 ( .A(n677), .B(n676), .Z(n718) );
  AND U750 ( .A(b[7]), .B(a[12]), .Z(n717) );
  XNOR U751 ( .A(n718), .B(n717), .Z(n719) );
  NAND U752 ( .A(b[0]), .B(a[20]), .Z(n678) );
  XNOR U753 ( .A(b[1]), .B(n678), .Z(n680) );
  NANDN U754 ( .A(b[0]), .B(a[19]), .Z(n679) );
  NAND U755 ( .A(n680), .B(n679), .Z(n720) );
  XNOR U756 ( .A(n719), .B(n720), .Z(n725) );
  XOR U757 ( .A(n726), .B(n725), .Z(n700) );
  NANDN U758 ( .A(n682), .B(n681), .Z(n686) );
  NANDN U759 ( .A(n684), .B(n683), .Z(n685) );
  AND U760 ( .A(n686), .B(n685), .Z(n699) );
  XNOR U761 ( .A(n700), .B(n699), .Z(n701) );
  NANDN U762 ( .A(n688), .B(n687), .Z(n692) );
  NAND U763 ( .A(n690), .B(n689), .Z(n691) );
  NAND U764 ( .A(n692), .B(n691), .Z(n702) );
  XNOR U765 ( .A(n701), .B(n702), .Z(n693) );
  XNOR U766 ( .A(n694), .B(n693), .Z(n695) );
  XNOR U767 ( .A(n696), .B(n695), .Z(n729) );
  XNOR U768 ( .A(sreg[268]), .B(n729), .Z(n730) );
  XNOR U769 ( .A(n731), .B(n730), .Z(c[268]) );
  NANDN U770 ( .A(n694), .B(n693), .Z(n698) );
  NANDN U771 ( .A(n696), .B(n695), .Z(n697) );
  AND U772 ( .A(n698), .B(n697), .Z(n742) );
  NANDN U773 ( .A(n700), .B(n699), .Z(n704) );
  NANDN U774 ( .A(n702), .B(n701), .Z(n703) );
  AND U775 ( .A(n704), .B(n703), .Z(n740) );
  NAND U776 ( .A(n26), .B(n705), .Z(n707) );
  XOR U777 ( .A(b[7]), .B(a[15]), .Z(n751) );
  NAND U778 ( .A(n10531), .B(n751), .Z(n706) );
  AND U779 ( .A(n707), .B(n706), .Z(n770) );
  NAND U780 ( .A(n23), .B(n708), .Z(n710) );
  XOR U781 ( .A(b[3]), .B(a[19]), .Z(n754) );
  NAND U782 ( .A(n24), .B(n754), .Z(n709) );
  NAND U783 ( .A(n710), .B(n709), .Z(n769) );
  XNOR U784 ( .A(n770), .B(n769), .Z(n772) );
  NAND U785 ( .A(b[0]), .B(a[21]), .Z(n711) );
  XNOR U786 ( .A(b[1]), .B(n711), .Z(n713) );
  NANDN U787 ( .A(b[0]), .B(a[20]), .Z(n712) );
  NAND U788 ( .A(n713), .B(n712), .Z(n766) );
  NAND U789 ( .A(n25), .B(n714), .Z(n716) );
  XOR U790 ( .A(b[5]), .B(a[17]), .Z(n760) );
  NAND U791 ( .A(n10456), .B(n760), .Z(n715) );
  AND U792 ( .A(n716), .B(n715), .Z(n764) );
  AND U793 ( .A(b[7]), .B(a[13]), .Z(n763) );
  XNOR U794 ( .A(n764), .B(n763), .Z(n765) );
  XNOR U795 ( .A(n766), .B(n765), .Z(n771) );
  XOR U796 ( .A(n772), .B(n771), .Z(n746) );
  NANDN U797 ( .A(n718), .B(n717), .Z(n722) );
  NANDN U798 ( .A(n720), .B(n719), .Z(n721) );
  AND U799 ( .A(n722), .B(n721), .Z(n745) );
  XNOR U800 ( .A(n746), .B(n745), .Z(n747) );
  NANDN U801 ( .A(n724), .B(n723), .Z(n728) );
  NAND U802 ( .A(n726), .B(n725), .Z(n727) );
  NAND U803 ( .A(n728), .B(n727), .Z(n748) );
  XNOR U804 ( .A(n747), .B(n748), .Z(n739) );
  XNOR U805 ( .A(n740), .B(n739), .Z(n741) );
  XNOR U806 ( .A(n742), .B(n741), .Z(n734) );
  XNOR U807 ( .A(sreg[269]), .B(n734), .Z(n736) );
  NANDN U808 ( .A(sreg[268]), .B(n729), .Z(n733) );
  NAND U809 ( .A(n731), .B(n730), .Z(n732) );
  NAND U810 ( .A(n733), .B(n732), .Z(n735) );
  XNOR U811 ( .A(n736), .B(n735), .Z(c[269]) );
  NANDN U812 ( .A(sreg[269]), .B(n734), .Z(n738) );
  NAND U813 ( .A(n736), .B(n735), .Z(n737) );
  AND U814 ( .A(n738), .B(n737), .Z(n777) );
  NANDN U815 ( .A(n740), .B(n739), .Z(n744) );
  NANDN U816 ( .A(n742), .B(n741), .Z(n743) );
  AND U817 ( .A(n744), .B(n743), .Z(n782) );
  NANDN U818 ( .A(n746), .B(n745), .Z(n750) );
  NANDN U819 ( .A(n748), .B(n747), .Z(n749) );
  AND U820 ( .A(n750), .B(n749), .Z(n781) );
  NAND U821 ( .A(n26), .B(n751), .Z(n753) );
  XOR U822 ( .A(b[7]), .B(a[16]), .Z(n792) );
  NAND U823 ( .A(n10531), .B(n792), .Z(n752) );
  AND U824 ( .A(n753), .B(n752), .Z(n811) );
  NAND U825 ( .A(n23), .B(n754), .Z(n756) );
  XOR U826 ( .A(b[3]), .B(a[20]), .Z(n795) );
  NAND U827 ( .A(n24), .B(n795), .Z(n755) );
  NAND U828 ( .A(n756), .B(n755), .Z(n810) );
  XNOR U829 ( .A(n811), .B(n810), .Z(n813) );
  NAND U830 ( .A(b[0]), .B(a[22]), .Z(n757) );
  XNOR U831 ( .A(b[1]), .B(n757), .Z(n759) );
  NANDN U832 ( .A(b[0]), .B(a[21]), .Z(n758) );
  NAND U833 ( .A(n759), .B(n758), .Z(n807) );
  NAND U834 ( .A(n25), .B(n760), .Z(n762) );
  XOR U835 ( .A(b[5]), .B(a[18]), .Z(n798) );
  NAND U836 ( .A(n10456), .B(n798), .Z(n761) );
  AND U837 ( .A(n762), .B(n761), .Z(n805) );
  AND U838 ( .A(b[7]), .B(a[14]), .Z(n804) );
  XNOR U839 ( .A(n805), .B(n804), .Z(n806) );
  XNOR U840 ( .A(n807), .B(n806), .Z(n812) );
  XOR U841 ( .A(n813), .B(n812), .Z(n787) );
  NANDN U842 ( .A(n764), .B(n763), .Z(n768) );
  NANDN U843 ( .A(n766), .B(n765), .Z(n767) );
  AND U844 ( .A(n768), .B(n767), .Z(n786) );
  XNOR U845 ( .A(n787), .B(n786), .Z(n788) );
  NANDN U846 ( .A(n770), .B(n769), .Z(n774) );
  NAND U847 ( .A(n772), .B(n771), .Z(n773) );
  NAND U848 ( .A(n774), .B(n773), .Z(n789) );
  XNOR U849 ( .A(n788), .B(n789), .Z(n780) );
  XOR U850 ( .A(n781), .B(n780), .Z(n783) );
  XOR U851 ( .A(n782), .B(n783), .Z(n775) );
  XNOR U852 ( .A(n775), .B(sreg[270]), .Z(n776) );
  XOR U853 ( .A(n777), .B(n776), .Z(c[270]) );
  NANDN U854 ( .A(n775), .B(sreg[270]), .Z(n779) );
  NAND U855 ( .A(n777), .B(n776), .Z(n778) );
  AND U856 ( .A(n779), .B(n778), .Z(n854) );
  NANDN U857 ( .A(n781), .B(n780), .Z(n785) );
  OR U858 ( .A(n783), .B(n782), .Z(n784) );
  AND U859 ( .A(n785), .B(n784), .Z(n819) );
  NANDN U860 ( .A(n787), .B(n786), .Z(n791) );
  NANDN U861 ( .A(n789), .B(n788), .Z(n790) );
  AND U862 ( .A(n791), .B(n790), .Z(n817) );
  NAND U863 ( .A(n26), .B(n792), .Z(n794) );
  XOR U864 ( .A(b[7]), .B(a[17]), .Z(n828) );
  NAND U865 ( .A(n10531), .B(n828), .Z(n793) );
  AND U866 ( .A(n794), .B(n793), .Z(n847) );
  NAND U867 ( .A(n23), .B(n795), .Z(n797) );
  XOR U868 ( .A(b[3]), .B(a[21]), .Z(n831) );
  NAND U869 ( .A(n24), .B(n831), .Z(n796) );
  NAND U870 ( .A(n797), .B(n796), .Z(n846) );
  XNOR U871 ( .A(n847), .B(n846), .Z(n849) );
  NAND U872 ( .A(n25), .B(n798), .Z(n800) );
  XOR U873 ( .A(b[5]), .B(a[19]), .Z(n837) );
  NAND U874 ( .A(n10456), .B(n837), .Z(n799) );
  AND U875 ( .A(n800), .B(n799), .Z(n841) );
  AND U876 ( .A(b[7]), .B(a[15]), .Z(n840) );
  XNOR U877 ( .A(n841), .B(n840), .Z(n842) );
  NAND U878 ( .A(b[0]), .B(a[23]), .Z(n801) );
  XNOR U879 ( .A(b[1]), .B(n801), .Z(n803) );
  NANDN U880 ( .A(b[0]), .B(a[22]), .Z(n802) );
  NAND U881 ( .A(n803), .B(n802), .Z(n843) );
  XNOR U882 ( .A(n842), .B(n843), .Z(n848) );
  XOR U883 ( .A(n849), .B(n848), .Z(n823) );
  NANDN U884 ( .A(n805), .B(n804), .Z(n809) );
  NANDN U885 ( .A(n807), .B(n806), .Z(n808) );
  AND U886 ( .A(n809), .B(n808), .Z(n822) );
  XNOR U887 ( .A(n823), .B(n822), .Z(n824) );
  NANDN U888 ( .A(n811), .B(n810), .Z(n815) );
  NAND U889 ( .A(n813), .B(n812), .Z(n814) );
  NAND U890 ( .A(n815), .B(n814), .Z(n825) );
  XNOR U891 ( .A(n824), .B(n825), .Z(n816) );
  XNOR U892 ( .A(n817), .B(n816), .Z(n818) );
  XNOR U893 ( .A(n819), .B(n818), .Z(n852) );
  XNOR U894 ( .A(sreg[271]), .B(n852), .Z(n853) );
  XNOR U895 ( .A(n854), .B(n853), .Z(c[271]) );
  NANDN U896 ( .A(n817), .B(n816), .Z(n821) );
  NANDN U897 ( .A(n819), .B(n818), .Z(n820) );
  AND U898 ( .A(n821), .B(n820), .Z(n865) );
  NANDN U899 ( .A(n823), .B(n822), .Z(n827) );
  NANDN U900 ( .A(n825), .B(n824), .Z(n826) );
  AND U901 ( .A(n827), .B(n826), .Z(n863) );
  NAND U902 ( .A(n26), .B(n828), .Z(n830) );
  XOR U903 ( .A(b[7]), .B(a[18]), .Z(n874) );
  NAND U904 ( .A(n10531), .B(n874), .Z(n829) );
  AND U905 ( .A(n830), .B(n829), .Z(n893) );
  NAND U906 ( .A(n23), .B(n831), .Z(n833) );
  XOR U907 ( .A(b[3]), .B(a[22]), .Z(n877) );
  NAND U908 ( .A(n24), .B(n877), .Z(n832) );
  NAND U909 ( .A(n833), .B(n832), .Z(n892) );
  XNOR U910 ( .A(n893), .B(n892), .Z(n895) );
  NAND U911 ( .A(b[0]), .B(a[24]), .Z(n834) );
  XNOR U912 ( .A(b[1]), .B(n834), .Z(n836) );
  NANDN U913 ( .A(b[0]), .B(a[23]), .Z(n835) );
  NAND U914 ( .A(n836), .B(n835), .Z(n889) );
  NAND U915 ( .A(n25), .B(n837), .Z(n839) );
  XOR U916 ( .A(b[5]), .B(a[20]), .Z(n883) );
  NAND U917 ( .A(n10456), .B(n883), .Z(n838) );
  AND U918 ( .A(n839), .B(n838), .Z(n887) );
  AND U919 ( .A(b[7]), .B(a[16]), .Z(n886) );
  XNOR U920 ( .A(n887), .B(n886), .Z(n888) );
  XNOR U921 ( .A(n889), .B(n888), .Z(n894) );
  XOR U922 ( .A(n895), .B(n894), .Z(n869) );
  NANDN U923 ( .A(n841), .B(n840), .Z(n845) );
  NANDN U924 ( .A(n843), .B(n842), .Z(n844) );
  AND U925 ( .A(n845), .B(n844), .Z(n868) );
  XNOR U926 ( .A(n869), .B(n868), .Z(n870) );
  NANDN U927 ( .A(n847), .B(n846), .Z(n851) );
  NAND U928 ( .A(n849), .B(n848), .Z(n850) );
  NAND U929 ( .A(n851), .B(n850), .Z(n871) );
  XNOR U930 ( .A(n870), .B(n871), .Z(n862) );
  XNOR U931 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U932 ( .A(n865), .B(n864), .Z(n857) );
  XNOR U933 ( .A(sreg[272]), .B(n857), .Z(n859) );
  NANDN U934 ( .A(sreg[271]), .B(n852), .Z(n856) );
  NAND U935 ( .A(n854), .B(n853), .Z(n855) );
  NAND U936 ( .A(n856), .B(n855), .Z(n858) );
  XNOR U937 ( .A(n859), .B(n858), .Z(c[272]) );
  NANDN U938 ( .A(sreg[272]), .B(n857), .Z(n861) );
  NAND U939 ( .A(n859), .B(n858), .Z(n860) );
  AND U940 ( .A(n861), .B(n860), .Z(n900) );
  NANDN U941 ( .A(n863), .B(n862), .Z(n867) );
  NANDN U942 ( .A(n865), .B(n864), .Z(n866) );
  AND U943 ( .A(n867), .B(n866), .Z(n905) );
  NANDN U944 ( .A(n869), .B(n868), .Z(n873) );
  NANDN U945 ( .A(n871), .B(n870), .Z(n872) );
  AND U946 ( .A(n873), .B(n872), .Z(n904) );
  NAND U947 ( .A(n26), .B(n874), .Z(n876) );
  XOR U948 ( .A(b[7]), .B(a[19]), .Z(n915) );
  NAND U949 ( .A(n10531), .B(n915), .Z(n875) );
  AND U950 ( .A(n876), .B(n875), .Z(n934) );
  NAND U951 ( .A(n23), .B(n877), .Z(n879) );
  XOR U952 ( .A(b[3]), .B(a[23]), .Z(n918) );
  NAND U953 ( .A(n24), .B(n918), .Z(n878) );
  NAND U954 ( .A(n879), .B(n878), .Z(n933) );
  XNOR U955 ( .A(n934), .B(n933), .Z(n936) );
  NAND U956 ( .A(b[0]), .B(a[25]), .Z(n880) );
  XNOR U957 ( .A(b[1]), .B(n880), .Z(n882) );
  NANDN U958 ( .A(b[0]), .B(a[24]), .Z(n881) );
  NAND U959 ( .A(n882), .B(n881), .Z(n930) );
  NAND U960 ( .A(n25), .B(n883), .Z(n885) );
  XOR U961 ( .A(b[5]), .B(a[21]), .Z(n924) );
  NAND U962 ( .A(n10456), .B(n924), .Z(n884) );
  AND U963 ( .A(n885), .B(n884), .Z(n928) );
  AND U964 ( .A(b[7]), .B(a[17]), .Z(n927) );
  XNOR U965 ( .A(n928), .B(n927), .Z(n929) );
  XNOR U966 ( .A(n930), .B(n929), .Z(n935) );
  XOR U967 ( .A(n936), .B(n935), .Z(n910) );
  NANDN U968 ( .A(n887), .B(n886), .Z(n891) );
  NANDN U969 ( .A(n889), .B(n888), .Z(n890) );
  AND U970 ( .A(n891), .B(n890), .Z(n909) );
  XNOR U971 ( .A(n910), .B(n909), .Z(n911) );
  NANDN U972 ( .A(n893), .B(n892), .Z(n897) );
  NAND U973 ( .A(n895), .B(n894), .Z(n896) );
  NAND U974 ( .A(n897), .B(n896), .Z(n912) );
  XNOR U975 ( .A(n911), .B(n912), .Z(n903) );
  XOR U976 ( .A(n904), .B(n903), .Z(n906) );
  XOR U977 ( .A(n905), .B(n906), .Z(n898) );
  XNOR U978 ( .A(n898), .B(sreg[273]), .Z(n899) );
  XOR U979 ( .A(n900), .B(n899), .Z(c[273]) );
  NANDN U980 ( .A(n898), .B(sreg[273]), .Z(n902) );
  NAND U981 ( .A(n900), .B(n899), .Z(n901) );
  AND U982 ( .A(n902), .B(n901), .Z(n977) );
  NANDN U983 ( .A(n904), .B(n903), .Z(n908) );
  OR U984 ( .A(n906), .B(n905), .Z(n907) );
  AND U985 ( .A(n908), .B(n907), .Z(n942) );
  NANDN U986 ( .A(n910), .B(n909), .Z(n914) );
  NANDN U987 ( .A(n912), .B(n911), .Z(n913) );
  AND U988 ( .A(n914), .B(n913), .Z(n940) );
  NAND U989 ( .A(n26), .B(n915), .Z(n917) );
  XOR U990 ( .A(b[7]), .B(a[20]), .Z(n951) );
  NAND U991 ( .A(n10531), .B(n951), .Z(n916) );
  AND U992 ( .A(n917), .B(n916), .Z(n970) );
  NAND U993 ( .A(n23), .B(n918), .Z(n920) );
  XOR U994 ( .A(b[3]), .B(a[24]), .Z(n954) );
  NAND U995 ( .A(n24), .B(n954), .Z(n919) );
  NAND U996 ( .A(n920), .B(n919), .Z(n969) );
  XNOR U997 ( .A(n970), .B(n969), .Z(n972) );
  NAND U998 ( .A(b[0]), .B(a[26]), .Z(n921) );
  XNOR U999 ( .A(b[1]), .B(n921), .Z(n923) );
  NANDN U1000 ( .A(b[0]), .B(a[25]), .Z(n922) );
  NAND U1001 ( .A(n923), .B(n922), .Z(n966) );
  NAND U1002 ( .A(n25), .B(n924), .Z(n926) );
  XOR U1003 ( .A(b[5]), .B(a[22]), .Z(n960) );
  NAND U1004 ( .A(n10456), .B(n960), .Z(n925) );
  AND U1005 ( .A(n926), .B(n925), .Z(n964) );
  AND U1006 ( .A(b[7]), .B(a[18]), .Z(n963) );
  XNOR U1007 ( .A(n964), .B(n963), .Z(n965) );
  XNOR U1008 ( .A(n966), .B(n965), .Z(n971) );
  XOR U1009 ( .A(n972), .B(n971), .Z(n946) );
  NANDN U1010 ( .A(n928), .B(n927), .Z(n932) );
  NANDN U1011 ( .A(n930), .B(n929), .Z(n931) );
  AND U1012 ( .A(n932), .B(n931), .Z(n945) );
  XNOR U1013 ( .A(n946), .B(n945), .Z(n947) );
  NANDN U1014 ( .A(n934), .B(n933), .Z(n938) );
  NAND U1015 ( .A(n936), .B(n935), .Z(n937) );
  NAND U1016 ( .A(n938), .B(n937), .Z(n948) );
  XNOR U1017 ( .A(n947), .B(n948), .Z(n939) );
  XNOR U1018 ( .A(n940), .B(n939), .Z(n941) );
  XNOR U1019 ( .A(n942), .B(n941), .Z(n975) );
  XNOR U1020 ( .A(sreg[274]), .B(n975), .Z(n976) );
  XNOR U1021 ( .A(n977), .B(n976), .Z(c[274]) );
  NANDN U1022 ( .A(n940), .B(n939), .Z(n944) );
  NANDN U1023 ( .A(n942), .B(n941), .Z(n943) );
  AND U1024 ( .A(n944), .B(n943), .Z(n988) );
  NANDN U1025 ( .A(n946), .B(n945), .Z(n950) );
  NANDN U1026 ( .A(n948), .B(n947), .Z(n949) );
  AND U1027 ( .A(n950), .B(n949), .Z(n986) );
  NAND U1028 ( .A(n26), .B(n951), .Z(n953) );
  XOR U1029 ( .A(b[7]), .B(a[21]), .Z(n997) );
  NAND U1030 ( .A(n10531), .B(n997), .Z(n952) );
  AND U1031 ( .A(n953), .B(n952), .Z(n1016) );
  NAND U1032 ( .A(n23), .B(n954), .Z(n956) );
  XOR U1033 ( .A(b[3]), .B(a[25]), .Z(n1000) );
  NAND U1034 ( .A(n24), .B(n1000), .Z(n955) );
  NAND U1035 ( .A(n956), .B(n955), .Z(n1015) );
  XNOR U1036 ( .A(n1016), .B(n1015), .Z(n1018) );
  NAND U1037 ( .A(b[0]), .B(a[27]), .Z(n957) );
  XNOR U1038 ( .A(b[1]), .B(n957), .Z(n959) );
  NANDN U1039 ( .A(b[0]), .B(a[26]), .Z(n958) );
  NAND U1040 ( .A(n959), .B(n958), .Z(n1012) );
  NAND U1041 ( .A(n25), .B(n960), .Z(n962) );
  XOR U1042 ( .A(b[5]), .B(a[23]), .Z(n1006) );
  NAND U1043 ( .A(n10456), .B(n1006), .Z(n961) );
  AND U1044 ( .A(n962), .B(n961), .Z(n1010) );
  AND U1045 ( .A(b[7]), .B(a[19]), .Z(n1009) );
  XNOR U1046 ( .A(n1010), .B(n1009), .Z(n1011) );
  XNOR U1047 ( .A(n1012), .B(n1011), .Z(n1017) );
  XOR U1048 ( .A(n1018), .B(n1017), .Z(n992) );
  NANDN U1049 ( .A(n964), .B(n963), .Z(n968) );
  NANDN U1050 ( .A(n966), .B(n965), .Z(n967) );
  AND U1051 ( .A(n968), .B(n967), .Z(n991) );
  XNOR U1052 ( .A(n992), .B(n991), .Z(n993) );
  NANDN U1053 ( .A(n970), .B(n969), .Z(n974) );
  NAND U1054 ( .A(n972), .B(n971), .Z(n973) );
  NAND U1055 ( .A(n974), .B(n973), .Z(n994) );
  XNOR U1056 ( .A(n993), .B(n994), .Z(n985) );
  XNOR U1057 ( .A(n986), .B(n985), .Z(n987) );
  XNOR U1058 ( .A(n988), .B(n987), .Z(n980) );
  XNOR U1059 ( .A(sreg[275]), .B(n980), .Z(n982) );
  NANDN U1060 ( .A(sreg[274]), .B(n975), .Z(n979) );
  NAND U1061 ( .A(n977), .B(n976), .Z(n978) );
  NAND U1062 ( .A(n979), .B(n978), .Z(n981) );
  XNOR U1063 ( .A(n982), .B(n981), .Z(c[275]) );
  NANDN U1064 ( .A(sreg[275]), .B(n980), .Z(n984) );
  NAND U1065 ( .A(n982), .B(n981), .Z(n983) );
  AND U1066 ( .A(n984), .B(n983), .Z(n1023) );
  NANDN U1067 ( .A(n986), .B(n985), .Z(n990) );
  NANDN U1068 ( .A(n988), .B(n987), .Z(n989) );
  AND U1069 ( .A(n990), .B(n989), .Z(n1028) );
  NANDN U1070 ( .A(n992), .B(n991), .Z(n996) );
  NANDN U1071 ( .A(n994), .B(n993), .Z(n995) );
  AND U1072 ( .A(n996), .B(n995), .Z(n1027) );
  NAND U1073 ( .A(n26), .B(n997), .Z(n999) );
  XOR U1074 ( .A(b[7]), .B(a[22]), .Z(n1038) );
  NAND U1075 ( .A(n10531), .B(n1038), .Z(n998) );
  AND U1076 ( .A(n999), .B(n998), .Z(n1057) );
  NAND U1077 ( .A(n23), .B(n1000), .Z(n1002) );
  XOR U1078 ( .A(b[3]), .B(a[26]), .Z(n1041) );
  NAND U1079 ( .A(n24), .B(n1041), .Z(n1001) );
  NAND U1080 ( .A(n1002), .B(n1001), .Z(n1056) );
  XNOR U1081 ( .A(n1057), .B(n1056), .Z(n1059) );
  NAND U1082 ( .A(b[0]), .B(a[28]), .Z(n1003) );
  XNOR U1083 ( .A(b[1]), .B(n1003), .Z(n1005) );
  NANDN U1084 ( .A(b[0]), .B(a[27]), .Z(n1004) );
  NAND U1085 ( .A(n1005), .B(n1004), .Z(n1053) );
  NAND U1086 ( .A(n25), .B(n1006), .Z(n1008) );
  XOR U1087 ( .A(b[5]), .B(a[24]), .Z(n1047) );
  NAND U1088 ( .A(n10456), .B(n1047), .Z(n1007) );
  AND U1089 ( .A(n1008), .B(n1007), .Z(n1051) );
  AND U1090 ( .A(b[7]), .B(a[20]), .Z(n1050) );
  XNOR U1091 ( .A(n1051), .B(n1050), .Z(n1052) );
  XNOR U1092 ( .A(n1053), .B(n1052), .Z(n1058) );
  XOR U1093 ( .A(n1059), .B(n1058), .Z(n1033) );
  NANDN U1094 ( .A(n1010), .B(n1009), .Z(n1014) );
  NANDN U1095 ( .A(n1012), .B(n1011), .Z(n1013) );
  AND U1096 ( .A(n1014), .B(n1013), .Z(n1032) );
  XNOR U1097 ( .A(n1033), .B(n1032), .Z(n1034) );
  NANDN U1098 ( .A(n1016), .B(n1015), .Z(n1020) );
  NAND U1099 ( .A(n1018), .B(n1017), .Z(n1019) );
  NAND U1100 ( .A(n1020), .B(n1019), .Z(n1035) );
  XNOR U1101 ( .A(n1034), .B(n1035), .Z(n1026) );
  XOR U1102 ( .A(n1027), .B(n1026), .Z(n1029) );
  XOR U1103 ( .A(n1028), .B(n1029), .Z(n1021) );
  XNOR U1104 ( .A(n1021), .B(sreg[276]), .Z(n1022) );
  XOR U1105 ( .A(n1023), .B(n1022), .Z(c[276]) );
  NANDN U1106 ( .A(n1021), .B(sreg[276]), .Z(n1025) );
  NAND U1107 ( .A(n1023), .B(n1022), .Z(n1024) );
  AND U1108 ( .A(n1025), .B(n1024), .Z(n1100) );
  NANDN U1109 ( .A(n1027), .B(n1026), .Z(n1031) );
  OR U1110 ( .A(n1029), .B(n1028), .Z(n1030) );
  AND U1111 ( .A(n1031), .B(n1030), .Z(n1065) );
  NANDN U1112 ( .A(n1033), .B(n1032), .Z(n1037) );
  NANDN U1113 ( .A(n1035), .B(n1034), .Z(n1036) );
  AND U1114 ( .A(n1037), .B(n1036), .Z(n1063) );
  NAND U1115 ( .A(n26), .B(n1038), .Z(n1040) );
  XOR U1116 ( .A(b[7]), .B(a[23]), .Z(n1074) );
  NAND U1117 ( .A(n10531), .B(n1074), .Z(n1039) );
  AND U1118 ( .A(n1040), .B(n1039), .Z(n1093) );
  NAND U1119 ( .A(n23), .B(n1041), .Z(n1043) );
  XOR U1120 ( .A(b[3]), .B(a[27]), .Z(n1077) );
  NAND U1121 ( .A(n24), .B(n1077), .Z(n1042) );
  NAND U1122 ( .A(n1043), .B(n1042), .Z(n1092) );
  XNOR U1123 ( .A(n1093), .B(n1092), .Z(n1095) );
  NAND U1124 ( .A(b[0]), .B(a[29]), .Z(n1044) );
  XNOR U1125 ( .A(b[1]), .B(n1044), .Z(n1046) );
  NANDN U1126 ( .A(b[0]), .B(a[28]), .Z(n1045) );
  NAND U1127 ( .A(n1046), .B(n1045), .Z(n1089) );
  NAND U1128 ( .A(n25), .B(n1047), .Z(n1049) );
  XOR U1129 ( .A(b[5]), .B(a[25]), .Z(n1083) );
  NAND U1130 ( .A(n10456), .B(n1083), .Z(n1048) );
  AND U1131 ( .A(n1049), .B(n1048), .Z(n1087) );
  AND U1132 ( .A(b[7]), .B(a[21]), .Z(n1086) );
  XNOR U1133 ( .A(n1087), .B(n1086), .Z(n1088) );
  XNOR U1134 ( .A(n1089), .B(n1088), .Z(n1094) );
  XOR U1135 ( .A(n1095), .B(n1094), .Z(n1069) );
  NANDN U1136 ( .A(n1051), .B(n1050), .Z(n1055) );
  NANDN U1137 ( .A(n1053), .B(n1052), .Z(n1054) );
  AND U1138 ( .A(n1055), .B(n1054), .Z(n1068) );
  XNOR U1139 ( .A(n1069), .B(n1068), .Z(n1070) );
  NANDN U1140 ( .A(n1057), .B(n1056), .Z(n1061) );
  NAND U1141 ( .A(n1059), .B(n1058), .Z(n1060) );
  NAND U1142 ( .A(n1061), .B(n1060), .Z(n1071) );
  XNOR U1143 ( .A(n1070), .B(n1071), .Z(n1062) );
  XNOR U1144 ( .A(n1063), .B(n1062), .Z(n1064) );
  XNOR U1145 ( .A(n1065), .B(n1064), .Z(n1098) );
  XNOR U1146 ( .A(sreg[277]), .B(n1098), .Z(n1099) );
  XNOR U1147 ( .A(n1100), .B(n1099), .Z(c[277]) );
  NANDN U1148 ( .A(n1063), .B(n1062), .Z(n1067) );
  NANDN U1149 ( .A(n1065), .B(n1064), .Z(n1066) );
  AND U1150 ( .A(n1067), .B(n1066), .Z(n1111) );
  NANDN U1151 ( .A(n1069), .B(n1068), .Z(n1073) );
  NANDN U1152 ( .A(n1071), .B(n1070), .Z(n1072) );
  AND U1153 ( .A(n1073), .B(n1072), .Z(n1109) );
  NAND U1154 ( .A(n26), .B(n1074), .Z(n1076) );
  XOR U1155 ( .A(b[7]), .B(a[24]), .Z(n1120) );
  NAND U1156 ( .A(n10531), .B(n1120), .Z(n1075) );
  AND U1157 ( .A(n1076), .B(n1075), .Z(n1139) );
  NAND U1158 ( .A(n23), .B(n1077), .Z(n1079) );
  XOR U1159 ( .A(b[3]), .B(a[28]), .Z(n1123) );
  NAND U1160 ( .A(n24), .B(n1123), .Z(n1078) );
  NAND U1161 ( .A(n1079), .B(n1078), .Z(n1138) );
  XNOR U1162 ( .A(n1139), .B(n1138), .Z(n1141) );
  NAND U1163 ( .A(b[0]), .B(a[30]), .Z(n1080) );
  XNOR U1164 ( .A(b[1]), .B(n1080), .Z(n1082) );
  NANDN U1165 ( .A(b[0]), .B(a[29]), .Z(n1081) );
  NAND U1166 ( .A(n1082), .B(n1081), .Z(n1135) );
  NAND U1167 ( .A(n25), .B(n1083), .Z(n1085) );
  XOR U1168 ( .A(b[5]), .B(a[26]), .Z(n1129) );
  NAND U1169 ( .A(n10456), .B(n1129), .Z(n1084) );
  AND U1170 ( .A(n1085), .B(n1084), .Z(n1133) );
  AND U1171 ( .A(b[7]), .B(a[22]), .Z(n1132) );
  XNOR U1172 ( .A(n1133), .B(n1132), .Z(n1134) );
  XNOR U1173 ( .A(n1135), .B(n1134), .Z(n1140) );
  XOR U1174 ( .A(n1141), .B(n1140), .Z(n1115) );
  NANDN U1175 ( .A(n1087), .B(n1086), .Z(n1091) );
  NANDN U1176 ( .A(n1089), .B(n1088), .Z(n1090) );
  AND U1177 ( .A(n1091), .B(n1090), .Z(n1114) );
  XNOR U1178 ( .A(n1115), .B(n1114), .Z(n1116) );
  NANDN U1179 ( .A(n1093), .B(n1092), .Z(n1097) );
  NAND U1180 ( .A(n1095), .B(n1094), .Z(n1096) );
  NAND U1181 ( .A(n1097), .B(n1096), .Z(n1117) );
  XNOR U1182 ( .A(n1116), .B(n1117), .Z(n1108) );
  XNOR U1183 ( .A(n1109), .B(n1108), .Z(n1110) );
  XNOR U1184 ( .A(n1111), .B(n1110), .Z(n1103) );
  XNOR U1185 ( .A(sreg[278]), .B(n1103), .Z(n1105) );
  NANDN U1186 ( .A(sreg[277]), .B(n1098), .Z(n1102) );
  NAND U1187 ( .A(n1100), .B(n1099), .Z(n1101) );
  NAND U1188 ( .A(n1102), .B(n1101), .Z(n1104) );
  XNOR U1189 ( .A(n1105), .B(n1104), .Z(c[278]) );
  NANDN U1190 ( .A(sreg[278]), .B(n1103), .Z(n1107) );
  NAND U1191 ( .A(n1105), .B(n1104), .Z(n1106) );
  AND U1192 ( .A(n1107), .B(n1106), .Z(n1146) );
  NANDN U1193 ( .A(n1109), .B(n1108), .Z(n1113) );
  NANDN U1194 ( .A(n1111), .B(n1110), .Z(n1112) );
  AND U1195 ( .A(n1113), .B(n1112), .Z(n1151) );
  NANDN U1196 ( .A(n1115), .B(n1114), .Z(n1119) );
  NANDN U1197 ( .A(n1117), .B(n1116), .Z(n1118) );
  AND U1198 ( .A(n1119), .B(n1118), .Z(n1150) );
  NAND U1199 ( .A(n26), .B(n1120), .Z(n1122) );
  XOR U1200 ( .A(b[7]), .B(a[25]), .Z(n1161) );
  NAND U1201 ( .A(n10531), .B(n1161), .Z(n1121) );
  AND U1202 ( .A(n1122), .B(n1121), .Z(n1180) );
  NAND U1203 ( .A(n23), .B(n1123), .Z(n1125) );
  XOR U1204 ( .A(b[3]), .B(a[29]), .Z(n1164) );
  NAND U1205 ( .A(n24), .B(n1164), .Z(n1124) );
  NAND U1206 ( .A(n1125), .B(n1124), .Z(n1179) );
  XNOR U1207 ( .A(n1180), .B(n1179), .Z(n1182) );
  NAND U1208 ( .A(b[0]), .B(a[31]), .Z(n1126) );
  XNOR U1209 ( .A(b[1]), .B(n1126), .Z(n1128) );
  NANDN U1210 ( .A(b[0]), .B(a[30]), .Z(n1127) );
  NAND U1211 ( .A(n1128), .B(n1127), .Z(n1176) );
  NAND U1212 ( .A(n25), .B(n1129), .Z(n1131) );
  XOR U1213 ( .A(b[5]), .B(a[27]), .Z(n1170) );
  NAND U1214 ( .A(n10456), .B(n1170), .Z(n1130) );
  AND U1215 ( .A(n1131), .B(n1130), .Z(n1174) );
  AND U1216 ( .A(b[7]), .B(a[23]), .Z(n1173) );
  XNOR U1217 ( .A(n1174), .B(n1173), .Z(n1175) );
  XNOR U1218 ( .A(n1176), .B(n1175), .Z(n1181) );
  XOR U1219 ( .A(n1182), .B(n1181), .Z(n1156) );
  NANDN U1220 ( .A(n1133), .B(n1132), .Z(n1137) );
  NANDN U1221 ( .A(n1135), .B(n1134), .Z(n1136) );
  AND U1222 ( .A(n1137), .B(n1136), .Z(n1155) );
  XNOR U1223 ( .A(n1156), .B(n1155), .Z(n1157) );
  NANDN U1224 ( .A(n1139), .B(n1138), .Z(n1143) );
  NAND U1225 ( .A(n1141), .B(n1140), .Z(n1142) );
  NAND U1226 ( .A(n1143), .B(n1142), .Z(n1158) );
  XNOR U1227 ( .A(n1157), .B(n1158), .Z(n1149) );
  XOR U1228 ( .A(n1150), .B(n1149), .Z(n1152) );
  XOR U1229 ( .A(n1151), .B(n1152), .Z(n1144) );
  XNOR U1230 ( .A(n1144), .B(sreg[279]), .Z(n1145) );
  XOR U1231 ( .A(n1146), .B(n1145), .Z(c[279]) );
  NANDN U1232 ( .A(n1144), .B(sreg[279]), .Z(n1148) );
  NAND U1233 ( .A(n1146), .B(n1145), .Z(n1147) );
  AND U1234 ( .A(n1148), .B(n1147), .Z(n1223) );
  NANDN U1235 ( .A(n1150), .B(n1149), .Z(n1154) );
  OR U1236 ( .A(n1152), .B(n1151), .Z(n1153) );
  AND U1237 ( .A(n1154), .B(n1153), .Z(n1188) );
  NANDN U1238 ( .A(n1156), .B(n1155), .Z(n1160) );
  NANDN U1239 ( .A(n1158), .B(n1157), .Z(n1159) );
  AND U1240 ( .A(n1160), .B(n1159), .Z(n1186) );
  NAND U1241 ( .A(n26), .B(n1161), .Z(n1163) );
  XOR U1242 ( .A(b[7]), .B(a[26]), .Z(n1197) );
  NAND U1243 ( .A(n10531), .B(n1197), .Z(n1162) );
  AND U1244 ( .A(n1163), .B(n1162), .Z(n1216) );
  NAND U1245 ( .A(n23), .B(n1164), .Z(n1166) );
  XOR U1246 ( .A(b[3]), .B(a[30]), .Z(n1200) );
  NAND U1247 ( .A(n24), .B(n1200), .Z(n1165) );
  NAND U1248 ( .A(n1166), .B(n1165), .Z(n1215) );
  XNOR U1249 ( .A(n1216), .B(n1215), .Z(n1218) );
  NAND U1250 ( .A(b[0]), .B(a[32]), .Z(n1167) );
  XNOR U1251 ( .A(b[1]), .B(n1167), .Z(n1169) );
  NANDN U1252 ( .A(b[0]), .B(a[31]), .Z(n1168) );
  NAND U1253 ( .A(n1169), .B(n1168), .Z(n1212) );
  NAND U1254 ( .A(n25), .B(n1170), .Z(n1172) );
  XOR U1255 ( .A(b[5]), .B(a[28]), .Z(n1206) );
  NAND U1256 ( .A(n10456), .B(n1206), .Z(n1171) );
  AND U1257 ( .A(n1172), .B(n1171), .Z(n1210) );
  AND U1258 ( .A(b[7]), .B(a[24]), .Z(n1209) );
  XNOR U1259 ( .A(n1210), .B(n1209), .Z(n1211) );
  XNOR U1260 ( .A(n1212), .B(n1211), .Z(n1217) );
  XOR U1261 ( .A(n1218), .B(n1217), .Z(n1192) );
  NANDN U1262 ( .A(n1174), .B(n1173), .Z(n1178) );
  NANDN U1263 ( .A(n1176), .B(n1175), .Z(n1177) );
  AND U1264 ( .A(n1178), .B(n1177), .Z(n1191) );
  XNOR U1265 ( .A(n1192), .B(n1191), .Z(n1193) );
  NANDN U1266 ( .A(n1180), .B(n1179), .Z(n1184) );
  NAND U1267 ( .A(n1182), .B(n1181), .Z(n1183) );
  NAND U1268 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U1269 ( .A(n1193), .B(n1194), .Z(n1185) );
  XNOR U1270 ( .A(n1186), .B(n1185), .Z(n1187) );
  XNOR U1271 ( .A(n1188), .B(n1187), .Z(n1221) );
  XNOR U1272 ( .A(sreg[280]), .B(n1221), .Z(n1222) );
  XNOR U1273 ( .A(n1223), .B(n1222), .Z(c[280]) );
  NANDN U1274 ( .A(n1186), .B(n1185), .Z(n1190) );
  NANDN U1275 ( .A(n1188), .B(n1187), .Z(n1189) );
  AND U1276 ( .A(n1190), .B(n1189), .Z(n1234) );
  NANDN U1277 ( .A(n1192), .B(n1191), .Z(n1196) );
  NANDN U1278 ( .A(n1194), .B(n1193), .Z(n1195) );
  AND U1279 ( .A(n1196), .B(n1195), .Z(n1232) );
  NAND U1280 ( .A(n26), .B(n1197), .Z(n1199) );
  XOR U1281 ( .A(b[7]), .B(a[27]), .Z(n1243) );
  NAND U1282 ( .A(n10531), .B(n1243), .Z(n1198) );
  AND U1283 ( .A(n1199), .B(n1198), .Z(n1262) );
  NAND U1284 ( .A(n23), .B(n1200), .Z(n1202) );
  XOR U1285 ( .A(b[3]), .B(a[31]), .Z(n1246) );
  NAND U1286 ( .A(n24), .B(n1246), .Z(n1201) );
  NAND U1287 ( .A(n1202), .B(n1201), .Z(n1261) );
  XNOR U1288 ( .A(n1262), .B(n1261), .Z(n1264) );
  NAND U1289 ( .A(b[0]), .B(a[33]), .Z(n1203) );
  XNOR U1290 ( .A(b[1]), .B(n1203), .Z(n1205) );
  NANDN U1291 ( .A(b[0]), .B(a[32]), .Z(n1204) );
  NAND U1292 ( .A(n1205), .B(n1204), .Z(n1258) );
  NAND U1293 ( .A(n25), .B(n1206), .Z(n1208) );
  XOR U1294 ( .A(b[5]), .B(a[29]), .Z(n1252) );
  NAND U1295 ( .A(n10456), .B(n1252), .Z(n1207) );
  AND U1296 ( .A(n1208), .B(n1207), .Z(n1256) );
  AND U1297 ( .A(b[7]), .B(a[25]), .Z(n1255) );
  XNOR U1298 ( .A(n1256), .B(n1255), .Z(n1257) );
  XNOR U1299 ( .A(n1258), .B(n1257), .Z(n1263) );
  XOR U1300 ( .A(n1264), .B(n1263), .Z(n1238) );
  NANDN U1301 ( .A(n1210), .B(n1209), .Z(n1214) );
  NANDN U1302 ( .A(n1212), .B(n1211), .Z(n1213) );
  AND U1303 ( .A(n1214), .B(n1213), .Z(n1237) );
  XNOR U1304 ( .A(n1238), .B(n1237), .Z(n1239) );
  NANDN U1305 ( .A(n1216), .B(n1215), .Z(n1220) );
  NAND U1306 ( .A(n1218), .B(n1217), .Z(n1219) );
  NAND U1307 ( .A(n1220), .B(n1219), .Z(n1240) );
  XNOR U1308 ( .A(n1239), .B(n1240), .Z(n1231) );
  XNOR U1309 ( .A(n1232), .B(n1231), .Z(n1233) );
  XNOR U1310 ( .A(n1234), .B(n1233), .Z(n1226) );
  XNOR U1311 ( .A(sreg[281]), .B(n1226), .Z(n1228) );
  NANDN U1312 ( .A(sreg[280]), .B(n1221), .Z(n1225) );
  NAND U1313 ( .A(n1223), .B(n1222), .Z(n1224) );
  NAND U1314 ( .A(n1225), .B(n1224), .Z(n1227) );
  XNOR U1315 ( .A(n1228), .B(n1227), .Z(c[281]) );
  NANDN U1316 ( .A(sreg[281]), .B(n1226), .Z(n1230) );
  NAND U1317 ( .A(n1228), .B(n1227), .Z(n1229) );
  AND U1318 ( .A(n1230), .B(n1229), .Z(n1269) );
  NANDN U1319 ( .A(n1232), .B(n1231), .Z(n1236) );
  NANDN U1320 ( .A(n1234), .B(n1233), .Z(n1235) );
  AND U1321 ( .A(n1236), .B(n1235), .Z(n1274) );
  NANDN U1322 ( .A(n1238), .B(n1237), .Z(n1242) );
  NANDN U1323 ( .A(n1240), .B(n1239), .Z(n1241) );
  AND U1324 ( .A(n1242), .B(n1241), .Z(n1273) );
  NAND U1325 ( .A(n26), .B(n1243), .Z(n1245) );
  XOR U1326 ( .A(b[7]), .B(a[28]), .Z(n1284) );
  NAND U1327 ( .A(n10531), .B(n1284), .Z(n1244) );
  AND U1328 ( .A(n1245), .B(n1244), .Z(n1303) );
  NAND U1329 ( .A(n23), .B(n1246), .Z(n1248) );
  XOR U1330 ( .A(b[3]), .B(a[32]), .Z(n1287) );
  NAND U1331 ( .A(n24), .B(n1287), .Z(n1247) );
  NAND U1332 ( .A(n1248), .B(n1247), .Z(n1302) );
  XNOR U1333 ( .A(n1303), .B(n1302), .Z(n1305) );
  NAND U1334 ( .A(b[0]), .B(a[34]), .Z(n1249) );
  XNOR U1335 ( .A(b[1]), .B(n1249), .Z(n1251) );
  NANDN U1336 ( .A(b[0]), .B(a[33]), .Z(n1250) );
  NAND U1337 ( .A(n1251), .B(n1250), .Z(n1299) );
  NAND U1338 ( .A(n25), .B(n1252), .Z(n1254) );
  XOR U1339 ( .A(b[5]), .B(a[30]), .Z(n1293) );
  NAND U1340 ( .A(n10456), .B(n1293), .Z(n1253) );
  AND U1341 ( .A(n1254), .B(n1253), .Z(n1297) );
  AND U1342 ( .A(b[7]), .B(a[26]), .Z(n1296) );
  XNOR U1343 ( .A(n1297), .B(n1296), .Z(n1298) );
  XNOR U1344 ( .A(n1299), .B(n1298), .Z(n1304) );
  XOR U1345 ( .A(n1305), .B(n1304), .Z(n1279) );
  NANDN U1346 ( .A(n1256), .B(n1255), .Z(n1260) );
  NANDN U1347 ( .A(n1258), .B(n1257), .Z(n1259) );
  AND U1348 ( .A(n1260), .B(n1259), .Z(n1278) );
  XNOR U1349 ( .A(n1279), .B(n1278), .Z(n1280) );
  NANDN U1350 ( .A(n1262), .B(n1261), .Z(n1266) );
  NAND U1351 ( .A(n1264), .B(n1263), .Z(n1265) );
  NAND U1352 ( .A(n1266), .B(n1265), .Z(n1281) );
  XNOR U1353 ( .A(n1280), .B(n1281), .Z(n1272) );
  XOR U1354 ( .A(n1273), .B(n1272), .Z(n1275) );
  XOR U1355 ( .A(n1274), .B(n1275), .Z(n1267) );
  XNOR U1356 ( .A(n1267), .B(sreg[282]), .Z(n1268) );
  XOR U1357 ( .A(n1269), .B(n1268), .Z(c[282]) );
  NANDN U1358 ( .A(n1267), .B(sreg[282]), .Z(n1271) );
  NAND U1359 ( .A(n1269), .B(n1268), .Z(n1270) );
  AND U1360 ( .A(n1271), .B(n1270), .Z(n1346) );
  NANDN U1361 ( .A(n1273), .B(n1272), .Z(n1277) );
  OR U1362 ( .A(n1275), .B(n1274), .Z(n1276) );
  AND U1363 ( .A(n1277), .B(n1276), .Z(n1311) );
  NANDN U1364 ( .A(n1279), .B(n1278), .Z(n1283) );
  NANDN U1365 ( .A(n1281), .B(n1280), .Z(n1282) );
  AND U1366 ( .A(n1283), .B(n1282), .Z(n1309) );
  NAND U1367 ( .A(n26), .B(n1284), .Z(n1286) );
  XOR U1368 ( .A(b[7]), .B(a[29]), .Z(n1320) );
  NAND U1369 ( .A(n10531), .B(n1320), .Z(n1285) );
  AND U1370 ( .A(n1286), .B(n1285), .Z(n1339) );
  NAND U1371 ( .A(n23), .B(n1287), .Z(n1289) );
  XOR U1372 ( .A(b[3]), .B(a[33]), .Z(n1323) );
  NAND U1373 ( .A(n24), .B(n1323), .Z(n1288) );
  NAND U1374 ( .A(n1289), .B(n1288), .Z(n1338) );
  XNOR U1375 ( .A(n1339), .B(n1338), .Z(n1341) );
  NAND U1376 ( .A(b[0]), .B(a[35]), .Z(n1290) );
  XNOR U1377 ( .A(b[1]), .B(n1290), .Z(n1292) );
  NANDN U1378 ( .A(b[0]), .B(a[34]), .Z(n1291) );
  NAND U1379 ( .A(n1292), .B(n1291), .Z(n1335) );
  NAND U1380 ( .A(n25), .B(n1293), .Z(n1295) );
  XOR U1381 ( .A(b[5]), .B(a[31]), .Z(n1329) );
  NAND U1382 ( .A(n10456), .B(n1329), .Z(n1294) );
  AND U1383 ( .A(n1295), .B(n1294), .Z(n1333) );
  AND U1384 ( .A(b[7]), .B(a[27]), .Z(n1332) );
  XNOR U1385 ( .A(n1333), .B(n1332), .Z(n1334) );
  XNOR U1386 ( .A(n1335), .B(n1334), .Z(n1340) );
  XOR U1387 ( .A(n1341), .B(n1340), .Z(n1315) );
  NANDN U1388 ( .A(n1297), .B(n1296), .Z(n1301) );
  NANDN U1389 ( .A(n1299), .B(n1298), .Z(n1300) );
  AND U1390 ( .A(n1301), .B(n1300), .Z(n1314) );
  XNOR U1391 ( .A(n1315), .B(n1314), .Z(n1316) );
  NANDN U1392 ( .A(n1303), .B(n1302), .Z(n1307) );
  NAND U1393 ( .A(n1305), .B(n1304), .Z(n1306) );
  NAND U1394 ( .A(n1307), .B(n1306), .Z(n1317) );
  XNOR U1395 ( .A(n1316), .B(n1317), .Z(n1308) );
  XNOR U1396 ( .A(n1309), .B(n1308), .Z(n1310) );
  XNOR U1397 ( .A(n1311), .B(n1310), .Z(n1344) );
  XNOR U1398 ( .A(sreg[283]), .B(n1344), .Z(n1345) );
  XNOR U1399 ( .A(n1346), .B(n1345), .Z(c[283]) );
  NANDN U1400 ( .A(n1309), .B(n1308), .Z(n1313) );
  NANDN U1401 ( .A(n1311), .B(n1310), .Z(n1312) );
  AND U1402 ( .A(n1313), .B(n1312), .Z(n1352) );
  NANDN U1403 ( .A(n1315), .B(n1314), .Z(n1319) );
  NANDN U1404 ( .A(n1317), .B(n1316), .Z(n1318) );
  AND U1405 ( .A(n1319), .B(n1318), .Z(n1350) );
  NAND U1406 ( .A(n26), .B(n1320), .Z(n1322) );
  XOR U1407 ( .A(b[7]), .B(a[30]), .Z(n1361) );
  NAND U1408 ( .A(n10531), .B(n1361), .Z(n1321) );
  AND U1409 ( .A(n1322), .B(n1321), .Z(n1380) );
  NAND U1410 ( .A(n23), .B(n1323), .Z(n1325) );
  XOR U1411 ( .A(b[3]), .B(a[34]), .Z(n1364) );
  NAND U1412 ( .A(n24), .B(n1364), .Z(n1324) );
  NAND U1413 ( .A(n1325), .B(n1324), .Z(n1379) );
  XNOR U1414 ( .A(n1380), .B(n1379), .Z(n1382) );
  NAND U1415 ( .A(b[0]), .B(a[36]), .Z(n1326) );
  XNOR U1416 ( .A(b[1]), .B(n1326), .Z(n1328) );
  NANDN U1417 ( .A(b[0]), .B(a[35]), .Z(n1327) );
  NAND U1418 ( .A(n1328), .B(n1327), .Z(n1376) );
  NAND U1419 ( .A(n25), .B(n1329), .Z(n1331) );
  XOR U1420 ( .A(b[5]), .B(a[32]), .Z(n1370) );
  NAND U1421 ( .A(n10456), .B(n1370), .Z(n1330) );
  AND U1422 ( .A(n1331), .B(n1330), .Z(n1374) );
  AND U1423 ( .A(b[7]), .B(a[28]), .Z(n1373) );
  XNOR U1424 ( .A(n1374), .B(n1373), .Z(n1375) );
  XNOR U1425 ( .A(n1376), .B(n1375), .Z(n1381) );
  XOR U1426 ( .A(n1382), .B(n1381), .Z(n1356) );
  NANDN U1427 ( .A(n1333), .B(n1332), .Z(n1337) );
  NANDN U1428 ( .A(n1335), .B(n1334), .Z(n1336) );
  AND U1429 ( .A(n1337), .B(n1336), .Z(n1355) );
  XNOR U1430 ( .A(n1356), .B(n1355), .Z(n1357) );
  NANDN U1431 ( .A(n1339), .B(n1338), .Z(n1343) );
  NAND U1432 ( .A(n1341), .B(n1340), .Z(n1342) );
  NAND U1433 ( .A(n1343), .B(n1342), .Z(n1358) );
  XNOR U1434 ( .A(n1357), .B(n1358), .Z(n1349) );
  XNOR U1435 ( .A(n1350), .B(n1349), .Z(n1351) );
  XNOR U1436 ( .A(n1352), .B(n1351), .Z(n1385) );
  XNOR U1437 ( .A(sreg[284]), .B(n1385), .Z(n1387) );
  NANDN U1438 ( .A(sreg[283]), .B(n1344), .Z(n1348) );
  NAND U1439 ( .A(n1346), .B(n1345), .Z(n1347) );
  NAND U1440 ( .A(n1348), .B(n1347), .Z(n1386) );
  XNOR U1441 ( .A(n1387), .B(n1386), .Z(c[284]) );
  NANDN U1442 ( .A(n1350), .B(n1349), .Z(n1354) );
  NANDN U1443 ( .A(n1352), .B(n1351), .Z(n1353) );
  AND U1444 ( .A(n1354), .B(n1353), .Z(n1393) );
  NANDN U1445 ( .A(n1356), .B(n1355), .Z(n1360) );
  NANDN U1446 ( .A(n1358), .B(n1357), .Z(n1359) );
  AND U1447 ( .A(n1360), .B(n1359), .Z(n1391) );
  NAND U1448 ( .A(n26), .B(n1361), .Z(n1363) );
  XOR U1449 ( .A(b[7]), .B(a[31]), .Z(n1402) );
  NAND U1450 ( .A(n10531), .B(n1402), .Z(n1362) );
  AND U1451 ( .A(n1363), .B(n1362), .Z(n1421) );
  NAND U1452 ( .A(n23), .B(n1364), .Z(n1366) );
  XOR U1453 ( .A(b[3]), .B(a[35]), .Z(n1405) );
  NAND U1454 ( .A(n24), .B(n1405), .Z(n1365) );
  NAND U1455 ( .A(n1366), .B(n1365), .Z(n1420) );
  XNOR U1456 ( .A(n1421), .B(n1420), .Z(n1423) );
  NAND U1457 ( .A(b[0]), .B(a[37]), .Z(n1367) );
  XNOR U1458 ( .A(b[1]), .B(n1367), .Z(n1369) );
  NANDN U1459 ( .A(b[0]), .B(a[36]), .Z(n1368) );
  NAND U1460 ( .A(n1369), .B(n1368), .Z(n1417) );
  NAND U1461 ( .A(n25), .B(n1370), .Z(n1372) );
  XOR U1462 ( .A(b[5]), .B(a[33]), .Z(n1411) );
  NAND U1463 ( .A(n10456), .B(n1411), .Z(n1371) );
  AND U1464 ( .A(n1372), .B(n1371), .Z(n1415) );
  AND U1465 ( .A(b[7]), .B(a[29]), .Z(n1414) );
  XNOR U1466 ( .A(n1415), .B(n1414), .Z(n1416) );
  XNOR U1467 ( .A(n1417), .B(n1416), .Z(n1422) );
  XOR U1468 ( .A(n1423), .B(n1422), .Z(n1397) );
  NANDN U1469 ( .A(n1374), .B(n1373), .Z(n1378) );
  NANDN U1470 ( .A(n1376), .B(n1375), .Z(n1377) );
  AND U1471 ( .A(n1378), .B(n1377), .Z(n1396) );
  XNOR U1472 ( .A(n1397), .B(n1396), .Z(n1398) );
  NANDN U1473 ( .A(n1380), .B(n1379), .Z(n1384) );
  NAND U1474 ( .A(n1382), .B(n1381), .Z(n1383) );
  NAND U1475 ( .A(n1384), .B(n1383), .Z(n1399) );
  XNOR U1476 ( .A(n1398), .B(n1399), .Z(n1390) );
  XNOR U1477 ( .A(n1391), .B(n1390), .Z(n1392) );
  XNOR U1478 ( .A(n1393), .B(n1392), .Z(n1426) );
  XNOR U1479 ( .A(sreg[285]), .B(n1426), .Z(n1428) );
  NANDN U1480 ( .A(sreg[284]), .B(n1385), .Z(n1389) );
  NAND U1481 ( .A(n1387), .B(n1386), .Z(n1388) );
  NAND U1482 ( .A(n1389), .B(n1388), .Z(n1427) );
  XNOR U1483 ( .A(n1428), .B(n1427), .Z(c[285]) );
  NANDN U1484 ( .A(n1391), .B(n1390), .Z(n1395) );
  NANDN U1485 ( .A(n1393), .B(n1392), .Z(n1394) );
  AND U1486 ( .A(n1395), .B(n1394), .Z(n1434) );
  NANDN U1487 ( .A(n1397), .B(n1396), .Z(n1401) );
  NANDN U1488 ( .A(n1399), .B(n1398), .Z(n1400) );
  AND U1489 ( .A(n1401), .B(n1400), .Z(n1432) );
  NAND U1490 ( .A(n26), .B(n1402), .Z(n1404) );
  XOR U1491 ( .A(b[7]), .B(a[32]), .Z(n1443) );
  NAND U1492 ( .A(n10531), .B(n1443), .Z(n1403) );
  AND U1493 ( .A(n1404), .B(n1403), .Z(n1462) );
  NAND U1494 ( .A(n23), .B(n1405), .Z(n1407) );
  XOR U1495 ( .A(b[3]), .B(a[36]), .Z(n1446) );
  NAND U1496 ( .A(n24), .B(n1446), .Z(n1406) );
  NAND U1497 ( .A(n1407), .B(n1406), .Z(n1461) );
  XNOR U1498 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U1499 ( .A(b[0]), .B(a[38]), .Z(n1408) );
  XNOR U1500 ( .A(b[1]), .B(n1408), .Z(n1410) );
  NANDN U1501 ( .A(b[0]), .B(a[37]), .Z(n1409) );
  NAND U1502 ( .A(n1410), .B(n1409), .Z(n1458) );
  NAND U1503 ( .A(n25), .B(n1411), .Z(n1413) );
  XOR U1504 ( .A(b[5]), .B(a[34]), .Z(n1452) );
  NAND U1505 ( .A(n10456), .B(n1452), .Z(n1412) );
  AND U1506 ( .A(n1413), .B(n1412), .Z(n1456) );
  AND U1507 ( .A(b[7]), .B(a[30]), .Z(n1455) );
  XNOR U1508 ( .A(n1456), .B(n1455), .Z(n1457) );
  XNOR U1509 ( .A(n1458), .B(n1457), .Z(n1463) );
  XOR U1510 ( .A(n1464), .B(n1463), .Z(n1438) );
  NANDN U1511 ( .A(n1415), .B(n1414), .Z(n1419) );
  NANDN U1512 ( .A(n1417), .B(n1416), .Z(n1418) );
  AND U1513 ( .A(n1419), .B(n1418), .Z(n1437) );
  XNOR U1514 ( .A(n1438), .B(n1437), .Z(n1439) );
  NANDN U1515 ( .A(n1421), .B(n1420), .Z(n1425) );
  NAND U1516 ( .A(n1423), .B(n1422), .Z(n1424) );
  NAND U1517 ( .A(n1425), .B(n1424), .Z(n1440) );
  XNOR U1518 ( .A(n1439), .B(n1440), .Z(n1431) );
  XNOR U1519 ( .A(n1432), .B(n1431), .Z(n1433) );
  XNOR U1520 ( .A(n1434), .B(n1433), .Z(n1467) );
  XNOR U1521 ( .A(sreg[286]), .B(n1467), .Z(n1469) );
  NANDN U1522 ( .A(sreg[285]), .B(n1426), .Z(n1430) );
  NAND U1523 ( .A(n1428), .B(n1427), .Z(n1429) );
  NAND U1524 ( .A(n1430), .B(n1429), .Z(n1468) );
  XNOR U1525 ( .A(n1469), .B(n1468), .Z(c[286]) );
  NANDN U1526 ( .A(n1432), .B(n1431), .Z(n1436) );
  NANDN U1527 ( .A(n1434), .B(n1433), .Z(n1435) );
  AND U1528 ( .A(n1436), .B(n1435), .Z(n1475) );
  NANDN U1529 ( .A(n1438), .B(n1437), .Z(n1442) );
  NANDN U1530 ( .A(n1440), .B(n1439), .Z(n1441) );
  AND U1531 ( .A(n1442), .B(n1441), .Z(n1473) );
  NAND U1532 ( .A(n26), .B(n1443), .Z(n1445) );
  XOR U1533 ( .A(b[7]), .B(a[33]), .Z(n1484) );
  NAND U1534 ( .A(n10531), .B(n1484), .Z(n1444) );
  AND U1535 ( .A(n1445), .B(n1444), .Z(n1503) );
  NAND U1536 ( .A(n23), .B(n1446), .Z(n1448) );
  XOR U1537 ( .A(b[3]), .B(a[37]), .Z(n1487) );
  NAND U1538 ( .A(n24), .B(n1487), .Z(n1447) );
  NAND U1539 ( .A(n1448), .B(n1447), .Z(n1502) );
  XNOR U1540 ( .A(n1503), .B(n1502), .Z(n1505) );
  NAND U1541 ( .A(b[0]), .B(a[39]), .Z(n1449) );
  XNOR U1542 ( .A(b[1]), .B(n1449), .Z(n1451) );
  NANDN U1543 ( .A(b[0]), .B(a[38]), .Z(n1450) );
  NAND U1544 ( .A(n1451), .B(n1450), .Z(n1499) );
  NAND U1545 ( .A(n25), .B(n1452), .Z(n1454) );
  XOR U1546 ( .A(b[5]), .B(a[35]), .Z(n1493) );
  NAND U1547 ( .A(n10456), .B(n1493), .Z(n1453) );
  AND U1548 ( .A(n1454), .B(n1453), .Z(n1497) );
  AND U1549 ( .A(b[7]), .B(a[31]), .Z(n1496) );
  XNOR U1550 ( .A(n1497), .B(n1496), .Z(n1498) );
  XNOR U1551 ( .A(n1499), .B(n1498), .Z(n1504) );
  XOR U1552 ( .A(n1505), .B(n1504), .Z(n1479) );
  NANDN U1553 ( .A(n1456), .B(n1455), .Z(n1460) );
  NANDN U1554 ( .A(n1458), .B(n1457), .Z(n1459) );
  AND U1555 ( .A(n1460), .B(n1459), .Z(n1478) );
  XNOR U1556 ( .A(n1479), .B(n1478), .Z(n1480) );
  NANDN U1557 ( .A(n1462), .B(n1461), .Z(n1466) );
  NAND U1558 ( .A(n1464), .B(n1463), .Z(n1465) );
  NAND U1559 ( .A(n1466), .B(n1465), .Z(n1481) );
  XNOR U1560 ( .A(n1480), .B(n1481), .Z(n1472) );
  XNOR U1561 ( .A(n1473), .B(n1472), .Z(n1474) );
  XNOR U1562 ( .A(n1475), .B(n1474), .Z(n1508) );
  XNOR U1563 ( .A(sreg[287]), .B(n1508), .Z(n1510) );
  NANDN U1564 ( .A(sreg[286]), .B(n1467), .Z(n1471) );
  NAND U1565 ( .A(n1469), .B(n1468), .Z(n1470) );
  NAND U1566 ( .A(n1471), .B(n1470), .Z(n1509) );
  XNOR U1567 ( .A(n1510), .B(n1509), .Z(c[287]) );
  NANDN U1568 ( .A(n1473), .B(n1472), .Z(n1477) );
  NANDN U1569 ( .A(n1475), .B(n1474), .Z(n1476) );
  AND U1570 ( .A(n1477), .B(n1476), .Z(n1516) );
  NANDN U1571 ( .A(n1479), .B(n1478), .Z(n1483) );
  NANDN U1572 ( .A(n1481), .B(n1480), .Z(n1482) );
  AND U1573 ( .A(n1483), .B(n1482), .Z(n1514) );
  NAND U1574 ( .A(n26), .B(n1484), .Z(n1486) );
  XOR U1575 ( .A(b[7]), .B(a[34]), .Z(n1525) );
  NAND U1576 ( .A(n10531), .B(n1525), .Z(n1485) );
  AND U1577 ( .A(n1486), .B(n1485), .Z(n1544) );
  NAND U1578 ( .A(n23), .B(n1487), .Z(n1489) );
  XOR U1579 ( .A(b[3]), .B(a[38]), .Z(n1528) );
  NAND U1580 ( .A(n24), .B(n1528), .Z(n1488) );
  NAND U1581 ( .A(n1489), .B(n1488), .Z(n1543) );
  XNOR U1582 ( .A(n1544), .B(n1543), .Z(n1546) );
  NAND U1583 ( .A(b[0]), .B(a[40]), .Z(n1490) );
  XNOR U1584 ( .A(b[1]), .B(n1490), .Z(n1492) );
  NANDN U1585 ( .A(b[0]), .B(a[39]), .Z(n1491) );
  NAND U1586 ( .A(n1492), .B(n1491), .Z(n1540) );
  NAND U1587 ( .A(n25), .B(n1493), .Z(n1495) );
  XOR U1588 ( .A(b[5]), .B(a[36]), .Z(n1531) );
  NAND U1589 ( .A(n10456), .B(n1531), .Z(n1494) );
  AND U1590 ( .A(n1495), .B(n1494), .Z(n1538) );
  AND U1591 ( .A(b[7]), .B(a[32]), .Z(n1537) );
  XNOR U1592 ( .A(n1538), .B(n1537), .Z(n1539) );
  XNOR U1593 ( .A(n1540), .B(n1539), .Z(n1545) );
  XOR U1594 ( .A(n1546), .B(n1545), .Z(n1520) );
  NANDN U1595 ( .A(n1497), .B(n1496), .Z(n1501) );
  NANDN U1596 ( .A(n1499), .B(n1498), .Z(n1500) );
  AND U1597 ( .A(n1501), .B(n1500), .Z(n1519) );
  XNOR U1598 ( .A(n1520), .B(n1519), .Z(n1521) );
  NANDN U1599 ( .A(n1503), .B(n1502), .Z(n1507) );
  NAND U1600 ( .A(n1505), .B(n1504), .Z(n1506) );
  NAND U1601 ( .A(n1507), .B(n1506), .Z(n1522) );
  XNOR U1602 ( .A(n1521), .B(n1522), .Z(n1513) );
  XNOR U1603 ( .A(n1514), .B(n1513), .Z(n1515) );
  XNOR U1604 ( .A(n1516), .B(n1515), .Z(n1549) );
  XNOR U1605 ( .A(sreg[288]), .B(n1549), .Z(n1551) );
  NANDN U1606 ( .A(sreg[287]), .B(n1508), .Z(n1512) );
  NAND U1607 ( .A(n1510), .B(n1509), .Z(n1511) );
  NAND U1608 ( .A(n1512), .B(n1511), .Z(n1550) );
  XNOR U1609 ( .A(n1551), .B(n1550), .Z(c[288]) );
  NANDN U1610 ( .A(n1514), .B(n1513), .Z(n1518) );
  NANDN U1611 ( .A(n1516), .B(n1515), .Z(n1517) );
  AND U1612 ( .A(n1518), .B(n1517), .Z(n1557) );
  NANDN U1613 ( .A(n1520), .B(n1519), .Z(n1524) );
  NANDN U1614 ( .A(n1522), .B(n1521), .Z(n1523) );
  AND U1615 ( .A(n1524), .B(n1523), .Z(n1555) );
  NAND U1616 ( .A(n26), .B(n1525), .Z(n1527) );
  XOR U1617 ( .A(b[7]), .B(a[35]), .Z(n1566) );
  NAND U1618 ( .A(n10531), .B(n1566), .Z(n1526) );
  AND U1619 ( .A(n1527), .B(n1526), .Z(n1585) );
  NAND U1620 ( .A(n23), .B(n1528), .Z(n1530) );
  XOR U1621 ( .A(b[3]), .B(a[39]), .Z(n1569) );
  NAND U1622 ( .A(n24), .B(n1569), .Z(n1529) );
  NAND U1623 ( .A(n1530), .B(n1529), .Z(n1584) );
  XNOR U1624 ( .A(n1585), .B(n1584), .Z(n1587) );
  NAND U1625 ( .A(n25), .B(n1531), .Z(n1533) );
  XOR U1626 ( .A(b[5]), .B(a[37]), .Z(n1575) );
  NAND U1627 ( .A(n10456), .B(n1575), .Z(n1532) );
  AND U1628 ( .A(n1533), .B(n1532), .Z(n1579) );
  AND U1629 ( .A(b[7]), .B(a[33]), .Z(n1578) );
  XNOR U1630 ( .A(n1579), .B(n1578), .Z(n1580) );
  NAND U1631 ( .A(b[0]), .B(a[41]), .Z(n1534) );
  XNOR U1632 ( .A(b[1]), .B(n1534), .Z(n1536) );
  NANDN U1633 ( .A(b[0]), .B(a[40]), .Z(n1535) );
  NAND U1634 ( .A(n1536), .B(n1535), .Z(n1581) );
  XNOR U1635 ( .A(n1580), .B(n1581), .Z(n1586) );
  XOR U1636 ( .A(n1587), .B(n1586), .Z(n1561) );
  NANDN U1637 ( .A(n1538), .B(n1537), .Z(n1542) );
  NANDN U1638 ( .A(n1540), .B(n1539), .Z(n1541) );
  AND U1639 ( .A(n1542), .B(n1541), .Z(n1560) );
  XNOR U1640 ( .A(n1561), .B(n1560), .Z(n1562) );
  NANDN U1641 ( .A(n1544), .B(n1543), .Z(n1548) );
  NAND U1642 ( .A(n1546), .B(n1545), .Z(n1547) );
  NAND U1643 ( .A(n1548), .B(n1547), .Z(n1563) );
  XNOR U1644 ( .A(n1562), .B(n1563), .Z(n1554) );
  XNOR U1645 ( .A(n1555), .B(n1554), .Z(n1556) );
  XNOR U1646 ( .A(n1557), .B(n1556), .Z(n1590) );
  XNOR U1647 ( .A(sreg[289]), .B(n1590), .Z(n1592) );
  NANDN U1648 ( .A(sreg[288]), .B(n1549), .Z(n1553) );
  NAND U1649 ( .A(n1551), .B(n1550), .Z(n1552) );
  NAND U1650 ( .A(n1553), .B(n1552), .Z(n1591) );
  XNOR U1651 ( .A(n1592), .B(n1591), .Z(c[289]) );
  NANDN U1652 ( .A(n1555), .B(n1554), .Z(n1559) );
  NANDN U1653 ( .A(n1557), .B(n1556), .Z(n1558) );
  AND U1654 ( .A(n1559), .B(n1558), .Z(n1598) );
  NANDN U1655 ( .A(n1561), .B(n1560), .Z(n1565) );
  NANDN U1656 ( .A(n1563), .B(n1562), .Z(n1564) );
  AND U1657 ( .A(n1565), .B(n1564), .Z(n1596) );
  NAND U1658 ( .A(n26), .B(n1566), .Z(n1568) );
  XOR U1659 ( .A(b[7]), .B(a[36]), .Z(n1607) );
  NAND U1660 ( .A(n10531), .B(n1607), .Z(n1567) );
  AND U1661 ( .A(n1568), .B(n1567), .Z(n1626) );
  NAND U1662 ( .A(n23), .B(n1569), .Z(n1571) );
  XOR U1663 ( .A(b[3]), .B(a[40]), .Z(n1610) );
  NAND U1664 ( .A(n24), .B(n1610), .Z(n1570) );
  NAND U1665 ( .A(n1571), .B(n1570), .Z(n1625) );
  XNOR U1666 ( .A(n1626), .B(n1625), .Z(n1628) );
  NAND U1667 ( .A(b[0]), .B(a[42]), .Z(n1572) );
  XNOR U1668 ( .A(b[1]), .B(n1572), .Z(n1574) );
  NANDN U1669 ( .A(b[0]), .B(a[41]), .Z(n1573) );
  NAND U1670 ( .A(n1574), .B(n1573), .Z(n1622) );
  NAND U1671 ( .A(n25), .B(n1575), .Z(n1577) );
  XOR U1672 ( .A(b[5]), .B(a[38]), .Z(n1613) );
  NAND U1673 ( .A(n10456), .B(n1613), .Z(n1576) );
  AND U1674 ( .A(n1577), .B(n1576), .Z(n1620) );
  AND U1675 ( .A(b[7]), .B(a[34]), .Z(n1619) );
  XNOR U1676 ( .A(n1620), .B(n1619), .Z(n1621) );
  XNOR U1677 ( .A(n1622), .B(n1621), .Z(n1627) );
  XOR U1678 ( .A(n1628), .B(n1627), .Z(n1602) );
  NANDN U1679 ( .A(n1579), .B(n1578), .Z(n1583) );
  NANDN U1680 ( .A(n1581), .B(n1580), .Z(n1582) );
  AND U1681 ( .A(n1583), .B(n1582), .Z(n1601) );
  XNOR U1682 ( .A(n1602), .B(n1601), .Z(n1603) );
  NANDN U1683 ( .A(n1585), .B(n1584), .Z(n1589) );
  NAND U1684 ( .A(n1587), .B(n1586), .Z(n1588) );
  NAND U1685 ( .A(n1589), .B(n1588), .Z(n1604) );
  XNOR U1686 ( .A(n1603), .B(n1604), .Z(n1595) );
  XNOR U1687 ( .A(n1596), .B(n1595), .Z(n1597) );
  XNOR U1688 ( .A(n1598), .B(n1597), .Z(n1631) );
  XNOR U1689 ( .A(sreg[290]), .B(n1631), .Z(n1633) );
  NANDN U1690 ( .A(sreg[289]), .B(n1590), .Z(n1594) );
  NAND U1691 ( .A(n1592), .B(n1591), .Z(n1593) );
  NAND U1692 ( .A(n1594), .B(n1593), .Z(n1632) );
  XNOR U1693 ( .A(n1633), .B(n1632), .Z(c[290]) );
  NANDN U1694 ( .A(n1596), .B(n1595), .Z(n1600) );
  NANDN U1695 ( .A(n1598), .B(n1597), .Z(n1599) );
  AND U1696 ( .A(n1600), .B(n1599), .Z(n1639) );
  NANDN U1697 ( .A(n1602), .B(n1601), .Z(n1606) );
  NANDN U1698 ( .A(n1604), .B(n1603), .Z(n1605) );
  AND U1699 ( .A(n1606), .B(n1605), .Z(n1637) );
  NAND U1700 ( .A(n26), .B(n1607), .Z(n1609) );
  XOR U1701 ( .A(b[7]), .B(a[37]), .Z(n1648) );
  NAND U1702 ( .A(n10531), .B(n1648), .Z(n1608) );
  AND U1703 ( .A(n1609), .B(n1608), .Z(n1667) );
  NAND U1704 ( .A(n23), .B(n1610), .Z(n1612) );
  XOR U1705 ( .A(b[3]), .B(a[41]), .Z(n1651) );
  NAND U1706 ( .A(n24), .B(n1651), .Z(n1611) );
  NAND U1707 ( .A(n1612), .B(n1611), .Z(n1666) );
  XNOR U1708 ( .A(n1667), .B(n1666), .Z(n1669) );
  NAND U1709 ( .A(n25), .B(n1613), .Z(n1615) );
  XOR U1710 ( .A(b[5]), .B(a[39]), .Z(n1657) );
  NAND U1711 ( .A(n10456), .B(n1657), .Z(n1614) );
  AND U1712 ( .A(n1615), .B(n1614), .Z(n1661) );
  AND U1713 ( .A(b[7]), .B(a[35]), .Z(n1660) );
  XNOR U1714 ( .A(n1661), .B(n1660), .Z(n1662) );
  NAND U1715 ( .A(b[0]), .B(a[43]), .Z(n1616) );
  XNOR U1716 ( .A(b[1]), .B(n1616), .Z(n1618) );
  NANDN U1717 ( .A(b[0]), .B(a[42]), .Z(n1617) );
  NAND U1718 ( .A(n1618), .B(n1617), .Z(n1663) );
  XNOR U1719 ( .A(n1662), .B(n1663), .Z(n1668) );
  XOR U1720 ( .A(n1669), .B(n1668), .Z(n1643) );
  NANDN U1721 ( .A(n1620), .B(n1619), .Z(n1624) );
  NANDN U1722 ( .A(n1622), .B(n1621), .Z(n1623) );
  AND U1723 ( .A(n1624), .B(n1623), .Z(n1642) );
  XNOR U1724 ( .A(n1643), .B(n1642), .Z(n1644) );
  NANDN U1725 ( .A(n1626), .B(n1625), .Z(n1630) );
  NAND U1726 ( .A(n1628), .B(n1627), .Z(n1629) );
  NAND U1727 ( .A(n1630), .B(n1629), .Z(n1645) );
  XNOR U1728 ( .A(n1644), .B(n1645), .Z(n1636) );
  XNOR U1729 ( .A(n1637), .B(n1636), .Z(n1638) );
  XNOR U1730 ( .A(n1639), .B(n1638), .Z(n1672) );
  XNOR U1731 ( .A(sreg[291]), .B(n1672), .Z(n1674) );
  NANDN U1732 ( .A(sreg[290]), .B(n1631), .Z(n1635) );
  NAND U1733 ( .A(n1633), .B(n1632), .Z(n1634) );
  NAND U1734 ( .A(n1635), .B(n1634), .Z(n1673) );
  XNOR U1735 ( .A(n1674), .B(n1673), .Z(c[291]) );
  NANDN U1736 ( .A(n1637), .B(n1636), .Z(n1641) );
  NANDN U1737 ( .A(n1639), .B(n1638), .Z(n1640) );
  AND U1738 ( .A(n1641), .B(n1640), .Z(n1680) );
  NANDN U1739 ( .A(n1643), .B(n1642), .Z(n1647) );
  NANDN U1740 ( .A(n1645), .B(n1644), .Z(n1646) );
  AND U1741 ( .A(n1647), .B(n1646), .Z(n1678) );
  NAND U1742 ( .A(n26), .B(n1648), .Z(n1650) );
  XOR U1743 ( .A(b[7]), .B(a[38]), .Z(n1689) );
  NAND U1744 ( .A(n10531), .B(n1689), .Z(n1649) );
  AND U1745 ( .A(n1650), .B(n1649), .Z(n1708) );
  NAND U1746 ( .A(n23), .B(n1651), .Z(n1653) );
  XOR U1747 ( .A(b[3]), .B(a[42]), .Z(n1692) );
  NAND U1748 ( .A(n24), .B(n1692), .Z(n1652) );
  NAND U1749 ( .A(n1653), .B(n1652), .Z(n1707) );
  XNOR U1750 ( .A(n1708), .B(n1707), .Z(n1710) );
  NAND U1751 ( .A(b[0]), .B(a[44]), .Z(n1654) );
  XNOR U1752 ( .A(b[1]), .B(n1654), .Z(n1656) );
  NANDN U1753 ( .A(b[0]), .B(a[43]), .Z(n1655) );
  NAND U1754 ( .A(n1656), .B(n1655), .Z(n1704) );
  NAND U1755 ( .A(n25), .B(n1657), .Z(n1659) );
  XOR U1756 ( .A(b[5]), .B(a[40]), .Z(n1698) );
  NAND U1757 ( .A(n10456), .B(n1698), .Z(n1658) );
  AND U1758 ( .A(n1659), .B(n1658), .Z(n1702) );
  AND U1759 ( .A(b[7]), .B(a[36]), .Z(n1701) );
  XNOR U1760 ( .A(n1702), .B(n1701), .Z(n1703) );
  XNOR U1761 ( .A(n1704), .B(n1703), .Z(n1709) );
  XOR U1762 ( .A(n1710), .B(n1709), .Z(n1684) );
  NANDN U1763 ( .A(n1661), .B(n1660), .Z(n1665) );
  NANDN U1764 ( .A(n1663), .B(n1662), .Z(n1664) );
  AND U1765 ( .A(n1665), .B(n1664), .Z(n1683) );
  XNOR U1766 ( .A(n1684), .B(n1683), .Z(n1685) );
  NANDN U1767 ( .A(n1667), .B(n1666), .Z(n1671) );
  NAND U1768 ( .A(n1669), .B(n1668), .Z(n1670) );
  NAND U1769 ( .A(n1671), .B(n1670), .Z(n1686) );
  XNOR U1770 ( .A(n1685), .B(n1686), .Z(n1677) );
  XNOR U1771 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U1772 ( .A(n1680), .B(n1679), .Z(n1713) );
  XNOR U1773 ( .A(sreg[292]), .B(n1713), .Z(n1715) );
  NANDN U1774 ( .A(sreg[291]), .B(n1672), .Z(n1676) );
  NAND U1775 ( .A(n1674), .B(n1673), .Z(n1675) );
  NAND U1776 ( .A(n1676), .B(n1675), .Z(n1714) );
  XNOR U1777 ( .A(n1715), .B(n1714), .Z(c[292]) );
  NANDN U1778 ( .A(n1678), .B(n1677), .Z(n1682) );
  NANDN U1779 ( .A(n1680), .B(n1679), .Z(n1681) );
  AND U1780 ( .A(n1682), .B(n1681), .Z(n1721) );
  NANDN U1781 ( .A(n1684), .B(n1683), .Z(n1688) );
  NANDN U1782 ( .A(n1686), .B(n1685), .Z(n1687) );
  AND U1783 ( .A(n1688), .B(n1687), .Z(n1719) );
  NAND U1784 ( .A(n26), .B(n1689), .Z(n1691) );
  XOR U1785 ( .A(b[7]), .B(a[39]), .Z(n1730) );
  NAND U1786 ( .A(n10531), .B(n1730), .Z(n1690) );
  AND U1787 ( .A(n1691), .B(n1690), .Z(n1749) );
  NAND U1788 ( .A(n23), .B(n1692), .Z(n1694) );
  XOR U1789 ( .A(b[3]), .B(a[43]), .Z(n1733) );
  NAND U1790 ( .A(n24), .B(n1733), .Z(n1693) );
  NAND U1791 ( .A(n1694), .B(n1693), .Z(n1748) );
  XNOR U1792 ( .A(n1749), .B(n1748), .Z(n1751) );
  NAND U1793 ( .A(b[0]), .B(a[45]), .Z(n1695) );
  XNOR U1794 ( .A(b[1]), .B(n1695), .Z(n1697) );
  NANDN U1795 ( .A(b[0]), .B(a[44]), .Z(n1696) );
  NAND U1796 ( .A(n1697), .B(n1696), .Z(n1745) );
  NAND U1797 ( .A(n25), .B(n1698), .Z(n1700) );
  XOR U1798 ( .A(b[5]), .B(a[41]), .Z(n1739) );
  NAND U1799 ( .A(n10456), .B(n1739), .Z(n1699) );
  AND U1800 ( .A(n1700), .B(n1699), .Z(n1743) );
  AND U1801 ( .A(b[7]), .B(a[37]), .Z(n1742) );
  XNOR U1802 ( .A(n1743), .B(n1742), .Z(n1744) );
  XNOR U1803 ( .A(n1745), .B(n1744), .Z(n1750) );
  XOR U1804 ( .A(n1751), .B(n1750), .Z(n1725) );
  NANDN U1805 ( .A(n1702), .B(n1701), .Z(n1706) );
  NANDN U1806 ( .A(n1704), .B(n1703), .Z(n1705) );
  AND U1807 ( .A(n1706), .B(n1705), .Z(n1724) );
  XNOR U1808 ( .A(n1725), .B(n1724), .Z(n1726) );
  NANDN U1809 ( .A(n1708), .B(n1707), .Z(n1712) );
  NAND U1810 ( .A(n1710), .B(n1709), .Z(n1711) );
  NAND U1811 ( .A(n1712), .B(n1711), .Z(n1727) );
  XNOR U1812 ( .A(n1726), .B(n1727), .Z(n1718) );
  XNOR U1813 ( .A(n1719), .B(n1718), .Z(n1720) );
  XNOR U1814 ( .A(n1721), .B(n1720), .Z(n1754) );
  XNOR U1815 ( .A(sreg[293]), .B(n1754), .Z(n1756) );
  NANDN U1816 ( .A(sreg[292]), .B(n1713), .Z(n1717) );
  NAND U1817 ( .A(n1715), .B(n1714), .Z(n1716) );
  NAND U1818 ( .A(n1717), .B(n1716), .Z(n1755) );
  XNOR U1819 ( .A(n1756), .B(n1755), .Z(c[293]) );
  NANDN U1820 ( .A(n1719), .B(n1718), .Z(n1723) );
  NANDN U1821 ( .A(n1721), .B(n1720), .Z(n1722) );
  AND U1822 ( .A(n1723), .B(n1722), .Z(n1762) );
  NANDN U1823 ( .A(n1725), .B(n1724), .Z(n1729) );
  NANDN U1824 ( .A(n1727), .B(n1726), .Z(n1728) );
  AND U1825 ( .A(n1729), .B(n1728), .Z(n1760) );
  NAND U1826 ( .A(n26), .B(n1730), .Z(n1732) );
  XOR U1827 ( .A(b[7]), .B(a[40]), .Z(n1771) );
  NAND U1828 ( .A(n10531), .B(n1771), .Z(n1731) );
  AND U1829 ( .A(n1732), .B(n1731), .Z(n1790) );
  NAND U1830 ( .A(n23), .B(n1733), .Z(n1735) );
  XOR U1831 ( .A(b[3]), .B(a[44]), .Z(n1774) );
  NAND U1832 ( .A(n24), .B(n1774), .Z(n1734) );
  NAND U1833 ( .A(n1735), .B(n1734), .Z(n1789) );
  XNOR U1834 ( .A(n1790), .B(n1789), .Z(n1792) );
  NAND U1835 ( .A(b[0]), .B(a[46]), .Z(n1736) );
  XNOR U1836 ( .A(b[1]), .B(n1736), .Z(n1738) );
  NANDN U1837 ( .A(b[0]), .B(a[45]), .Z(n1737) );
  NAND U1838 ( .A(n1738), .B(n1737), .Z(n1786) );
  NAND U1839 ( .A(n25), .B(n1739), .Z(n1741) );
  XOR U1840 ( .A(b[5]), .B(a[42]), .Z(n1780) );
  NAND U1841 ( .A(n10456), .B(n1780), .Z(n1740) );
  AND U1842 ( .A(n1741), .B(n1740), .Z(n1784) );
  AND U1843 ( .A(b[7]), .B(a[38]), .Z(n1783) );
  XNOR U1844 ( .A(n1784), .B(n1783), .Z(n1785) );
  XNOR U1845 ( .A(n1786), .B(n1785), .Z(n1791) );
  XOR U1846 ( .A(n1792), .B(n1791), .Z(n1766) );
  NANDN U1847 ( .A(n1743), .B(n1742), .Z(n1747) );
  NANDN U1848 ( .A(n1745), .B(n1744), .Z(n1746) );
  AND U1849 ( .A(n1747), .B(n1746), .Z(n1765) );
  XNOR U1850 ( .A(n1766), .B(n1765), .Z(n1767) );
  NANDN U1851 ( .A(n1749), .B(n1748), .Z(n1753) );
  NAND U1852 ( .A(n1751), .B(n1750), .Z(n1752) );
  NAND U1853 ( .A(n1753), .B(n1752), .Z(n1768) );
  XNOR U1854 ( .A(n1767), .B(n1768), .Z(n1759) );
  XNOR U1855 ( .A(n1760), .B(n1759), .Z(n1761) );
  XNOR U1856 ( .A(n1762), .B(n1761), .Z(n1795) );
  XNOR U1857 ( .A(sreg[294]), .B(n1795), .Z(n1797) );
  NANDN U1858 ( .A(sreg[293]), .B(n1754), .Z(n1758) );
  NAND U1859 ( .A(n1756), .B(n1755), .Z(n1757) );
  NAND U1860 ( .A(n1758), .B(n1757), .Z(n1796) );
  XNOR U1861 ( .A(n1797), .B(n1796), .Z(c[294]) );
  NANDN U1862 ( .A(n1760), .B(n1759), .Z(n1764) );
  NANDN U1863 ( .A(n1762), .B(n1761), .Z(n1763) );
  AND U1864 ( .A(n1764), .B(n1763), .Z(n1803) );
  NANDN U1865 ( .A(n1766), .B(n1765), .Z(n1770) );
  NANDN U1866 ( .A(n1768), .B(n1767), .Z(n1769) );
  AND U1867 ( .A(n1770), .B(n1769), .Z(n1801) );
  NAND U1868 ( .A(n26), .B(n1771), .Z(n1773) );
  XOR U1869 ( .A(b[7]), .B(a[41]), .Z(n1812) );
  NAND U1870 ( .A(n10531), .B(n1812), .Z(n1772) );
  AND U1871 ( .A(n1773), .B(n1772), .Z(n1831) );
  NAND U1872 ( .A(n23), .B(n1774), .Z(n1776) );
  XOR U1873 ( .A(b[3]), .B(a[45]), .Z(n1815) );
  NAND U1874 ( .A(n24), .B(n1815), .Z(n1775) );
  NAND U1875 ( .A(n1776), .B(n1775), .Z(n1830) );
  XNOR U1876 ( .A(n1831), .B(n1830), .Z(n1833) );
  NAND U1877 ( .A(b[0]), .B(a[47]), .Z(n1777) );
  XNOR U1878 ( .A(b[1]), .B(n1777), .Z(n1779) );
  NANDN U1879 ( .A(b[0]), .B(a[46]), .Z(n1778) );
  NAND U1880 ( .A(n1779), .B(n1778), .Z(n1827) );
  NAND U1881 ( .A(n25), .B(n1780), .Z(n1782) );
  XOR U1882 ( .A(b[5]), .B(a[43]), .Z(n1821) );
  NAND U1883 ( .A(n10456), .B(n1821), .Z(n1781) );
  AND U1884 ( .A(n1782), .B(n1781), .Z(n1825) );
  AND U1885 ( .A(b[7]), .B(a[39]), .Z(n1824) );
  XNOR U1886 ( .A(n1825), .B(n1824), .Z(n1826) );
  XNOR U1887 ( .A(n1827), .B(n1826), .Z(n1832) );
  XOR U1888 ( .A(n1833), .B(n1832), .Z(n1807) );
  NANDN U1889 ( .A(n1784), .B(n1783), .Z(n1788) );
  NANDN U1890 ( .A(n1786), .B(n1785), .Z(n1787) );
  AND U1891 ( .A(n1788), .B(n1787), .Z(n1806) );
  XNOR U1892 ( .A(n1807), .B(n1806), .Z(n1808) );
  NANDN U1893 ( .A(n1790), .B(n1789), .Z(n1794) );
  NAND U1894 ( .A(n1792), .B(n1791), .Z(n1793) );
  NAND U1895 ( .A(n1794), .B(n1793), .Z(n1809) );
  XNOR U1896 ( .A(n1808), .B(n1809), .Z(n1800) );
  XNOR U1897 ( .A(n1801), .B(n1800), .Z(n1802) );
  XNOR U1898 ( .A(n1803), .B(n1802), .Z(n1836) );
  XNOR U1899 ( .A(sreg[295]), .B(n1836), .Z(n1838) );
  NANDN U1900 ( .A(sreg[294]), .B(n1795), .Z(n1799) );
  NAND U1901 ( .A(n1797), .B(n1796), .Z(n1798) );
  NAND U1902 ( .A(n1799), .B(n1798), .Z(n1837) );
  XNOR U1903 ( .A(n1838), .B(n1837), .Z(c[295]) );
  NANDN U1904 ( .A(n1801), .B(n1800), .Z(n1805) );
  NANDN U1905 ( .A(n1803), .B(n1802), .Z(n1804) );
  AND U1906 ( .A(n1805), .B(n1804), .Z(n1844) );
  NANDN U1907 ( .A(n1807), .B(n1806), .Z(n1811) );
  NANDN U1908 ( .A(n1809), .B(n1808), .Z(n1810) );
  AND U1909 ( .A(n1811), .B(n1810), .Z(n1842) );
  NAND U1910 ( .A(n26), .B(n1812), .Z(n1814) );
  XOR U1911 ( .A(b[7]), .B(a[42]), .Z(n1853) );
  NAND U1912 ( .A(n10531), .B(n1853), .Z(n1813) );
  AND U1913 ( .A(n1814), .B(n1813), .Z(n1872) );
  NAND U1914 ( .A(n23), .B(n1815), .Z(n1817) );
  XOR U1915 ( .A(b[3]), .B(a[46]), .Z(n1856) );
  NAND U1916 ( .A(n24), .B(n1856), .Z(n1816) );
  NAND U1917 ( .A(n1817), .B(n1816), .Z(n1871) );
  XNOR U1918 ( .A(n1872), .B(n1871), .Z(n1874) );
  NAND U1919 ( .A(b[0]), .B(a[48]), .Z(n1818) );
  XNOR U1920 ( .A(b[1]), .B(n1818), .Z(n1820) );
  NANDN U1921 ( .A(b[0]), .B(a[47]), .Z(n1819) );
  NAND U1922 ( .A(n1820), .B(n1819), .Z(n1868) );
  NAND U1923 ( .A(n25), .B(n1821), .Z(n1823) );
  XOR U1924 ( .A(b[5]), .B(a[44]), .Z(n1862) );
  NAND U1925 ( .A(n10456), .B(n1862), .Z(n1822) );
  AND U1926 ( .A(n1823), .B(n1822), .Z(n1866) );
  AND U1927 ( .A(b[7]), .B(a[40]), .Z(n1865) );
  XNOR U1928 ( .A(n1866), .B(n1865), .Z(n1867) );
  XNOR U1929 ( .A(n1868), .B(n1867), .Z(n1873) );
  XOR U1930 ( .A(n1874), .B(n1873), .Z(n1848) );
  NANDN U1931 ( .A(n1825), .B(n1824), .Z(n1829) );
  NANDN U1932 ( .A(n1827), .B(n1826), .Z(n1828) );
  AND U1933 ( .A(n1829), .B(n1828), .Z(n1847) );
  XNOR U1934 ( .A(n1848), .B(n1847), .Z(n1849) );
  NANDN U1935 ( .A(n1831), .B(n1830), .Z(n1835) );
  NAND U1936 ( .A(n1833), .B(n1832), .Z(n1834) );
  NAND U1937 ( .A(n1835), .B(n1834), .Z(n1850) );
  XNOR U1938 ( .A(n1849), .B(n1850), .Z(n1841) );
  XNOR U1939 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U1940 ( .A(n1844), .B(n1843), .Z(n1877) );
  XNOR U1941 ( .A(sreg[296]), .B(n1877), .Z(n1879) );
  NANDN U1942 ( .A(sreg[295]), .B(n1836), .Z(n1840) );
  NAND U1943 ( .A(n1838), .B(n1837), .Z(n1839) );
  NAND U1944 ( .A(n1840), .B(n1839), .Z(n1878) );
  XNOR U1945 ( .A(n1879), .B(n1878), .Z(c[296]) );
  NANDN U1946 ( .A(n1842), .B(n1841), .Z(n1846) );
  NANDN U1947 ( .A(n1844), .B(n1843), .Z(n1845) );
  AND U1948 ( .A(n1846), .B(n1845), .Z(n1885) );
  NANDN U1949 ( .A(n1848), .B(n1847), .Z(n1852) );
  NANDN U1950 ( .A(n1850), .B(n1849), .Z(n1851) );
  AND U1951 ( .A(n1852), .B(n1851), .Z(n1883) );
  NAND U1952 ( .A(n26), .B(n1853), .Z(n1855) );
  XOR U1953 ( .A(b[7]), .B(a[43]), .Z(n1894) );
  NAND U1954 ( .A(n10531), .B(n1894), .Z(n1854) );
  AND U1955 ( .A(n1855), .B(n1854), .Z(n1913) );
  NAND U1956 ( .A(n23), .B(n1856), .Z(n1858) );
  XOR U1957 ( .A(b[3]), .B(a[47]), .Z(n1897) );
  NAND U1958 ( .A(n24), .B(n1897), .Z(n1857) );
  NAND U1959 ( .A(n1858), .B(n1857), .Z(n1912) );
  XNOR U1960 ( .A(n1913), .B(n1912), .Z(n1915) );
  NAND U1961 ( .A(b[0]), .B(a[49]), .Z(n1859) );
  XNOR U1962 ( .A(b[1]), .B(n1859), .Z(n1861) );
  NANDN U1963 ( .A(b[0]), .B(a[48]), .Z(n1860) );
  NAND U1964 ( .A(n1861), .B(n1860), .Z(n1909) );
  NAND U1965 ( .A(n25), .B(n1862), .Z(n1864) );
  XOR U1966 ( .A(b[5]), .B(a[45]), .Z(n1900) );
  NAND U1967 ( .A(n10456), .B(n1900), .Z(n1863) );
  AND U1968 ( .A(n1864), .B(n1863), .Z(n1907) );
  AND U1969 ( .A(b[7]), .B(a[41]), .Z(n1906) );
  XNOR U1970 ( .A(n1907), .B(n1906), .Z(n1908) );
  XNOR U1971 ( .A(n1909), .B(n1908), .Z(n1914) );
  XOR U1972 ( .A(n1915), .B(n1914), .Z(n1889) );
  NANDN U1973 ( .A(n1866), .B(n1865), .Z(n1870) );
  NANDN U1974 ( .A(n1868), .B(n1867), .Z(n1869) );
  AND U1975 ( .A(n1870), .B(n1869), .Z(n1888) );
  XNOR U1976 ( .A(n1889), .B(n1888), .Z(n1890) );
  NANDN U1977 ( .A(n1872), .B(n1871), .Z(n1876) );
  NAND U1978 ( .A(n1874), .B(n1873), .Z(n1875) );
  NAND U1979 ( .A(n1876), .B(n1875), .Z(n1891) );
  XNOR U1980 ( .A(n1890), .B(n1891), .Z(n1882) );
  XNOR U1981 ( .A(n1883), .B(n1882), .Z(n1884) );
  XNOR U1982 ( .A(n1885), .B(n1884), .Z(n1918) );
  XNOR U1983 ( .A(sreg[297]), .B(n1918), .Z(n1920) );
  NANDN U1984 ( .A(sreg[296]), .B(n1877), .Z(n1881) );
  NAND U1985 ( .A(n1879), .B(n1878), .Z(n1880) );
  NAND U1986 ( .A(n1881), .B(n1880), .Z(n1919) );
  XNOR U1987 ( .A(n1920), .B(n1919), .Z(c[297]) );
  NANDN U1988 ( .A(n1883), .B(n1882), .Z(n1887) );
  NANDN U1989 ( .A(n1885), .B(n1884), .Z(n1886) );
  AND U1990 ( .A(n1887), .B(n1886), .Z(n1926) );
  NANDN U1991 ( .A(n1889), .B(n1888), .Z(n1893) );
  NANDN U1992 ( .A(n1891), .B(n1890), .Z(n1892) );
  AND U1993 ( .A(n1893), .B(n1892), .Z(n1924) );
  NAND U1994 ( .A(n26), .B(n1894), .Z(n1896) );
  XOR U1995 ( .A(b[7]), .B(a[44]), .Z(n1935) );
  NAND U1996 ( .A(n10531), .B(n1935), .Z(n1895) );
  AND U1997 ( .A(n1896), .B(n1895), .Z(n1954) );
  NAND U1998 ( .A(n23), .B(n1897), .Z(n1899) );
  XOR U1999 ( .A(b[3]), .B(a[48]), .Z(n1938) );
  NAND U2000 ( .A(n24), .B(n1938), .Z(n1898) );
  NAND U2001 ( .A(n1899), .B(n1898), .Z(n1953) );
  XNOR U2002 ( .A(n1954), .B(n1953), .Z(n1956) );
  NAND U2003 ( .A(n25), .B(n1900), .Z(n1902) );
  XOR U2004 ( .A(b[5]), .B(a[46]), .Z(n1944) );
  NAND U2005 ( .A(n10456), .B(n1944), .Z(n1901) );
  AND U2006 ( .A(n1902), .B(n1901), .Z(n1948) );
  AND U2007 ( .A(b[7]), .B(a[42]), .Z(n1947) );
  XNOR U2008 ( .A(n1948), .B(n1947), .Z(n1949) );
  NAND U2009 ( .A(b[0]), .B(a[50]), .Z(n1903) );
  XNOR U2010 ( .A(b[1]), .B(n1903), .Z(n1905) );
  NANDN U2011 ( .A(b[0]), .B(a[49]), .Z(n1904) );
  NAND U2012 ( .A(n1905), .B(n1904), .Z(n1950) );
  XNOR U2013 ( .A(n1949), .B(n1950), .Z(n1955) );
  XOR U2014 ( .A(n1956), .B(n1955), .Z(n1930) );
  NANDN U2015 ( .A(n1907), .B(n1906), .Z(n1911) );
  NANDN U2016 ( .A(n1909), .B(n1908), .Z(n1910) );
  AND U2017 ( .A(n1911), .B(n1910), .Z(n1929) );
  XNOR U2018 ( .A(n1930), .B(n1929), .Z(n1931) );
  NANDN U2019 ( .A(n1913), .B(n1912), .Z(n1917) );
  NAND U2020 ( .A(n1915), .B(n1914), .Z(n1916) );
  NAND U2021 ( .A(n1917), .B(n1916), .Z(n1932) );
  XNOR U2022 ( .A(n1931), .B(n1932), .Z(n1923) );
  XNOR U2023 ( .A(n1924), .B(n1923), .Z(n1925) );
  XNOR U2024 ( .A(n1926), .B(n1925), .Z(n1959) );
  XNOR U2025 ( .A(sreg[298]), .B(n1959), .Z(n1961) );
  NANDN U2026 ( .A(sreg[297]), .B(n1918), .Z(n1922) );
  NAND U2027 ( .A(n1920), .B(n1919), .Z(n1921) );
  NAND U2028 ( .A(n1922), .B(n1921), .Z(n1960) );
  XNOR U2029 ( .A(n1961), .B(n1960), .Z(c[298]) );
  NANDN U2030 ( .A(n1924), .B(n1923), .Z(n1928) );
  NANDN U2031 ( .A(n1926), .B(n1925), .Z(n1927) );
  AND U2032 ( .A(n1928), .B(n1927), .Z(n1967) );
  NANDN U2033 ( .A(n1930), .B(n1929), .Z(n1934) );
  NANDN U2034 ( .A(n1932), .B(n1931), .Z(n1933) );
  AND U2035 ( .A(n1934), .B(n1933), .Z(n1965) );
  NAND U2036 ( .A(n26), .B(n1935), .Z(n1937) );
  XOR U2037 ( .A(b[7]), .B(a[45]), .Z(n1976) );
  NAND U2038 ( .A(n10531), .B(n1976), .Z(n1936) );
  AND U2039 ( .A(n1937), .B(n1936), .Z(n1995) );
  NAND U2040 ( .A(n23), .B(n1938), .Z(n1940) );
  XOR U2041 ( .A(b[3]), .B(a[49]), .Z(n1979) );
  NAND U2042 ( .A(n24), .B(n1979), .Z(n1939) );
  NAND U2043 ( .A(n1940), .B(n1939), .Z(n1994) );
  XNOR U2044 ( .A(n1995), .B(n1994), .Z(n1997) );
  NAND U2045 ( .A(b[0]), .B(a[51]), .Z(n1941) );
  XNOR U2046 ( .A(b[1]), .B(n1941), .Z(n1943) );
  NANDN U2047 ( .A(b[0]), .B(a[50]), .Z(n1942) );
  NAND U2048 ( .A(n1943), .B(n1942), .Z(n1991) );
  NAND U2049 ( .A(n25), .B(n1944), .Z(n1946) );
  XOR U2050 ( .A(b[5]), .B(a[47]), .Z(n1985) );
  NAND U2051 ( .A(n10456), .B(n1985), .Z(n1945) );
  AND U2052 ( .A(n1946), .B(n1945), .Z(n1989) );
  AND U2053 ( .A(b[7]), .B(a[43]), .Z(n1988) );
  XNOR U2054 ( .A(n1989), .B(n1988), .Z(n1990) );
  XNOR U2055 ( .A(n1991), .B(n1990), .Z(n1996) );
  XOR U2056 ( .A(n1997), .B(n1996), .Z(n1971) );
  NANDN U2057 ( .A(n1948), .B(n1947), .Z(n1952) );
  NANDN U2058 ( .A(n1950), .B(n1949), .Z(n1951) );
  AND U2059 ( .A(n1952), .B(n1951), .Z(n1970) );
  XNOR U2060 ( .A(n1971), .B(n1970), .Z(n1972) );
  NANDN U2061 ( .A(n1954), .B(n1953), .Z(n1958) );
  NAND U2062 ( .A(n1956), .B(n1955), .Z(n1957) );
  NAND U2063 ( .A(n1958), .B(n1957), .Z(n1973) );
  XNOR U2064 ( .A(n1972), .B(n1973), .Z(n1964) );
  XNOR U2065 ( .A(n1965), .B(n1964), .Z(n1966) );
  XNOR U2066 ( .A(n1967), .B(n1966), .Z(n2000) );
  XNOR U2067 ( .A(sreg[299]), .B(n2000), .Z(n2002) );
  NANDN U2068 ( .A(sreg[298]), .B(n1959), .Z(n1963) );
  NAND U2069 ( .A(n1961), .B(n1960), .Z(n1962) );
  NAND U2070 ( .A(n1963), .B(n1962), .Z(n2001) );
  XNOR U2071 ( .A(n2002), .B(n2001), .Z(c[299]) );
  NANDN U2072 ( .A(n1965), .B(n1964), .Z(n1969) );
  NANDN U2073 ( .A(n1967), .B(n1966), .Z(n1968) );
  AND U2074 ( .A(n1969), .B(n1968), .Z(n2008) );
  NANDN U2075 ( .A(n1971), .B(n1970), .Z(n1975) );
  NANDN U2076 ( .A(n1973), .B(n1972), .Z(n1974) );
  AND U2077 ( .A(n1975), .B(n1974), .Z(n2006) );
  NAND U2078 ( .A(n26), .B(n1976), .Z(n1978) );
  XOR U2079 ( .A(b[7]), .B(a[46]), .Z(n2017) );
  NAND U2080 ( .A(n10531), .B(n2017), .Z(n1977) );
  AND U2081 ( .A(n1978), .B(n1977), .Z(n2036) );
  NAND U2082 ( .A(n23), .B(n1979), .Z(n1981) );
  XOR U2083 ( .A(b[3]), .B(a[50]), .Z(n2020) );
  NAND U2084 ( .A(n24), .B(n2020), .Z(n1980) );
  NAND U2085 ( .A(n1981), .B(n1980), .Z(n2035) );
  XNOR U2086 ( .A(n2036), .B(n2035), .Z(n2038) );
  NAND U2087 ( .A(b[0]), .B(a[52]), .Z(n1982) );
  XNOR U2088 ( .A(b[1]), .B(n1982), .Z(n1984) );
  NANDN U2089 ( .A(b[0]), .B(a[51]), .Z(n1983) );
  NAND U2090 ( .A(n1984), .B(n1983), .Z(n2032) );
  NAND U2091 ( .A(n25), .B(n1985), .Z(n1987) );
  XOR U2092 ( .A(b[5]), .B(a[48]), .Z(n2026) );
  NAND U2093 ( .A(n10456), .B(n2026), .Z(n1986) );
  AND U2094 ( .A(n1987), .B(n1986), .Z(n2030) );
  AND U2095 ( .A(b[7]), .B(a[44]), .Z(n2029) );
  XNOR U2096 ( .A(n2030), .B(n2029), .Z(n2031) );
  XNOR U2097 ( .A(n2032), .B(n2031), .Z(n2037) );
  XOR U2098 ( .A(n2038), .B(n2037), .Z(n2012) );
  NANDN U2099 ( .A(n1989), .B(n1988), .Z(n1993) );
  NANDN U2100 ( .A(n1991), .B(n1990), .Z(n1992) );
  AND U2101 ( .A(n1993), .B(n1992), .Z(n2011) );
  XNOR U2102 ( .A(n2012), .B(n2011), .Z(n2013) );
  NANDN U2103 ( .A(n1995), .B(n1994), .Z(n1999) );
  NAND U2104 ( .A(n1997), .B(n1996), .Z(n1998) );
  NAND U2105 ( .A(n1999), .B(n1998), .Z(n2014) );
  XNOR U2106 ( .A(n2013), .B(n2014), .Z(n2005) );
  XNOR U2107 ( .A(n2006), .B(n2005), .Z(n2007) );
  XNOR U2108 ( .A(n2008), .B(n2007), .Z(n2041) );
  XNOR U2109 ( .A(sreg[300]), .B(n2041), .Z(n2043) );
  NANDN U2110 ( .A(sreg[299]), .B(n2000), .Z(n2004) );
  NAND U2111 ( .A(n2002), .B(n2001), .Z(n2003) );
  NAND U2112 ( .A(n2004), .B(n2003), .Z(n2042) );
  XNOR U2113 ( .A(n2043), .B(n2042), .Z(c[300]) );
  NANDN U2114 ( .A(n2006), .B(n2005), .Z(n2010) );
  NANDN U2115 ( .A(n2008), .B(n2007), .Z(n2009) );
  AND U2116 ( .A(n2010), .B(n2009), .Z(n2049) );
  NANDN U2117 ( .A(n2012), .B(n2011), .Z(n2016) );
  NANDN U2118 ( .A(n2014), .B(n2013), .Z(n2015) );
  AND U2119 ( .A(n2016), .B(n2015), .Z(n2047) );
  NAND U2120 ( .A(n26), .B(n2017), .Z(n2019) );
  XOR U2121 ( .A(b[7]), .B(a[47]), .Z(n2058) );
  NAND U2122 ( .A(n10531), .B(n2058), .Z(n2018) );
  AND U2123 ( .A(n2019), .B(n2018), .Z(n2077) );
  NAND U2124 ( .A(n23), .B(n2020), .Z(n2022) );
  XOR U2125 ( .A(b[3]), .B(a[51]), .Z(n2061) );
  NAND U2126 ( .A(n24), .B(n2061), .Z(n2021) );
  NAND U2127 ( .A(n2022), .B(n2021), .Z(n2076) );
  XNOR U2128 ( .A(n2077), .B(n2076), .Z(n2079) );
  NAND U2129 ( .A(b[0]), .B(a[53]), .Z(n2023) );
  XNOR U2130 ( .A(b[1]), .B(n2023), .Z(n2025) );
  NANDN U2131 ( .A(b[0]), .B(a[52]), .Z(n2024) );
  NAND U2132 ( .A(n2025), .B(n2024), .Z(n2073) );
  NAND U2133 ( .A(n25), .B(n2026), .Z(n2028) );
  XOR U2134 ( .A(b[5]), .B(a[49]), .Z(n2064) );
  NAND U2135 ( .A(n10456), .B(n2064), .Z(n2027) );
  AND U2136 ( .A(n2028), .B(n2027), .Z(n2071) );
  AND U2137 ( .A(b[7]), .B(a[45]), .Z(n2070) );
  XNOR U2138 ( .A(n2071), .B(n2070), .Z(n2072) );
  XNOR U2139 ( .A(n2073), .B(n2072), .Z(n2078) );
  XOR U2140 ( .A(n2079), .B(n2078), .Z(n2053) );
  NANDN U2141 ( .A(n2030), .B(n2029), .Z(n2034) );
  NANDN U2142 ( .A(n2032), .B(n2031), .Z(n2033) );
  AND U2143 ( .A(n2034), .B(n2033), .Z(n2052) );
  XNOR U2144 ( .A(n2053), .B(n2052), .Z(n2054) );
  NANDN U2145 ( .A(n2036), .B(n2035), .Z(n2040) );
  NAND U2146 ( .A(n2038), .B(n2037), .Z(n2039) );
  NAND U2147 ( .A(n2040), .B(n2039), .Z(n2055) );
  XNOR U2148 ( .A(n2054), .B(n2055), .Z(n2046) );
  XNOR U2149 ( .A(n2047), .B(n2046), .Z(n2048) );
  XNOR U2150 ( .A(n2049), .B(n2048), .Z(n2082) );
  XNOR U2151 ( .A(sreg[301]), .B(n2082), .Z(n2084) );
  NANDN U2152 ( .A(sreg[300]), .B(n2041), .Z(n2045) );
  NAND U2153 ( .A(n2043), .B(n2042), .Z(n2044) );
  NAND U2154 ( .A(n2045), .B(n2044), .Z(n2083) );
  XNOR U2155 ( .A(n2084), .B(n2083), .Z(c[301]) );
  NANDN U2156 ( .A(n2047), .B(n2046), .Z(n2051) );
  NANDN U2157 ( .A(n2049), .B(n2048), .Z(n2050) );
  AND U2158 ( .A(n2051), .B(n2050), .Z(n2090) );
  NANDN U2159 ( .A(n2053), .B(n2052), .Z(n2057) );
  NANDN U2160 ( .A(n2055), .B(n2054), .Z(n2056) );
  AND U2161 ( .A(n2057), .B(n2056), .Z(n2088) );
  NAND U2162 ( .A(n26), .B(n2058), .Z(n2060) );
  XOR U2163 ( .A(b[7]), .B(a[48]), .Z(n2099) );
  NAND U2164 ( .A(n10531), .B(n2099), .Z(n2059) );
  AND U2165 ( .A(n2060), .B(n2059), .Z(n2118) );
  NAND U2166 ( .A(n23), .B(n2061), .Z(n2063) );
  XOR U2167 ( .A(b[3]), .B(a[52]), .Z(n2102) );
  NAND U2168 ( .A(n24), .B(n2102), .Z(n2062) );
  NAND U2169 ( .A(n2063), .B(n2062), .Z(n2117) );
  XNOR U2170 ( .A(n2118), .B(n2117), .Z(n2120) );
  NAND U2171 ( .A(n25), .B(n2064), .Z(n2066) );
  XOR U2172 ( .A(b[5]), .B(a[50]), .Z(n2105) );
  NAND U2173 ( .A(n10456), .B(n2105), .Z(n2065) );
  AND U2174 ( .A(n2066), .B(n2065), .Z(n2112) );
  AND U2175 ( .A(b[7]), .B(a[46]), .Z(n2111) );
  XNOR U2176 ( .A(n2112), .B(n2111), .Z(n2113) );
  NAND U2177 ( .A(b[0]), .B(a[54]), .Z(n2067) );
  XNOR U2178 ( .A(b[1]), .B(n2067), .Z(n2069) );
  NANDN U2179 ( .A(b[0]), .B(a[53]), .Z(n2068) );
  NAND U2180 ( .A(n2069), .B(n2068), .Z(n2114) );
  XNOR U2181 ( .A(n2113), .B(n2114), .Z(n2119) );
  XOR U2182 ( .A(n2120), .B(n2119), .Z(n2094) );
  NANDN U2183 ( .A(n2071), .B(n2070), .Z(n2075) );
  NANDN U2184 ( .A(n2073), .B(n2072), .Z(n2074) );
  AND U2185 ( .A(n2075), .B(n2074), .Z(n2093) );
  XNOR U2186 ( .A(n2094), .B(n2093), .Z(n2095) );
  NANDN U2187 ( .A(n2077), .B(n2076), .Z(n2081) );
  NAND U2188 ( .A(n2079), .B(n2078), .Z(n2080) );
  NAND U2189 ( .A(n2081), .B(n2080), .Z(n2096) );
  XNOR U2190 ( .A(n2095), .B(n2096), .Z(n2087) );
  XNOR U2191 ( .A(n2088), .B(n2087), .Z(n2089) );
  XNOR U2192 ( .A(n2090), .B(n2089), .Z(n2123) );
  XNOR U2193 ( .A(sreg[302]), .B(n2123), .Z(n2125) );
  NANDN U2194 ( .A(sreg[301]), .B(n2082), .Z(n2086) );
  NAND U2195 ( .A(n2084), .B(n2083), .Z(n2085) );
  NAND U2196 ( .A(n2086), .B(n2085), .Z(n2124) );
  XNOR U2197 ( .A(n2125), .B(n2124), .Z(c[302]) );
  NANDN U2198 ( .A(n2088), .B(n2087), .Z(n2092) );
  NANDN U2199 ( .A(n2090), .B(n2089), .Z(n2091) );
  AND U2200 ( .A(n2092), .B(n2091), .Z(n2131) );
  NANDN U2201 ( .A(n2094), .B(n2093), .Z(n2098) );
  NANDN U2202 ( .A(n2096), .B(n2095), .Z(n2097) );
  AND U2203 ( .A(n2098), .B(n2097), .Z(n2129) );
  NAND U2204 ( .A(n26), .B(n2099), .Z(n2101) );
  XOR U2205 ( .A(b[7]), .B(a[49]), .Z(n2140) );
  NAND U2206 ( .A(n10531), .B(n2140), .Z(n2100) );
  AND U2207 ( .A(n2101), .B(n2100), .Z(n2159) );
  NAND U2208 ( .A(n23), .B(n2102), .Z(n2104) );
  XOR U2209 ( .A(b[3]), .B(a[53]), .Z(n2143) );
  NAND U2210 ( .A(n24), .B(n2143), .Z(n2103) );
  NAND U2211 ( .A(n2104), .B(n2103), .Z(n2158) );
  XNOR U2212 ( .A(n2159), .B(n2158), .Z(n2161) );
  NAND U2213 ( .A(n25), .B(n2105), .Z(n2107) );
  XOR U2214 ( .A(b[5]), .B(a[51]), .Z(n2149) );
  NAND U2215 ( .A(n10456), .B(n2149), .Z(n2106) );
  AND U2216 ( .A(n2107), .B(n2106), .Z(n2153) );
  AND U2217 ( .A(b[7]), .B(a[47]), .Z(n2152) );
  XNOR U2218 ( .A(n2153), .B(n2152), .Z(n2154) );
  NAND U2219 ( .A(b[0]), .B(a[55]), .Z(n2108) );
  XNOR U2220 ( .A(b[1]), .B(n2108), .Z(n2110) );
  NANDN U2221 ( .A(b[0]), .B(a[54]), .Z(n2109) );
  NAND U2222 ( .A(n2110), .B(n2109), .Z(n2155) );
  XNOR U2223 ( .A(n2154), .B(n2155), .Z(n2160) );
  XOR U2224 ( .A(n2161), .B(n2160), .Z(n2135) );
  NANDN U2225 ( .A(n2112), .B(n2111), .Z(n2116) );
  NANDN U2226 ( .A(n2114), .B(n2113), .Z(n2115) );
  AND U2227 ( .A(n2116), .B(n2115), .Z(n2134) );
  XNOR U2228 ( .A(n2135), .B(n2134), .Z(n2136) );
  NANDN U2229 ( .A(n2118), .B(n2117), .Z(n2122) );
  NAND U2230 ( .A(n2120), .B(n2119), .Z(n2121) );
  NAND U2231 ( .A(n2122), .B(n2121), .Z(n2137) );
  XNOR U2232 ( .A(n2136), .B(n2137), .Z(n2128) );
  XNOR U2233 ( .A(n2129), .B(n2128), .Z(n2130) );
  XNOR U2234 ( .A(n2131), .B(n2130), .Z(n2164) );
  XNOR U2235 ( .A(sreg[303]), .B(n2164), .Z(n2166) );
  NANDN U2236 ( .A(sreg[302]), .B(n2123), .Z(n2127) );
  NAND U2237 ( .A(n2125), .B(n2124), .Z(n2126) );
  NAND U2238 ( .A(n2127), .B(n2126), .Z(n2165) );
  XNOR U2239 ( .A(n2166), .B(n2165), .Z(c[303]) );
  NANDN U2240 ( .A(n2129), .B(n2128), .Z(n2133) );
  NANDN U2241 ( .A(n2131), .B(n2130), .Z(n2132) );
  AND U2242 ( .A(n2133), .B(n2132), .Z(n2172) );
  NANDN U2243 ( .A(n2135), .B(n2134), .Z(n2139) );
  NANDN U2244 ( .A(n2137), .B(n2136), .Z(n2138) );
  AND U2245 ( .A(n2139), .B(n2138), .Z(n2170) );
  NAND U2246 ( .A(n26), .B(n2140), .Z(n2142) );
  XOR U2247 ( .A(b[7]), .B(a[50]), .Z(n2181) );
  NAND U2248 ( .A(n10531), .B(n2181), .Z(n2141) );
  AND U2249 ( .A(n2142), .B(n2141), .Z(n2200) );
  NAND U2250 ( .A(n23), .B(n2143), .Z(n2145) );
  XOR U2251 ( .A(b[3]), .B(a[54]), .Z(n2184) );
  NAND U2252 ( .A(n24), .B(n2184), .Z(n2144) );
  NAND U2253 ( .A(n2145), .B(n2144), .Z(n2199) );
  XNOR U2254 ( .A(n2200), .B(n2199), .Z(n2202) );
  NAND U2255 ( .A(b[0]), .B(a[56]), .Z(n2146) );
  XNOR U2256 ( .A(b[1]), .B(n2146), .Z(n2148) );
  NANDN U2257 ( .A(b[0]), .B(a[55]), .Z(n2147) );
  NAND U2258 ( .A(n2148), .B(n2147), .Z(n2196) );
  NAND U2259 ( .A(n25), .B(n2149), .Z(n2151) );
  XOR U2260 ( .A(b[5]), .B(a[52]), .Z(n2190) );
  NAND U2261 ( .A(n10456), .B(n2190), .Z(n2150) );
  AND U2262 ( .A(n2151), .B(n2150), .Z(n2194) );
  AND U2263 ( .A(b[7]), .B(a[48]), .Z(n2193) );
  XNOR U2264 ( .A(n2194), .B(n2193), .Z(n2195) );
  XNOR U2265 ( .A(n2196), .B(n2195), .Z(n2201) );
  XOR U2266 ( .A(n2202), .B(n2201), .Z(n2176) );
  NANDN U2267 ( .A(n2153), .B(n2152), .Z(n2157) );
  NANDN U2268 ( .A(n2155), .B(n2154), .Z(n2156) );
  AND U2269 ( .A(n2157), .B(n2156), .Z(n2175) );
  XNOR U2270 ( .A(n2176), .B(n2175), .Z(n2177) );
  NANDN U2271 ( .A(n2159), .B(n2158), .Z(n2163) );
  NAND U2272 ( .A(n2161), .B(n2160), .Z(n2162) );
  NAND U2273 ( .A(n2163), .B(n2162), .Z(n2178) );
  XNOR U2274 ( .A(n2177), .B(n2178), .Z(n2169) );
  XNOR U2275 ( .A(n2170), .B(n2169), .Z(n2171) );
  XNOR U2276 ( .A(n2172), .B(n2171), .Z(n2205) );
  XNOR U2277 ( .A(sreg[304]), .B(n2205), .Z(n2207) );
  NANDN U2278 ( .A(sreg[303]), .B(n2164), .Z(n2168) );
  NAND U2279 ( .A(n2166), .B(n2165), .Z(n2167) );
  NAND U2280 ( .A(n2168), .B(n2167), .Z(n2206) );
  XNOR U2281 ( .A(n2207), .B(n2206), .Z(c[304]) );
  NANDN U2282 ( .A(n2170), .B(n2169), .Z(n2174) );
  NANDN U2283 ( .A(n2172), .B(n2171), .Z(n2173) );
  AND U2284 ( .A(n2174), .B(n2173), .Z(n2213) );
  NANDN U2285 ( .A(n2176), .B(n2175), .Z(n2180) );
  NANDN U2286 ( .A(n2178), .B(n2177), .Z(n2179) );
  AND U2287 ( .A(n2180), .B(n2179), .Z(n2211) );
  NAND U2288 ( .A(n26), .B(n2181), .Z(n2183) );
  XOR U2289 ( .A(b[7]), .B(a[51]), .Z(n2222) );
  NAND U2290 ( .A(n10531), .B(n2222), .Z(n2182) );
  AND U2291 ( .A(n2183), .B(n2182), .Z(n2241) );
  NAND U2292 ( .A(n23), .B(n2184), .Z(n2186) );
  XOR U2293 ( .A(b[3]), .B(a[55]), .Z(n2225) );
  NAND U2294 ( .A(n24), .B(n2225), .Z(n2185) );
  NAND U2295 ( .A(n2186), .B(n2185), .Z(n2240) );
  XNOR U2296 ( .A(n2241), .B(n2240), .Z(n2243) );
  NAND U2297 ( .A(b[0]), .B(a[57]), .Z(n2187) );
  XNOR U2298 ( .A(b[1]), .B(n2187), .Z(n2189) );
  NANDN U2299 ( .A(b[0]), .B(a[56]), .Z(n2188) );
  NAND U2300 ( .A(n2189), .B(n2188), .Z(n2237) );
  NAND U2301 ( .A(n25), .B(n2190), .Z(n2192) );
  XOR U2302 ( .A(b[5]), .B(a[53]), .Z(n2228) );
  NAND U2303 ( .A(n10456), .B(n2228), .Z(n2191) );
  AND U2304 ( .A(n2192), .B(n2191), .Z(n2235) );
  AND U2305 ( .A(b[7]), .B(a[49]), .Z(n2234) );
  XNOR U2306 ( .A(n2235), .B(n2234), .Z(n2236) );
  XNOR U2307 ( .A(n2237), .B(n2236), .Z(n2242) );
  XOR U2308 ( .A(n2243), .B(n2242), .Z(n2217) );
  NANDN U2309 ( .A(n2194), .B(n2193), .Z(n2198) );
  NANDN U2310 ( .A(n2196), .B(n2195), .Z(n2197) );
  AND U2311 ( .A(n2198), .B(n2197), .Z(n2216) );
  XNOR U2312 ( .A(n2217), .B(n2216), .Z(n2218) );
  NANDN U2313 ( .A(n2200), .B(n2199), .Z(n2204) );
  NAND U2314 ( .A(n2202), .B(n2201), .Z(n2203) );
  NAND U2315 ( .A(n2204), .B(n2203), .Z(n2219) );
  XNOR U2316 ( .A(n2218), .B(n2219), .Z(n2210) );
  XNOR U2317 ( .A(n2211), .B(n2210), .Z(n2212) );
  XNOR U2318 ( .A(n2213), .B(n2212), .Z(n2246) );
  XNOR U2319 ( .A(sreg[305]), .B(n2246), .Z(n2248) );
  NANDN U2320 ( .A(sreg[304]), .B(n2205), .Z(n2209) );
  NAND U2321 ( .A(n2207), .B(n2206), .Z(n2208) );
  NAND U2322 ( .A(n2209), .B(n2208), .Z(n2247) );
  XNOR U2323 ( .A(n2248), .B(n2247), .Z(c[305]) );
  NANDN U2324 ( .A(n2211), .B(n2210), .Z(n2215) );
  NANDN U2325 ( .A(n2213), .B(n2212), .Z(n2214) );
  AND U2326 ( .A(n2215), .B(n2214), .Z(n2254) );
  NANDN U2327 ( .A(n2217), .B(n2216), .Z(n2221) );
  NANDN U2328 ( .A(n2219), .B(n2218), .Z(n2220) );
  AND U2329 ( .A(n2221), .B(n2220), .Z(n2252) );
  NAND U2330 ( .A(n26), .B(n2222), .Z(n2224) );
  XOR U2331 ( .A(b[7]), .B(a[52]), .Z(n2263) );
  NAND U2332 ( .A(n10531), .B(n2263), .Z(n2223) );
  AND U2333 ( .A(n2224), .B(n2223), .Z(n2282) );
  NAND U2334 ( .A(n23), .B(n2225), .Z(n2227) );
  XOR U2335 ( .A(b[3]), .B(a[56]), .Z(n2266) );
  NAND U2336 ( .A(n24), .B(n2266), .Z(n2226) );
  NAND U2337 ( .A(n2227), .B(n2226), .Z(n2281) );
  XNOR U2338 ( .A(n2282), .B(n2281), .Z(n2284) );
  NAND U2339 ( .A(n25), .B(n2228), .Z(n2230) );
  XOR U2340 ( .A(b[5]), .B(a[54]), .Z(n2272) );
  NAND U2341 ( .A(n10456), .B(n2272), .Z(n2229) );
  AND U2342 ( .A(n2230), .B(n2229), .Z(n2276) );
  AND U2343 ( .A(b[7]), .B(a[50]), .Z(n2275) );
  XNOR U2344 ( .A(n2276), .B(n2275), .Z(n2277) );
  NAND U2345 ( .A(b[0]), .B(a[58]), .Z(n2231) );
  XNOR U2346 ( .A(b[1]), .B(n2231), .Z(n2233) );
  NANDN U2347 ( .A(b[0]), .B(a[57]), .Z(n2232) );
  NAND U2348 ( .A(n2233), .B(n2232), .Z(n2278) );
  XNOR U2349 ( .A(n2277), .B(n2278), .Z(n2283) );
  XOR U2350 ( .A(n2284), .B(n2283), .Z(n2258) );
  NANDN U2351 ( .A(n2235), .B(n2234), .Z(n2239) );
  NANDN U2352 ( .A(n2237), .B(n2236), .Z(n2238) );
  AND U2353 ( .A(n2239), .B(n2238), .Z(n2257) );
  XNOR U2354 ( .A(n2258), .B(n2257), .Z(n2259) );
  NANDN U2355 ( .A(n2241), .B(n2240), .Z(n2245) );
  NAND U2356 ( .A(n2243), .B(n2242), .Z(n2244) );
  NAND U2357 ( .A(n2245), .B(n2244), .Z(n2260) );
  XNOR U2358 ( .A(n2259), .B(n2260), .Z(n2251) );
  XNOR U2359 ( .A(n2252), .B(n2251), .Z(n2253) );
  XNOR U2360 ( .A(n2254), .B(n2253), .Z(n2287) );
  XNOR U2361 ( .A(sreg[306]), .B(n2287), .Z(n2289) );
  NANDN U2362 ( .A(sreg[305]), .B(n2246), .Z(n2250) );
  NAND U2363 ( .A(n2248), .B(n2247), .Z(n2249) );
  NAND U2364 ( .A(n2250), .B(n2249), .Z(n2288) );
  XNOR U2365 ( .A(n2289), .B(n2288), .Z(c[306]) );
  NANDN U2366 ( .A(n2252), .B(n2251), .Z(n2256) );
  NANDN U2367 ( .A(n2254), .B(n2253), .Z(n2255) );
  AND U2368 ( .A(n2256), .B(n2255), .Z(n2295) );
  NANDN U2369 ( .A(n2258), .B(n2257), .Z(n2262) );
  NANDN U2370 ( .A(n2260), .B(n2259), .Z(n2261) );
  AND U2371 ( .A(n2262), .B(n2261), .Z(n2293) );
  NAND U2372 ( .A(n26), .B(n2263), .Z(n2265) );
  XOR U2373 ( .A(b[7]), .B(a[53]), .Z(n2304) );
  NAND U2374 ( .A(n10531), .B(n2304), .Z(n2264) );
  AND U2375 ( .A(n2265), .B(n2264), .Z(n2323) );
  NAND U2376 ( .A(n23), .B(n2266), .Z(n2268) );
  XOR U2377 ( .A(b[3]), .B(a[57]), .Z(n2307) );
  NAND U2378 ( .A(n24), .B(n2307), .Z(n2267) );
  NAND U2379 ( .A(n2268), .B(n2267), .Z(n2322) );
  XNOR U2380 ( .A(n2323), .B(n2322), .Z(n2325) );
  NAND U2381 ( .A(b[0]), .B(a[59]), .Z(n2269) );
  XNOR U2382 ( .A(b[1]), .B(n2269), .Z(n2271) );
  NANDN U2383 ( .A(b[0]), .B(a[58]), .Z(n2270) );
  NAND U2384 ( .A(n2271), .B(n2270), .Z(n2319) );
  NAND U2385 ( .A(n25), .B(n2272), .Z(n2274) );
  XOR U2386 ( .A(b[5]), .B(a[55]), .Z(n2313) );
  NAND U2387 ( .A(n10456), .B(n2313), .Z(n2273) );
  AND U2388 ( .A(n2274), .B(n2273), .Z(n2317) );
  AND U2389 ( .A(b[7]), .B(a[51]), .Z(n2316) );
  XNOR U2390 ( .A(n2317), .B(n2316), .Z(n2318) );
  XNOR U2391 ( .A(n2319), .B(n2318), .Z(n2324) );
  XOR U2392 ( .A(n2325), .B(n2324), .Z(n2299) );
  NANDN U2393 ( .A(n2276), .B(n2275), .Z(n2280) );
  NANDN U2394 ( .A(n2278), .B(n2277), .Z(n2279) );
  AND U2395 ( .A(n2280), .B(n2279), .Z(n2298) );
  XNOR U2396 ( .A(n2299), .B(n2298), .Z(n2300) );
  NANDN U2397 ( .A(n2282), .B(n2281), .Z(n2286) );
  NAND U2398 ( .A(n2284), .B(n2283), .Z(n2285) );
  NAND U2399 ( .A(n2286), .B(n2285), .Z(n2301) );
  XNOR U2400 ( .A(n2300), .B(n2301), .Z(n2292) );
  XNOR U2401 ( .A(n2293), .B(n2292), .Z(n2294) );
  XNOR U2402 ( .A(n2295), .B(n2294), .Z(n2328) );
  XNOR U2403 ( .A(sreg[307]), .B(n2328), .Z(n2330) );
  NANDN U2404 ( .A(sreg[306]), .B(n2287), .Z(n2291) );
  NAND U2405 ( .A(n2289), .B(n2288), .Z(n2290) );
  NAND U2406 ( .A(n2291), .B(n2290), .Z(n2329) );
  XNOR U2407 ( .A(n2330), .B(n2329), .Z(c[307]) );
  NANDN U2408 ( .A(n2293), .B(n2292), .Z(n2297) );
  NANDN U2409 ( .A(n2295), .B(n2294), .Z(n2296) );
  AND U2410 ( .A(n2297), .B(n2296), .Z(n2336) );
  NANDN U2411 ( .A(n2299), .B(n2298), .Z(n2303) );
  NANDN U2412 ( .A(n2301), .B(n2300), .Z(n2302) );
  AND U2413 ( .A(n2303), .B(n2302), .Z(n2334) );
  NAND U2414 ( .A(n26), .B(n2304), .Z(n2306) );
  XOR U2415 ( .A(b[7]), .B(a[54]), .Z(n2345) );
  NAND U2416 ( .A(n10531), .B(n2345), .Z(n2305) );
  AND U2417 ( .A(n2306), .B(n2305), .Z(n2364) );
  NAND U2418 ( .A(n23), .B(n2307), .Z(n2309) );
  XOR U2419 ( .A(b[3]), .B(a[58]), .Z(n2348) );
  NAND U2420 ( .A(n24), .B(n2348), .Z(n2308) );
  NAND U2421 ( .A(n2309), .B(n2308), .Z(n2363) );
  XNOR U2422 ( .A(n2364), .B(n2363), .Z(n2366) );
  NAND U2423 ( .A(b[0]), .B(a[60]), .Z(n2310) );
  XNOR U2424 ( .A(b[1]), .B(n2310), .Z(n2312) );
  NANDN U2425 ( .A(b[0]), .B(a[59]), .Z(n2311) );
  NAND U2426 ( .A(n2312), .B(n2311), .Z(n2360) );
  NAND U2427 ( .A(n25), .B(n2313), .Z(n2315) );
  XOR U2428 ( .A(b[5]), .B(a[56]), .Z(n2354) );
  NAND U2429 ( .A(n10456), .B(n2354), .Z(n2314) );
  AND U2430 ( .A(n2315), .B(n2314), .Z(n2358) );
  AND U2431 ( .A(b[7]), .B(a[52]), .Z(n2357) );
  XNOR U2432 ( .A(n2358), .B(n2357), .Z(n2359) );
  XNOR U2433 ( .A(n2360), .B(n2359), .Z(n2365) );
  XOR U2434 ( .A(n2366), .B(n2365), .Z(n2340) );
  NANDN U2435 ( .A(n2317), .B(n2316), .Z(n2321) );
  NANDN U2436 ( .A(n2319), .B(n2318), .Z(n2320) );
  AND U2437 ( .A(n2321), .B(n2320), .Z(n2339) );
  XNOR U2438 ( .A(n2340), .B(n2339), .Z(n2341) );
  NANDN U2439 ( .A(n2323), .B(n2322), .Z(n2327) );
  NAND U2440 ( .A(n2325), .B(n2324), .Z(n2326) );
  NAND U2441 ( .A(n2327), .B(n2326), .Z(n2342) );
  XNOR U2442 ( .A(n2341), .B(n2342), .Z(n2333) );
  XNOR U2443 ( .A(n2334), .B(n2333), .Z(n2335) );
  XNOR U2444 ( .A(n2336), .B(n2335), .Z(n2369) );
  XNOR U2445 ( .A(sreg[308]), .B(n2369), .Z(n2371) );
  NANDN U2446 ( .A(sreg[307]), .B(n2328), .Z(n2332) );
  NAND U2447 ( .A(n2330), .B(n2329), .Z(n2331) );
  NAND U2448 ( .A(n2332), .B(n2331), .Z(n2370) );
  XNOR U2449 ( .A(n2371), .B(n2370), .Z(c[308]) );
  NANDN U2450 ( .A(n2334), .B(n2333), .Z(n2338) );
  NANDN U2451 ( .A(n2336), .B(n2335), .Z(n2337) );
  AND U2452 ( .A(n2338), .B(n2337), .Z(n2377) );
  NANDN U2453 ( .A(n2340), .B(n2339), .Z(n2344) );
  NANDN U2454 ( .A(n2342), .B(n2341), .Z(n2343) );
  AND U2455 ( .A(n2344), .B(n2343), .Z(n2375) );
  NAND U2456 ( .A(n26), .B(n2345), .Z(n2347) );
  XOR U2457 ( .A(b[7]), .B(a[55]), .Z(n2386) );
  NAND U2458 ( .A(n10531), .B(n2386), .Z(n2346) );
  AND U2459 ( .A(n2347), .B(n2346), .Z(n2405) );
  NAND U2460 ( .A(n23), .B(n2348), .Z(n2350) );
  XOR U2461 ( .A(b[3]), .B(a[59]), .Z(n2389) );
  NAND U2462 ( .A(n24), .B(n2389), .Z(n2349) );
  NAND U2463 ( .A(n2350), .B(n2349), .Z(n2404) );
  XNOR U2464 ( .A(n2405), .B(n2404), .Z(n2407) );
  NAND U2465 ( .A(b[0]), .B(a[61]), .Z(n2351) );
  XNOR U2466 ( .A(b[1]), .B(n2351), .Z(n2353) );
  NANDN U2467 ( .A(b[0]), .B(a[60]), .Z(n2352) );
  NAND U2468 ( .A(n2353), .B(n2352), .Z(n2401) );
  NAND U2469 ( .A(n25), .B(n2354), .Z(n2356) );
  XOR U2470 ( .A(b[5]), .B(a[57]), .Z(n2395) );
  NAND U2471 ( .A(n10456), .B(n2395), .Z(n2355) );
  AND U2472 ( .A(n2356), .B(n2355), .Z(n2399) );
  AND U2473 ( .A(b[7]), .B(a[53]), .Z(n2398) );
  XNOR U2474 ( .A(n2399), .B(n2398), .Z(n2400) );
  XNOR U2475 ( .A(n2401), .B(n2400), .Z(n2406) );
  XOR U2476 ( .A(n2407), .B(n2406), .Z(n2381) );
  NANDN U2477 ( .A(n2358), .B(n2357), .Z(n2362) );
  NANDN U2478 ( .A(n2360), .B(n2359), .Z(n2361) );
  AND U2479 ( .A(n2362), .B(n2361), .Z(n2380) );
  XNOR U2480 ( .A(n2381), .B(n2380), .Z(n2382) );
  NANDN U2481 ( .A(n2364), .B(n2363), .Z(n2368) );
  NAND U2482 ( .A(n2366), .B(n2365), .Z(n2367) );
  NAND U2483 ( .A(n2368), .B(n2367), .Z(n2383) );
  XNOR U2484 ( .A(n2382), .B(n2383), .Z(n2374) );
  XNOR U2485 ( .A(n2375), .B(n2374), .Z(n2376) );
  XNOR U2486 ( .A(n2377), .B(n2376), .Z(n2410) );
  XNOR U2487 ( .A(sreg[309]), .B(n2410), .Z(n2412) );
  NANDN U2488 ( .A(sreg[308]), .B(n2369), .Z(n2373) );
  NAND U2489 ( .A(n2371), .B(n2370), .Z(n2372) );
  NAND U2490 ( .A(n2373), .B(n2372), .Z(n2411) );
  XNOR U2491 ( .A(n2412), .B(n2411), .Z(c[309]) );
  NANDN U2492 ( .A(n2375), .B(n2374), .Z(n2379) );
  NANDN U2493 ( .A(n2377), .B(n2376), .Z(n2378) );
  AND U2494 ( .A(n2379), .B(n2378), .Z(n2418) );
  NANDN U2495 ( .A(n2381), .B(n2380), .Z(n2385) );
  NANDN U2496 ( .A(n2383), .B(n2382), .Z(n2384) );
  AND U2497 ( .A(n2385), .B(n2384), .Z(n2416) );
  NAND U2498 ( .A(n26), .B(n2386), .Z(n2388) );
  XOR U2499 ( .A(b[7]), .B(a[56]), .Z(n2427) );
  NAND U2500 ( .A(n10531), .B(n2427), .Z(n2387) );
  AND U2501 ( .A(n2388), .B(n2387), .Z(n2446) );
  NAND U2502 ( .A(n23), .B(n2389), .Z(n2391) );
  XOR U2503 ( .A(b[3]), .B(a[60]), .Z(n2430) );
  NAND U2504 ( .A(n24), .B(n2430), .Z(n2390) );
  NAND U2505 ( .A(n2391), .B(n2390), .Z(n2445) );
  XNOR U2506 ( .A(n2446), .B(n2445), .Z(n2448) );
  NAND U2507 ( .A(b[0]), .B(a[62]), .Z(n2392) );
  XNOR U2508 ( .A(b[1]), .B(n2392), .Z(n2394) );
  NANDN U2509 ( .A(b[0]), .B(a[61]), .Z(n2393) );
  NAND U2510 ( .A(n2394), .B(n2393), .Z(n2442) );
  NAND U2511 ( .A(n25), .B(n2395), .Z(n2397) );
  XOR U2512 ( .A(b[5]), .B(a[58]), .Z(n2436) );
  NAND U2513 ( .A(n10456), .B(n2436), .Z(n2396) );
  AND U2514 ( .A(n2397), .B(n2396), .Z(n2440) );
  AND U2515 ( .A(b[7]), .B(a[54]), .Z(n2439) );
  XNOR U2516 ( .A(n2440), .B(n2439), .Z(n2441) );
  XNOR U2517 ( .A(n2442), .B(n2441), .Z(n2447) );
  XOR U2518 ( .A(n2448), .B(n2447), .Z(n2422) );
  NANDN U2519 ( .A(n2399), .B(n2398), .Z(n2403) );
  NANDN U2520 ( .A(n2401), .B(n2400), .Z(n2402) );
  AND U2521 ( .A(n2403), .B(n2402), .Z(n2421) );
  XNOR U2522 ( .A(n2422), .B(n2421), .Z(n2423) );
  NANDN U2523 ( .A(n2405), .B(n2404), .Z(n2409) );
  NAND U2524 ( .A(n2407), .B(n2406), .Z(n2408) );
  NAND U2525 ( .A(n2409), .B(n2408), .Z(n2424) );
  XNOR U2526 ( .A(n2423), .B(n2424), .Z(n2415) );
  XNOR U2527 ( .A(n2416), .B(n2415), .Z(n2417) );
  XNOR U2528 ( .A(n2418), .B(n2417), .Z(n2451) );
  XNOR U2529 ( .A(sreg[310]), .B(n2451), .Z(n2453) );
  NANDN U2530 ( .A(sreg[309]), .B(n2410), .Z(n2414) );
  NAND U2531 ( .A(n2412), .B(n2411), .Z(n2413) );
  NAND U2532 ( .A(n2414), .B(n2413), .Z(n2452) );
  XNOR U2533 ( .A(n2453), .B(n2452), .Z(c[310]) );
  NANDN U2534 ( .A(n2416), .B(n2415), .Z(n2420) );
  NANDN U2535 ( .A(n2418), .B(n2417), .Z(n2419) );
  AND U2536 ( .A(n2420), .B(n2419), .Z(n2459) );
  NANDN U2537 ( .A(n2422), .B(n2421), .Z(n2426) );
  NANDN U2538 ( .A(n2424), .B(n2423), .Z(n2425) );
  AND U2539 ( .A(n2426), .B(n2425), .Z(n2457) );
  NAND U2540 ( .A(n26), .B(n2427), .Z(n2429) );
  XOR U2541 ( .A(b[7]), .B(a[57]), .Z(n2468) );
  NAND U2542 ( .A(n10531), .B(n2468), .Z(n2428) );
  AND U2543 ( .A(n2429), .B(n2428), .Z(n2487) );
  NAND U2544 ( .A(n23), .B(n2430), .Z(n2432) );
  XOR U2545 ( .A(b[3]), .B(a[61]), .Z(n2471) );
  NAND U2546 ( .A(n24), .B(n2471), .Z(n2431) );
  NAND U2547 ( .A(n2432), .B(n2431), .Z(n2486) );
  XNOR U2548 ( .A(n2487), .B(n2486), .Z(n2489) );
  NAND U2549 ( .A(b[0]), .B(a[63]), .Z(n2433) );
  XNOR U2550 ( .A(b[1]), .B(n2433), .Z(n2435) );
  NANDN U2551 ( .A(b[0]), .B(a[62]), .Z(n2434) );
  NAND U2552 ( .A(n2435), .B(n2434), .Z(n2483) );
  NAND U2553 ( .A(n25), .B(n2436), .Z(n2438) );
  XOR U2554 ( .A(b[5]), .B(a[59]), .Z(n2474) );
  NAND U2555 ( .A(n10456), .B(n2474), .Z(n2437) );
  AND U2556 ( .A(n2438), .B(n2437), .Z(n2481) );
  AND U2557 ( .A(b[7]), .B(a[55]), .Z(n2480) );
  XNOR U2558 ( .A(n2481), .B(n2480), .Z(n2482) );
  XNOR U2559 ( .A(n2483), .B(n2482), .Z(n2488) );
  XOR U2560 ( .A(n2489), .B(n2488), .Z(n2463) );
  NANDN U2561 ( .A(n2440), .B(n2439), .Z(n2444) );
  NANDN U2562 ( .A(n2442), .B(n2441), .Z(n2443) );
  AND U2563 ( .A(n2444), .B(n2443), .Z(n2462) );
  XNOR U2564 ( .A(n2463), .B(n2462), .Z(n2464) );
  NANDN U2565 ( .A(n2446), .B(n2445), .Z(n2450) );
  NAND U2566 ( .A(n2448), .B(n2447), .Z(n2449) );
  NAND U2567 ( .A(n2450), .B(n2449), .Z(n2465) );
  XNOR U2568 ( .A(n2464), .B(n2465), .Z(n2456) );
  XNOR U2569 ( .A(n2457), .B(n2456), .Z(n2458) );
  XNOR U2570 ( .A(n2459), .B(n2458), .Z(n2492) );
  XNOR U2571 ( .A(sreg[311]), .B(n2492), .Z(n2494) );
  NANDN U2572 ( .A(sreg[310]), .B(n2451), .Z(n2455) );
  NAND U2573 ( .A(n2453), .B(n2452), .Z(n2454) );
  NAND U2574 ( .A(n2455), .B(n2454), .Z(n2493) );
  XNOR U2575 ( .A(n2494), .B(n2493), .Z(c[311]) );
  NANDN U2576 ( .A(n2457), .B(n2456), .Z(n2461) );
  NANDN U2577 ( .A(n2459), .B(n2458), .Z(n2460) );
  AND U2578 ( .A(n2461), .B(n2460), .Z(n2500) );
  NANDN U2579 ( .A(n2463), .B(n2462), .Z(n2467) );
  NANDN U2580 ( .A(n2465), .B(n2464), .Z(n2466) );
  AND U2581 ( .A(n2467), .B(n2466), .Z(n2498) );
  NAND U2582 ( .A(n26), .B(n2468), .Z(n2470) );
  XOR U2583 ( .A(b[7]), .B(a[58]), .Z(n2509) );
  NAND U2584 ( .A(n10531), .B(n2509), .Z(n2469) );
  AND U2585 ( .A(n2470), .B(n2469), .Z(n2528) );
  NAND U2586 ( .A(n23), .B(n2471), .Z(n2473) );
  XOR U2587 ( .A(b[3]), .B(a[62]), .Z(n2512) );
  NAND U2588 ( .A(n24), .B(n2512), .Z(n2472) );
  NAND U2589 ( .A(n2473), .B(n2472), .Z(n2527) );
  XNOR U2590 ( .A(n2528), .B(n2527), .Z(n2530) );
  NAND U2591 ( .A(n25), .B(n2474), .Z(n2476) );
  XOR U2592 ( .A(b[5]), .B(a[60]), .Z(n2518) );
  NAND U2593 ( .A(n10456), .B(n2518), .Z(n2475) );
  AND U2594 ( .A(n2476), .B(n2475), .Z(n2522) );
  AND U2595 ( .A(b[7]), .B(a[56]), .Z(n2521) );
  XNOR U2596 ( .A(n2522), .B(n2521), .Z(n2523) );
  NAND U2597 ( .A(b[0]), .B(a[64]), .Z(n2477) );
  XNOR U2598 ( .A(b[1]), .B(n2477), .Z(n2479) );
  NANDN U2599 ( .A(b[0]), .B(a[63]), .Z(n2478) );
  NAND U2600 ( .A(n2479), .B(n2478), .Z(n2524) );
  XNOR U2601 ( .A(n2523), .B(n2524), .Z(n2529) );
  XOR U2602 ( .A(n2530), .B(n2529), .Z(n2504) );
  NANDN U2603 ( .A(n2481), .B(n2480), .Z(n2485) );
  NANDN U2604 ( .A(n2483), .B(n2482), .Z(n2484) );
  AND U2605 ( .A(n2485), .B(n2484), .Z(n2503) );
  XNOR U2606 ( .A(n2504), .B(n2503), .Z(n2505) );
  NANDN U2607 ( .A(n2487), .B(n2486), .Z(n2491) );
  NAND U2608 ( .A(n2489), .B(n2488), .Z(n2490) );
  NAND U2609 ( .A(n2491), .B(n2490), .Z(n2506) );
  XNOR U2610 ( .A(n2505), .B(n2506), .Z(n2497) );
  XNOR U2611 ( .A(n2498), .B(n2497), .Z(n2499) );
  XNOR U2612 ( .A(n2500), .B(n2499), .Z(n2533) );
  XNOR U2613 ( .A(sreg[312]), .B(n2533), .Z(n2535) );
  NANDN U2614 ( .A(sreg[311]), .B(n2492), .Z(n2496) );
  NAND U2615 ( .A(n2494), .B(n2493), .Z(n2495) );
  NAND U2616 ( .A(n2496), .B(n2495), .Z(n2534) );
  XNOR U2617 ( .A(n2535), .B(n2534), .Z(c[312]) );
  NANDN U2618 ( .A(n2498), .B(n2497), .Z(n2502) );
  NANDN U2619 ( .A(n2500), .B(n2499), .Z(n2501) );
  AND U2620 ( .A(n2502), .B(n2501), .Z(n2541) );
  NANDN U2621 ( .A(n2504), .B(n2503), .Z(n2508) );
  NANDN U2622 ( .A(n2506), .B(n2505), .Z(n2507) );
  AND U2623 ( .A(n2508), .B(n2507), .Z(n2539) );
  NAND U2624 ( .A(n26), .B(n2509), .Z(n2511) );
  XOR U2625 ( .A(b[7]), .B(a[59]), .Z(n2550) );
  NAND U2626 ( .A(n10531), .B(n2550), .Z(n2510) );
  AND U2627 ( .A(n2511), .B(n2510), .Z(n2569) );
  NAND U2628 ( .A(n23), .B(n2512), .Z(n2514) );
  XOR U2629 ( .A(b[3]), .B(a[63]), .Z(n2553) );
  NAND U2630 ( .A(n24), .B(n2553), .Z(n2513) );
  NAND U2631 ( .A(n2514), .B(n2513), .Z(n2568) );
  XNOR U2632 ( .A(n2569), .B(n2568), .Z(n2571) );
  NAND U2633 ( .A(b[0]), .B(a[65]), .Z(n2515) );
  XNOR U2634 ( .A(b[1]), .B(n2515), .Z(n2517) );
  NANDN U2635 ( .A(b[0]), .B(a[64]), .Z(n2516) );
  NAND U2636 ( .A(n2517), .B(n2516), .Z(n2565) );
  NAND U2637 ( .A(n25), .B(n2518), .Z(n2520) );
  XOR U2638 ( .A(b[5]), .B(a[61]), .Z(n2559) );
  NAND U2639 ( .A(n10456), .B(n2559), .Z(n2519) );
  AND U2640 ( .A(n2520), .B(n2519), .Z(n2563) );
  AND U2641 ( .A(b[7]), .B(a[57]), .Z(n2562) );
  XNOR U2642 ( .A(n2563), .B(n2562), .Z(n2564) );
  XNOR U2643 ( .A(n2565), .B(n2564), .Z(n2570) );
  XOR U2644 ( .A(n2571), .B(n2570), .Z(n2545) );
  NANDN U2645 ( .A(n2522), .B(n2521), .Z(n2526) );
  NANDN U2646 ( .A(n2524), .B(n2523), .Z(n2525) );
  AND U2647 ( .A(n2526), .B(n2525), .Z(n2544) );
  XNOR U2648 ( .A(n2545), .B(n2544), .Z(n2546) );
  NANDN U2649 ( .A(n2528), .B(n2527), .Z(n2532) );
  NAND U2650 ( .A(n2530), .B(n2529), .Z(n2531) );
  NAND U2651 ( .A(n2532), .B(n2531), .Z(n2547) );
  XNOR U2652 ( .A(n2546), .B(n2547), .Z(n2538) );
  XNOR U2653 ( .A(n2539), .B(n2538), .Z(n2540) );
  XNOR U2654 ( .A(n2541), .B(n2540), .Z(n2574) );
  XNOR U2655 ( .A(sreg[313]), .B(n2574), .Z(n2576) );
  NANDN U2656 ( .A(sreg[312]), .B(n2533), .Z(n2537) );
  NAND U2657 ( .A(n2535), .B(n2534), .Z(n2536) );
  NAND U2658 ( .A(n2537), .B(n2536), .Z(n2575) );
  XNOR U2659 ( .A(n2576), .B(n2575), .Z(c[313]) );
  NANDN U2660 ( .A(n2539), .B(n2538), .Z(n2543) );
  NANDN U2661 ( .A(n2541), .B(n2540), .Z(n2542) );
  AND U2662 ( .A(n2543), .B(n2542), .Z(n2582) );
  NANDN U2663 ( .A(n2545), .B(n2544), .Z(n2549) );
  NANDN U2664 ( .A(n2547), .B(n2546), .Z(n2548) );
  AND U2665 ( .A(n2549), .B(n2548), .Z(n2580) );
  NAND U2666 ( .A(n26), .B(n2550), .Z(n2552) );
  XOR U2667 ( .A(b[7]), .B(a[60]), .Z(n2591) );
  NAND U2668 ( .A(n10531), .B(n2591), .Z(n2551) );
  AND U2669 ( .A(n2552), .B(n2551), .Z(n2610) );
  NAND U2670 ( .A(n23), .B(n2553), .Z(n2555) );
  XOR U2671 ( .A(b[3]), .B(a[64]), .Z(n2594) );
  NAND U2672 ( .A(n24), .B(n2594), .Z(n2554) );
  NAND U2673 ( .A(n2555), .B(n2554), .Z(n2609) );
  XNOR U2674 ( .A(n2610), .B(n2609), .Z(n2612) );
  NAND U2675 ( .A(b[0]), .B(a[66]), .Z(n2556) );
  XNOR U2676 ( .A(b[1]), .B(n2556), .Z(n2558) );
  NANDN U2677 ( .A(b[0]), .B(a[65]), .Z(n2557) );
  NAND U2678 ( .A(n2558), .B(n2557), .Z(n2606) );
  NAND U2679 ( .A(n25), .B(n2559), .Z(n2561) );
  XOR U2680 ( .A(b[5]), .B(a[62]), .Z(n2597) );
  NAND U2681 ( .A(n10456), .B(n2597), .Z(n2560) );
  AND U2682 ( .A(n2561), .B(n2560), .Z(n2604) );
  AND U2683 ( .A(b[7]), .B(a[58]), .Z(n2603) );
  XNOR U2684 ( .A(n2604), .B(n2603), .Z(n2605) );
  XNOR U2685 ( .A(n2606), .B(n2605), .Z(n2611) );
  XOR U2686 ( .A(n2612), .B(n2611), .Z(n2586) );
  NANDN U2687 ( .A(n2563), .B(n2562), .Z(n2567) );
  NANDN U2688 ( .A(n2565), .B(n2564), .Z(n2566) );
  AND U2689 ( .A(n2567), .B(n2566), .Z(n2585) );
  XNOR U2690 ( .A(n2586), .B(n2585), .Z(n2587) );
  NANDN U2691 ( .A(n2569), .B(n2568), .Z(n2573) );
  NAND U2692 ( .A(n2571), .B(n2570), .Z(n2572) );
  NAND U2693 ( .A(n2573), .B(n2572), .Z(n2588) );
  XNOR U2694 ( .A(n2587), .B(n2588), .Z(n2579) );
  XNOR U2695 ( .A(n2580), .B(n2579), .Z(n2581) );
  XNOR U2696 ( .A(n2582), .B(n2581), .Z(n2615) );
  XNOR U2697 ( .A(sreg[314]), .B(n2615), .Z(n2617) );
  NANDN U2698 ( .A(sreg[313]), .B(n2574), .Z(n2578) );
  NAND U2699 ( .A(n2576), .B(n2575), .Z(n2577) );
  NAND U2700 ( .A(n2578), .B(n2577), .Z(n2616) );
  XNOR U2701 ( .A(n2617), .B(n2616), .Z(c[314]) );
  NANDN U2702 ( .A(n2580), .B(n2579), .Z(n2584) );
  NANDN U2703 ( .A(n2582), .B(n2581), .Z(n2583) );
  AND U2704 ( .A(n2584), .B(n2583), .Z(n2623) );
  NANDN U2705 ( .A(n2586), .B(n2585), .Z(n2590) );
  NANDN U2706 ( .A(n2588), .B(n2587), .Z(n2589) );
  AND U2707 ( .A(n2590), .B(n2589), .Z(n2621) );
  NAND U2708 ( .A(n26), .B(n2591), .Z(n2593) );
  XOR U2709 ( .A(b[7]), .B(a[61]), .Z(n2632) );
  NAND U2710 ( .A(n10531), .B(n2632), .Z(n2592) );
  AND U2711 ( .A(n2593), .B(n2592), .Z(n2651) );
  NAND U2712 ( .A(n23), .B(n2594), .Z(n2596) );
  XOR U2713 ( .A(b[3]), .B(a[65]), .Z(n2635) );
  NAND U2714 ( .A(n24), .B(n2635), .Z(n2595) );
  NAND U2715 ( .A(n2596), .B(n2595), .Z(n2650) );
  XNOR U2716 ( .A(n2651), .B(n2650), .Z(n2653) );
  NAND U2717 ( .A(n25), .B(n2597), .Z(n2599) );
  XOR U2718 ( .A(b[5]), .B(a[63]), .Z(n2641) );
  NAND U2719 ( .A(n10456), .B(n2641), .Z(n2598) );
  AND U2720 ( .A(n2599), .B(n2598), .Z(n2645) );
  AND U2721 ( .A(b[7]), .B(a[59]), .Z(n2644) );
  XNOR U2722 ( .A(n2645), .B(n2644), .Z(n2646) );
  NAND U2723 ( .A(b[0]), .B(a[67]), .Z(n2600) );
  XNOR U2724 ( .A(b[1]), .B(n2600), .Z(n2602) );
  NANDN U2725 ( .A(b[0]), .B(a[66]), .Z(n2601) );
  NAND U2726 ( .A(n2602), .B(n2601), .Z(n2647) );
  XNOR U2727 ( .A(n2646), .B(n2647), .Z(n2652) );
  XOR U2728 ( .A(n2653), .B(n2652), .Z(n2627) );
  NANDN U2729 ( .A(n2604), .B(n2603), .Z(n2608) );
  NANDN U2730 ( .A(n2606), .B(n2605), .Z(n2607) );
  AND U2731 ( .A(n2608), .B(n2607), .Z(n2626) );
  XNOR U2732 ( .A(n2627), .B(n2626), .Z(n2628) );
  NANDN U2733 ( .A(n2610), .B(n2609), .Z(n2614) );
  NAND U2734 ( .A(n2612), .B(n2611), .Z(n2613) );
  NAND U2735 ( .A(n2614), .B(n2613), .Z(n2629) );
  XNOR U2736 ( .A(n2628), .B(n2629), .Z(n2620) );
  XNOR U2737 ( .A(n2621), .B(n2620), .Z(n2622) );
  XNOR U2738 ( .A(n2623), .B(n2622), .Z(n2656) );
  XNOR U2739 ( .A(sreg[315]), .B(n2656), .Z(n2658) );
  NANDN U2740 ( .A(sreg[314]), .B(n2615), .Z(n2619) );
  NAND U2741 ( .A(n2617), .B(n2616), .Z(n2618) );
  NAND U2742 ( .A(n2619), .B(n2618), .Z(n2657) );
  XNOR U2743 ( .A(n2658), .B(n2657), .Z(c[315]) );
  NANDN U2744 ( .A(n2621), .B(n2620), .Z(n2625) );
  NANDN U2745 ( .A(n2623), .B(n2622), .Z(n2624) );
  AND U2746 ( .A(n2625), .B(n2624), .Z(n2664) );
  NANDN U2747 ( .A(n2627), .B(n2626), .Z(n2631) );
  NANDN U2748 ( .A(n2629), .B(n2628), .Z(n2630) );
  AND U2749 ( .A(n2631), .B(n2630), .Z(n2662) );
  NAND U2750 ( .A(n26), .B(n2632), .Z(n2634) );
  XOR U2751 ( .A(b[7]), .B(a[62]), .Z(n2673) );
  NAND U2752 ( .A(n10531), .B(n2673), .Z(n2633) );
  AND U2753 ( .A(n2634), .B(n2633), .Z(n2692) );
  NAND U2754 ( .A(n23), .B(n2635), .Z(n2637) );
  XOR U2755 ( .A(b[3]), .B(a[66]), .Z(n2676) );
  NAND U2756 ( .A(n24), .B(n2676), .Z(n2636) );
  NAND U2757 ( .A(n2637), .B(n2636), .Z(n2691) );
  XNOR U2758 ( .A(n2692), .B(n2691), .Z(n2694) );
  NAND U2759 ( .A(b[0]), .B(a[68]), .Z(n2638) );
  XNOR U2760 ( .A(b[1]), .B(n2638), .Z(n2640) );
  NANDN U2761 ( .A(b[0]), .B(a[67]), .Z(n2639) );
  NAND U2762 ( .A(n2640), .B(n2639), .Z(n2688) );
  NAND U2763 ( .A(n25), .B(n2641), .Z(n2643) );
  XOR U2764 ( .A(b[5]), .B(a[64]), .Z(n2682) );
  NAND U2765 ( .A(n10456), .B(n2682), .Z(n2642) );
  AND U2766 ( .A(n2643), .B(n2642), .Z(n2686) );
  AND U2767 ( .A(b[7]), .B(a[60]), .Z(n2685) );
  XNOR U2768 ( .A(n2686), .B(n2685), .Z(n2687) );
  XNOR U2769 ( .A(n2688), .B(n2687), .Z(n2693) );
  XOR U2770 ( .A(n2694), .B(n2693), .Z(n2668) );
  NANDN U2771 ( .A(n2645), .B(n2644), .Z(n2649) );
  NANDN U2772 ( .A(n2647), .B(n2646), .Z(n2648) );
  AND U2773 ( .A(n2649), .B(n2648), .Z(n2667) );
  XNOR U2774 ( .A(n2668), .B(n2667), .Z(n2669) );
  NANDN U2775 ( .A(n2651), .B(n2650), .Z(n2655) );
  NAND U2776 ( .A(n2653), .B(n2652), .Z(n2654) );
  NAND U2777 ( .A(n2655), .B(n2654), .Z(n2670) );
  XNOR U2778 ( .A(n2669), .B(n2670), .Z(n2661) );
  XNOR U2779 ( .A(n2662), .B(n2661), .Z(n2663) );
  XNOR U2780 ( .A(n2664), .B(n2663), .Z(n2697) );
  XNOR U2781 ( .A(sreg[316]), .B(n2697), .Z(n2699) );
  NANDN U2782 ( .A(sreg[315]), .B(n2656), .Z(n2660) );
  NAND U2783 ( .A(n2658), .B(n2657), .Z(n2659) );
  NAND U2784 ( .A(n2660), .B(n2659), .Z(n2698) );
  XNOR U2785 ( .A(n2699), .B(n2698), .Z(c[316]) );
  NANDN U2786 ( .A(n2662), .B(n2661), .Z(n2666) );
  NANDN U2787 ( .A(n2664), .B(n2663), .Z(n2665) );
  AND U2788 ( .A(n2666), .B(n2665), .Z(n2709) );
  NANDN U2789 ( .A(n2668), .B(n2667), .Z(n2672) );
  NANDN U2790 ( .A(n2670), .B(n2669), .Z(n2671) );
  AND U2791 ( .A(n2672), .B(n2671), .Z(n2708) );
  NAND U2792 ( .A(n26), .B(n2673), .Z(n2675) );
  XOR U2793 ( .A(b[7]), .B(a[63]), .Z(n2719) );
  NAND U2794 ( .A(n10531), .B(n2719), .Z(n2674) );
  AND U2795 ( .A(n2675), .B(n2674), .Z(n2738) );
  NAND U2796 ( .A(n23), .B(n2676), .Z(n2678) );
  XOR U2797 ( .A(b[3]), .B(a[67]), .Z(n2722) );
  NAND U2798 ( .A(n24), .B(n2722), .Z(n2677) );
  NAND U2799 ( .A(n2678), .B(n2677), .Z(n2737) );
  XNOR U2800 ( .A(n2738), .B(n2737), .Z(n2740) );
  NAND U2801 ( .A(b[0]), .B(a[69]), .Z(n2679) );
  XNOR U2802 ( .A(b[1]), .B(n2679), .Z(n2681) );
  NANDN U2803 ( .A(b[0]), .B(a[68]), .Z(n2680) );
  NAND U2804 ( .A(n2681), .B(n2680), .Z(n2734) );
  NAND U2805 ( .A(n25), .B(n2682), .Z(n2684) );
  XOR U2806 ( .A(b[5]), .B(a[65]), .Z(n2725) );
  NAND U2807 ( .A(n10456), .B(n2725), .Z(n2683) );
  AND U2808 ( .A(n2684), .B(n2683), .Z(n2732) );
  AND U2809 ( .A(b[7]), .B(a[61]), .Z(n2731) );
  XNOR U2810 ( .A(n2732), .B(n2731), .Z(n2733) );
  XNOR U2811 ( .A(n2734), .B(n2733), .Z(n2739) );
  XOR U2812 ( .A(n2740), .B(n2739), .Z(n2714) );
  NANDN U2813 ( .A(n2686), .B(n2685), .Z(n2690) );
  NANDN U2814 ( .A(n2688), .B(n2687), .Z(n2689) );
  AND U2815 ( .A(n2690), .B(n2689), .Z(n2713) );
  XNOR U2816 ( .A(n2714), .B(n2713), .Z(n2715) );
  NANDN U2817 ( .A(n2692), .B(n2691), .Z(n2696) );
  NAND U2818 ( .A(n2694), .B(n2693), .Z(n2695) );
  NAND U2819 ( .A(n2696), .B(n2695), .Z(n2716) );
  XNOR U2820 ( .A(n2715), .B(n2716), .Z(n2707) );
  XOR U2821 ( .A(n2708), .B(n2707), .Z(n2710) );
  XOR U2822 ( .A(n2709), .B(n2710), .Z(n2702) );
  XNOR U2823 ( .A(n2702), .B(sreg[317]), .Z(n2704) );
  NANDN U2824 ( .A(sreg[316]), .B(n2697), .Z(n2701) );
  NAND U2825 ( .A(n2699), .B(n2698), .Z(n2700) );
  AND U2826 ( .A(n2701), .B(n2700), .Z(n2703) );
  XOR U2827 ( .A(n2704), .B(n2703), .Z(c[317]) );
  NANDN U2828 ( .A(n2702), .B(sreg[317]), .Z(n2706) );
  NAND U2829 ( .A(n2704), .B(n2703), .Z(n2705) );
  AND U2830 ( .A(n2706), .B(n2705), .Z(n2781) );
  NANDN U2831 ( .A(n2708), .B(n2707), .Z(n2712) );
  OR U2832 ( .A(n2710), .B(n2709), .Z(n2711) );
  AND U2833 ( .A(n2712), .B(n2711), .Z(n2746) );
  NANDN U2834 ( .A(n2714), .B(n2713), .Z(n2718) );
  NANDN U2835 ( .A(n2716), .B(n2715), .Z(n2717) );
  AND U2836 ( .A(n2718), .B(n2717), .Z(n2744) );
  NAND U2837 ( .A(n26), .B(n2719), .Z(n2721) );
  XOR U2838 ( .A(b[7]), .B(a[64]), .Z(n2755) );
  NAND U2839 ( .A(n10531), .B(n2755), .Z(n2720) );
  AND U2840 ( .A(n2721), .B(n2720), .Z(n2774) );
  NAND U2841 ( .A(n23), .B(n2722), .Z(n2724) );
  XOR U2842 ( .A(b[3]), .B(a[68]), .Z(n2758) );
  NAND U2843 ( .A(n24), .B(n2758), .Z(n2723) );
  NAND U2844 ( .A(n2724), .B(n2723), .Z(n2773) );
  XNOR U2845 ( .A(n2774), .B(n2773), .Z(n2776) );
  NAND U2846 ( .A(n25), .B(n2725), .Z(n2727) );
  XOR U2847 ( .A(b[5]), .B(a[66]), .Z(n2764) );
  NAND U2848 ( .A(n10456), .B(n2764), .Z(n2726) );
  AND U2849 ( .A(n2727), .B(n2726), .Z(n2768) );
  AND U2850 ( .A(b[7]), .B(a[62]), .Z(n2767) );
  XNOR U2851 ( .A(n2768), .B(n2767), .Z(n2769) );
  NAND U2852 ( .A(b[0]), .B(a[70]), .Z(n2728) );
  XNOR U2853 ( .A(b[1]), .B(n2728), .Z(n2730) );
  NANDN U2854 ( .A(b[0]), .B(a[69]), .Z(n2729) );
  NAND U2855 ( .A(n2730), .B(n2729), .Z(n2770) );
  XNOR U2856 ( .A(n2769), .B(n2770), .Z(n2775) );
  XOR U2857 ( .A(n2776), .B(n2775), .Z(n2750) );
  NANDN U2858 ( .A(n2732), .B(n2731), .Z(n2736) );
  NANDN U2859 ( .A(n2734), .B(n2733), .Z(n2735) );
  AND U2860 ( .A(n2736), .B(n2735), .Z(n2749) );
  XNOR U2861 ( .A(n2750), .B(n2749), .Z(n2751) );
  NANDN U2862 ( .A(n2738), .B(n2737), .Z(n2742) );
  NAND U2863 ( .A(n2740), .B(n2739), .Z(n2741) );
  NAND U2864 ( .A(n2742), .B(n2741), .Z(n2752) );
  XNOR U2865 ( .A(n2751), .B(n2752), .Z(n2743) );
  XNOR U2866 ( .A(n2744), .B(n2743), .Z(n2745) );
  XNOR U2867 ( .A(n2746), .B(n2745), .Z(n2779) );
  XNOR U2868 ( .A(sreg[318]), .B(n2779), .Z(n2780) );
  XNOR U2869 ( .A(n2781), .B(n2780), .Z(c[318]) );
  NANDN U2870 ( .A(n2744), .B(n2743), .Z(n2748) );
  NANDN U2871 ( .A(n2746), .B(n2745), .Z(n2747) );
  AND U2872 ( .A(n2748), .B(n2747), .Z(n2787) );
  NANDN U2873 ( .A(n2750), .B(n2749), .Z(n2754) );
  NANDN U2874 ( .A(n2752), .B(n2751), .Z(n2753) );
  AND U2875 ( .A(n2754), .B(n2753), .Z(n2785) );
  NAND U2876 ( .A(n26), .B(n2755), .Z(n2757) );
  XOR U2877 ( .A(b[7]), .B(a[65]), .Z(n2796) );
  NAND U2878 ( .A(n10531), .B(n2796), .Z(n2756) );
  AND U2879 ( .A(n2757), .B(n2756), .Z(n2815) );
  NAND U2880 ( .A(n23), .B(n2758), .Z(n2760) );
  XOR U2881 ( .A(b[3]), .B(a[69]), .Z(n2799) );
  NAND U2882 ( .A(n24), .B(n2799), .Z(n2759) );
  NAND U2883 ( .A(n2760), .B(n2759), .Z(n2814) );
  XNOR U2884 ( .A(n2815), .B(n2814), .Z(n2817) );
  NAND U2885 ( .A(b[0]), .B(a[71]), .Z(n2761) );
  XNOR U2886 ( .A(b[1]), .B(n2761), .Z(n2763) );
  NANDN U2887 ( .A(b[0]), .B(a[70]), .Z(n2762) );
  NAND U2888 ( .A(n2763), .B(n2762), .Z(n2811) );
  NAND U2889 ( .A(n25), .B(n2764), .Z(n2766) );
  XOR U2890 ( .A(b[5]), .B(a[67]), .Z(n2802) );
  NAND U2891 ( .A(n10456), .B(n2802), .Z(n2765) );
  AND U2892 ( .A(n2766), .B(n2765), .Z(n2809) );
  AND U2893 ( .A(b[7]), .B(a[63]), .Z(n2808) );
  XNOR U2894 ( .A(n2809), .B(n2808), .Z(n2810) );
  XNOR U2895 ( .A(n2811), .B(n2810), .Z(n2816) );
  XOR U2896 ( .A(n2817), .B(n2816), .Z(n2791) );
  NANDN U2897 ( .A(n2768), .B(n2767), .Z(n2772) );
  NANDN U2898 ( .A(n2770), .B(n2769), .Z(n2771) );
  AND U2899 ( .A(n2772), .B(n2771), .Z(n2790) );
  XNOR U2900 ( .A(n2791), .B(n2790), .Z(n2792) );
  NANDN U2901 ( .A(n2774), .B(n2773), .Z(n2778) );
  NAND U2902 ( .A(n2776), .B(n2775), .Z(n2777) );
  NAND U2903 ( .A(n2778), .B(n2777), .Z(n2793) );
  XNOR U2904 ( .A(n2792), .B(n2793), .Z(n2784) );
  XNOR U2905 ( .A(n2785), .B(n2784), .Z(n2786) );
  XNOR U2906 ( .A(n2787), .B(n2786), .Z(n2820) );
  XNOR U2907 ( .A(sreg[319]), .B(n2820), .Z(n2822) );
  NANDN U2908 ( .A(sreg[318]), .B(n2779), .Z(n2783) );
  NAND U2909 ( .A(n2781), .B(n2780), .Z(n2782) );
  NAND U2910 ( .A(n2783), .B(n2782), .Z(n2821) );
  XNOR U2911 ( .A(n2822), .B(n2821), .Z(c[319]) );
  NANDN U2912 ( .A(n2785), .B(n2784), .Z(n2789) );
  NANDN U2913 ( .A(n2787), .B(n2786), .Z(n2788) );
  AND U2914 ( .A(n2789), .B(n2788), .Z(n2828) );
  NANDN U2915 ( .A(n2791), .B(n2790), .Z(n2795) );
  NANDN U2916 ( .A(n2793), .B(n2792), .Z(n2794) );
  AND U2917 ( .A(n2795), .B(n2794), .Z(n2826) );
  NAND U2918 ( .A(n26), .B(n2796), .Z(n2798) );
  XOR U2919 ( .A(b[7]), .B(a[66]), .Z(n2837) );
  NAND U2920 ( .A(n10531), .B(n2837), .Z(n2797) );
  AND U2921 ( .A(n2798), .B(n2797), .Z(n2856) );
  NAND U2922 ( .A(n23), .B(n2799), .Z(n2801) );
  XOR U2923 ( .A(b[3]), .B(a[70]), .Z(n2840) );
  NAND U2924 ( .A(n24), .B(n2840), .Z(n2800) );
  NAND U2925 ( .A(n2801), .B(n2800), .Z(n2855) );
  XNOR U2926 ( .A(n2856), .B(n2855), .Z(n2858) );
  NAND U2927 ( .A(n25), .B(n2802), .Z(n2804) );
  XOR U2928 ( .A(b[5]), .B(a[68]), .Z(n2846) );
  NAND U2929 ( .A(n10456), .B(n2846), .Z(n2803) );
  AND U2930 ( .A(n2804), .B(n2803), .Z(n2850) );
  AND U2931 ( .A(b[7]), .B(a[64]), .Z(n2849) );
  XNOR U2932 ( .A(n2850), .B(n2849), .Z(n2851) );
  NAND U2933 ( .A(b[0]), .B(a[72]), .Z(n2805) );
  XNOR U2934 ( .A(b[1]), .B(n2805), .Z(n2807) );
  NANDN U2935 ( .A(b[0]), .B(a[71]), .Z(n2806) );
  NAND U2936 ( .A(n2807), .B(n2806), .Z(n2852) );
  XNOR U2937 ( .A(n2851), .B(n2852), .Z(n2857) );
  XOR U2938 ( .A(n2858), .B(n2857), .Z(n2832) );
  NANDN U2939 ( .A(n2809), .B(n2808), .Z(n2813) );
  NANDN U2940 ( .A(n2811), .B(n2810), .Z(n2812) );
  AND U2941 ( .A(n2813), .B(n2812), .Z(n2831) );
  XNOR U2942 ( .A(n2832), .B(n2831), .Z(n2833) );
  NANDN U2943 ( .A(n2815), .B(n2814), .Z(n2819) );
  NAND U2944 ( .A(n2817), .B(n2816), .Z(n2818) );
  NAND U2945 ( .A(n2819), .B(n2818), .Z(n2834) );
  XNOR U2946 ( .A(n2833), .B(n2834), .Z(n2825) );
  XNOR U2947 ( .A(n2826), .B(n2825), .Z(n2827) );
  XNOR U2948 ( .A(n2828), .B(n2827), .Z(n2861) );
  XNOR U2949 ( .A(sreg[320]), .B(n2861), .Z(n2863) );
  NANDN U2950 ( .A(sreg[319]), .B(n2820), .Z(n2824) );
  NAND U2951 ( .A(n2822), .B(n2821), .Z(n2823) );
  NAND U2952 ( .A(n2824), .B(n2823), .Z(n2862) );
  XNOR U2953 ( .A(n2863), .B(n2862), .Z(c[320]) );
  NANDN U2954 ( .A(n2826), .B(n2825), .Z(n2830) );
  NANDN U2955 ( .A(n2828), .B(n2827), .Z(n2829) );
  AND U2956 ( .A(n2830), .B(n2829), .Z(n2869) );
  NANDN U2957 ( .A(n2832), .B(n2831), .Z(n2836) );
  NANDN U2958 ( .A(n2834), .B(n2833), .Z(n2835) );
  AND U2959 ( .A(n2836), .B(n2835), .Z(n2867) );
  NAND U2960 ( .A(n26), .B(n2837), .Z(n2839) );
  XOR U2961 ( .A(b[7]), .B(a[67]), .Z(n2878) );
  NAND U2962 ( .A(n10531), .B(n2878), .Z(n2838) );
  AND U2963 ( .A(n2839), .B(n2838), .Z(n2897) );
  NAND U2964 ( .A(n23), .B(n2840), .Z(n2842) );
  XOR U2965 ( .A(b[3]), .B(a[71]), .Z(n2881) );
  NAND U2966 ( .A(n24), .B(n2881), .Z(n2841) );
  NAND U2967 ( .A(n2842), .B(n2841), .Z(n2896) );
  XNOR U2968 ( .A(n2897), .B(n2896), .Z(n2899) );
  NAND U2969 ( .A(b[0]), .B(a[73]), .Z(n2843) );
  XNOR U2970 ( .A(b[1]), .B(n2843), .Z(n2845) );
  NANDN U2971 ( .A(b[0]), .B(a[72]), .Z(n2844) );
  NAND U2972 ( .A(n2845), .B(n2844), .Z(n2893) );
  NAND U2973 ( .A(n25), .B(n2846), .Z(n2848) );
  XOR U2974 ( .A(b[5]), .B(a[69]), .Z(n2887) );
  NAND U2975 ( .A(n10456), .B(n2887), .Z(n2847) );
  AND U2976 ( .A(n2848), .B(n2847), .Z(n2891) );
  AND U2977 ( .A(b[7]), .B(a[65]), .Z(n2890) );
  XNOR U2978 ( .A(n2891), .B(n2890), .Z(n2892) );
  XNOR U2979 ( .A(n2893), .B(n2892), .Z(n2898) );
  XOR U2980 ( .A(n2899), .B(n2898), .Z(n2873) );
  NANDN U2981 ( .A(n2850), .B(n2849), .Z(n2854) );
  NANDN U2982 ( .A(n2852), .B(n2851), .Z(n2853) );
  AND U2983 ( .A(n2854), .B(n2853), .Z(n2872) );
  XNOR U2984 ( .A(n2873), .B(n2872), .Z(n2874) );
  NANDN U2985 ( .A(n2856), .B(n2855), .Z(n2860) );
  NAND U2986 ( .A(n2858), .B(n2857), .Z(n2859) );
  NAND U2987 ( .A(n2860), .B(n2859), .Z(n2875) );
  XNOR U2988 ( .A(n2874), .B(n2875), .Z(n2866) );
  XNOR U2989 ( .A(n2867), .B(n2866), .Z(n2868) );
  XNOR U2990 ( .A(n2869), .B(n2868), .Z(n2902) );
  XNOR U2991 ( .A(sreg[321]), .B(n2902), .Z(n2904) );
  NANDN U2992 ( .A(sreg[320]), .B(n2861), .Z(n2865) );
  NAND U2993 ( .A(n2863), .B(n2862), .Z(n2864) );
  NAND U2994 ( .A(n2865), .B(n2864), .Z(n2903) );
  XNOR U2995 ( .A(n2904), .B(n2903), .Z(c[321]) );
  NANDN U2996 ( .A(n2867), .B(n2866), .Z(n2871) );
  NANDN U2997 ( .A(n2869), .B(n2868), .Z(n2870) );
  AND U2998 ( .A(n2871), .B(n2870), .Z(n2910) );
  NANDN U2999 ( .A(n2873), .B(n2872), .Z(n2877) );
  NANDN U3000 ( .A(n2875), .B(n2874), .Z(n2876) );
  AND U3001 ( .A(n2877), .B(n2876), .Z(n2908) );
  NAND U3002 ( .A(n26), .B(n2878), .Z(n2880) );
  XOR U3003 ( .A(b[7]), .B(a[68]), .Z(n2919) );
  NAND U3004 ( .A(n10531), .B(n2919), .Z(n2879) );
  AND U3005 ( .A(n2880), .B(n2879), .Z(n2938) );
  NAND U3006 ( .A(n23), .B(n2881), .Z(n2883) );
  XOR U3007 ( .A(b[3]), .B(a[72]), .Z(n2922) );
  NAND U3008 ( .A(n24), .B(n2922), .Z(n2882) );
  NAND U3009 ( .A(n2883), .B(n2882), .Z(n2937) );
  XNOR U3010 ( .A(n2938), .B(n2937), .Z(n2940) );
  NAND U3011 ( .A(b[0]), .B(a[74]), .Z(n2884) );
  XNOR U3012 ( .A(b[1]), .B(n2884), .Z(n2886) );
  NANDN U3013 ( .A(b[0]), .B(a[73]), .Z(n2885) );
  NAND U3014 ( .A(n2886), .B(n2885), .Z(n2934) );
  NAND U3015 ( .A(n25), .B(n2887), .Z(n2889) );
  XOR U3016 ( .A(b[5]), .B(a[70]), .Z(n2928) );
  NAND U3017 ( .A(n10456), .B(n2928), .Z(n2888) );
  AND U3018 ( .A(n2889), .B(n2888), .Z(n2932) );
  AND U3019 ( .A(b[7]), .B(a[66]), .Z(n2931) );
  XNOR U3020 ( .A(n2932), .B(n2931), .Z(n2933) );
  XNOR U3021 ( .A(n2934), .B(n2933), .Z(n2939) );
  XOR U3022 ( .A(n2940), .B(n2939), .Z(n2914) );
  NANDN U3023 ( .A(n2891), .B(n2890), .Z(n2895) );
  NANDN U3024 ( .A(n2893), .B(n2892), .Z(n2894) );
  AND U3025 ( .A(n2895), .B(n2894), .Z(n2913) );
  XNOR U3026 ( .A(n2914), .B(n2913), .Z(n2915) );
  NANDN U3027 ( .A(n2897), .B(n2896), .Z(n2901) );
  NAND U3028 ( .A(n2899), .B(n2898), .Z(n2900) );
  NAND U3029 ( .A(n2901), .B(n2900), .Z(n2916) );
  XNOR U3030 ( .A(n2915), .B(n2916), .Z(n2907) );
  XNOR U3031 ( .A(n2908), .B(n2907), .Z(n2909) );
  XNOR U3032 ( .A(n2910), .B(n2909), .Z(n2943) );
  XNOR U3033 ( .A(sreg[322]), .B(n2943), .Z(n2945) );
  NANDN U3034 ( .A(sreg[321]), .B(n2902), .Z(n2906) );
  NAND U3035 ( .A(n2904), .B(n2903), .Z(n2905) );
  NAND U3036 ( .A(n2906), .B(n2905), .Z(n2944) );
  XNOR U3037 ( .A(n2945), .B(n2944), .Z(c[322]) );
  NANDN U3038 ( .A(n2908), .B(n2907), .Z(n2912) );
  NANDN U3039 ( .A(n2910), .B(n2909), .Z(n2911) );
  AND U3040 ( .A(n2912), .B(n2911), .Z(n2951) );
  NANDN U3041 ( .A(n2914), .B(n2913), .Z(n2918) );
  NANDN U3042 ( .A(n2916), .B(n2915), .Z(n2917) );
  AND U3043 ( .A(n2918), .B(n2917), .Z(n2949) );
  NAND U3044 ( .A(n26), .B(n2919), .Z(n2921) );
  XOR U3045 ( .A(b[7]), .B(a[69]), .Z(n2960) );
  NAND U3046 ( .A(n10531), .B(n2960), .Z(n2920) );
  AND U3047 ( .A(n2921), .B(n2920), .Z(n2979) );
  NAND U3048 ( .A(n23), .B(n2922), .Z(n2924) );
  XOR U3049 ( .A(b[3]), .B(a[73]), .Z(n2963) );
  NAND U3050 ( .A(n24), .B(n2963), .Z(n2923) );
  NAND U3051 ( .A(n2924), .B(n2923), .Z(n2978) );
  XNOR U3052 ( .A(n2979), .B(n2978), .Z(n2981) );
  NAND U3053 ( .A(b[0]), .B(a[75]), .Z(n2925) );
  XNOR U3054 ( .A(b[1]), .B(n2925), .Z(n2927) );
  NANDN U3055 ( .A(b[0]), .B(a[74]), .Z(n2926) );
  NAND U3056 ( .A(n2927), .B(n2926), .Z(n2975) );
  NAND U3057 ( .A(n25), .B(n2928), .Z(n2930) );
  XOR U3058 ( .A(b[5]), .B(a[71]), .Z(n2969) );
  NAND U3059 ( .A(n10456), .B(n2969), .Z(n2929) );
  AND U3060 ( .A(n2930), .B(n2929), .Z(n2973) );
  AND U3061 ( .A(b[7]), .B(a[67]), .Z(n2972) );
  XNOR U3062 ( .A(n2973), .B(n2972), .Z(n2974) );
  XNOR U3063 ( .A(n2975), .B(n2974), .Z(n2980) );
  XOR U3064 ( .A(n2981), .B(n2980), .Z(n2955) );
  NANDN U3065 ( .A(n2932), .B(n2931), .Z(n2936) );
  NANDN U3066 ( .A(n2934), .B(n2933), .Z(n2935) );
  AND U3067 ( .A(n2936), .B(n2935), .Z(n2954) );
  XNOR U3068 ( .A(n2955), .B(n2954), .Z(n2956) );
  NANDN U3069 ( .A(n2938), .B(n2937), .Z(n2942) );
  NAND U3070 ( .A(n2940), .B(n2939), .Z(n2941) );
  NAND U3071 ( .A(n2942), .B(n2941), .Z(n2957) );
  XNOR U3072 ( .A(n2956), .B(n2957), .Z(n2948) );
  XNOR U3073 ( .A(n2949), .B(n2948), .Z(n2950) );
  XNOR U3074 ( .A(n2951), .B(n2950), .Z(n2984) );
  XNOR U3075 ( .A(sreg[323]), .B(n2984), .Z(n2986) );
  NANDN U3076 ( .A(sreg[322]), .B(n2943), .Z(n2947) );
  NAND U3077 ( .A(n2945), .B(n2944), .Z(n2946) );
  NAND U3078 ( .A(n2947), .B(n2946), .Z(n2985) );
  XNOR U3079 ( .A(n2986), .B(n2985), .Z(c[323]) );
  NANDN U3080 ( .A(n2949), .B(n2948), .Z(n2953) );
  NANDN U3081 ( .A(n2951), .B(n2950), .Z(n2952) );
  AND U3082 ( .A(n2953), .B(n2952), .Z(n2992) );
  NANDN U3083 ( .A(n2955), .B(n2954), .Z(n2959) );
  NANDN U3084 ( .A(n2957), .B(n2956), .Z(n2958) );
  AND U3085 ( .A(n2959), .B(n2958), .Z(n2990) );
  NAND U3086 ( .A(n26), .B(n2960), .Z(n2962) );
  XOR U3087 ( .A(b[7]), .B(a[70]), .Z(n3001) );
  NAND U3088 ( .A(n10531), .B(n3001), .Z(n2961) );
  AND U3089 ( .A(n2962), .B(n2961), .Z(n3020) );
  NAND U3090 ( .A(n23), .B(n2963), .Z(n2965) );
  XOR U3091 ( .A(b[3]), .B(a[74]), .Z(n3004) );
  NAND U3092 ( .A(n24), .B(n3004), .Z(n2964) );
  NAND U3093 ( .A(n2965), .B(n2964), .Z(n3019) );
  XNOR U3094 ( .A(n3020), .B(n3019), .Z(n3022) );
  NAND U3095 ( .A(b[0]), .B(a[76]), .Z(n2966) );
  XNOR U3096 ( .A(b[1]), .B(n2966), .Z(n2968) );
  NANDN U3097 ( .A(b[0]), .B(a[75]), .Z(n2967) );
  NAND U3098 ( .A(n2968), .B(n2967), .Z(n3016) );
  NAND U3099 ( .A(n25), .B(n2969), .Z(n2971) );
  XOR U3100 ( .A(b[5]), .B(a[72]), .Z(n3010) );
  NAND U3101 ( .A(n10456), .B(n3010), .Z(n2970) );
  AND U3102 ( .A(n2971), .B(n2970), .Z(n3014) );
  AND U3103 ( .A(b[7]), .B(a[68]), .Z(n3013) );
  XNOR U3104 ( .A(n3014), .B(n3013), .Z(n3015) );
  XNOR U3105 ( .A(n3016), .B(n3015), .Z(n3021) );
  XOR U3106 ( .A(n3022), .B(n3021), .Z(n2996) );
  NANDN U3107 ( .A(n2973), .B(n2972), .Z(n2977) );
  NANDN U3108 ( .A(n2975), .B(n2974), .Z(n2976) );
  AND U3109 ( .A(n2977), .B(n2976), .Z(n2995) );
  XNOR U3110 ( .A(n2996), .B(n2995), .Z(n2997) );
  NANDN U3111 ( .A(n2979), .B(n2978), .Z(n2983) );
  NAND U3112 ( .A(n2981), .B(n2980), .Z(n2982) );
  NAND U3113 ( .A(n2983), .B(n2982), .Z(n2998) );
  XNOR U3114 ( .A(n2997), .B(n2998), .Z(n2989) );
  XNOR U3115 ( .A(n2990), .B(n2989), .Z(n2991) );
  XNOR U3116 ( .A(n2992), .B(n2991), .Z(n3025) );
  XNOR U3117 ( .A(sreg[324]), .B(n3025), .Z(n3027) );
  NANDN U3118 ( .A(sreg[323]), .B(n2984), .Z(n2988) );
  NAND U3119 ( .A(n2986), .B(n2985), .Z(n2987) );
  NAND U3120 ( .A(n2988), .B(n2987), .Z(n3026) );
  XNOR U3121 ( .A(n3027), .B(n3026), .Z(c[324]) );
  NANDN U3122 ( .A(n2990), .B(n2989), .Z(n2994) );
  NANDN U3123 ( .A(n2992), .B(n2991), .Z(n2993) );
  AND U3124 ( .A(n2994), .B(n2993), .Z(n3033) );
  NANDN U3125 ( .A(n2996), .B(n2995), .Z(n3000) );
  NANDN U3126 ( .A(n2998), .B(n2997), .Z(n2999) );
  AND U3127 ( .A(n3000), .B(n2999), .Z(n3031) );
  NAND U3128 ( .A(n26), .B(n3001), .Z(n3003) );
  XOR U3129 ( .A(b[7]), .B(a[71]), .Z(n3042) );
  NAND U3130 ( .A(n10531), .B(n3042), .Z(n3002) );
  AND U3131 ( .A(n3003), .B(n3002), .Z(n3061) );
  NAND U3132 ( .A(n23), .B(n3004), .Z(n3006) );
  XOR U3133 ( .A(b[3]), .B(a[75]), .Z(n3045) );
  NAND U3134 ( .A(n24), .B(n3045), .Z(n3005) );
  NAND U3135 ( .A(n3006), .B(n3005), .Z(n3060) );
  XNOR U3136 ( .A(n3061), .B(n3060), .Z(n3063) );
  NAND U3137 ( .A(b[0]), .B(a[77]), .Z(n3007) );
  XNOR U3138 ( .A(b[1]), .B(n3007), .Z(n3009) );
  NANDN U3139 ( .A(b[0]), .B(a[76]), .Z(n3008) );
  NAND U3140 ( .A(n3009), .B(n3008), .Z(n3057) );
  NAND U3141 ( .A(n25), .B(n3010), .Z(n3012) );
  XOR U3142 ( .A(b[5]), .B(a[73]), .Z(n3051) );
  NAND U3143 ( .A(n10456), .B(n3051), .Z(n3011) );
  AND U3144 ( .A(n3012), .B(n3011), .Z(n3055) );
  AND U3145 ( .A(b[7]), .B(a[69]), .Z(n3054) );
  XNOR U3146 ( .A(n3055), .B(n3054), .Z(n3056) );
  XNOR U3147 ( .A(n3057), .B(n3056), .Z(n3062) );
  XOR U3148 ( .A(n3063), .B(n3062), .Z(n3037) );
  NANDN U3149 ( .A(n3014), .B(n3013), .Z(n3018) );
  NANDN U3150 ( .A(n3016), .B(n3015), .Z(n3017) );
  AND U3151 ( .A(n3018), .B(n3017), .Z(n3036) );
  XNOR U3152 ( .A(n3037), .B(n3036), .Z(n3038) );
  NANDN U3153 ( .A(n3020), .B(n3019), .Z(n3024) );
  NAND U3154 ( .A(n3022), .B(n3021), .Z(n3023) );
  NAND U3155 ( .A(n3024), .B(n3023), .Z(n3039) );
  XNOR U3156 ( .A(n3038), .B(n3039), .Z(n3030) );
  XNOR U3157 ( .A(n3031), .B(n3030), .Z(n3032) );
  XNOR U3158 ( .A(n3033), .B(n3032), .Z(n3066) );
  XNOR U3159 ( .A(sreg[325]), .B(n3066), .Z(n3068) );
  NANDN U3160 ( .A(sreg[324]), .B(n3025), .Z(n3029) );
  NAND U3161 ( .A(n3027), .B(n3026), .Z(n3028) );
  NAND U3162 ( .A(n3029), .B(n3028), .Z(n3067) );
  XNOR U3163 ( .A(n3068), .B(n3067), .Z(c[325]) );
  NANDN U3164 ( .A(n3031), .B(n3030), .Z(n3035) );
  NANDN U3165 ( .A(n3033), .B(n3032), .Z(n3034) );
  AND U3166 ( .A(n3035), .B(n3034), .Z(n3074) );
  NANDN U3167 ( .A(n3037), .B(n3036), .Z(n3041) );
  NANDN U3168 ( .A(n3039), .B(n3038), .Z(n3040) );
  AND U3169 ( .A(n3041), .B(n3040), .Z(n3072) );
  NAND U3170 ( .A(n26), .B(n3042), .Z(n3044) );
  XOR U3171 ( .A(b[7]), .B(a[72]), .Z(n3083) );
  NAND U3172 ( .A(n10531), .B(n3083), .Z(n3043) );
  AND U3173 ( .A(n3044), .B(n3043), .Z(n3102) );
  NAND U3174 ( .A(n23), .B(n3045), .Z(n3047) );
  XOR U3175 ( .A(b[3]), .B(a[76]), .Z(n3086) );
  NAND U3176 ( .A(n24), .B(n3086), .Z(n3046) );
  NAND U3177 ( .A(n3047), .B(n3046), .Z(n3101) );
  XNOR U3178 ( .A(n3102), .B(n3101), .Z(n3104) );
  NAND U3179 ( .A(b[0]), .B(a[78]), .Z(n3048) );
  XNOR U3180 ( .A(b[1]), .B(n3048), .Z(n3050) );
  NANDN U3181 ( .A(b[0]), .B(a[77]), .Z(n3049) );
  NAND U3182 ( .A(n3050), .B(n3049), .Z(n3098) );
  NAND U3183 ( .A(n25), .B(n3051), .Z(n3053) );
  XOR U3184 ( .A(b[5]), .B(a[74]), .Z(n3089) );
  NAND U3185 ( .A(n10456), .B(n3089), .Z(n3052) );
  AND U3186 ( .A(n3053), .B(n3052), .Z(n3096) );
  AND U3187 ( .A(b[7]), .B(a[70]), .Z(n3095) );
  XNOR U3188 ( .A(n3096), .B(n3095), .Z(n3097) );
  XNOR U3189 ( .A(n3098), .B(n3097), .Z(n3103) );
  XOR U3190 ( .A(n3104), .B(n3103), .Z(n3078) );
  NANDN U3191 ( .A(n3055), .B(n3054), .Z(n3059) );
  NANDN U3192 ( .A(n3057), .B(n3056), .Z(n3058) );
  AND U3193 ( .A(n3059), .B(n3058), .Z(n3077) );
  XNOR U3194 ( .A(n3078), .B(n3077), .Z(n3079) );
  NANDN U3195 ( .A(n3061), .B(n3060), .Z(n3065) );
  NAND U3196 ( .A(n3063), .B(n3062), .Z(n3064) );
  NAND U3197 ( .A(n3065), .B(n3064), .Z(n3080) );
  XNOR U3198 ( .A(n3079), .B(n3080), .Z(n3071) );
  XNOR U3199 ( .A(n3072), .B(n3071), .Z(n3073) );
  XNOR U3200 ( .A(n3074), .B(n3073), .Z(n3107) );
  XNOR U3201 ( .A(sreg[326]), .B(n3107), .Z(n3109) );
  NANDN U3202 ( .A(sreg[325]), .B(n3066), .Z(n3070) );
  NAND U3203 ( .A(n3068), .B(n3067), .Z(n3069) );
  NAND U3204 ( .A(n3070), .B(n3069), .Z(n3108) );
  XNOR U3205 ( .A(n3109), .B(n3108), .Z(c[326]) );
  NANDN U3206 ( .A(n3072), .B(n3071), .Z(n3076) );
  NANDN U3207 ( .A(n3074), .B(n3073), .Z(n3075) );
  AND U3208 ( .A(n3076), .B(n3075), .Z(n3115) );
  NANDN U3209 ( .A(n3078), .B(n3077), .Z(n3082) );
  NANDN U3210 ( .A(n3080), .B(n3079), .Z(n3081) );
  AND U3211 ( .A(n3082), .B(n3081), .Z(n3113) );
  NAND U3212 ( .A(n26), .B(n3083), .Z(n3085) );
  XOR U3213 ( .A(b[7]), .B(a[73]), .Z(n3124) );
  NAND U3214 ( .A(n10531), .B(n3124), .Z(n3084) );
  AND U3215 ( .A(n3085), .B(n3084), .Z(n3143) );
  NAND U3216 ( .A(n23), .B(n3086), .Z(n3088) );
  XOR U3217 ( .A(b[3]), .B(a[77]), .Z(n3127) );
  NAND U3218 ( .A(n24), .B(n3127), .Z(n3087) );
  NAND U3219 ( .A(n3088), .B(n3087), .Z(n3142) );
  XNOR U3220 ( .A(n3143), .B(n3142), .Z(n3145) );
  NAND U3221 ( .A(n25), .B(n3089), .Z(n3091) );
  XOR U3222 ( .A(b[5]), .B(a[75]), .Z(n3133) );
  NAND U3223 ( .A(n10456), .B(n3133), .Z(n3090) );
  AND U3224 ( .A(n3091), .B(n3090), .Z(n3137) );
  AND U3225 ( .A(b[7]), .B(a[71]), .Z(n3136) );
  XNOR U3226 ( .A(n3137), .B(n3136), .Z(n3138) );
  NAND U3227 ( .A(b[0]), .B(a[79]), .Z(n3092) );
  XNOR U3228 ( .A(b[1]), .B(n3092), .Z(n3094) );
  NANDN U3229 ( .A(b[0]), .B(a[78]), .Z(n3093) );
  NAND U3230 ( .A(n3094), .B(n3093), .Z(n3139) );
  XNOR U3231 ( .A(n3138), .B(n3139), .Z(n3144) );
  XOR U3232 ( .A(n3145), .B(n3144), .Z(n3119) );
  NANDN U3233 ( .A(n3096), .B(n3095), .Z(n3100) );
  NANDN U3234 ( .A(n3098), .B(n3097), .Z(n3099) );
  AND U3235 ( .A(n3100), .B(n3099), .Z(n3118) );
  XNOR U3236 ( .A(n3119), .B(n3118), .Z(n3120) );
  NANDN U3237 ( .A(n3102), .B(n3101), .Z(n3106) );
  NAND U3238 ( .A(n3104), .B(n3103), .Z(n3105) );
  NAND U3239 ( .A(n3106), .B(n3105), .Z(n3121) );
  XNOR U3240 ( .A(n3120), .B(n3121), .Z(n3112) );
  XNOR U3241 ( .A(n3113), .B(n3112), .Z(n3114) );
  XNOR U3242 ( .A(n3115), .B(n3114), .Z(n3148) );
  XNOR U3243 ( .A(sreg[327]), .B(n3148), .Z(n3150) );
  NANDN U3244 ( .A(sreg[326]), .B(n3107), .Z(n3111) );
  NAND U3245 ( .A(n3109), .B(n3108), .Z(n3110) );
  NAND U3246 ( .A(n3111), .B(n3110), .Z(n3149) );
  XNOR U3247 ( .A(n3150), .B(n3149), .Z(c[327]) );
  NANDN U3248 ( .A(n3113), .B(n3112), .Z(n3117) );
  NANDN U3249 ( .A(n3115), .B(n3114), .Z(n3116) );
  AND U3250 ( .A(n3117), .B(n3116), .Z(n3156) );
  NANDN U3251 ( .A(n3119), .B(n3118), .Z(n3123) );
  NANDN U3252 ( .A(n3121), .B(n3120), .Z(n3122) );
  AND U3253 ( .A(n3123), .B(n3122), .Z(n3154) );
  NAND U3254 ( .A(n26), .B(n3124), .Z(n3126) );
  XOR U3255 ( .A(b[7]), .B(a[74]), .Z(n3165) );
  NAND U3256 ( .A(n10531), .B(n3165), .Z(n3125) );
  AND U3257 ( .A(n3126), .B(n3125), .Z(n3184) );
  NAND U3258 ( .A(n23), .B(n3127), .Z(n3129) );
  XOR U3259 ( .A(b[3]), .B(a[78]), .Z(n3168) );
  NAND U3260 ( .A(n24), .B(n3168), .Z(n3128) );
  NAND U3261 ( .A(n3129), .B(n3128), .Z(n3183) );
  XNOR U3262 ( .A(n3184), .B(n3183), .Z(n3186) );
  NAND U3263 ( .A(b[0]), .B(a[80]), .Z(n3130) );
  XNOR U3264 ( .A(b[1]), .B(n3130), .Z(n3132) );
  NANDN U3265 ( .A(b[0]), .B(a[79]), .Z(n3131) );
  NAND U3266 ( .A(n3132), .B(n3131), .Z(n3180) );
  NAND U3267 ( .A(n25), .B(n3133), .Z(n3135) );
  XOR U3268 ( .A(b[5]), .B(a[76]), .Z(n3174) );
  NAND U3269 ( .A(n10456), .B(n3174), .Z(n3134) );
  AND U3270 ( .A(n3135), .B(n3134), .Z(n3178) );
  AND U3271 ( .A(b[7]), .B(a[72]), .Z(n3177) );
  XNOR U3272 ( .A(n3178), .B(n3177), .Z(n3179) );
  XNOR U3273 ( .A(n3180), .B(n3179), .Z(n3185) );
  XOR U3274 ( .A(n3186), .B(n3185), .Z(n3160) );
  NANDN U3275 ( .A(n3137), .B(n3136), .Z(n3141) );
  NANDN U3276 ( .A(n3139), .B(n3138), .Z(n3140) );
  AND U3277 ( .A(n3141), .B(n3140), .Z(n3159) );
  XNOR U3278 ( .A(n3160), .B(n3159), .Z(n3161) );
  NANDN U3279 ( .A(n3143), .B(n3142), .Z(n3147) );
  NAND U3280 ( .A(n3145), .B(n3144), .Z(n3146) );
  NAND U3281 ( .A(n3147), .B(n3146), .Z(n3162) );
  XNOR U3282 ( .A(n3161), .B(n3162), .Z(n3153) );
  XNOR U3283 ( .A(n3154), .B(n3153), .Z(n3155) );
  XNOR U3284 ( .A(n3156), .B(n3155), .Z(n3189) );
  XNOR U3285 ( .A(sreg[328]), .B(n3189), .Z(n3191) );
  NANDN U3286 ( .A(sreg[327]), .B(n3148), .Z(n3152) );
  NAND U3287 ( .A(n3150), .B(n3149), .Z(n3151) );
  NAND U3288 ( .A(n3152), .B(n3151), .Z(n3190) );
  XNOR U3289 ( .A(n3191), .B(n3190), .Z(c[328]) );
  NANDN U3290 ( .A(n3154), .B(n3153), .Z(n3158) );
  NANDN U3291 ( .A(n3156), .B(n3155), .Z(n3157) );
  AND U3292 ( .A(n3158), .B(n3157), .Z(n3197) );
  NANDN U3293 ( .A(n3160), .B(n3159), .Z(n3164) );
  NANDN U3294 ( .A(n3162), .B(n3161), .Z(n3163) );
  AND U3295 ( .A(n3164), .B(n3163), .Z(n3195) );
  NAND U3296 ( .A(n26), .B(n3165), .Z(n3167) );
  XOR U3297 ( .A(b[7]), .B(a[75]), .Z(n3206) );
  NAND U3298 ( .A(n10531), .B(n3206), .Z(n3166) );
  AND U3299 ( .A(n3167), .B(n3166), .Z(n3225) );
  NAND U3300 ( .A(n23), .B(n3168), .Z(n3170) );
  XOR U3301 ( .A(b[3]), .B(a[79]), .Z(n3209) );
  NAND U3302 ( .A(n24), .B(n3209), .Z(n3169) );
  NAND U3303 ( .A(n3170), .B(n3169), .Z(n3224) );
  XNOR U3304 ( .A(n3225), .B(n3224), .Z(n3227) );
  NAND U3305 ( .A(b[0]), .B(a[81]), .Z(n3171) );
  XNOR U3306 ( .A(b[1]), .B(n3171), .Z(n3173) );
  NANDN U3307 ( .A(b[0]), .B(a[80]), .Z(n3172) );
  NAND U3308 ( .A(n3173), .B(n3172), .Z(n3221) );
  NAND U3309 ( .A(n25), .B(n3174), .Z(n3176) );
  XOR U3310 ( .A(b[5]), .B(a[77]), .Z(n3215) );
  NAND U3311 ( .A(n10456), .B(n3215), .Z(n3175) );
  AND U3312 ( .A(n3176), .B(n3175), .Z(n3219) );
  AND U3313 ( .A(b[7]), .B(a[73]), .Z(n3218) );
  XNOR U3314 ( .A(n3219), .B(n3218), .Z(n3220) );
  XNOR U3315 ( .A(n3221), .B(n3220), .Z(n3226) );
  XOR U3316 ( .A(n3227), .B(n3226), .Z(n3201) );
  NANDN U3317 ( .A(n3178), .B(n3177), .Z(n3182) );
  NANDN U3318 ( .A(n3180), .B(n3179), .Z(n3181) );
  AND U3319 ( .A(n3182), .B(n3181), .Z(n3200) );
  XNOR U3320 ( .A(n3201), .B(n3200), .Z(n3202) );
  NANDN U3321 ( .A(n3184), .B(n3183), .Z(n3188) );
  NAND U3322 ( .A(n3186), .B(n3185), .Z(n3187) );
  NAND U3323 ( .A(n3188), .B(n3187), .Z(n3203) );
  XNOR U3324 ( .A(n3202), .B(n3203), .Z(n3194) );
  XNOR U3325 ( .A(n3195), .B(n3194), .Z(n3196) );
  XNOR U3326 ( .A(n3197), .B(n3196), .Z(n3230) );
  XNOR U3327 ( .A(sreg[329]), .B(n3230), .Z(n3232) );
  NANDN U3328 ( .A(sreg[328]), .B(n3189), .Z(n3193) );
  NAND U3329 ( .A(n3191), .B(n3190), .Z(n3192) );
  NAND U3330 ( .A(n3193), .B(n3192), .Z(n3231) );
  XNOR U3331 ( .A(n3232), .B(n3231), .Z(c[329]) );
  NANDN U3332 ( .A(n3195), .B(n3194), .Z(n3199) );
  NANDN U3333 ( .A(n3197), .B(n3196), .Z(n3198) );
  AND U3334 ( .A(n3199), .B(n3198), .Z(n3238) );
  NANDN U3335 ( .A(n3201), .B(n3200), .Z(n3205) );
  NANDN U3336 ( .A(n3203), .B(n3202), .Z(n3204) );
  AND U3337 ( .A(n3205), .B(n3204), .Z(n3236) );
  NAND U3338 ( .A(n26), .B(n3206), .Z(n3208) );
  XOR U3339 ( .A(b[7]), .B(a[76]), .Z(n3247) );
  NAND U3340 ( .A(n10531), .B(n3247), .Z(n3207) );
  AND U3341 ( .A(n3208), .B(n3207), .Z(n3266) );
  NAND U3342 ( .A(n23), .B(n3209), .Z(n3211) );
  XOR U3343 ( .A(b[3]), .B(a[80]), .Z(n3250) );
  NAND U3344 ( .A(n24), .B(n3250), .Z(n3210) );
  NAND U3345 ( .A(n3211), .B(n3210), .Z(n3265) );
  XNOR U3346 ( .A(n3266), .B(n3265), .Z(n3268) );
  NAND U3347 ( .A(b[0]), .B(a[82]), .Z(n3212) );
  XNOR U3348 ( .A(b[1]), .B(n3212), .Z(n3214) );
  NANDN U3349 ( .A(b[0]), .B(a[81]), .Z(n3213) );
  NAND U3350 ( .A(n3214), .B(n3213), .Z(n3262) );
  NAND U3351 ( .A(n25), .B(n3215), .Z(n3217) );
  XOR U3352 ( .A(b[5]), .B(a[78]), .Z(n3256) );
  NAND U3353 ( .A(n10456), .B(n3256), .Z(n3216) );
  AND U3354 ( .A(n3217), .B(n3216), .Z(n3260) );
  AND U3355 ( .A(b[7]), .B(a[74]), .Z(n3259) );
  XNOR U3356 ( .A(n3260), .B(n3259), .Z(n3261) );
  XNOR U3357 ( .A(n3262), .B(n3261), .Z(n3267) );
  XOR U3358 ( .A(n3268), .B(n3267), .Z(n3242) );
  NANDN U3359 ( .A(n3219), .B(n3218), .Z(n3223) );
  NANDN U3360 ( .A(n3221), .B(n3220), .Z(n3222) );
  AND U3361 ( .A(n3223), .B(n3222), .Z(n3241) );
  XNOR U3362 ( .A(n3242), .B(n3241), .Z(n3243) );
  NANDN U3363 ( .A(n3225), .B(n3224), .Z(n3229) );
  NAND U3364 ( .A(n3227), .B(n3226), .Z(n3228) );
  NAND U3365 ( .A(n3229), .B(n3228), .Z(n3244) );
  XNOR U3366 ( .A(n3243), .B(n3244), .Z(n3235) );
  XNOR U3367 ( .A(n3236), .B(n3235), .Z(n3237) );
  XNOR U3368 ( .A(n3238), .B(n3237), .Z(n3271) );
  XNOR U3369 ( .A(sreg[330]), .B(n3271), .Z(n3273) );
  NANDN U3370 ( .A(sreg[329]), .B(n3230), .Z(n3234) );
  NAND U3371 ( .A(n3232), .B(n3231), .Z(n3233) );
  NAND U3372 ( .A(n3234), .B(n3233), .Z(n3272) );
  XNOR U3373 ( .A(n3273), .B(n3272), .Z(c[330]) );
  NANDN U3374 ( .A(n3236), .B(n3235), .Z(n3240) );
  NANDN U3375 ( .A(n3238), .B(n3237), .Z(n3239) );
  AND U3376 ( .A(n3240), .B(n3239), .Z(n3279) );
  NANDN U3377 ( .A(n3242), .B(n3241), .Z(n3246) );
  NANDN U3378 ( .A(n3244), .B(n3243), .Z(n3245) );
  AND U3379 ( .A(n3246), .B(n3245), .Z(n3277) );
  NAND U3380 ( .A(n26), .B(n3247), .Z(n3249) );
  XOR U3381 ( .A(b[7]), .B(a[77]), .Z(n3288) );
  NAND U3382 ( .A(n10531), .B(n3288), .Z(n3248) );
  AND U3383 ( .A(n3249), .B(n3248), .Z(n3307) );
  NAND U3384 ( .A(n23), .B(n3250), .Z(n3252) );
  XOR U3385 ( .A(b[3]), .B(a[81]), .Z(n3291) );
  NAND U3386 ( .A(n24), .B(n3291), .Z(n3251) );
  NAND U3387 ( .A(n3252), .B(n3251), .Z(n3306) );
  XNOR U3388 ( .A(n3307), .B(n3306), .Z(n3309) );
  NAND U3389 ( .A(b[0]), .B(a[83]), .Z(n3253) );
  XNOR U3390 ( .A(b[1]), .B(n3253), .Z(n3255) );
  NANDN U3391 ( .A(b[0]), .B(a[82]), .Z(n3254) );
  NAND U3392 ( .A(n3255), .B(n3254), .Z(n3303) );
  NAND U3393 ( .A(n25), .B(n3256), .Z(n3258) );
  XOR U3394 ( .A(b[5]), .B(a[79]), .Z(n3297) );
  NAND U3395 ( .A(n10456), .B(n3297), .Z(n3257) );
  AND U3396 ( .A(n3258), .B(n3257), .Z(n3301) );
  AND U3397 ( .A(b[7]), .B(a[75]), .Z(n3300) );
  XNOR U3398 ( .A(n3301), .B(n3300), .Z(n3302) );
  XNOR U3399 ( .A(n3303), .B(n3302), .Z(n3308) );
  XOR U3400 ( .A(n3309), .B(n3308), .Z(n3283) );
  NANDN U3401 ( .A(n3260), .B(n3259), .Z(n3264) );
  NANDN U3402 ( .A(n3262), .B(n3261), .Z(n3263) );
  AND U3403 ( .A(n3264), .B(n3263), .Z(n3282) );
  XNOR U3404 ( .A(n3283), .B(n3282), .Z(n3284) );
  NANDN U3405 ( .A(n3266), .B(n3265), .Z(n3270) );
  NAND U3406 ( .A(n3268), .B(n3267), .Z(n3269) );
  NAND U3407 ( .A(n3270), .B(n3269), .Z(n3285) );
  XNOR U3408 ( .A(n3284), .B(n3285), .Z(n3276) );
  XNOR U3409 ( .A(n3277), .B(n3276), .Z(n3278) );
  XNOR U3410 ( .A(n3279), .B(n3278), .Z(n3312) );
  XNOR U3411 ( .A(sreg[331]), .B(n3312), .Z(n3314) );
  NANDN U3412 ( .A(sreg[330]), .B(n3271), .Z(n3275) );
  NAND U3413 ( .A(n3273), .B(n3272), .Z(n3274) );
  NAND U3414 ( .A(n3275), .B(n3274), .Z(n3313) );
  XNOR U3415 ( .A(n3314), .B(n3313), .Z(c[331]) );
  NANDN U3416 ( .A(n3277), .B(n3276), .Z(n3281) );
  NANDN U3417 ( .A(n3279), .B(n3278), .Z(n3280) );
  AND U3418 ( .A(n3281), .B(n3280), .Z(n3320) );
  NANDN U3419 ( .A(n3283), .B(n3282), .Z(n3287) );
  NANDN U3420 ( .A(n3285), .B(n3284), .Z(n3286) );
  AND U3421 ( .A(n3287), .B(n3286), .Z(n3318) );
  NAND U3422 ( .A(n26), .B(n3288), .Z(n3290) );
  XOR U3423 ( .A(b[7]), .B(a[78]), .Z(n3329) );
  NAND U3424 ( .A(n10531), .B(n3329), .Z(n3289) );
  AND U3425 ( .A(n3290), .B(n3289), .Z(n3348) );
  NAND U3426 ( .A(n23), .B(n3291), .Z(n3293) );
  XOR U3427 ( .A(b[3]), .B(a[82]), .Z(n3332) );
  NAND U3428 ( .A(n24), .B(n3332), .Z(n3292) );
  NAND U3429 ( .A(n3293), .B(n3292), .Z(n3347) );
  XNOR U3430 ( .A(n3348), .B(n3347), .Z(n3350) );
  NAND U3431 ( .A(b[0]), .B(a[84]), .Z(n3294) );
  XNOR U3432 ( .A(b[1]), .B(n3294), .Z(n3296) );
  NANDN U3433 ( .A(b[0]), .B(a[83]), .Z(n3295) );
  NAND U3434 ( .A(n3296), .B(n3295), .Z(n3344) );
  NAND U3435 ( .A(n25), .B(n3297), .Z(n3299) );
  XOR U3436 ( .A(b[5]), .B(a[80]), .Z(n3338) );
  NAND U3437 ( .A(n10456), .B(n3338), .Z(n3298) );
  AND U3438 ( .A(n3299), .B(n3298), .Z(n3342) );
  AND U3439 ( .A(b[7]), .B(a[76]), .Z(n3341) );
  XNOR U3440 ( .A(n3342), .B(n3341), .Z(n3343) );
  XNOR U3441 ( .A(n3344), .B(n3343), .Z(n3349) );
  XOR U3442 ( .A(n3350), .B(n3349), .Z(n3324) );
  NANDN U3443 ( .A(n3301), .B(n3300), .Z(n3305) );
  NANDN U3444 ( .A(n3303), .B(n3302), .Z(n3304) );
  AND U3445 ( .A(n3305), .B(n3304), .Z(n3323) );
  XNOR U3446 ( .A(n3324), .B(n3323), .Z(n3325) );
  NANDN U3447 ( .A(n3307), .B(n3306), .Z(n3311) );
  NAND U3448 ( .A(n3309), .B(n3308), .Z(n3310) );
  NAND U3449 ( .A(n3311), .B(n3310), .Z(n3326) );
  XNOR U3450 ( .A(n3325), .B(n3326), .Z(n3317) );
  XNOR U3451 ( .A(n3318), .B(n3317), .Z(n3319) );
  XNOR U3452 ( .A(n3320), .B(n3319), .Z(n3353) );
  XNOR U3453 ( .A(sreg[332]), .B(n3353), .Z(n3355) );
  NANDN U3454 ( .A(sreg[331]), .B(n3312), .Z(n3316) );
  NAND U3455 ( .A(n3314), .B(n3313), .Z(n3315) );
  NAND U3456 ( .A(n3316), .B(n3315), .Z(n3354) );
  XNOR U3457 ( .A(n3355), .B(n3354), .Z(c[332]) );
  NANDN U3458 ( .A(n3318), .B(n3317), .Z(n3322) );
  NANDN U3459 ( .A(n3320), .B(n3319), .Z(n3321) );
  AND U3460 ( .A(n3322), .B(n3321), .Z(n3361) );
  NANDN U3461 ( .A(n3324), .B(n3323), .Z(n3328) );
  NANDN U3462 ( .A(n3326), .B(n3325), .Z(n3327) );
  AND U3463 ( .A(n3328), .B(n3327), .Z(n3359) );
  NAND U3464 ( .A(n26), .B(n3329), .Z(n3331) );
  XOR U3465 ( .A(b[7]), .B(a[79]), .Z(n3370) );
  NAND U3466 ( .A(n10531), .B(n3370), .Z(n3330) );
  AND U3467 ( .A(n3331), .B(n3330), .Z(n3389) );
  NAND U3468 ( .A(n23), .B(n3332), .Z(n3334) );
  XOR U3469 ( .A(b[3]), .B(a[83]), .Z(n3373) );
  NAND U3470 ( .A(n24), .B(n3373), .Z(n3333) );
  NAND U3471 ( .A(n3334), .B(n3333), .Z(n3388) );
  XNOR U3472 ( .A(n3389), .B(n3388), .Z(n3391) );
  NAND U3473 ( .A(b[0]), .B(a[85]), .Z(n3335) );
  XNOR U3474 ( .A(b[1]), .B(n3335), .Z(n3337) );
  NANDN U3475 ( .A(b[0]), .B(a[84]), .Z(n3336) );
  NAND U3476 ( .A(n3337), .B(n3336), .Z(n3385) );
  NAND U3477 ( .A(n25), .B(n3338), .Z(n3340) );
  XOR U3478 ( .A(b[5]), .B(a[81]), .Z(n3379) );
  NAND U3479 ( .A(n10456), .B(n3379), .Z(n3339) );
  AND U3480 ( .A(n3340), .B(n3339), .Z(n3383) );
  AND U3481 ( .A(b[7]), .B(a[77]), .Z(n3382) );
  XNOR U3482 ( .A(n3383), .B(n3382), .Z(n3384) );
  XNOR U3483 ( .A(n3385), .B(n3384), .Z(n3390) );
  XOR U3484 ( .A(n3391), .B(n3390), .Z(n3365) );
  NANDN U3485 ( .A(n3342), .B(n3341), .Z(n3346) );
  NANDN U3486 ( .A(n3344), .B(n3343), .Z(n3345) );
  AND U3487 ( .A(n3346), .B(n3345), .Z(n3364) );
  XNOR U3488 ( .A(n3365), .B(n3364), .Z(n3366) );
  NANDN U3489 ( .A(n3348), .B(n3347), .Z(n3352) );
  NAND U3490 ( .A(n3350), .B(n3349), .Z(n3351) );
  NAND U3491 ( .A(n3352), .B(n3351), .Z(n3367) );
  XNOR U3492 ( .A(n3366), .B(n3367), .Z(n3358) );
  XNOR U3493 ( .A(n3359), .B(n3358), .Z(n3360) );
  XNOR U3494 ( .A(n3361), .B(n3360), .Z(n3394) );
  XNOR U3495 ( .A(sreg[333]), .B(n3394), .Z(n3396) );
  NANDN U3496 ( .A(sreg[332]), .B(n3353), .Z(n3357) );
  NAND U3497 ( .A(n3355), .B(n3354), .Z(n3356) );
  NAND U3498 ( .A(n3357), .B(n3356), .Z(n3395) );
  XNOR U3499 ( .A(n3396), .B(n3395), .Z(c[333]) );
  NANDN U3500 ( .A(n3359), .B(n3358), .Z(n3363) );
  NANDN U3501 ( .A(n3361), .B(n3360), .Z(n3362) );
  AND U3502 ( .A(n3363), .B(n3362), .Z(n3402) );
  NANDN U3503 ( .A(n3365), .B(n3364), .Z(n3369) );
  NANDN U3504 ( .A(n3367), .B(n3366), .Z(n3368) );
  AND U3505 ( .A(n3369), .B(n3368), .Z(n3400) );
  NAND U3506 ( .A(n26), .B(n3370), .Z(n3372) );
  XOR U3507 ( .A(b[7]), .B(a[80]), .Z(n3411) );
  NAND U3508 ( .A(n10531), .B(n3411), .Z(n3371) );
  AND U3509 ( .A(n3372), .B(n3371), .Z(n3430) );
  NAND U3510 ( .A(n23), .B(n3373), .Z(n3375) );
  XOR U3511 ( .A(b[3]), .B(a[84]), .Z(n3414) );
  NAND U3512 ( .A(n24), .B(n3414), .Z(n3374) );
  NAND U3513 ( .A(n3375), .B(n3374), .Z(n3429) );
  XNOR U3514 ( .A(n3430), .B(n3429), .Z(n3432) );
  NAND U3515 ( .A(b[0]), .B(a[86]), .Z(n3376) );
  XNOR U3516 ( .A(b[1]), .B(n3376), .Z(n3378) );
  NANDN U3517 ( .A(b[0]), .B(a[85]), .Z(n3377) );
  NAND U3518 ( .A(n3378), .B(n3377), .Z(n3426) );
  NAND U3519 ( .A(n25), .B(n3379), .Z(n3381) );
  XOR U3520 ( .A(b[5]), .B(a[82]), .Z(n3417) );
  NAND U3521 ( .A(n10456), .B(n3417), .Z(n3380) );
  AND U3522 ( .A(n3381), .B(n3380), .Z(n3424) );
  AND U3523 ( .A(b[7]), .B(a[78]), .Z(n3423) );
  XNOR U3524 ( .A(n3424), .B(n3423), .Z(n3425) );
  XNOR U3525 ( .A(n3426), .B(n3425), .Z(n3431) );
  XOR U3526 ( .A(n3432), .B(n3431), .Z(n3406) );
  NANDN U3527 ( .A(n3383), .B(n3382), .Z(n3387) );
  NANDN U3528 ( .A(n3385), .B(n3384), .Z(n3386) );
  AND U3529 ( .A(n3387), .B(n3386), .Z(n3405) );
  XNOR U3530 ( .A(n3406), .B(n3405), .Z(n3407) );
  NANDN U3531 ( .A(n3389), .B(n3388), .Z(n3393) );
  NAND U3532 ( .A(n3391), .B(n3390), .Z(n3392) );
  NAND U3533 ( .A(n3393), .B(n3392), .Z(n3408) );
  XNOR U3534 ( .A(n3407), .B(n3408), .Z(n3399) );
  XNOR U3535 ( .A(n3400), .B(n3399), .Z(n3401) );
  XNOR U3536 ( .A(n3402), .B(n3401), .Z(n3435) );
  XNOR U3537 ( .A(sreg[334]), .B(n3435), .Z(n3437) );
  NANDN U3538 ( .A(sreg[333]), .B(n3394), .Z(n3398) );
  NAND U3539 ( .A(n3396), .B(n3395), .Z(n3397) );
  NAND U3540 ( .A(n3398), .B(n3397), .Z(n3436) );
  XNOR U3541 ( .A(n3437), .B(n3436), .Z(c[334]) );
  NANDN U3542 ( .A(n3400), .B(n3399), .Z(n3404) );
  NANDN U3543 ( .A(n3402), .B(n3401), .Z(n3403) );
  AND U3544 ( .A(n3404), .B(n3403), .Z(n3443) );
  NANDN U3545 ( .A(n3406), .B(n3405), .Z(n3410) );
  NANDN U3546 ( .A(n3408), .B(n3407), .Z(n3409) );
  AND U3547 ( .A(n3410), .B(n3409), .Z(n3441) );
  NAND U3548 ( .A(n26), .B(n3411), .Z(n3413) );
  XOR U3549 ( .A(b[7]), .B(a[81]), .Z(n3452) );
  NAND U3550 ( .A(n10531), .B(n3452), .Z(n3412) );
  AND U3551 ( .A(n3413), .B(n3412), .Z(n3471) );
  NAND U3552 ( .A(n23), .B(n3414), .Z(n3416) );
  XOR U3553 ( .A(b[3]), .B(a[85]), .Z(n3455) );
  NAND U3554 ( .A(n24), .B(n3455), .Z(n3415) );
  NAND U3555 ( .A(n3416), .B(n3415), .Z(n3470) );
  XNOR U3556 ( .A(n3471), .B(n3470), .Z(n3473) );
  NAND U3557 ( .A(n25), .B(n3417), .Z(n3419) );
  XOR U3558 ( .A(b[5]), .B(a[83]), .Z(n3461) );
  NAND U3559 ( .A(n10456), .B(n3461), .Z(n3418) );
  AND U3560 ( .A(n3419), .B(n3418), .Z(n3465) );
  AND U3561 ( .A(b[7]), .B(a[79]), .Z(n3464) );
  XNOR U3562 ( .A(n3465), .B(n3464), .Z(n3466) );
  NAND U3563 ( .A(b[0]), .B(a[87]), .Z(n3420) );
  XNOR U3564 ( .A(b[1]), .B(n3420), .Z(n3422) );
  NANDN U3565 ( .A(b[0]), .B(a[86]), .Z(n3421) );
  NAND U3566 ( .A(n3422), .B(n3421), .Z(n3467) );
  XNOR U3567 ( .A(n3466), .B(n3467), .Z(n3472) );
  XOR U3568 ( .A(n3473), .B(n3472), .Z(n3447) );
  NANDN U3569 ( .A(n3424), .B(n3423), .Z(n3428) );
  NANDN U3570 ( .A(n3426), .B(n3425), .Z(n3427) );
  AND U3571 ( .A(n3428), .B(n3427), .Z(n3446) );
  XNOR U3572 ( .A(n3447), .B(n3446), .Z(n3448) );
  NANDN U3573 ( .A(n3430), .B(n3429), .Z(n3434) );
  NAND U3574 ( .A(n3432), .B(n3431), .Z(n3433) );
  NAND U3575 ( .A(n3434), .B(n3433), .Z(n3449) );
  XNOR U3576 ( .A(n3448), .B(n3449), .Z(n3440) );
  XNOR U3577 ( .A(n3441), .B(n3440), .Z(n3442) );
  XNOR U3578 ( .A(n3443), .B(n3442), .Z(n3476) );
  XNOR U3579 ( .A(sreg[335]), .B(n3476), .Z(n3478) );
  NANDN U3580 ( .A(sreg[334]), .B(n3435), .Z(n3439) );
  NAND U3581 ( .A(n3437), .B(n3436), .Z(n3438) );
  NAND U3582 ( .A(n3439), .B(n3438), .Z(n3477) );
  XNOR U3583 ( .A(n3478), .B(n3477), .Z(c[335]) );
  NANDN U3584 ( .A(n3441), .B(n3440), .Z(n3445) );
  NANDN U3585 ( .A(n3443), .B(n3442), .Z(n3444) );
  AND U3586 ( .A(n3445), .B(n3444), .Z(n3484) );
  NANDN U3587 ( .A(n3447), .B(n3446), .Z(n3451) );
  NANDN U3588 ( .A(n3449), .B(n3448), .Z(n3450) );
  AND U3589 ( .A(n3451), .B(n3450), .Z(n3482) );
  NAND U3590 ( .A(n26), .B(n3452), .Z(n3454) );
  XOR U3591 ( .A(b[7]), .B(a[82]), .Z(n3493) );
  NAND U3592 ( .A(n10531), .B(n3493), .Z(n3453) );
  AND U3593 ( .A(n3454), .B(n3453), .Z(n3512) );
  NAND U3594 ( .A(n23), .B(n3455), .Z(n3457) );
  XOR U3595 ( .A(b[3]), .B(a[86]), .Z(n3496) );
  NAND U3596 ( .A(n24), .B(n3496), .Z(n3456) );
  NAND U3597 ( .A(n3457), .B(n3456), .Z(n3511) );
  XNOR U3598 ( .A(n3512), .B(n3511), .Z(n3514) );
  NAND U3599 ( .A(b[0]), .B(a[88]), .Z(n3458) );
  XNOR U3600 ( .A(b[1]), .B(n3458), .Z(n3460) );
  NANDN U3601 ( .A(b[0]), .B(a[87]), .Z(n3459) );
  NAND U3602 ( .A(n3460), .B(n3459), .Z(n3508) );
  NAND U3603 ( .A(n25), .B(n3461), .Z(n3463) );
  XOR U3604 ( .A(b[5]), .B(a[84]), .Z(n3502) );
  NAND U3605 ( .A(n10456), .B(n3502), .Z(n3462) );
  AND U3606 ( .A(n3463), .B(n3462), .Z(n3506) );
  AND U3607 ( .A(b[7]), .B(a[80]), .Z(n3505) );
  XNOR U3608 ( .A(n3506), .B(n3505), .Z(n3507) );
  XNOR U3609 ( .A(n3508), .B(n3507), .Z(n3513) );
  XOR U3610 ( .A(n3514), .B(n3513), .Z(n3488) );
  NANDN U3611 ( .A(n3465), .B(n3464), .Z(n3469) );
  NANDN U3612 ( .A(n3467), .B(n3466), .Z(n3468) );
  AND U3613 ( .A(n3469), .B(n3468), .Z(n3487) );
  XNOR U3614 ( .A(n3488), .B(n3487), .Z(n3489) );
  NANDN U3615 ( .A(n3471), .B(n3470), .Z(n3475) );
  NAND U3616 ( .A(n3473), .B(n3472), .Z(n3474) );
  NAND U3617 ( .A(n3475), .B(n3474), .Z(n3490) );
  XNOR U3618 ( .A(n3489), .B(n3490), .Z(n3481) );
  XNOR U3619 ( .A(n3482), .B(n3481), .Z(n3483) );
  XNOR U3620 ( .A(n3484), .B(n3483), .Z(n3517) );
  XNOR U3621 ( .A(sreg[336]), .B(n3517), .Z(n3519) );
  NANDN U3622 ( .A(sreg[335]), .B(n3476), .Z(n3480) );
  NAND U3623 ( .A(n3478), .B(n3477), .Z(n3479) );
  NAND U3624 ( .A(n3480), .B(n3479), .Z(n3518) );
  XNOR U3625 ( .A(n3519), .B(n3518), .Z(c[336]) );
  NANDN U3626 ( .A(n3482), .B(n3481), .Z(n3486) );
  NANDN U3627 ( .A(n3484), .B(n3483), .Z(n3485) );
  AND U3628 ( .A(n3486), .B(n3485), .Z(n3525) );
  NANDN U3629 ( .A(n3488), .B(n3487), .Z(n3492) );
  NANDN U3630 ( .A(n3490), .B(n3489), .Z(n3491) );
  AND U3631 ( .A(n3492), .B(n3491), .Z(n3523) );
  NAND U3632 ( .A(n26), .B(n3493), .Z(n3495) );
  XOR U3633 ( .A(b[7]), .B(a[83]), .Z(n3534) );
  NAND U3634 ( .A(n10531), .B(n3534), .Z(n3494) );
  AND U3635 ( .A(n3495), .B(n3494), .Z(n3553) );
  NAND U3636 ( .A(n23), .B(n3496), .Z(n3498) );
  XOR U3637 ( .A(b[3]), .B(a[87]), .Z(n3537) );
  NAND U3638 ( .A(n24), .B(n3537), .Z(n3497) );
  NAND U3639 ( .A(n3498), .B(n3497), .Z(n3552) );
  XNOR U3640 ( .A(n3553), .B(n3552), .Z(n3555) );
  NAND U3641 ( .A(b[0]), .B(a[89]), .Z(n3499) );
  XNOR U3642 ( .A(b[1]), .B(n3499), .Z(n3501) );
  NANDN U3643 ( .A(b[0]), .B(a[88]), .Z(n3500) );
  NAND U3644 ( .A(n3501), .B(n3500), .Z(n3549) );
  NAND U3645 ( .A(n25), .B(n3502), .Z(n3504) );
  XOR U3646 ( .A(b[5]), .B(a[85]), .Z(n3543) );
  NAND U3647 ( .A(n10456), .B(n3543), .Z(n3503) );
  AND U3648 ( .A(n3504), .B(n3503), .Z(n3547) );
  AND U3649 ( .A(b[7]), .B(a[81]), .Z(n3546) );
  XNOR U3650 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U3651 ( .A(n3549), .B(n3548), .Z(n3554) );
  XOR U3652 ( .A(n3555), .B(n3554), .Z(n3529) );
  NANDN U3653 ( .A(n3506), .B(n3505), .Z(n3510) );
  NANDN U3654 ( .A(n3508), .B(n3507), .Z(n3509) );
  AND U3655 ( .A(n3510), .B(n3509), .Z(n3528) );
  XNOR U3656 ( .A(n3529), .B(n3528), .Z(n3530) );
  NANDN U3657 ( .A(n3512), .B(n3511), .Z(n3516) );
  NAND U3658 ( .A(n3514), .B(n3513), .Z(n3515) );
  NAND U3659 ( .A(n3516), .B(n3515), .Z(n3531) );
  XNOR U3660 ( .A(n3530), .B(n3531), .Z(n3522) );
  XNOR U3661 ( .A(n3523), .B(n3522), .Z(n3524) );
  XNOR U3662 ( .A(n3525), .B(n3524), .Z(n3558) );
  XNOR U3663 ( .A(sreg[337]), .B(n3558), .Z(n3560) );
  NANDN U3664 ( .A(sreg[336]), .B(n3517), .Z(n3521) );
  NAND U3665 ( .A(n3519), .B(n3518), .Z(n3520) );
  NAND U3666 ( .A(n3521), .B(n3520), .Z(n3559) );
  XNOR U3667 ( .A(n3560), .B(n3559), .Z(c[337]) );
  NANDN U3668 ( .A(n3523), .B(n3522), .Z(n3527) );
  NANDN U3669 ( .A(n3525), .B(n3524), .Z(n3526) );
  AND U3670 ( .A(n3527), .B(n3526), .Z(n3566) );
  NANDN U3671 ( .A(n3529), .B(n3528), .Z(n3533) );
  NANDN U3672 ( .A(n3531), .B(n3530), .Z(n3532) );
  AND U3673 ( .A(n3533), .B(n3532), .Z(n3564) );
  NAND U3674 ( .A(n26), .B(n3534), .Z(n3536) );
  XOR U3675 ( .A(b[7]), .B(a[84]), .Z(n3575) );
  NAND U3676 ( .A(n10531), .B(n3575), .Z(n3535) );
  AND U3677 ( .A(n3536), .B(n3535), .Z(n3594) );
  NAND U3678 ( .A(n23), .B(n3537), .Z(n3539) );
  XOR U3679 ( .A(b[3]), .B(a[88]), .Z(n3578) );
  NAND U3680 ( .A(n24), .B(n3578), .Z(n3538) );
  NAND U3681 ( .A(n3539), .B(n3538), .Z(n3593) );
  XNOR U3682 ( .A(n3594), .B(n3593), .Z(n3596) );
  NAND U3683 ( .A(b[0]), .B(a[90]), .Z(n3540) );
  XNOR U3684 ( .A(b[1]), .B(n3540), .Z(n3542) );
  NANDN U3685 ( .A(b[0]), .B(a[89]), .Z(n3541) );
  NAND U3686 ( .A(n3542), .B(n3541), .Z(n3590) );
  NAND U3687 ( .A(n25), .B(n3543), .Z(n3545) );
  XOR U3688 ( .A(b[5]), .B(a[86]), .Z(n3584) );
  NAND U3689 ( .A(n10456), .B(n3584), .Z(n3544) );
  AND U3690 ( .A(n3545), .B(n3544), .Z(n3588) );
  AND U3691 ( .A(b[7]), .B(a[82]), .Z(n3587) );
  XNOR U3692 ( .A(n3588), .B(n3587), .Z(n3589) );
  XNOR U3693 ( .A(n3590), .B(n3589), .Z(n3595) );
  XOR U3694 ( .A(n3596), .B(n3595), .Z(n3570) );
  NANDN U3695 ( .A(n3547), .B(n3546), .Z(n3551) );
  NANDN U3696 ( .A(n3549), .B(n3548), .Z(n3550) );
  AND U3697 ( .A(n3551), .B(n3550), .Z(n3569) );
  XNOR U3698 ( .A(n3570), .B(n3569), .Z(n3571) );
  NANDN U3699 ( .A(n3553), .B(n3552), .Z(n3557) );
  NAND U3700 ( .A(n3555), .B(n3554), .Z(n3556) );
  NAND U3701 ( .A(n3557), .B(n3556), .Z(n3572) );
  XNOR U3702 ( .A(n3571), .B(n3572), .Z(n3563) );
  XNOR U3703 ( .A(n3564), .B(n3563), .Z(n3565) );
  XNOR U3704 ( .A(n3566), .B(n3565), .Z(n3599) );
  XNOR U3705 ( .A(sreg[338]), .B(n3599), .Z(n3601) );
  NANDN U3706 ( .A(sreg[337]), .B(n3558), .Z(n3562) );
  NAND U3707 ( .A(n3560), .B(n3559), .Z(n3561) );
  NAND U3708 ( .A(n3562), .B(n3561), .Z(n3600) );
  XNOR U3709 ( .A(n3601), .B(n3600), .Z(c[338]) );
  NANDN U3710 ( .A(n3564), .B(n3563), .Z(n3568) );
  NANDN U3711 ( .A(n3566), .B(n3565), .Z(n3567) );
  AND U3712 ( .A(n3568), .B(n3567), .Z(n3607) );
  NANDN U3713 ( .A(n3570), .B(n3569), .Z(n3574) );
  NANDN U3714 ( .A(n3572), .B(n3571), .Z(n3573) );
  AND U3715 ( .A(n3574), .B(n3573), .Z(n3605) );
  NAND U3716 ( .A(n26), .B(n3575), .Z(n3577) );
  XOR U3717 ( .A(b[7]), .B(a[85]), .Z(n3616) );
  NAND U3718 ( .A(n10531), .B(n3616), .Z(n3576) );
  AND U3719 ( .A(n3577), .B(n3576), .Z(n3635) );
  NAND U3720 ( .A(n23), .B(n3578), .Z(n3580) );
  XOR U3721 ( .A(b[3]), .B(a[89]), .Z(n3619) );
  NAND U3722 ( .A(n24), .B(n3619), .Z(n3579) );
  NAND U3723 ( .A(n3580), .B(n3579), .Z(n3634) );
  XNOR U3724 ( .A(n3635), .B(n3634), .Z(n3637) );
  NAND U3725 ( .A(b[0]), .B(a[91]), .Z(n3581) );
  XNOR U3726 ( .A(b[1]), .B(n3581), .Z(n3583) );
  NANDN U3727 ( .A(b[0]), .B(a[90]), .Z(n3582) );
  NAND U3728 ( .A(n3583), .B(n3582), .Z(n3631) );
  NAND U3729 ( .A(n25), .B(n3584), .Z(n3586) );
  XOR U3730 ( .A(b[5]), .B(a[87]), .Z(n3622) );
  NAND U3731 ( .A(n10456), .B(n3622), .Z(n3585) );
  AND U3732 ( .A(n3586), .B(n3585), .Z(n3629) );
  AND U3733 ( .A(b[7]), .B(a[83]), .Z(n3628) );
  XNOR U3734 ( .A(n3629), .B(n3628), .Z(n3630) );
  XNOR U3735 ( .A(n3631), .B(n3630), .Z(n3636) );
  XOR U3736 ( .A(n3637), .B(n3636), .Z(n3611) );
  NANDN U3737 ( .A(n3588), .B(n3587), .Z(n3592) );
  NANDN U3738 ( .A(n3590), .B(n3589), .Z(n3591) );
  AND U3739 ( .A(n3592), .B(n3591), .Z(n3610) );
  XNOR U3740 ( .A(n3611), .B(n3610), .Z(n3612) );
  NANDN U3741 ( .A(n3594), .B(n3593), .Z(n3598) );
  NAND U3742 ( .A(n3596), .B(n3595), .Z(n3597) );
  NAND U3743 ( .A(n3598), .B(n3597), .Z(n3613) );
  XNOR U3744 ( .A(n3612), .B(n3613), .Z(n3604) );
  XNOR U3745 ( .A(n3605), .B(n3604), .Z(n3606) );
  XNOR U3746 ( .A(n3607), .B(n3606), .Z(n3640) );
  XNOR U3747 ( .A(sreg[339]), .B(n3640), .Z(n3642) );
  NANDN U3748 ( .A(sreg[338]), .B(n3599), .Z(n3603) );
  NAND U3749 ( .A(n3601), .B(n3600), .Z(n3602) );
  NAND U3750 ( .A(n3603), .B(n3602), .Z(n3641) );
  XNOR U3751 ( .A(n3642), .B(n3641), .Z(c[339]) );
  NANDN U3752 ( .A(n3605), .B(n3604), .Z(n3609) );
  NANDN U3753 ( .A(n3607), .B(n3606), .Z(n3608) );
  AND U3754 ( .A(n3609), .B(n3608), .Z(n3648) );
  NANDN U3755 ( .A(n3611), .B(n3610), .Z(n3615) );
  NANDN U3756 ( .A(n3613), .B(n3612), .Z(n3614) );
  AND U3757 ( .A(n3615), .B(n3614), .Z(n3646) );
  NAND U3758 ( .A(n26), .B(n3616), .Z(n3618) );
  XOR U3759 ( .A(b[7]), .B(a[86]), .Z(n3657) );
  NAND U3760 ( .A(n10531), .B(n3657), .Z(n3617) );
  AND U3761 ( .A(n3618), .B(n3617), .Z(n3676) );
  NAND U3762 ( .A(n23), .B(n3619), .Z(n3621) );
  XOR U3763 ( .A(b[3]), .B(a[90]), .Z(n3660) );
  NAND U3764 ( .A(n24), .B(n3660), .Z(n3620) );
  NAND U3765 ( .A(n3621), .B(n3620), .Z(n3675) );
  XNOR U3766 ( .A(n3676), .B(n3675), .Z(n3678) );
  NAND U3767 ( .A(n25), .B(n3622), .Z(n3624) );
  XOR U3768 ( .A(b[5]), .B(a[88]), .Z(n3666) );
  NAND U3769 ( .A(n10456), .B(n3666), .Z(n3623) );
  AND U3770 ( .A(n3624), .B(n3623), .Z(n3670) );
  AND U3771 ( .A(b[7]), .B(a[84]), .Z(n3669) );
  XNOR U3772 ( .A(n3670), .B(n3669), .Z(n3671) );
  NAND U3773 ( .A(b[0]), .B(a[92]), .Z(n3625) );
  XNOR U3774 ( .A(b[1]), .B(n3625), .Z(n3627) );
  NANDN U3775 ( .A(b[0]), .B(a[91]), .Z(n3626) );
  NAND U3776 ( .A(n3627), .B(n3626), .Z(n3672) );
  XNOR U3777 ( .A(n3671), .B(n3672), .Z(n3677) );
  XOR U3778 ( .A(n3678), .B(n3677), .Z(n3652) );
  NANDN U3779 ( .A(n3629), .B(n3628), .Z(n3633) );
  NANDN U3780 ( .A(n3631), .B(n3630), .Z(n3632) );
  AND U3781 ( .A(n3633), .B(n3632), .Z(n3651) );
  XNOR U3782 ( .A(n3652), .B(n3651), .Z(n3653) );
  NANDN U3783 ( .A(n3635), .B(n3634), .Z(n3639) );
  NAND U3784 ( .A(n3637), .B(n3636), .Z(n3638) );
  NAND U3785 ( .A(n3639), .B(n3638), .Z(n3654) );
  XNOR U3786 ( .A(n3653), .B(n3654), .Z(n3645) );
  XNOR U3787 ( .A(n3646), .B(n3645), .Z(n3647) );
  XNOR U3788 ( .A(n3648), .B(n3647), .Z(n3681) );
  XNOR U3789 ( .A(sreg[340]), .B(n3681), .Z(n3683) );
  NANDN U3790 ( .A(sreg[339]), .B(n3640), .Z(n3644) );
  NAND U3791 ( .A(n3642), .B(n3641), .Z(n3643) );
  NAND U3792 ( .A(n3644), .B(n3643), .Z(n3682) );
  XNOR U3793 ( .A(n3683), .B(n3682), .Z(c[340]) );
  NANDN U3794 ( .A(n3646), .B(n3645), .Z(n3650) );
  NANDN U3795 ( .A(n3648), .B(n3647), .Z(n3649) );
  AND U3796 ( .A(n3650), .B(n3649), .Z(n3689) );
  NANDN U3797 ( .A(n3652), .B(n3651), .Z(n3656) );
  NANDN U3798 ( .A(n3654), .B(n3653), .Z(n3655) );
  AND U3799 ( .A(n3656), .B(n3655), .Z(n3687) );
  NAND U3800 ( .A(n26), .B(n3657), .Z(n3659) );
  XOR U3801 ( .A(b[7]), .B(a[87]), .Z(n3698) );
  NAND U3802 ( .A(n10531), .B(n3698), .Z(n3658) );
  AND U3803 ( .A(n3659), .B(n3658), .Z(n3717) );
  NAND U3804 ( .A(n23), .B(n3660), .Z(n3662) );
  XOR U3805 ( .A(b[3]), .B(a[91]), .Z(n3701) );
  NAND U3806 ( .A(n24), .B(n3701), .Z(n3661) );
  NAND U3807 ( .A(n3662), .B(n3661), .Z(n3716) );
  XNOR U3808 ( .A(n3717), .B(n3716), .Z(n3719) );
  NAND U3809 ( .A(b[0]), .B(a[93]), .Z(n3663) );
  XNOR U3810 ( .A(b[1]), .B(n3663), .Z(n3665) );
  NANDN U3811 ( .A(b[0]), .B(a[92]), .Z(n3664) );
  NAND U3812 ( .A(n3665), .B(n3664), .Z(n3713) );
  NAND U3813 ( .A(n25), .B(n3666), .Z(n3668) );
  XOR U3814 ( .A(b[5]), .B(a[89]), .Z(n3707) );
  NAND U3815 ( .A(n10456), .B(n3707), .Z(n3667) );
  AND U3816 ( .A(n3668), .B(n3667), .Z(n3711) );
  AND U3817 ( .A(b[7]), .B(a[85]), .Z(n3710) );
  XNOR U3818 ( .A(n3711), .B(n3710), .Z(n3712) );
  XNOR U3819 ( .A(n3713), .B(n3712), .Z(n3718) );
  XOR U3820 ( .A(n3719), .B(n3718), .Z(n3693) );
  NANDN U3821 ( .A(n3670), .B(n3669), .Z(n3674) );
  NANDN U3822 ( .A(n3672), .B(n3671), .Z(n3673) );
  AND U3823 ( .A(n3674), .B(n3673), .Z(n3692) );
  XNOR U3824 ( .A(n3693), .B(n3692), .Z(n3694) );
  NANDN U3825 ( .A(n3676), .B(n3675), .Z(n3680) );
  NAND U3826 ( .A(n3678), .B(n3677), .Z(n3679) );
  NAND U3827 ( .A(n3680), .B(n3679), .Z(n3695) );
  XNOR U3828 ( .A(n3694), .B(n3695), .Z(n3686) );
  XNOR U3829 ( .A(n3687), .B(n3686), .Z(n3688) );
  XNOR U3830 ( .A(n3689), .B(n3688), .Z(n3722) );
  XNOR U3831 ( .A(sreg[341]), .B(n3722), .Z(n3724) );
  NANDN U3832 ( .A(sreg[340]), .B(n3681), .Z(n3685) );
  NAND U3833 ( .A(n3683), .B(n3682), .Z(n3684) );
  NAND U3834 ( .A(n3685), .B(n3684), .Z(n3723) );
  XNOR U3835 ( .A(n3724), .B(n3723), .Z(c[341]) );
  NANDN U3836 ( .A(n3687), .B(n3686), .Z(n3691) );
  NANDN U3837 ( .A(n3689), .B(n3688), .Z(n3690) );
  AND U3838 ( .A(n3691), .B(n3690), .Z(n3730) );
  NANDN U3839 ( .A(n3693), .B(n3692), .Z(n3697) );
  NANDN U3840 ( .A(n3695), .B(n3694), .Z(n3696) );
  AND U3841 ( .A(n3697), .B(n3696), .Z(n3728) );
  NAND U3842 ( .A(n26), .B(n3698), .Z(n3700) );
  XOR U3843 ( .A(b[7]), .B(a[88]), .Z(n3739) );
  NAND U3844 ( .A(n10531), .B(n3739), .Z(n3699) );
  AND U3845 ( .A(n3700), .B(n3699), .Z(n3758) );
  NAND U3846 ( .A(n23), .B(n3701), .Z(n3703) );
  XOR U3847 ( .A(b[3]), .B(a[92]), .Z(n3742) );
  NAND U3848 ( .A(n24), .B(n3742), .Z(n3702) );
  NAND U3849 ( .A(n3703), .B(n3702), .Z(n3757) );
  XNOR U3850 ( .A(n3758), .B(n3757), .Z(n3760) );
  NAND U3851 ( .A(b[0]), .B(a[94]), .Z(n3704) );
  XNOR U3852 ( .A(b[1]), .B(n3704), .Z(n3706) );
  NANDN U3853 ( .A(b[0]), .B(a[93]), .Z(n3705) );
  NAND U3854 ( .A(n3706), .B(n3705), .Z(n3754) );
  NAND U3855 ( .A(n25), .B(n3707), .Z(n3709) );
  XOR U3856 ( .A(b[5]), .B(a[90]), .Z(n3748) );
  NAND U3857 ( .A(n10456), .B(n3748), .Z(n3708) );
  AND U3858 ( .A(n3709), .B(n3708), .Z(n3752) );
  AND U3859 ( .A(b[7]), .B(a[86]), .Z(n3751) );
  XNOR U3860 ( .A(n3752), .B(n3751), .Z(n3753) );
  XNOR U3861 ( .A(n3754), .B(n3753), .Z(n3759) );
  XOR U3862 ( .A(n3760), .B(n3759), .Z(n3734) );
  NANDN U3863 ( .A(n3711), .B(n3710), .Z(n3715) );
  NANDN U3864 ( .A(n3713), .B(n3712), .Z(n3714) );
  AND U3865 ( .A(n3715), .B(n3714), .Z(n3733) );
  XNOR U3866 ( .A(n3734), .B(n3733), .Z(n3735) );
  NANDN U3867 ( .A(n3717), .B(n3716), .Z(n3721) );
  NAND U3868 ( .A(n3719), .B(n3718), .Z(n3720) );
  NAND U3869 ( .A(n3721), .B(n3720), .Z(n3736) );
  XNOR U3870 ( .A(n3735), .B(n3736), .Z(n3727) );
  XNOR U3871 ( .A(n3728), .B(n3727), .Z(n3729) );
  XNOR U3872 ( .A(n3730), .B(n3729), .Z(n3763) );
  XNOR U3873 ( .A(sreg[342]), .B(n3763), .Z(n3765) );
  NANDN U3874 ( .A(sreg[341]), .B(n3722), .Z(n3726) );
  NAND U3875 ( .A(n3724), .B(n3723), .Z(n3725) );
  NAND U3876 ( .A(n3726), .B(n3725), .Z(n3764) );
  XNOR U3877 ( .A(n3765), .B(n3764), .Z(c[342]) );
  NANDN U3878 ( .A(n3728), .B(n3727), .Z(n3732) );
  NANDN U3879 ( .A(n3730), .B(n3729), .Z(n3731) );
  AND U3880 ( .A(n3732), .B(n3731), .Z(n3771) );
  NANDN U3881 ( .A(n3734), .B(n3733), .Z(n3738) );
  NANDN U3882 ( .A(n3736), .B(n3735), .Z(n3737) );
  AND U3883 ( .A(n3738), .B(n3737), .Z(n3769) );
  NAND U3884 ( .A(n26), .B(n3739), .Z(n3741) );
  XOR U3885 ( .A(b[7]), .B(a[89]), .Z(n3780) );
  NAND U3886 ( .A(n10531), .B(n3780), .Z(n3740) );
  AND U3887 ( .A(n3741), .B(n3740), .Z(n3799) );
  NAND U3888 ( .A(n23), .B(n3742), .Z(n3744) );
  XOR U3889 ( .A(b[3]), .B(a[93]), .Z(n3783) );
  NAND U3890 ( .A(n24), .B(n3783), .Z(n3743) );
  NAND U3891 ( .A(n3744), .B(n3743), .Z(n3798) );
  XNOR U3892 ( .A(n3799), .B(n3798), .Z(n3801) );
  NAND U3893 ( .A(b[0]), .B(a[95]), .Z(n3745) );
  XNOR U3894 ( .A(b[1]), .B(n3745), .Z(n3747) );
  NANDN U3895 ( .A(b[0]), .B(a[94]), .Z(n3746) );
  NAND U3896 ( .A(n3747), .B(n3746), .Z(n3795) );
  NAND U3897 ( .A(n25), .B(n3748), .Z(n3750) );
  XOR U3898 ( .A(b[5]), .B(a[91]), .Z(n3786) );
  NAND U3899 ( .A(n10456), .B(n3786), .Z(n3749) );
  AND U3900 ( .A(n3750), .B(n3749), .Z(n3793) );
  AND U3901 ( .A(b[7]), .B(a[87]), .Z(n3792) );
  XNOR U3902 ( .A(n3793), .B(n3792), .Z(n3794) );
  XNOR U3903 ( .A(n3795), .B(n3794), .Z(n3800) );
  XOR U3904 ( .A(n3801), .B(n3800), .Z(n3775) );
  NANDN U3905 ( .A(n3752), .B(n3751), .Z(n3756) );
  NANDN U3906 ( .A(n3754), .B(n3753), .Z(n3755) );
  AND U3907 ( .A(n3756), .B(n3755), .Z(n3774) );
  XNOR U3908 ( .A(n3775), .B(n3774), .Z(n3776) );
  NANDN U3909 ( .A(n3758), .B(n3757), .Z(n3762) );
  NAND U3910 ( .A(n3760), .B(n3759), .Z(n3761) );
  NAND U3911 ( .A(n3762), .B(n3761), .Z(n3777) );
  XNOR U3912 ( .A(n3776), .B(n3777), .Z(n3768) );
  XNOR U3913 ( .A(n3769), .B(n3768), .Z(n3770) );
  XNOR U3914 ( .A(n3771), .B(n3770), .Z(n3804) );
  XNOR U3915 ( .A(sreg[343]), .B(n3804), .Z(n3806) );
  NANDN U3916 ( .A(sreg[342]), .B(n3763), .Z(n3767) );
  NAND U3917 ( .A(n3765), .B(n3764), .Z(n3766) );
  NAND U3918 ( .A(n3767), .B(n3766), .Z(n3805) );
  XNOR U3919 ( .A(n3806), .B(n3805), .Z(c[343]) );
  NANDN U3920 ( .A(n3769), .B(n3768), .Z(n3773) );
  NANDN U3921 ( .A(n3771), .B(n3770), .Z(n3772) );
  AND U3922 ( .A(n3773), .B(n3772), .Z(n3812) );
  NANDN U3923 ( .A(n3775), .B(n3774), .Z(n3779) );
  NANDN U3924 ( .A(n3777), .B(n3776), .Z(n3778) );
  AND U3925 ( .A(n3779), .B(n3778), .Z(n3810) );
  NAND U3926 ( .A(n26), .B(n3780), .Z(n3782) );
  XOR U3927 ( .A(b[7]), .B(a[90]), .Z(n3821) );
  NAND U3928 ( .A(n10531), .B(n3821), .Z(n3781) );
  AND U3929 ( .A(n3782), .B(n3781), .Z(n3840) );
  NAND U3930 ( .A(n23), .B(n3783), .Z(n3785) );
  XOR U3931 ( .A(b[3]), .B(a[94]), .Z(n3824) );
  NAND U3932 ( .A(n24), .B(n3824), .Z(n3784) );
  NAND U3933 ( .A(n3785), .B(n3784), .Z(n3839) );
  XNOR U3934 ( .A(n3840), .B(n3839), .Z(n3842) );
  NAND U3935 ( .A(n25), .B(n3786), .Z(n3788) );
  XOR U3936 ( .A(b[5]), .B(a[92]), .Z(n3830) );
  NAND U3937 ( .A(n10456), .B(n3830), .Z(n3787) );
  AND U3938 ( .A(n3788), .B(n3787), .Z(n3834) );
  AND U3939 ( .A(b[7]), .B(a[88]), .Z(n3833) );
  XNOR U3940 ( .A(n3834), .B(n3833), .Z(n3835) );
  NAND U3941 ( .A(b[0]), .B(a[96]), .Z(n3789) );
  XNOR U3942 ( .A(b[1]), .B(n3789), .Z(n3791) );
  NANDN U3943 ( .A(b[0]), .B(a[95]), .Z(n3790) );
  NAND U3944 ( .A(n3791), .B(n3790), .Z(n3836) );
  XNOR U3945 ( .A(n3835), .B(n3836), .Z(n3841) );
  XOR U3946 ( .A(n3842), .B(n3841), .Z(n3816) );
  NANDN U3947 ( .A(n3793), .B(n3792), .Z(n3797) );
  NANDN U3948 ( .A(n3795), .B(n3794), .Z(n3796) );
  AND U3949 ( .A(n3797), .B(n3796), .Z(n3815) );
  XNOR U3950 ( .A(n3816), .B(n3815), .Z(n3817) );
  NANDN U3951 ( .A(n3799), .B(n3798), .Z(n3803) );
  NAND U3952 ( .A(n3801), .B(n3800), .Z(n3802) );
  NAND U3953 ( .A(n3803), .B(n3802), .Z(n3818) );
  XNOR U3954 ( .A(n3817), .B(n3818), .Z(n3809) );
  XNOR U3955 ( .A(n3810), .B(n3809), .Z(n3811) );
  XNOR U3956 ( .A(n3812), .B(n3811), .Z(n3845) );
  XNOR U3957 ( .A(sreg[344]), .B(n3845), .Z(n3847) );
  NANDN U3958 ( .A(sreg[343]), .B(n3804), .Z(n3808) );
  NAND U3959 ( .A(n3806), .B(n3805), .Z(n3807) );
  NAND U3960 ( .A(n3808), .B(n3807), .Z(n3846) );
  XNOR U3961 ( .A(n3847), .B(n3846), .Z(c[344]) );
  NANDN U3962 ( .A(n3810), .B(n3809), .Z(n3814) );
  NANDN U3963 ( .A(n3812), .B(n3811), .Z(n3813) );
  AND U3964 ( .A(n3814), .B(n3813), .Z(n3853) );
  NANDN U3965 ( .A(n3816), .B(n3815), .Z(n3820) );
  NANDN U3966 ( .A(n3818), .B(n3817), .Z(n3819) );
  AND U3967 ( .A(n3820), .B(n3819), .Z(n3851) );
  NAND U3968 ( .A(n26), .B(n3821), .Z(n3823) );
  XOR U3969 ( .A(b[7]), .B(a[91]), .Z(n3862) );
  NAND U3970 ( .A(n10531), .B(n3862), .Z(n3822) );
  AND U3971 ( .A(n3823), .B(n3822), .Z(n3881) );
  NAND U3972 ( .A(n23), .B(n3824), .Z(n3826) );
  XOR U3973 ( .A(b[3]), .B(a[95]), .Z(n3865) );
  NAND U3974 ( .A(n24), .B(n3865), .Z(n3825) );
  NAND U3975 ( .A(n3826), .B(n3825), .Z(n3880) );
  XNOR U3976 ( .A(n3881), .B(n3880), .Z(n3883) );
  NAND U3977 ( .A(b[0]), .B(a[97]), .Z(n3827) );
  XNOR U3978 ( .A(b[1]), .B(n3827), .Z(n3829) );
  NANDN U3979 ( .A(b[0]), .B(a[96]), .Z(n3828) );
  NAND U3980 ( .A(n3829), .B(n3828), .Z(n3877) );
  NAND U3981 ( .A(n25), .B(n3830), .Z(n3832) );
  XOR U3982 ( .A(b[5]), .B(a[93]), .Z(n3868) );
  NAND U3983 ( .A(n10456), .B(n3868), .Z(n3831) );
  AND U3984 ( .A(n3832), .B(n3831), .Z(n3875) );
  AND U3985 ( .A(b[7]), .B(a[89]), .Z(n3874) );
  XNOR U3986 ( .A(n3875), .B(n3874), .Z(n3876) );
  XNOR U3987 ( .A(n3877), .B(n3876), .Z(n3882) );
  XOR U3988 ( .A(n3883), .B(n3882), .Z(n3857) );
  NANDN U3989 ( .A(n3834), .B(n3833), .Z(n3838) );
  NANDN U3990 ( .A(n3836), .B(n3835), .Z(n3837) );
  AND U3991 ( .A(n3838), .B(n3837), .Z(n3856) );
  XNOR U3992 ( .A(n3857), .B(n3856), .Z(n3858) );
  NANDN U3993 ( .A(n3840), .B(n3839), .Z(n3844) );
  NAND U3994 ( .A(n3842), .B(n3841), .Z(n3843) );
  NAND U3995 ( .A(n3844), .B(n3843), .Z(n3859) );
  XNOR U3996 ( .A(n3858), .B(n3859), .Z(n3850) );
  XNOR U3997 ( .A(n3851), .B(n3850), .Z(n3852) );
  XNOR U3998 ( .A(n3853), .B(n3852), .Z(n3886) );
  XNOR U3999 ( .A(sreg[345]), .B(n3886), .Z(n3888) );
  NANDN U4000 ( .A(sreg[344]), .B(n3845), .Z(n3849) );
  NAND U4001 ( .A(n3847), .B(n3846), .Z(n3848) );
  NAND U4002 ( .A(n3849), .B(n3848), .Z(n3887) );
  XNOR U4003 ( .A(n3888), .B(n3887), .Z(c[345]) );
  NANDN U4004 ( .A(n3851), .B(n3850), .Z(n3855) );
  NANDN U4005 ( .A(n3853), .B(n3852), .Z(n3854) );
  AND U4006 ( .A(n3855), .B(n3854), .Z(n3894) );
  NANDN U4007 ( .A(n3857), .B(n3856), .Z(n3861) );
  NANDN U4008 ( .A(n3859), .B(n3858), .Z(n3860) );
  AND U4009 ( .A(n3861), .B(n3860), .Z(n3892) );
  NAND U4010 ( .A(n26), .B(n3862), .Z(n3864) );
  XOR U4011 ( .A(b[7]), .B(a[92]), .Z(n3903) );
  NAND U4012 ( .A(n10531), .B(n3903), .Z(n3863) );
  AND U4013 ( .A(n3864), .B(n3863), .Z(n3922) );
  NAND U4014 ( .A(n23), .B(n3865), .Z(n3867) );
  XOR U4015 ( .A(b[3]), .B(a[96]), .Z(n3906) );
  NAND U4016 ( .A(n24), .B(n3906), .Z(n3866) );
  NAND U4017 ( .A(n3867), .B(n3866), .Z(n3921) );
  XNOR U4018 ( .A(n3922), .B(n3921), .Z(n3924) );
  NAND U4019 ( .A(n25), .B(n3868), .Z(n3870) );
  XOR U4020 ( .A(b[5]), .B(a[94]), .Z(n3912) );
  NAND U4021 ( .A(n10456), .B(n3912), .Z(n3869) );
  AND U4022 ( .A(n3870), .B(n3869), .Z(n3916) );
  AND U4023 ( .A(b[7]), .B(a[90]), .Z(n3915) );
  XNOR U4024 ( .A(n3916), .B(n3915), .Z(n3917) );
  NAND U4025 ( .A(b[0]), .B(a[98]), .Z(n3871) );
  XNOR U4026 ( .A(b[1]), .B(n3871), .Z(n3873) );
  NANDN U4027 ( .A(b[0]), .B(a[97]), .Z(n3872) );
  NAND U4028 ( .A(n3873), .B(n3872), .Z(n3918) );
  XNOR U4029 ( .A(n3917), .B(n3918), .Z(n3923) );
  XOR U4030 ( .A(n3924), .B(n3923), .Z(n3898) );
  NANDN U4031 ( .A(n3875), .B(n3874), .Z(n3879) );
  NANDN U4032 ( .A(n3877), .B(n3876), .Z(n3878) );
  AND U4033 ( .A(n3879), .B(n3878), .Z(n3897) );
  XNOR U4034 ( .A(n3898), .B(n3897), .Z(n3899) );
  NANDN U4035 ( .A(n3881), .B(n3880), .Z(n3885) );
  NAND U4036 ( .A(n3883), .B(n3882), .Z(n3884) );
  NAND U4037 ( .A(n3885), .B(n3884), .Z(n3900) );
  XNOR U4038 ( .A(n3899), .B(n3900), .Z(n3891) );
  XNOR U4039 ( .A(n3892), .B(n3891), .Z(n3893) );
  XNOR U4040 ( .A(n3894), .B(n3893), .Z(n3927) );
  XNOR U4041 ( .A(sreg[346]), .B(n3927), .Z(n3929) );
  NANDN U4042 ( .A(sreg[345]), .B(n3886), .Z(n3890) );
  NAND U4043 ( .A(n3888), .B(n3887), .Z(n3889) );
  NAND U4044 ( .A(n3890), .B(n3889), .Z(n3928) );
  XNOR U4045 ( .A(n3929), .B(n3928), .Z(c[346]) );
  NANDN U4046 ( .A(n3892), .B(n3891), .Z(n3896) );
  NANDN U4047 ( .A(n3894), .B(n3893), .Z(n3895) );
  AND U4048 ( .A(n3896), .B(n3895), .Z(n3935) );
  NANDN U4049 ( .A(n3898), .B(n3897), .Z(n3902) );
  NANDN U4050 ( .A(n3900), .B(n3899), .Z(n3901) );
  AND U4051 ( .A(n3902), .B(n3901), .Z(n3933) );
  NAND U4052 ( .A(n26), .B(n3903), .Z(n3905) );
  XOR U4053 ( .A(b[7]), .B(a[93]), .Z(n3944) );
  NAND U4054 ( .A(n10531), .B(n3944), .Z(n3904) );
  AND U4055 ( .A(n3905), .B(n3904), .Z(n3963) );
  NAND U4056 ( .A(n23), .B(n3906), .Z(n3908) );
  XOR U4057 ( .A(b[3]), .B(a[97]), .Z(n3947) );
  NAND U4058 ( .A(n24), .B(n3947), .Z(n3907) );
  NAND U4059 ( .A(n3908), .B(n3907), .Z(n3962) );
  XNOR U4060 ( .A(n3963), .B(n3962), .Z(n3965) );
  NAND U4061 ( .A(b[0]), .B(a[99]), .Z(n3909) );
  XNOR U4062 ( .A(b[1]), .B(n3909), .Z(n3911) );
  NANDN U4063 ( .A(b[0]), .B(a[98]), .Z(n3910) );
  NAND U4064 ( .A(n3911), .B(n3910), .Z(n3959) );
  NAND U4065 ( .A(n25), .B(n3912), .Z(n3914) );
  XOR U4066 ( .A(b[5]), .B(a[95]), .Z(n3953) );
  NAND U4067 ( .A(n10456), .B(n3953), .Z(n3913) );
  AND U4068 ( .A(n3914), .B(n3913), .Z(n3957) );
  AND U4069 ( .A(b[7]), .B(a[91]), .Z(n3956) );
  XNOR U4070 ( .A(n3957), .B(n3956), .Z(n3958) );
  XNOR U4071 ( .A(n3959), .B(n3958), .Z(n3964) );
  XOR U4072 ( .A(n3965), .B(n3964), .Z(n3939) );
  NANDN U4073 ( .A(n3916), .B(n3915), .Z(n3920) );
  NANDN U4074 ( .A(n3918), .B(n3917), .Z(n3919) );
  AND U4075 ( .A(n3920), .B(n3919), .Z(n3938) );
  XNOR U4076 ( .A(n3939), .B(n3938), .Z(n3940) );
  NANDN U4077 ( .A(n3922), .B(n3921), .Z(n3926) );
  NAND U4078 ( .A(n3924), .B(n3923), .Z(n3925) );
  NAND U4079 ( .A(n3926), .B(n3925), .Z(n3941) );
  XNOR U4080 ( .A(n3940), .B(n3941), .Z(n3932) );
  XNOR U4081 ( .A(n3933), .B(n3932), .Z(n3934) );
  XNOR U4082 ( .A(n3935), .B(n3934), .Z(n3968) );
  XNOR U4083 ( .A(sreg[347]), .B(n3968), .Z(n3970) );
  NANDN U4084 ( .A(sreg[346]), .B(n3927), .Z(n3931) );
  NAND U4085 ( .A(n3929), .B(n3928), .Z(n3930) );
  NAND U4086 ( .A(n3931), .B(n3930), .Z(n3969) );
  XNOR U4087 ( .A(n3970), .B(n3969), .Z(c[347]) );
  NANDN U4088 ( .A(n3933), .B(n3932), .Z(n3937) );
  NANDN U4089 ( .A(n3935), .B(n3934), .Z(n3936) );
  AND U4090 ( .A(n3937), .B(n3936), .Z(n3976) );
  NANDN U4091 ( .A(n3939), .B(n3938), .Z(n3943) );
  NANDN U4092 ( .A(n3941), .B(n3940), .Z(n3942) );
  AND U4093 ( .A(n3943), .B(n3942), .Z(n3974) );
  NAND U4094 ( .A(n26), .B(n3944), .Z(n3946) );
  XOR U4095 ( .A(b[7]), .B(a[94]), .Z(n3985) );
  NAND U4096 ( .A(n10531), .B(n3985), .Z(n3945) );
  AND U4097 ( .A(n3946), .B(n3945), .Z(n4004) );
  NAND U4098 ( .A(n23), .B(n3947), .Z(n3949) );
  XOR U4099 ( .A(b[3]), .B(a[98]), .Z(n3988) );
  NAND U4100 ( .A(n24), .B(n3988), .Z(n3948) );
  NAND U4101 ( .A(n3949), .B(n3948), .Z(n4003) );
  XNOR U4102 ( .A(n4004), .B(n4003), .Z(n4006) );
  NAND U4103 ( .A(b[0]), .B(a[100]), .Z(n3950) );
  XNOR U4104 ( .A(b[1]), .B(n3950), .Z(n3952) );
  NANDN U4105 ( .A(b[0]), .B(a[99]), .Z(n3951) );
  NAND U4106 ( .A(n3952), .B(n3951), .Z(n4000) );
  NAND U4107 ( .A(n25), .B(n3953), .Z(n3955) );
  XOR U4108 ( .A(b[5]), .B(a[96]), .Z(n3994) );
  NAND U4109 ( .A(n10456), .B(n3994), .Z(n3954) );
  AND U4110 ( .A(n3955), .B(n3954), .Z(n3998) );
  AND U4111 ( .A(b[7]), .B(a[92]), .Z(n3997) );
  XNOR U4112 ( .A(n3998), .B(n3997), .Z(n3999) );
  XNOR U4113 ( .A(n4000), .B(n3999), .Z(n4005) );
  XOR U4114 ( .A(n4006), .B(n4005), .Z(n3980) );
  NANDN U4115 ( .A(n3957), .B(n3956), .Z(n3961) );
  NANDN U4116 ( .A(n3959), .B(n3958), .Z(n3960) );
  AND U4117 ( .A(n3961), .B(n3960), .Z(n3979) );
  XNOR U4118 ( .A(n3980), .B(n3979), .Z(n3981) );
  NANDN U4119 ( .A(n3963), .B(n3962), .Z(n3967) );
  NAND U4120 ( .A(n3965), .B(n3964), .Z(n3966) );
  NAND U4121 ( .A(n3967), .B(n3966), .Z(n3982) );
  XNOR U4122 ( .A(n3981), .B(n3982), .Z(n3973) );
  XNOR U4123 ( .A(n3974), .B(n3973), .Z(n3975) );
  XNOR U4124 ( .A(n3976), .B(n3975), .Z(n4009) );
  XNOR U4125 ( .A(sreg[348]), .B(n4009), .Z(n4011) );
  NANDN U4126 ( .A(sreg[347]), .B(n3968), .Z(n3972) );
  NAND U4127 ( .A(n3970), .B(n3969), .Z(n3971) );
  NAND U4128 ( .A(n3972), .B(n3971), .Z(n4010) );
  XNOR U4129 ( .A(n4011), .B(n4010), .Z(c[348]) );
  NANDN U4130 ( .A(n3974), .B(n3973), .Z(n3978) );
  NANDN U4131 ( .A(n3976), .B(n3975), .Z(n3977) );
  AND U4132 ( .A(n3978), .B(n3977), .Z(n4017) );
  NANDN U4133 ( .A(n3980), .B(n3979), .Z(n3984) );
  NANDN U4134 ( .A(n3982), .B(n3981), .Z(n3983) );
  AND U4135 ( .A(n3984), .B(n3983), .Z(n4015) );
  NAND U4136 ( .A(n26), .B(n3985), .Z(n3987) );
  XOR U4137 ( .A(b[7]), .B(a[95]), .Z(n4026) );
  NAND U4138 ( .A(n10531), .B(n4026), .Z(n3986) );
  AND U4139 ( .A(n3987), .B(n3986), .Z(n4045) );
  NAND U4140 ( .A(n23), .B(n3988), .Z(n3990) );
  XOR U4141 ( .A(b[3]), .B(a[99]), .Z(n4029) );
  NAND U4142 ( .A(n24), .B(n4029), .Z(n3989) );
  NAND U4143 ( .A(n3990), .B(n3989), .Z(n4044) );
  XNOR U4144 ( .A(n4045), .B(n4044), .Z(n4047) );
  NAND U4145 ( .A(b[0]), .B(a[101]), .Z(n3991) );
  XNOR U4146 ( .A(b[1]), .B(n3991), .Z(n3993) );
  NANDN U4147 ( .A(b[0]), .B(a[100]), .Z(n3992) );
  NAND U4148 ( .A(n3993), .B(n3992), .Z(n4041) );
  NAND U4149 ( .A(n25), .B(n3994), .Z(n3996) );
  XOR U4150 ( .A(b[5]), .B(a[97]), .Z(n4035) );
  NAND U4151 ( .A(n10456), .B(n4035), .Z(n3995) );
  AND U4152 ( .A(n3996), .B(n3995), .Z(n4039) );
  AND U4153 ( .A(b[7]), .B(a[93]), .Z(n4038) );
  XNOR U4154 ( .A(n4039), .B(n4038), .Z(n4040) );
  XNOR U4155 ( .A(n4041), .B(n4040), .Z(n4046) );
  XOR U4156 ( .A(n4047), .B(n4046), .Z(n4021) );
  NANDN U4157 ( .A(n3998), .B(n3997), .Z(n4002) );
  NANDN U4158 ( .A(n4000), .B(n3999), .Z(n4001) );
  AND U4159 ( .A(n4002), .B(n4001), .Z(n4020) );
  XNOR U4160 ( .A(n4021), .B(n4020), .Z(n4022) );
  NANDN U4161 ( .A(n4004), .B(n4003), .Z(n4008) );
  NAND U4162 ( .A(n4006), .B(n4005), .Z(n4007) );
  NAND U4163 ( .A(n4008), .B(n4007), .Z(n4023) );
  XNOR U4164 ( .A(n4022), .B(n4023), .Z(n4014) );
  XNOR U4165 ( .A(n4015), .B(n4014), .Z(n4016) );
  XNOR U4166 ( .A(n4017), .B(n4016), .Z(n4050) );
  XNOR U4167 ( .A(sreg[349]), .B(n4050), .Z(n4052) );
  NANDN U4168 ( .A(sreg[348]), .B(n4009), .Z(n4013) );
  NAND U4169 ( .A(n4011), .B(n4010), .Z(n4012) );
  NAND U4170 ( .A(n4013), .B(n4012), .Z(n4051) );
  XNOR U4171 ( .A(n4052), .B(n4051), .Z(c[349]) );
  NANDN U4172 ( .A(n4015), .B(n4014), .Z(n4019) );
  NANDN U4173 ( .A(n4017), .B(n4016), .Z(n4018) );
  AND U4174 ( .A(n4019), .B(n4018), .Z(n4058) );
  NANDN U4175 ( .A(n4021), .B(n4020), .Z(n4025) );
  NANDN U4176 ( .A(n4023), .B(n4022), .Z(n4024) );
  AND U4177 ( .A(n4025), .B(n4024), .Z(n4056) );
  NAND U4178 ( .A(n26), .B(n4026), .Z(n4028) );
  XOR U4179 ( .A(b[7]), .B(a[96]), .Z(n4067) );
  NAND U4180 ( .A(n10531), .B(n4067), .Z(n4027) );
  AND U4181 ( .A(n4028), .B(n4027), .Z(n4086) );
  NAND U4182 ( .A(n23), .B(n4029), .Z(n4031) );
  XOR U4183 ( .A(b[3]), .B(a[100]), .Z(n4070) );
  NAND U4184 ( .A(n24), .B(n4070), .Z(n4030) );
  NAND U4185 ( .A(n4031), .B(n4030), .Z(n4085) );
  XNOR U4186 ( .A(n4086), .B(n4085), .Z(n4088) );
  NAND U4187 ( .A(b[0]), .B(a[102]), .Z(n4032) );
  XNOR U4188 ( .A(b[1]), .B(n4032), .Z(n4034) );
  NANDN U4189 ( .A(b[0]), .B(a[101]), .Z(n4033) );
  NAND U4190 ( .A(n4034), .B(n4033), .Z(n4082) );
  NAND U4191 ( .A(n25), .B(n4035), .Z(n4037) );
  XOR U4192 ( .A(b[5]), .B(a[98]), .Z(n4076) );
  NAND U4193 ( .A(n10456), .B(n4076), .Z(n4036) );
  AND U4194 ( .A(n4037), .B(n4036), .Z(n4080) );
  AND U4195 ( .A(b[7]), .B(a[94]), .Z(n4079) );
  XNOR U4196 ( .A(n4080), .B(n4079), .Z(n4081) );
  XNOR U4197 ( .A(n4082), .B(n4081), .Z(n4087) );
  XOR U4198 ( .A(n4088), .B(n4087), .Z(n4062) );
  NANDN U4199 ( .A(n4039), .B(n4038), .Z(n4043) );
  NANDN U4200 ( .A(n4041), .B(n4040), .Z(n4042) );
  AND U4201 ( .A(n4043), .B(n4042), .Z(n4061) );
  XNOR U4202 ( .A(n4062), .B(n4061), .Z(n4063) );
  NANDN U4203 ( .A(n4045), .B(n4044), .Z(n4049) );
  NAND U4204 ( .A(n4047), .B(n4046), .Z(n4048) );
  NAND U4205 ( .A(n4049), .B(n4048), .Z(n4064) );
  XNOR U4206 ( .A(n4063), .B(n4064), .Z(n4055) );
  XNOR U4207 ( .A(n4056), .B(n4055), .Z(n4057) );
  XNOR U4208 ( .A(n4058), .B(n4057), .Z(n4091) );
  XNOR U4209 ( .A(sreg[350]), .B(n4091), .Z(n4093) );
  NANDN U4210 ( .A(sreg[349]), .B(n4050), .Z(n4054) );
  NAND U4211 ( .A(n4052), .B(n4051), .Z(n4053) );
  NAND U4212 ( .A(n4054), .B(n4053), .Z(n4092) );
  XNOR U4213 ( .A(n4093), .B(n4092), .Z(c[350]) );
  NANDN U4214 ( .A(n4056), .B(n4055), .Z(n4060) );
  NANDN U4215 ( .A(n4058), .B(n4057), .Z(n4059) );
  AND U4216 ( .A(n4060), .B(n4059), .Z(n4099) );
  NANDN U4217 ( .A(n4062), .B(n4061), .Z(n4066) );
  NANDN U4218 ( .A(n4064), .B(n4063), .Z(n4065) );
  AND U4219 ( .A(n4066), .B(n4065), .Z(n4097) );
  NAND U4220 ( .A(n26), .B(n4067), .Z(n4069) );
  XOR U4221 ( .A(b[7]), .B(a[97]), .Z(n4108) );
  NAND U4222 ( .A(n10531), .B(n4108), .Z(n4068) );
  AND U4223 ( .A(n4069), .B(n4068), .Z(n4127) );
  NAND U4224 ( .A(n23), .B(n4070), .Z(n4072) );
  XOR U4225 ( .A(b[3]), .B(a[101]), .Z(n4111) );
  NAND U4226 ( .A(n24), .B(n4111), .Z(n4071) );
  NAND U4227 ( .A(n4072), .B(n4071), .Z(n4126) );
  XNOR U4228 ( .A(n4127), .B(n4126), .Z(n4129) );
  NAND U4229 ( .A(b[0]), .B(a[103]), .Z(n4073) );
  XNOR U4230 ( .A(b[1]), .B(n4073), .Z(n4075) );
  NANDN U4231 ( .A(b[0]), .B(a[102]), .Z(n4074) );
  NAND U4232 ( .A(n4075), .B(n4074), .Z(n4123) );
  NAND U4233 ( .A(n25), .B(n4076), .Z(n4078) );
  XOR U4234 ( .A(b[5]), .B(a[99]), .Z(n4117) );
  NAND U4235 ( .A(n10456), .B(n4117), .Z(n4077) );
  AND U4236 ( .A(n4078), .B(n4077), .Z(n4121) );
  AND U4237 ( .A(b[7]), .B(a[95]), .Z(n4120) );
  XNOR U4238 ( .A(n4121), .B(n4120), .Z(n4122) );
  XNOR U4239 ( .A(n4123), .B(n4122), .Z(n4128) );
  XOR U4240 ( .A(n4129), .B(n4128), .Z(n4103) );
  NANDN U4241 ( .A(n4080), .B(n4079), .Z(n4084) );
  NANDN U4242 ( .A(n4082), .B(n4081), .Z(n4083) );
  AND U4243 ( .A(n4084), .B(n4083), .Z(n4102) );
  XNOR U4244 ( .A(n4103), .B(n4102), .Z(n4104) );
  NANDN U4245 ( .A(n4086), .B(n4085), .Z(n4090) );
  NAND U4246 ( .A(n4088), .B(n4087), .Z(n4089) );
  NAND U4247 ( .A(n4090), .B(n4089), .Z(n4105) );
  XNOR U4248 ( .A(n4104), .B(n4105), .Z(n4096) );
  XNOR U4249 ( .A(n4097), .B(n4096), .Z(n4098) );
  XNOR U4250 ( .A(n4099), .B(n4098), .Z(n4132) );
  XNOR U4251 ( .A(sreg[351]), .B(n4132), .Z(n4134) );
  NANDN U4252 ( .A(sreg[350]), .B(n4091), .Z(n4095) );
  NAND U4253 ( .A(n4093), .B(n4092), .Z(n4094) );
  NAND U4254 ( .A(n4095), .B(n4094), .Z(n4133) );
  XNOR U4255 ( .A(n4134), .B(n4133), .Z(c[351]) );
  NANDN U4256 ( .A(n4097), .B(n4096), .Z(n4101) );
  NANDN U4257 ( .A(n4099), .B(n4098), .Z(n4100) );
  AND U4258 ( .A(n4101), .B(n4100), .Z(n4140) );
  NANDN U4259 ( .A(n4103), .B(n4102), .Z(n4107) );
  NANDN U4260 ( .A(n4105), .B(n4104), .Z(n4106) );
  AND U4261 ( .A(n4107), .B(n4106), .Z(n4138) );
  NAND U4262 ( .A(n26), .B(n4108), .Z(n4110) );
  XOR U4263 ( .A(b[7]), .B(a[98]), .Z(n4149) );
  NAND U4264 ( .A(n10531), .B(n4149), .Z(n4109) );
  AND U4265 ( .A(n4110), .B(n4109), .Z(n4168) );
  NAND U4266 ( .A(n23), .B(n4111), .Z(n4113) );
  XOR U4267 ( .A(b[3]), .B(a[102]), .Z(n4152) );
  NAND U4268 ( .A(n24), .B(n4152), .Z(n4112) );
  NAND U4269 ( .A(n4113), .B(n4112), .Z(n4167) );
  XNOR U4270 ( .A(n4168), .B(n4167), .Z(n4170) );
  NAND U4271 ( .A(b[0]), .B(a[104]), .Z(n4114) );
  XNOR U4272 ( .A(b[1]), .B(n4114), .Z(n4116) );
  NANDN U4273 ( .A(b[0]), .B(a[103]), .Z(n4115) );
  NAND U4274 ( .A(n4116), .B(n4115), .Z(n4164) );
  NAND U4275 ( .A(n25), .B(n4117), .Z(n4119) );
  XOR U4276 ( .A(b[5]), .B(a[100]), .Z(n4158) );
  NAND U4277 ( .A(n10456), .B(n4158), .Z(n4118) );
  AND U4278 ( .A(n4119), .B(n4118), .Z(n4162) );
  AND U4279 ( .A(b[7]), .B(a[96]), .Z(n4161) );
  XNOR U4280 ( .A(n4162), .B(n4161), .Z(n4163) );
  XNOR U4281 ( .A(n4164), .B(n4163), .Z(n4169) );
  XOR U4282 ( .A(n4170), .B(n4169), .Z(n4144) );
  NANDN U4283 ( .A(n4121), .B(n4120), .Z(n4125) );
  NANDN U4284 ( .A(n4123), .B(n4122), .Z(n4124) );
  AND U4285 ( .A(n4125), .B(n4124), .Z(n4143) );
  XNOR U4286 ( .A(n4144), .B(n4143), .Z(n4145) );
  NANDN U4287 ( .A(n4127), .B(n4126), .Z(n4131) );
  NAND U4288 ( .A(n4129), .B(n4128), .Z(n4130) );
  NAND U4289 ( .A(n4131), .B(n4130), .Z(n4146) );
  XNOR U4290 ( .A(n4145), .B(n4146), .Z(n4137) );
  XNOR U4291 ( .A(n4138), .B(n4137), .Z(n4139) );
  XNOR U4292 ( .A(n4140), .B(n4139), .Z(n4173) );
  XNOR U4293 ( .A(sreg[352]), .B(n4173), .Z(n4175) );
  NANDN U4294 ( .A(sreg[351]), .B(n4132), .Z(n4136) );
  NAND U4295 ( .A(n4134), .B(n4133), .Z(n4135) );
  NAND U4296 ( .A(n4136), .B(n4135), .Z(n4174) );
  XNOR U4297 ( .A(n4175), .B(n4174), .Z(c[352]) );
  NANDN U4298 ( .A(n4138), .B(n4137), .Z(n4142) );
  NANDN U4299 ( .A(n4140), .B(n4139), .Z(n4141) );
  AND U4300 ( .A(n4142), .B(n4141), .Z(n4181) );
  NANDN U4301 ( .A(n4144), .B(n4143), .Z(n4148) );
  NANDN U4302 ( .A(n4146), .B(n4145), .Z(n4147) );
  AND U4303 ( .A(n4148), .B(n4147), .Z(n4179) );
  NAND U4304 ( .A(n26), .B(n4149), .Z(n4151) );
  XOR U4305 ( .A(b[7]), .B(a[99]), .Z(n4190) );
  NAND U4306 ( .A(n10531), .B(n4190), .Z(n4150) );
  AND U4307 ( .A(n4151), .B(n4150), .Z(n4209) );
  NAND U4308 ( .A(n23), .B(n4152), .Z(n4154) );
  XOR U4309 ( .A(b[3]), .B(a[103]), .Z(n4193) );
  NAND U4310 ( .A(n24), .B(n4193), .Z(n4153) );
  NAND U4311 ( .A(n4154), .B(n4153), .Z(n4208) );
  XNOR U4312 ( .A(n4209), .B(n4208), .Z(n4211) );
  NAND U4313 ( .A(b[0]), .B(a[105]), .Z(n4155) );
  XNOR U4314 ( .A(b[1]), .B(n4155), .Z(n4157) );
  NANDN U4315 ( .A(b[0]), .B(a[104]), .Z(n4156) );
  NAND U4316 ( .A(n4157), .B(n4156), .Z(n4205) );
  NAND U4317 ( .A(n25), .B(n4158), .Z(n4160) );
  XOR U4318 ( .A(b[5]), .B(a[101]), .Z(n4199) );
  NAND U4319 ( .A(n10456), .B(n4199), .Z(n4159) );
  AND U4320 ( .A(n4160), .B(n4159), .Z(n4203) );
  AND U4321 ( .A(b[7]), .B(a[97]), .Z(n4202) );
  XNOR U4322 ( .A(n4203), .B(n4202), .Z(n4204) );
  XNOR U4323 ( .A(n4205), .B(n4204), .Z(n4210) );
  XOR U4324 ( .A(n4211), .B(n4210), .Z(n4185) );
  NANDN U4325 ( .A(n4162), .B(n4161), .Z(n4166) );
  NANDN U4326 ( .A(n4164), .B(n4163), .Z(n4165) );
  AND U4327 ( .A(n4166), .B(n4165), .Z(n4184) );
  XNOR U4328 ( .A(n4185), .B(n4184), .Z(n4186) );
  NANDN U4329 ( .A(n4168), .B(n4167), .Z(n4172) );
  NAND U4330 ( .A(n4170), .B(n4169), .Z(n4171) );
  NAND U4331 ( .A(n4172), .B(n4171), .Z(n4187) );
  XNOR U4332 ( .A(n4186), .B(n4187), .Z(n4178) );
  XNOR U4333 ( .A(n4179), .B(n4178), .Z(n4180) );
  XNOR U4334 ( .A(n4181), .B(n4180), .Z(n4214) );
  XNOR U4335 ( .A(sreg[353]), .B(n4214), .Z(n4216) );
  NANDN U4336 ( .A(sreg[352]), .B(n4173), .Z(n4177) );
  NAND U4337 ( .A(n4175), .B(n4174), .Z(n4176) );
  NAND U4338 ( .A(n4177), .B(n4176), .Z(n4215) );
  XNOR U4339 ( .A(n4216), .B(n4215), .Z(c[353]) );
  NANDN U4340 ( .A(n4179), .B(n4178), .Z(n4183) );
  NANDN U4341 ( .A(n4181), .B(n4180), .Z(n4182) );
  AND U4342 ( .A(n4183), .B(n4182), .Z(n4222) );
  NANDN U4343 ( .A(n4185), .B(n4184), .Z(n4189) );
  NANDN U4344 ( .A(n4187), .B(n4186), .Z(n4188) );
  AND U4345 ( .A(n4189), .B(n4188), .Z(n4220) );
  NAND U4346 ( .A(n26), .B(n4190), .Z(n4192) );
  XOR U4347 ( .A(b[7]), .B(a[100]), .Z(n4231) );
  NAND U4348 ( .A(n10531), .B(n4231), .Z(n4191) );
  AND U4349 ( .A(n4192), .B(n4191), .Z(n4250) );
  NAND U4350 ( .A(n23), .B(n4193), .Z(n4195) );
  XOR U4351 ( .A(b[3]), .B(a[104]), .Z(n4234) );
  NAND U4352 ( .A(n24), .B(n4234), .Z(n4194) );
  NAND U4353 ( .A(n4195), .B(n4194), .Z(n4249) );
  XNOR U4354 ( .A(n4250), .B(n4249), .Z(n4252) );
  NAND U4355 ( .A(b[0]), .B(a[106]), .Z(n4196) );
  XNOR U4356 ( .A(b[1]), .B(n4196), .Z(n4198) );
  NANDN U4357 ( .A(b[0]), .B(a[105]), .Z(n4197) );
  NAND U4358 ( .A(n4198), .B(n4197), .Z(n4246) );
  NAND U4359 ( .A(n25), .B(n4199), .Z(n4201) );
  XOR U4360 ( .A(b[5]), .B(a[102]), .Z(n4240) );
  NAND U4361 ( .A(n10456), .B(n4240), .Z(n4200) );
  AND U4362 ( .A(n4201), .B(n4200), .Z(n4244) );
  AND U4363 ( .A(b[7]), .B(a[98]), .Z(n4243) );
  XNOR U4364 ( .A(n4244), .B(n4243), .Z(n4245) );
  XNOR U4365 ( .A(n4246), .B(n4245), .Z(n4251) );
  XOR U4366 ( .A(n4252), .B(n4251), .Z(n4226) );
  NANDN U4367 ( .A(n4203), .B(n4202), .Z(n4207) );
  NANDN U4368 ( .A(n4205), .B(n4204), .Z(n4206) );
  AND U4369 ( .A(n4207), .B(n4206), .Z(n4225) );
  XNOR U4370 ( .A(n4226), .B(n4225), .Z(n4227) );
  NANDN U4371 ( .A(n4209), .B(n4208), .Z(n4213) );
  NAND U4372 ( .A(n4211), .B(n4210), .Z(n4212) );
  NAND U4373 ( .A(n4213), .B(n4212), .Z(n4228) );
  XNOR U4374 ( .A(n4227), .B(n4228), .Z(n4219) );
  XNOR U4375 ( .A(n4220), .B(n4219), .Z(n4221) );
  XNOR U4376 ( .A(n4222), .B(n4221), .Z(n4255) );
  XNOR U4377 ( .A(sreg[354]), .B(n4255), .Z(n4257) );
  NANDN U4378 ( .A(sreg[353]), .B(n4214), .Z(n4218) );
  NAND U4379 ( .A(n4216), .B(n4215), .Z(n4217) );
  NAND U4380 ( .A(n4218), .B(n4217), .Z(n4256) );
  XNOR U4381 ( .A(n4257), .B(n4256), .Z(c[354]) );
  NANDN U4382 ( .A(n4220), .B(n4219), .Z(n4224) );
  NANDN U4383 ( .A(n4222), .B(n4221), .Z(n4223) );
  AND U4384 ( .A(n4224), .B(n4223), .Z(n4263) );
  NANDN U4385 ( .A(n4226), .B(n4225), .Z(n4230) );
  NANDN U4386 ( .A(n4228), .B(n4227), .Z(n4229) );
  AND U4387 ( .A(n4230), .B(n4229), .Z(n4261) );
  NAND U4388 ( .A(n26), .B(n4231), .Z(n4233) );
  XOR U4389 ( .A(b[7]), .B(a[101]), .Z(n4272) );
  NAND U4390 ( .A(n10531), .B(n4272), .Z(n4232) );
  AND U4391 ( .A(n4233), .B(n4232), .Z(n4291) );
  NAND U4392 ( .A(n23), .B(n4234), .Z(n4236) );
  XOR U4393 ( .A(b[3]), .B(a[105]), .Z(n4275) );
  NAND U4394 ( .A(n24), .B(n4275), .Z(n4235) );
  NAND U4395 ( .A(n4236), .B(n4235), .Z(n4290) );
  XNOR U4396 ( .A(n4291), .B(n4290), .Z(n4293) );
  NAND U4397 ( .A(b[0]), .B(a[107]), .Z(n4237) );
  XNOR U4398 ( .A(b[1]), .B(n4237), .Z(n4239) );
  NANDN U4399 ( .A(b[0]), .B(a[106]), .Z(n4238) );
  NAND U4400 ( .A(n4239), .B(n4238), .Z(n4287) );
  NAND U4401 ( .A(n25), .B(n4240), .Z(n4242) );
  XOR U4402 ( .A(b[5]), .B(a[103]), .Z(n4281) );
  NAND U4403 ( .A(n10456), .B(n4281), .Z(n4241) );
  AND U4404 ( .A(n4242), .B(n4241), .Z(n4285) );
  AND U4405 ( .A(b[7]), .B(a[99]), .Z(n4284) );
  XNOR U4406 ( .A(n4285), .B(n4284), .Z(n4286) );
  XNOR U4407 ( .A(n4287), .B(n4286), .Z(n4292) );
  XOR U4408 ( .A(n4293), .B(n4292), .Z(n4267) );
  NANDN U4409 ( .A(n4244), .B(n4243), .Z(n4248) );
  NANDN U4410 ( .A(n4246), .B(n4245), .Z(n4247) );
  AND U4411 ( .A(n4248), .B(n4247), .Z(n4266) );
  XNOR U4412 ( .A(n4267), .B(n4266), .Z(n4268) );
  NANDN U4413 ( .A(n4250), .B(n4249), .Z(n4254) );
  NAND U4414 ( .A(n4252), .B(n4251), .Z(n4253) );
  NAND U4415 ( .A(n4254), .B(n4253), .Z(n4269) );
  XNOR U4416 ( .A(n4268), .B(n4269), .Z(n4260) );
  XNOR U4417 ( .A(n4261), .B(n4260), .Z(n4262) );
  XNOR U4418 ( .A(n4263), .B(n4262), .Z(n4296) );
  XNOR U4419 ( .A(sreg[355]), .B(n4296), .Z(n4298) );
  NANDN U4420 ( .A(sreg[354]), .B(n4255), .Z(n4259) );
  NAND U4421 ( .A(n4257), .B(n4256), .Z(n4258) );
  NAND U4422 ( .A(n4259), .B(n4258), .Z(n4297) );
  XNOR U4423 ( .A(n4298), .B(n4297), .Z(c[355]) );
  NANDN U4424 ( .A(n4261), .B(n4260), .Z(n4265) );
  NANDN U4425 ( .A(n4263), .B(n4262), .Z(n4264) );
  AND U4426 ( .A(n4265), .B(n4264), .Z(n4304) );
  NANDN U4427 ( .A(n4267), .B(n4266), .Z(n4271) );
  NANDN U4428 ( .A(n4269), .B(n4268), .Z(n4270) );
  AND U4429 ( .A(n4271), .B(n4270), .Z(n4302) );
  NAND U4430 ( .A(n26), .B(n4272), .Z(n4274) );
  XOR U4431 ( .A(b[7]), .B(a[102]), .Z(n4313) );
  NAND U4432 ( .A(n10531), .B(n4313), .Z(n4273) );
  AND U4433 ( .A(n4274), .B(n4273), .Z(n4332) );
  NAND U4434 ( .A(n23), .B(n4275), .Z(n4277) );
  XOR U4435 ( .A(b[3]), .B(a[106]), .Z(n4316) );
  NAND U4436 ( .A(n24), .B(n4316), .Z(n4276) );
  NAND U4437 ( .A(n4277), .B(n4276), .Z(n4331) );
  XNOR U4438 ( .A(n4332), .B(n4331), .Z(n4334) );
  NAND U4439 ( .A(b[0]), .B(a[108]), .Z(n4278) );
  XNOR U4440 ( .A(b[1]), .B(n4278), .Z(n4280) );
  NANDN U4441 ( .A(b[0]), .B(a[107]), .Z(n4279) );
  NAND U4442 ( .A(n4280), .B(n4279), .Z(n4328) );
  NAND U4443 ( .A(n25), .B(n4281), .Z(n4283) );
  XOR U4444 ( .A(b[5]), .B(a[104]), .Z(n4322) );
  NAND U4445 ( .A(n10456), .B(n4322), .Z(n4282) );
  AND U4446 ( .A(n4283), .B(n4282), .Z(n4326) );
  AND U4447 ( .A(b[7]), .B(a[100]), .Z(n4325) );
  XNOR U4448 ( .A(n4326), .B(n4325), .Z(n4327) );
  XNOR U4449 ( .A(n4328), .B(n4327), .Z(n4333) );
  XOR U4450 ( .A(n4334), .B(n4333), .Z(n4308) );
  NANDN U4451 ( .A(n4285), .B(n4284), .Z(n4289) );
  NANDN U4452 ( .A(n4287), .B(n4286), .Z(n4288) );
  AND U4453 ( .A(n4289), .B(n4288), .Z(n4307) );
  XNOR U4454 ( .A(n4308), .B(n4307), .Z(n4309) );
  NANDN U4455 ( .A(n4291), .B(n4290), .Z(n4295) );
  NAND U4456 ( .A(n4293), .B(n4292), .Z(n4294) );
  NAND U4457 ( .A(n4295), .B(n4294), .Z(n4310) );
  XNOR U4458 ( .A(n4309), .B(n4310), .Z(n4301) );
  XNOR U4459 ( .A(n4302), .B(n4301), .Z(n4303) );
  XNOR U4460 ( .A(n4304), .B(n4303), .Z(n4337) );
  XNOR U4461 ( .A(sreg[356]), .B(n4337), .Z(n4339) );
  NANDN U4462 ( .A(sreg[355]), .B(n4296), .Z(n4300) );
  NAND U4463 ( .A(n4298), .B(n4297), .Z(n4299) );
  NAND U4464 ( .A(n4300), .B(n4299), .Z(n4338) );
  XNOR U4465 ( .A(n4339), .B(n4338), .Z(c[356]) );
  NANDN U4466 ( .A(n4302), .B(n4301), .Z(n4306) );
  NANDN U4467 ( .A(n4304), .B(n4303), .Z(n4305) );
  AND U4468 ( .A(n4306), .B(n4305), .Z(n4345) );
  NANDN U4469 ( .A(n4308), .B(n4307), .Z(n4312) );
  NANDN U4470 ( .A(n4310), .B(n4309), .Z(n4311) );
  AND U4471 ( .A(n4312), .B(n4311), .Z(n4343) );
  NAND U4472 ( .A(n26), .B(n4313), .Z(n4315) );
  XOR U4473 ( .A(b[7]), .B(a[103]), .Z(n4354) );
  NAND U4474 ( .A(n10531), .B(n4354), .Z(n4314) );
  AND U4475 ( .A(n4315), .B(n4314), .Z(n4373) );
  NAND U4476 ( .A(n23), .B(n4316), .Z(n4318) );
  XOR U4477 ( .A(b[3]), .B(a[107]), .Z(n4357) );
  NAND U4478 ( .A(n24), .B(n4357), .Z(n4317) );
  NAND U4479 ( .A(n4318), .B(n4317), .Z(n4372) );
  XNOR U4480 ( .A(n4373), .B(n4372), .Z(n4375) );
  NAND U4481 ( .A(b[0]), .B(a[109]), .Z(n4319) );
  XNOR U4482 ( .A(b[1]), .B(n4319), .Z(n4321) );
  NANDN U4483 ( .A(b[0]), .B(a[108]), .Z(n4320) );
  NAND U4484 ( .A(n4321), .B(n4320), .Z(n4369) );
  NAND U4485 ( .A(n25), .B(n4322), .Z(n4324) );
  XOR U4486 ( .A(b[5]), .B(a[105]), .Z(n4363) );
  NAND U4487 ( .A(n10456), .B(n4363), .Z(n4323) );
  AND U4488 ( .A(n4324), .B(n4323), .Z(n4367) );
  AND U4489 ( .A(b[7]), .B(a[101]), .Z(n4366) );
  XNOR U4490 ( .A(n4367), .B(n4366), .Z(n4368) );
  XNOR U4491 ( .A(n4369), .B(n4368), .Z(n4374) );
  XOR U4492 ( .A(n4375), .B(n4374), .Z(n4349) );
  NANDN U4493 ( .A(n4326), .B(n4325), .Z(n4330) );
  NANDN U4494 ( .A(n4328), .B(n4327), .Z(n4329) );
  AND U4495 ( .A(n4330), .B(n4329), .Z(n4348) );
  XNOR U4496 ( .A(n4349), .B(n4348), .Z(n4350) );
  NANDN U4497 ( .A(n4332), .B(n4331), .Z(n4336) );
  NAND U4498 ( .A(n4334), .B(n4333), .Z(n4335) );
  NAND U4499 ( .A(n4336), .B(n4335), .Z(n4351) );
  XNOR U4500 ( .A(n4350), .B(n4351), .Z(n4342) );
  XNOR U4501 ( .A(n4343), .B(n4342), .Z(n4344) );
  XNOR U4502 ( .A(n4345), .B(n4344), .Z(n4378) );
  XNOR U4503 ( .A(sreg[357]), .B(n4378), .Z(n4380) );
  NANDN U4504 ( .A(sreg[356]), .B(n4337), .Z(n4341) );
  NAND U4505 ( .A(n4339), .B(n4338), .Z(n4340) );
  NAND U4506 ( .A(n4341), .B(n4340), .Z(n4379) );
  XNOR U4507 ( .A(n4380), .B(n4379), .Z(c[357]) );
  NANDN U4508 ( .A(n4343), .B(n4342), .Z(n4347) );
  NANDN U4509 ( .A(n4345), .B(n4344), .Z(n4346) );
  AND U4510 ( .A(n4347), .B(n4346), .Z(n4386) );
  NANDN U4511 ( .A(n4349), .B(n4348), .Z(n4353) );
  NANDN U4512 ( .A(n4351), .B(n4350), .Z(n4352) );
  AND U4513 ( .A(n4353), .B(n4352), .Z(n4384) );
  NAND U4514 ( .A(n26), .B(n4354), .Z(n4356) );
  XOR U4515 ( .A(b[7]), .B(a[104]), .Z(n4395) );
  NAND U4516 ( .A(n10531), .B(n4395), .Z(n4355) );
  AND U4517 ( .A(n4356), .B(n4355), .Z(n4414) );
  NAND U4518 ( .A(n23), .B(n4357), .Z(n4359) );
  XOR U4519 ( .A(b[3]), .B(a[108]), .Z(n4398) );
  NAND U4520 ( .A(n24), .B(n4398), .Z(n4358) );
  NAND U4521 ( .A(n4359), .B(n4358), .Z(n4413) );
  XNOR U4522 ( .A(n4414), .B(n4413), .Z(n4416) );
  NAND U4523 ( .A(b[0]), .B(a[110]), .Z(n4360) );
  XNOR U4524 ( .A(b[1]), .B(n4360), .Z(n4362) );
  NANDN U4525 ( .A(b[0]), .B(a[109]), .Z(n4361) );
  NAND U4526 ( .A(n4362), .B(n4361), .Z(n4410) );
  NAND U4527 ( .A(n25), .B(n4363), .Z(n4365) );
  XOR U4528 ( .A(b[5]), .B(a[106]), .Z(n4404) );
  NAND U4529 ( .A(n10456), .B(n4404), .Z(n4364) );
  AND U4530 ( .A(n4365), .B(n4364), .Z(n4408) );
  AND U4531 ( .A(b[7]), .B(a[102]), .Z(n4407) );
  XNOR U4532 ( .A(n4408), .B(n4407), .Z(n4409) );
  XNOR U4533 ( .A(n4410), .B(n4409), .Z(n4415) );
  XOR U4534 ( .A(n4416), .B(n4415), .Z(n4390) );
  NANDN U4535 ( .A(n4367), .B(n4366), .Z(n4371) );
  NANDN U4536 ( .A(n4369), .B(n4368), .Z(n4370) );
  AND U4537 ( .A(n4371), .B(n4370), .Z(n4389) );
  XNOR U4538 ( .A(n4390), .B(n4389), .Z(n4391) );
  NANDN U4539 ( .A(n4373), .B(n4372), .Z(n4377) );
  NAND U4540 ( .A(n4375), .B(n4374), .Z(n4376) );
  NAND U4541 ( .A(n4377), .B(n4376), .Z(n4392) );
  XNOR U4542 ( .A(n4391), .B(n4392), .Z(n4383) );
  XNOR U4543 ( .A(n4384), .B(n4383), .Z(n4385) );
  XNOR U4544 ( .A(n4386), .B(n4385), .Z(n4419) );
  XNOR U4545 ( .A(sreg[358]), .B(n4419), .Z(n4421) );
  NANDN U4546 ( .A(sreg[357]), .B(n4378), .Z(n4382) );
  NAND U4547 ( .A(n4380), .B(n4379), .Z(n4381) );
  NAND U4548 ( .A(n4382), .B(n4381), .Z(n4420) );
  XNOR U4549 ( .A(n4421), .B(n4420), .Z(c[358]) );
  NANDN U4550 ( .A(n4384), .B(n4383), .Z(n4388) );
  NANDN U4551 ( .A(n4386), .B(n4385), .Z(n4387) );
  AND U4552 ( .A(n4388), .B(n4387), .Z(n4427) );
  NANDN U4553 ( .A(n4390), .B(n4389), .Z(n4394) );
  NANDN U4554 ( .A(n4392), .B(n4391), .Z(n4393) );
  AND U4555 ( .A(n4394), .B(n4393), .Z(n4425) );
  NAND U4556 ( .A(n26), .B(n4395), .Z(n4397) );
  XOR U4557 ( .A(b[7]), .B(a[105]), .Z(n4436) );
  NAND U4558 ( .A(n10531), .B(n4436), .Z(n4396) );
  AND U4559 ( .A(n4397), .B(n4396), .Z(n4455) );
  NAND U4560 ( .A(n23), .B(n4398), .Z(n4400) );
  XOR U4561 ( .A(b[3]), .B(a[109]), .Z(n4439) );
  NAND U4562 ( .A(n24), .B(n4439), .Z(n4399) );
  NAND U4563 ( .A(n4400), .B(n4399), .Z(n4454) );
  XNOR U4564 ( .A(n4455), .B(n4454), .Z(n4457) );
  NAND U4565 ( .A(b[0]), .B(a[111]), .Z(n4401) );
  XNOR U4566 ( .A(b[1]), .B(n4401), .Z(n4403) );
  NANDN U4567 ( .A(b[0]), .B(a[110]), .Z(n4402) );
  NAND U4568 ( .A(n4403), .B(n4402), .Z(n4451) );
  NAND U4569 ( .A(n25), .B(n4404), .Z(n4406) );
  XOR U4570 ( .A(b[5]), .B(a[107]), .Z(n4445) );
  NAND U4571 ( .A(n10456), .B(n4445), .Z(n4405) );
  AND U4572 ( .A(n4406), .B(n4405), .Z(n4449) );
  AND U4573 ( .A(b[7]), .B(a[103]), .Z(n4448) );
  XNOR U4574 ( .A(n4449), .B(n4448), .Z(n4450) );
  XNOR U4575 ( .A(n4451), .B(n4450), .Z(n4456) );
  XOR U4576 ( .A(n4457), .B(n4456), .Z(n4431) );
  NANDN U4577 ( .A(n4408), .B(n4407), .Z(n4412) );
  NANDN U4578 ( .A(n4410), .B(n4409), .Z(n4411) );
  AND U4579 ( .A(n4412), .B(n4411), .Z(n4430) );
  XNOR U4580 ( .A(n4431), .B(n4430), .Z(n4432) );
  NANDN U4581 ( .A(n4414), .B(n4413), .Z(n4418) );
  NAND U4582 ( .A(n4416), .B(n4415), .Z(n4417) );
  NAND U4583 ( .A(n4418), .B(n4417), .Z(n4433) );
  XNOR U4584 ( .A(n4432), .B(n4433), .Z(n4424) );
  XNOR U4585 ( .A(n4425), .B(n4424), .Z(n4426) );
  XNOR U4586 ( .A(n4427), .B(n4426), .Z(n4460) );
  XNOR U4587 ( .A(sreg[359]), .B(n4460), .Z(n4462) );
  NANDN U4588 ( .A(sreg[358]), .B(n4419), .Z(n4423) );
  NAND U4589 ( .A(n4421), .B(n4420), .Z(n4422) );
  NAND U4590 ( .A(n4423), .B(n4422), .Z(n4461) );
  XNOR U4591 ( .A(n4462), .B(n4461), .Z(c[359]) );
  NANDN U4592 ( .A(n4425), .B(n4424), .Z(n4429) );
  NANDN U4593 ( .A(n4427), .B(n4426), .Z(n4428) );
  AND U4594 ( .A(n4429), .B(n4428), .Z(n4468) );
  NANDN U4595 ( .A(n4431), .B(n4430), .Z(n4435) );
  NANDN U4596 ( .A(n4433), .B(n4432), .Z(n4434) );
  AND U4597 ( .A(n4435), .B(n4434), .Z(n4466) );
  NAND U4598 ( .A(n26), .B(n4436), .Z(n4438) );
  XOR U4599 ( .A(b[7]), .B(a[106]), .Z(n4477) );
  NAND U4600 ( .A(n10531), .B(n4477), .Z(n4437) );
  AND U4601 ( .A(n4438), .B(n4437), .Z(n4496) );
  NAND U4602 ( .A(n23), .B(n4439), .Z(n4441) );
  XOR U4603 ( .A(b[3]), .B(a[110]), .Z(n4480) );
  NAND U4604 ( .A(n24), .B(n4480), .Z(n4440) );
  NAND U4605 ( .A(n4441), .B(n4440), .Z(n4495) );
  XNOR U4606 ( .A(n4496), .B(n4495), .Z(n4498) );
  NAND U4607 ( .A(b[0]), .B(a[112]), .Z(n4442) );
  XNOR U4608 ( .A(b[1]), .B(n4442), .Z(n4444) );
  NANDN U4609 ( .A(b[0]), .B(a[111]), .Z(n4443) );
  NAND U4610 ( .A(n4444), .B(n4443), .Z(n4492) );
  NAND U4611 ( .A(n25), .B(n4445), .Z(n4447) );
  XOR U4612 ( .A(b[5]), .B(a[108]), .Z(n4486) );
  NAND U4613 ( .A(n10456), .B(n4486), .Z(n4446) );
  AND U4614 ( .A(n4447), .B(n4446), .Z(n4490) );
  AND U4615 ( .A(b[7]), .B(a[104]), .Z(n4489) );
  XNOR U4616 ( .A(n4490), .B(n4489), .Z(n4491) );
  XNOR U4617 ( .A(n4492), .B(n4491), .Z(n4497) );
  XOR U4618 ( .A(n4498), .B(n4497), .Z(n4472) );
  NANDN U4619 ( .A(n4449), .B(n4448), .Z(n4453) );
  NANDN U4620 ( .A(n4451), .B(n4450), .Z(n4452) );
  AND U4621 ( .A(n4453), .B(n4452), .Z(n4471) );
  XNOR U4622 ( .A(n4472), .B(n4471), .Z(n4473) );
  NANDN U4623 ( .A(n4455), .B(n4454), .Z(n4459) );
  NAND U4624 ( .A(n4457), .B(n4456), .Z(n4458) );
  NAND U4625 ( .A(n4459), .B(n4458), .Z(n4474) );
  XNOR U4626 ( .A(n4473), .B(n4474), .Z(n4465) );
  XNOR U4627 ( .A(n4466), .B(n4465), .Z(n4467) );
  XNOR U4628 ( .A(n4468), .B(n4467), .Z(n4501) );
  XNOR U4629 ( .A(sreg[360]), .B(n4501), .Z(n4503) );
  NANDN U4630 ( .A(sreg[359]), .B(n4460), .Z(n4464) );
  NAND U4631 ( .A(n4462), .B(n4461), .Z(n4463) );
  NAND U4632 ( .A(n4464), .B(n4463), .Z(n4502) );
  XNOR U4633 ( .A(n4503), .B(n4502), .Z(c[360]) );
  NANDN U4634 ( .A(n4466), .B(n4465), .Z(n4470) );
  NANDN U4635 ( .A(n4468), .B(n4467), .Z(n4469) );
  AND U4636 ( .A(n4470), .B(n4469), .Z(n4509) );
  NANDN U4637 ( .A(n4472), .B(n4471), .Z(n4476) );
  NANDN U4638 ( .A(n4474), .B(n4473), .Z(n4475) );
  AND U4639 ( .A(n4476), .B(n4475), .Z(n4507) );
  NAND U4640 ( .A(n26), .B(n4477), .Z(n4479) );
  XOR U4641 ( .A(b[7]), .B(a[107]), .Z(n4518) );
  NAND U4642 ( .A(n10531), .B(n4518), .Z(n4478) );
  AND U4643 ( .A(n4479), .B(n4478), .Z(n4537) );
  NAND U4644 ( .A(n23), .B(n4480), .Z(n4482) );
  XOR U4645 ( .A(b[3]), .B(a[111]), .Z(n4521) );
  NAND U4646 ( .A(n24), .B(n4521), .Z(n4481) );
  NAND U4647 ( .A(n4482), .B(n4481), .Z(n4536) );
  XNOR U4648 ( .A(n4537), .B(n4536), .Z(n4539) );
  NAND U4649 ( .A(b[0]), .B(a[113]), .Z(n4483) );
  XNOR U4650 ( .A(b[1]), .B(n4483), .Z(n4485) );
  NANDN U4651 ( .A(b[0]), .B(a[112]), .Z(n4484) );
  NAND U4652 ( .A(n4485), .B(n4484), .Z(n4533) );
  NAND U4653 ( .A(n25), .B(n4486), .Z(n4488) );
  XOR U4654 ( .A(b[5]), .B(a[109]), .Z(n4527) );
  NAND U4655 ( .A(n10456), .B(n4527), .Z(n4487) );
  AND U4656 ( .A(n4488), .B(n4487), .Z(n4531) );
  AND U4657 ( .A(b[7]), .B(a[105]), .Z(n4530) );
  XNOR U4658 ( .A(n4531), .B(n4530), .Z(n4532) );
  XNOR U4659 ( .A(n4533), .B(n4532), .Z(n4538) );
  XOR U4660 ( .A(n4539), .B(n4538), .Z(n4513) );
  NANDN U4661 ( .A(n4490), .B(n4489), .Z(n4494) );
  NANDN U4662 ( .A(n4492), .B(n4491), .Z(n4493) );
  AND U4663 ( .A(n4494), .B(n4493), .Z(n4512) );
  XNOR U4664 ( .A(n4513), .B(n4512), .Z(n4514) );
  NANDN U4665 ( .A(n4496), .B(n4495), .Z(n4500) );
  NAND U4666 ( .A(n4498), .B(n4497), .Z(n4499) );
  NAND U4667 ( .A(n4500), .B(n4499), .Z(n4515) );
  XNOR U4668 ( .A(n4514), .B(n4515), .Z(n4506) );
  XNOR U4669 ( .A(n4507), .B(n4506), .Z(n4508) );
  XNOR U4670 ( .A(n4509), .B(n4508), .Z(n4542) );
  XNOR U4671 ( .A(sreg[361]), .B(n4542), .Z(n4544) );
  NANDN U4672 ( .A(sreg[360]), .B(n4501), .Z(n4505) );
  NAND U4673 ( .A(n4503), .B(n4502), .Z(n4504) );
  NAND U4674 ( .A(n4505), .B(n4504), .Z(n4543) );
  XNOR U4675 ( .A(n4544), .B(n4543), .Z(c[361]) );
  NANDN U4676 ( .A(n4507), .B(n4506), .Z(n4511) );
  NANDN U4677 ( .A(n4509), .B(n4508), .Z(n4510) );
  AND U4678 ( .A(n4511), .B(n4510), .Z(n4550) );
  NANDN U4679 ( .A(n4513), .B(n4512), .Z(n4517) );
  NANDN U4680 ( .A(n4515), .B(n4514), .Z(n4516) );
  AND U4681 ( .A(n4517), .B(n4516), .Z(n4548) );
  NAND U4682 ( .A(n26), .B(n4518), .Z(n4520) );
  XOR U4683 ( .A(b[7]), .B(a[108]), .Z(n4559) );
  NAND U4684 ( .A(n10531), .B(n4559), .Z(n4519) );
  AND U4685 ( .A(n4520), .B(n4519), .Z(n4578) );
  NAND U4686 ( .A(n23), .B(n4521), .Z(n4523) );
  XOR U4687 ( .A(b[3]), .B(a[112]), .Z(n4562) );
  NAND U4688 ( .A(n24), .B(n4562), .Z(n4522) );
  NAND U4689 ( .A(n4523), .B(n4522), .Z(n4577) );
  XNOR U4690 ( .A(n4578), .B(n4577), .Z(n4580) );
  NAND U4691 ( .A(b[0]), .B(a[114]), .Z(n4524) );
  XNOR U4692 ( .A(b[1]), .B(n4524), .Z(n4526) );
  NANDN U4693 ( .A(b[0]), .B(a[113]), .Z(n4525) );
  NAND U4694 ( .A(n4526), .B(n4525), .Z(n4574) );
  NAND U4695 ( .A(n25), .B(n4527), .Z(n4529) );
  XOR U4696 ( .A(b[5]), .B(a[110]), .Z(n4568) );
  NAND U4697 ( .A(n10456), .B(n4568), .Z(n4528) );
  AND U4698 ( .A(n4529), .B(n4528), .Z(n4572) );
  AND U4699 ( .A(b[7]), .B(a[106]), .Z(n4571) );
  XNOR U4700 ( .A(n4572), .B(n4571), .Z(n4573) );
  XNOR U4701 ( .A(n4574), .B(n4573), .Z(n4579) );
  XOR U4702 ( .A(n4580), .B(n4579), .Z(n4554) );
  NANDN U4703 ( .A(n4531), .B(n4530), .Z(n4535) );
  NANDN U4704 ( .A(n4533), .B(n4532), .Z(n4534) );
  AND U4705 ( .A(n4535), .B(n4534), .Z(n4553) );
  XNOR U4706 ( .A(n4554), .B(n4553), .Z(n4555) );
  NANDN U4707 ( .A(n4537), .B(n4536), .Z(n4541) );
  NAND U4708 ( .A(n4539), .B(n4538), .Z(n4540) );
  NAND U4709 ( .A(n4541), .B(n4540), .Z(n4556) );
  XNOR U4710 ( .A(n4555), .B(n4556), .Z(n4547) );
  XNOR U4711 ( .A(n4548), .B(n4547), .Z(n4549) );
  XNOR U4712 ( .A(n4550), .B(n4549), .Z(n4583) );
  XNOR U4713 ( .A(sreg[362]), .B(n4583), .Z(n4585) );
  NANDN U4714 ( .A(sreg[361]), .B(n4542), .Z(n4546) );
  NAND U4715 ( .A(n4544), .B(n4543), .Z(n4545) );
  NAND U4716 ( .A(n4546), .B(n4545), .Z(n4584) );
  XNOR U4717 ( .A(n4585), .B(n4584), .Z(c[362]) );
  NANDN U4718 ( .A(n4548), .B(n4547), .Z(n4552) );
  NANDN U4719 ( .A(n4550), .B(n4549), .Z(n4551) );
  AND U4720 ( .A(n4552), .B(n4551), .Z(n4591) );
  NANDN U4721 ( .A(n4554), .B(n4553), .Z(n4558) );
  NANDN U4722 ( .A(n4556), .B(n4555), .Z(n4557) );
  AND U4723 ( .A(n4558), .B(n4557), .Z(n4589) );
  NAND U4724 ( .A(n26), .B(n4559), .Z(n4561) );
  XOR U4725 ( .A(b[7]), .B(a[109]), .Z(n4600) );
  NAND U4726 ( .A(n10531), .B(n4600), .Z(n4560) );
  AND U4727 ( .A(n4561), .B(n4560), .Z(n4619) );
  NAND U4728 ( .A(n23), .B(n4562), .Z(n4564) );
  XOR U4729 ( .A(b[3]), .B(a[113]), .Z(n4603) );
  NAND U4730 ( .A(n24), .B(n4603), .Z(n4563) );
  NAND U4731 ( .A(n4564), .B(n4563), .Z(n4618) );
  XNOR U4732 ( .A(n4619), .B(n4618), .Z(n4621) );
  NAND U4733 ( .A(b[0]), .B(a[115]), .Z(n4565) );
  XNOR U4734 ( .A(b[1]), .B(n4565), .Z(n4567) );
  NANDN U4735 ( .A(b[0]), .B(a[114]), .Z(n4566) );
  NAND U4736 ( .A(n4567), .B(n4566), .Z(n4615) );
  NAND U4737 ( .A(n25), .B(n4568), .Z(n4570) );
  XOR U4738 ( .A(b[5]), .B(a[111]), .Z(n4606) );
  NAND U4739 ( .A(n10456), .B(n4606), .Z(n4569) );
  AND U4740 ( .A(n4570), .B(n4569), .Z(n4613) );
  AND U4741 ( .A(b[7]), .B(a[107]), .Z(n4612) );
  XNOR U4742 ( .A(n4613), .B(n4612), .Z(n4614) );
  XNOR U4743 ( .A(n4615), .B(n4614), .Z(n4620) );
  XOR U4744 ( .A(n4621), .B(n4620), .Z(n4595) );
  NANDN U4745 ( .A(n4572), .B(n4571), .Z(n4576) );
  NANDN U4746 ( .A(n4574), .B(n4573), .Z(n4575) );
  AND U4747 ( .A(n4576), .B(n4575), .Z(n4594) );
  XNOR U4748 ( .A(n4595), .B(n4594), .Z(n4596) );
  NANDN U4749 ( .A(n4578), .B(n4577), .Z(n4582) );
  NAND U4750 ( .A(n4580), .B(n4579), .Z(n4581) );
  NAND U4751 ( .A(n4582), .B(n4581), .Z(n4597) );
  XNOR U4752 ( .A(n4596), .B(n4597), .Z(n4588) );
  XNOR U4753 ( .A(n4589), .B(n4588), .Z(n4590) );
  XNOR U4754 ( .A(n4591), .B(n4590), .Z(n4624) );
  XNOR U4755 ( .A(sreg[363]), .B(n4624), .Z(n4626) );
  NANDN U4756 ( .A(sreg[362]), .B(n4583), .Z(n4587) );
  NAND U4757 ( .A(n4585), .B(n4584), .Z(n4586) );
  NAND U4758 ( .A(n4587), .B(n4586), .Z(n4625) );
  XNOR U4759 ( .A(n4626), .B(n4625), .Z(c[363]) );
  NANDN U4760 ( .A(n4589), .B(n4588), .Z(n4593) );
  NANDN U4761 ( .A(n4591), .B(n4590), .Z(n4592) );
  AND U4762 ( .A(n4593), .B(n4592), .Z(n4632) );
  NANDN U4763 ( .A(n4595), .B(n4594), .Z(n4599) );
  NANDN U4764 ( .A(n4597), .B(n4596), .Z(n4598) );
  AND U4765 ( .A(n4599), .B(n4598), .Z(n4630) );
  NAND U4766 ( .A(n26), .B(n4600), .Z(n4602) );
  XOR U4767 ( .A(b[7]), .B(a[110]), .Z(n4641) );
  NAND U4768 ( .A(n10531), .B(n4641), .Z(n4601) );
  AND U4769 ( .A(n4602), .B(n4601), .Z(n4660) );
  NAND U4770 ( .A(n23), .B(n4603), .Z(n4605) );
  XOR U4771 ( .A(b[3]), .B(a[114]), .Z(n4644) );
  NAND U4772 ( .A(n24), .B(n4644), .Z(n4604) );
  NAND U4773 ( .A(n4605), .B(n4604), .Z(n4659) );
  XNOR U4774 ( .A(n4660), .B(n4659), .Z(n4662) );
  NAND U4775 ( .A(n25), .B(n4606), .Z(n4608) );
  XOR U4776 ( .A(b[5]), .B(a[112]), .Z(n4650) );
  NAND U4777 ( .A(n10456), .B(n4650), .Z(n4607) );
  AND U4778 ( .A(n4608), .B(n4607), .Z(n4654) );
  AND U4779 ( .A(b[7]), .B(a[108]), .Z(n4653) );
  XNOR U4780 ( .A(n4654), .B(n4653), .Z(n4655) );
  NAND U4781 ( .A(b[0]), .B(a[116]), .Z(n4609) );
  XNOR U4782 ( .A(b[1]), .B(n4609), .Z(n4611) );
  NANDN U4783 ( .A(b[0]), .B(a[115]), .Z(n4610) );
  NAND U4784 ( .A(n4611), .B(n4610), .Z(n4656) );
  XNOR U4785 ( .A(n4655), .B(n4656), .Z(n4661) );
  XOR U4786 ( .A(n4662), .B(n4661), .Z(n4636) );
  NANDN U4787 ( .A(n4613), .B(n4612), .Z(n4617) );
  NANDN U4788 ( .A(n4615), .B(n4614), .Z(n4616) );
  AND U4789 ( .A(n4617), .B(n4616), .Z(n4635) );
  XNOR U4790 ( .A(n4636), .B(n4635), .Z(n4637) );
  NANDN U4791 ( .A(n4619), .B(n4618), .Z(n4623) );
  NAND U4792 ( .A(n4621), .B(n4620), .Z(n4622) );
  NAND U4793 ( .A(n4623), .B(n4622), .Z(n4638) );
  XNOR U4794 ( .A(n4637), .B(n4638), .Z(n4629) );
  XNOR U4795 ( .A(n4630), .B(n4629), .Z(n4631) );
  XNOR U4796 ( .A(n4632), .B(n4631), .Z(n4665) );
  XNOR U4797 ( .A(sreg[364]), .B(n4665), .Z(n4667) );
  NANDN U4798 ( .A(sreg[363]), .B(n4624), .Z(n4628) );
  NAND U4799 ( .A(n4626), .B(n4625), .Z(n4627) );
  NAND U4800 ( .A(n4628), .B(n4627), .Z(n4666) );
  XNOR U4801 ( .A(n4667), .B(n4666), .Z(c[364]) );
  NANDN U4802 ( .A(n4630), .B(n4629), .Z(n4634) );
  NANDN U4803 ( .A(n4632), .B(n4631), .Z(n4633) );
  AND U4804 ( .A(n4634), .B(n4633), .Z(n4673) );
  NANDN U4805 ( .A(n4636), .B(n4635), .Z(n4640) );
  NANDN U4806 ( .A(n4638), .B(n4637), .Z(n4639) );
  AND U4807 ( .A(n4640), .B(n4639), .Z(n4671) );
  NAND U4808 ( .A(n26), .B(n4641), .Z(n4643) );
  XOR U4809 ( .A(b[7]), .B(a[111]), .Z(n4682) );
  NAND U4810 ( .A(n10531), .B(n4682), .Z(n4642) );
  AND U4811 ( .A(n4643), .B(n4642), .Z(n4701) );
  NAND U4812 ( .A(n23), .B(n4644), .Z(n4646) );
  XOR U4813 ( .A(b[3]), .B(a[115]), .Z(n4685) );
  NAND U4814 ( .A(n24), .B(n4685), .Z(n4645) );
  NAND U4815 ( .A(n4646), .B(n4645), .Z(n4700) );
  XNOR U4816 ( .A(n4701), .B(n4700), .Z(n4703) );
  NAND U4817 ( .A(b[0]), .B(a[117]), .Z(n4647) );
  XNOR U4818 ( .A(b[1]), .B(n4647), .Z(n4649) );
  NANDN U4819 ( .A(b[0]), .B(a[116]), .Z(n4648) );
  NAND U4820 ( .A(n4649), .B(n4648), .Z(n4697) );
  NAND U4821 ( .A(n25), .B(n4650), .Z(n4652) );
  XOR U4822 ( .A(b[5]), .B(a[113]), .Z(n4691) );
  NAND U4823 ( .A(n10456), .B(n4691), .Z(n4651) );
  AND U4824 ( .A(n4652), .B(n4651), .Z(n4695) );
  AND U4825 ( .A(b[7]), .B(a[109]), .Z(n4694) );
  XNOR U4826 ( .A(n4695), .B(n4694), .Z(n4696) );
  XNOR U4827 ( .A(n4697), .B(n4696), .Z(n4702) );
  XOR U4828 ( .A(n4703), .B(n4702), .Z(n4677) );
  NANDN U4829 ( .A(n4654), .B(n4653), .Z(n4658) );
  NANDN U4830 ( .A(n4656), .B(n4655), .Z(n4657) );
  AND U4831 ( .A(n4658), .B(n4657), .Z(n4676) );
  XNOR U4832 ( .A(n4677), .B(n4676), .Z(n4678) );
  NANDN U4833 ( .A(n4660), .B(n4659), .Z(n4664) );
  NAND U4834 ( .A(n4662), .B(n4661), .Z(n4663) );
  NAND U4835 ( .A(n4664), .B(n4663), .Z(n4679) );
  XNOR U4836 ( .A(n4678), .B(n4679), .Z(n4670) );
  XNOR U4837 ( .A(n4671), .B(n4670), .Z(n4672) );
  XNOR U4838 ( .A(n4673), .B(n4672), .Z(n4706) );
  XNOR U4839 ( .A(sreg[365]), .B(n4706), .Z(n4708) );
  NANDN U4840 ( .A(sreg[364]), .B(n4665), .Z(n4669) );
  NAND U4841 ( .A(n4667), .B(n4666), .Z(n4668) );
  NAND U4842 ( .A(n4669), .B(n4668), .Z(n4707) );
  XNOR U4843 ( .A(n4708), .B(n4707), .Z(c[365]) );
  NANDN U4844 ( .A(n4671), .B(n4670), .Z(n4675) );
  NANDN U4845 ( .A(n4673), .B(n4672), .Z(n4674) );
  AND U4846 ( .A(n4675), .B(n4674), .Z(n4714) );
  NANDN U4847 ( .A(n4677), .B(n4676), .Z(n4681) );
  NANDN U4848 ( .A(n4679), .B(n4678), .Z(n4680) );
  AND U4849 ( .A(n4681), .B(n4680), .Z(n4712) );
  NAND U4850 ( .A(n26), .B(n4682), .Z(n4684) );
  XOR U4851 ( .A(b[7]), .B(a[112]), .Z(n4723) );
  NAND U4852 ( .A(n10531), .B(n4723), .Z(n4683) );
  AND U4853 ( .A(n4684), .B(n4683), .Z(n4742) );
  NAND U4854 ( .A(n23), .B(n4685), .Z(n4687) );
  XOR U4855 ( .A(b[3]), .B(a[116]), .Z(n4726) );
  NAND U4856 ( .A(n24), .B(n4726), .Z(n4686) );
  NAND U4857 ( .A(n4687), .B(n4686), .Z(n4741) );
  XNOR U4858 ( .A(n4742), .B(n4741), .Z(n4744) );
  NAND U4859 ( .A(b[0]), .B(a[118]), .Z(n4688) );
  XNOR U4860 ( .A(b[1]), .B(n4688), .Z(n4690) );
  NANDN U4861 ( .A(b[0]), .B(a[117]), .Z(n4689) );
  NAND U4862 ( .A(n4690), .B(n4689), .Z(n4738) );
  NAND U4863 ( .A(n25), .B(n4691), .Z(n4693) );
  XOR U4864 ( .A(b[5]), .B(a[114]), .Z(n4729) );
  NAND U4865 ( .A(n10456), .B(n4729), .Z(n4692) );
  AND U4866 ( .A(n4693), .B(n4692), .Z(n4736) );
  AND U4867 ( .A(b[7]), .B(a[110]), .Z(n4735) );
  XNOR U4868 ( .A(n4736), .B(n4735), .Z(n4737) );
  XNOR U4869 ( .A(n4738), .B(n4737), .Z(n4743) );
  XOR U4870 ( .A(n4744), .B(n4743), .Z(n4718) );
  NANDN U4871 ( .A(n4695), .B(n4694), .Z(n4699) );
  NANDN U4872 ( .A(n4697), .B(n4696), .Z(n4698) );
  AND U4873 ( .A(n4699), .B(n4698), .Z(n4717) );
  XNOR U4874 ( .A(n4718), .B(n4717), .Z(n4719) );
  NANDN U4875 ( .A(n4701), .B(n4700), .Z(n4705) );
  NAND U4876 ( .A(n4703), .B(n4702), .Z(n4704) );
  NAND U4877 ( .A(n4705), .B(n4704), .Z(n4720) );
  XNOR U4878 ( .A(n4719), .B(n4720), .Z(n4711) );
  XNOR U4879 ( .A(n4712), .B(n4711), .Z(n4713) );
  XNOR U4880 ( .A(n4714), .B(n4713), .Z(n4747) );
  XNOR U4881 ( .A(sreg[366]), .B(n4747), .Z(n4749) );
  NANDN U4882 ( .A(sreg[365]), .B(n4706), .Z(n4710) );
  NAND U4883 ( .A(n4708), .B(n4707), .Z(n4709) );
  NAND U4884 ( .A(n4710), .B(n4709), .Z(n4748) );
  XNOR U4885 ( .A(n4749), .B(n4748), .Z(c[366]) );
  NANDN U4886 ( .A(n4712), .B(n4711), .Z(n4716) );
  NANDN U4887 ( .A(n4714), .B(n4713), .Z(n4715) );
  AND U4888 ( .A(n4716), .B(n4715), .Z(n4755) );
  NANDN U4889 ( .A(n4718), .B(n4717), .Z(n4722) );
  NANDN U4890 ( .A(n4720), .B(n4719), .Z(n4721) );
  AND U4891 ( .A(n4722), .B(n4721), .Z(n4753) );
  NAND U4892 ( .A(n26), .B(n4723), .Z(n4725) );
  XOR U4893 ( .A(b[7]), .B(a[113]), .Z(n4764) );
  NAND U4894 ( .A(n10531), .B(n4764), .Z(n4724) );
  AND U4895 ( .A(n4725), .B(n4724), .Z(n4783) );
  NAND U4896 ( .A(n23), .B(n4726), .Z(n4728) );
  XOR U4897 ( .A(b[3]), .B(a[117]), .Z(n4767) );
  NAND U4898 ( .A(n24), .B(n4767), .Z(n4727) );
  NAND U4899 ( .A(n4728), .B(n4727), .Z(n4782) );
  XNOR U4900 ( .A(n4783), .B(n4782), .Z(n4785) );
  NAND U4901 ( .A(n25), .B(n4729), .Z(n4731) );
  XOR U4902 ( .A(b[5]), .B(a[115]), .Z(n4773) );
  NAND U4903 ( .A(n10456), .B(n4773), .Z(n4730) );
  AND U4904 ( .A(n4731), .B(n4730), .Z(n4777) );
  AND U4905 ( .A(b[7]), .B(a[111]), .Z(n4776) );
  XNOR U4906 ( .A(n4777), .B(n4776), .Z(n4778) );
  NAND U4907 ( .A(b[0]), .B(a[119]), .Z(n4732) );
  XNOR U4908 ( .A(b[1]), .B(n4732), .Z(n4734) );
  NANDN U4909 ( .A(b[0]), .B(a[118]), .Z(n4733) );
  NAND U4910 ( .A(n4734), .B(n4733), .Z(n4779) );
  XNOR U4911 ( .A(n4778), .B(n4779), .Z(n4784) );
  XOR U4912 ( .A(n4785), .B(n4784), .Z(n4759) );
  NANDN U4913 ( .A(n4736), .B(n4735), .Z(n4740) );
  NANDN U4914 ( .A(n4738), .B(n4737), .Z(n4739) );
  AND U4915 ( .A(n4740), .B(n4739), .Z(n4758) );
  XNOR U4916 ( .A(n4759), .B(n4758), .Z(n4760) );
  NANDN U4917 ( .A(n4742), .B(n4741), .Z(n4746) );
  NAND U4918 ( .A(n4744), .B(n4743), .Z(n4745) );
  NAND U4919 ( .A(n4746), .B(n4745), .Z(n4761) );
  XNOR U4920 ( .A(n4760), .B(n4761), .Z(n4752) );
  XNOR U4921 ( .A(n4753), .B(n4752), .Z(n4754) );
  XNOR U4922 ( .A(n4755), .B(n4754), .Z(n4788) );
  XNOR U4923 ( .A(sreg[367]), .B(n4788), .Z(n4790) );
  NANDN U4924 ( .A(sreg[366]), .B(n4747), .Z(n4751) );
  NAND U4925 ( .A(n4749), .B(n4748), .Z(n4750) );
  NAND U4926 ( .A(n4751), .B(n4750), .Z(n4789) );
  XNOR U4927 ( .A(n4790), .B(n4789), .Z(c[367]) );
  NANDN U4928 ( .A(n4753), .B(n4752), .Z(n4757) );
  NANDN U4929 ( .A(n4755), .B(n4754), .Z(n4756) );
  AND U4930 ( .A(n4757), .B(n4756), .Z(n4796) );
  NANDN U4931 ( .A(n4759), .B(n4758), .Z(n4763) );
  NANDN U4932 ( .A(n4761), .B(n4760), .Z(n4762) );
  AND U4933 ( .A(n4763), .B(n4762), .Z(n4794) );
  NAND U4934 ( .A(n26), .B(n4764), .Z(n4766) );
  XOR U4935 ( .A(b[7]), .B(a[114]), .Z(n4805) );
  NAND U4936 ( .A(n10531), .B(n4805), .Z(n4765) );
  AND U4937 ( .A(n4766), .B(n4765), .Z(n4824) );
  NAND U4938 ( .A(n23), .B(n4767), .Z(n4769) );
  XOR U4939 ( .A(b[3]), .B(a[118]), .Z(n4808) );
  NAND U4940 ( .A(n24), .B(n4808), .Z(n4768) );
  NAND U4941 ( .A(n4769), .B(n4768), .Z(n4823) );
  XNOR U4942 ( .A(n4824), .B(n4823), .Z(n4826) );
  NAND U4943 ( .A(b[0]), .B(a[120]), .Z(n4770) );
  XNOR U4944 ( .A(b[1]), .B(n4770), .Z(n4772) );
  NANDN U4945 ( .A(b[0]), .B(a[119]), .Z(n4771) );
  NAND U4946 ( .A(n4772), .B(n4771), .Z(n4820) );
  NAND U4947 ( .A(n25), .B(n4773), .Z(n4775) );
  XOR U4948 ( .A(b[5]), .B(a[116]), .Z(n4814) );
  NAND U4949 ( .A(n10456), .B(n4814), .Z(n4774) );
  AND U4950 ( .A(n4775), .B(n4774), .Z(n4818) );
  AND U4951 ( .A(b[7]), .B(a[112]), .Z(n4817) );
  XNOR U4952 ( .A(n4818), .B(n4817), .Z(n4819) );
  XNOR U4953 ( .A(n4820), .B(n4819), .Z(n4825) );
  XOR U4954 ( .A(n4826), .B(n4825), .Z(n4800) );
  NANDN U4955 ( .A(n4777), .B(n4776), .Z(n4781) );
  NANDN U4956 ( .A(n4779), .B(n4778), .Z(n4780) );
  AND U4957 ( .A(n4781), .B(n4780), .Z(n4799) );
  XNOR U4958 ( .A(n4800), .B(n4799), .Z(n4801) );
  NANDN U4959 ( .A(n4783), .B(n4782), .Z(n4787) );
  NAND U4960 ( .A(n4785), .B(n4784), .Z(n4786) );
  NAND U4961 ( .A(n4787), .B(n4786), .Z(n4802) );
  XNOR U4962 ( .A(n4801), .B(n4802), .Z(n4793) );
  XNOR U4963 ( .A(n4794), .B(n4793), .Z(n4795) );
  XNOR U4964 ( .A(n4796), .B(n4795), .Z(n4829) );
  XNOR U4965 ( .A(sreg[368]), .B(n4829), .Z(n4831) );
  NANDN U4966 ( .A(sreg[367]), .B(n4788), .Z(n4792) );
  NAND U4967 ( .A(n4790), .B(n4789), .Z(n4791) );
  NAND U4968 ( .A(n4792), .B(n4791), .Z(n4830) );
  XNOR U4969 ( .A(n4831), .B(n4830), .Z(c[368]) );
  NANDN U4970 ( .A(n4794), .B(n4793), .Z(n4798) );
  NANDN U4971 ( .A(n4796), .B(n4795), .Z(n4797) );
  AND U4972 ( .A(n4798), .B(n4797), .Z(n4837) );
  NANDN U4973 ( .A(n4800), .B(n4799), .Z(n4804) );
  NANDN U4974 ( .A(n4802), .B(n4801), .Z(n4803) );
  AND U4975 ( .A(n4804), .B(n4803), .Z(n4835) );
  NAND U4976 ( .A(n26), .B(n4805), .Z(n4807) );
  XOR U4977 ( .A(b[7]), .B(a[115]), .Z(n4846) );
  NAND U4978 ( .A(n10531), .B(n4846), .Z(n4806) );
  AND U4979 ( .A(n4807), .B(n4806), .Z(n4865) );
  NAND U4980 ( .A(n23), .B(n4808), .Z(n4810) );
  XOR U4981 ( .A(b[3]), .B(a[119]), .Z(n4849) );
  NAND U4982 ( .A(n24), .B(n4849), .Z(n4809) );
  NAND U4983 ( .A(n4810), .B(n4809), .Z(n4864) );
  XNOR U4984 ( .A(n4865), .B(n4864), .Z(n4867) );
  NAND U4985 ( .A(b[0]), .B(a[121]), .Z(n4811) );
  XNOR U4986 ( .A(b[1]), .B(n4811), .Z(n4813) );
  NANDN U4987 ( .A(b[0]), .B(a[120]), .Z(n4812) );
  NAND U4988 ( .A(n4813), .B(n4812), .Z(n4861) );
  NAND U4989 ( .A(n25), .B(n4814), .Z(n4816) );
  XOR U4990 ( .A(b[5]), .B(a[117]), .Z(n4855) );
  NAND U4991 ( .A(n10456), .B(n4855), .Z(n4815) );
  AND U4992 ( .A(n4816), .B(n4815), .Z(n4859) );
  AND U4993 ( .A(b[7]), .B(a[113]), .Z(n4858) );
  XNOR U4994 ( .A(n4859), .B(n4858), .Z(n4860) );
  XNOR U4995 ( .A(n4861), .B(n4860), .Z(n4866) );
  XOR U4996 ( .A(n4867), .B(n4866), .Z(n4841) );
  NANDN U4997 ( .A(n4818), .B(n4817), .Z(n4822) );
  NANDN U4998 ( .A(n4820), .B(n4819), .Z(n4821) );
  AND U4999 ( .A(n4822), .B(n4821), .Z(n4840) );
  XNOR U5000 ( .A(n4841), .B(n4840), .Z(n4842) );
  NANDN U5001 ( .A(n4824), .B(n4823), .Z(n4828) );
  NAND U5002 ( .A(n4826), .B(n4825), .Z(n4827) );
  NAND U5003 ( .A(n4828), .B(n4827), .Z(n4843) );
  XNOR U5004 ( .A(n4842), .B(n4843), .Z(n4834) );
  XNOR U5005 ( .A(n4835), .B(n4834), .Z(n4836) );
  XNOR U5006 ( .A(n4837), .B(n4836), .Z(n4870) );
  XNOR U5007 ( .A(sreg[369]), .B(n4870), .Z(n4872) );
  NANDN U5008 ( .A(sreg[368]), .B(n4829), .Z(n4833) );
  NAND U5009 ( .A(n4831), .B(n4830), .Z(n4832) );
  NAND U5010 ( .A(n4833), .B(n4832), .Z(n4871) );
  XNOR U5011 ( .A(n4872), .B(n4871), .Z(c[369]) );
  NANDN U5012 ( .A(n4835), .B(n4834), .Z(n4839) );
  NANDN U5013 ( .A(n4837), .B(n4836), .Z(n4838) );
  AND U5014 ( .A(n4839), .B(n4838), .Z(n4878) );
  NANDN U5015 ( .A(n4841), .B(n4840), .Z(n4845) );
  NANDN U5016 ( .A(n4843), .B(n4842), .Z(n4844) );
  AND U5017 ( .A(n4845), .B(n4844), .Z(n4876) );
  NAND U5018 ( .A(n26), .B(n4846), .Z(n4848) );
  XOR U5019 ( .A(b[7]), .B(a[116]), .Z(n4887) );
  NAND U5020 ( .A(n10531), .B(n4887), .Z(n4847) );
  AND U5021 ( .A(n4848), .B(n4847), .Z(n4906) );
  NAND U5022 ( .A(n23), .B(n4849), .Z(n4851) );
  XOR U5023 ( .A(b[3]), .B(a[120]), .Z(n4890) );
  NAND U5024 ( .A(n24), .B(n4890), .Z(n4850) );
  NAND U5025 ( .A(n4851), .B(n4850), .Z(n4905) );
  XNOR U5026 ( .A(n4906), .B(n4905), .Z(n4908) );
  NAND U5027 ( .A(b[0]), .B(a[122]), .Z(n4852) );
  XNOR U5028 ( .A(b[1]), .B(n4852), .Z(n4854) );
  NANDN U5029 ( .A(b[0]), .B(a[121]), .Z(n4853) );
  NAND U5030 ( .A(n4854), .B(n4853), .Z(n4902) );
  NAND U5031 ( .A(n25), .B(n4855), .Z(n4857) );
  XOR U5032 ( .A(b[5]), .B(a[118]), .Z(n4896) );
  NAND U5033 ( .A(n10456), .B(n4896), .Z(n4856) );
  AND U5034 ( .A(n4857), .B(n4856), .Z(n4900) );
  AND U5035 ( .A(b[7]), .B(a[114]), .Z(n4899) );
  XNOR U5036 ( .A(n4900), .B(n4899), .Z(n4901) );
  XNOR U5037 ( .A(n4902), .B(n4901), .Z(n4907) );
  XOR U5038 ( .A(n4908), .B(n4907), .Z(n4882) );
  NANDN U5039 ( .A(n4859), .B(n4858), .Z(n4863) );
  NANDN U5040 ( .A(n4861), .B(n4860), .Z(n4862) );
  AND U5041 ( .A(n4863), .B(n4862), .Z(n4881) );
  XNOR U5042 ( .A(n4882), .B(n4881), .Z(n4883) );
  NANDN U5043 ( .A(n4865), .B(n4864), .Z(n4869) );
  NAND U5044 ( .A(n4867), .B(n4866), .Z(n4868) );
  NAND U5045 ( .A(n4869), .B(n4868), .Z(n4884) );
  XNOR U5046 ( .A(n4883), .B(n4884), .Z(n4875) );
  XNOR U5047 ( .A(n4876), .B(n4875), .Z(n4877) );
  XNOR U5048 ( .A(n4878), .B(n4877), .Z(n4911) );
  XNOR U5049 ( .A(sreg[370]), .B(n4911), .Z(n4913) );
  NANDN U5050 ( .A(sreg[369]), .B(n4870), .Z(n4874) );
  NAND U5051 ( .A(n4872), .B(n4871), .Z(n4873) );
  NAND U5052 ( .A(n4874), .B(n4873), .Z(n4912) );
  XNOR U5053 ( .A(n4913), .B(n4912), .Z(c[370]) );
  NANDN U5054 ( .A(n4876), .B(n4875), .Z(n4880) );
  NANDN U5055 ( .A(n4878), .B(n4877), .Z(n4879) );
  AND U5056 ( .A(n4880), .B(n4879), .Z(n4919) );
  NANDN U5057 ( .A(n4882), .B(n4881), .Z(n4886) );
  NANDN U5058 ( .A(n4884), .B(n4883), .Z(n4885) );
  AND U5059 ( .A(n4886), .B(n4885), .Z(n4917) );
  NAND U5060 ( .A(n26), .B(n4887), .Z(n4889) );
  XOR U5061 ( .A(b[7]), .B(a[117]), .Z(n4928) );
  NAND U5062 ( .A(n10531), .B(n4928), .Z(n4888) );
  AND U5063 ( .A(n4889), .B(n4888), .Z(n4947) );
  NAND U5064 ( .A(n23), .B(n4890), .Z(n4892) );
  XOR U5065 ( .A(b[3]), .B(a[121]), .Z(n4931) );
  NAND U5066 ( .A(n24), .B(n4931), .Z(n4891) );
  NAND U5067 ( .A(n4892), .B(n4891), .Z(n4946) );
  XNOR U5068 ( .A(n4947), .B(n4946), .Z(n4949) );
  NAND U5069 ( .A(b[0]), .B(a[123]), .Z(n4893) );
  XNOR U5070 ( .A(b[1]), .B(n4893), .Z(n4895) );
  NANDN U5071 ( .A(b[0]), .B(a[122]), .Z(n4894) );
  NAND U5072 ( .A(n4895), .B(n4894), .Z(n4943) );
  NAND U5073 ( .A(n25), .B(n4896), .Z(n4898) );
  XOR U5074 ( .A(b[5]), .B(a[119]), .Z(n4934) );
  NAND U5075 ( .A(n10456), .B(n4934), .Z(n4897) );
  AND U5076 ( .A(n4898), .B(n4897), .Z(n4941) );
  AND U5077 ( .A(b[7]), .B(a[115]), .Z(n4940) );
  XNOR U5078 ( .A(n4941), .B(n4940), .Z(n4942) );
  XNOR U5079 ( .A(n4943), .B(n4942), .Z(n4948) );
  XOR U5080 ( .A(n4949), .B(n4948), .Z(n4923) );
  NANDN U5081 ( .A(n4900), .B(n4899), .Z(n4904) );
  NANDN U5082 ( .A(n4902), .B(n4901), .Z(n4903) );
  AND U5083 ( .A(n4904), .B(n4903), .Z(n4922) );
  XNOR U5084 ( .A(n4923), .B(n4922), .Z(n4924) );
  NANDN U5085 ( .A(n4906), .B(n4905), .Z(n4910) );
  NAND U5086 ( .A(n4908), .B(n4907), .Z(n4909) );
  NAND U5087 ( .A(n4910), .B(n4909), .Z(n4925) );
  XNOR U5088 ( .A(n4924), .B(n4925), .Z(n4916) );
  XNOR U5089 ( .A(n4917), .B(n4916), .Z(n4918) );
  XNOR U5090 ( .A(n4919), .B(n4918), .Z(n4952) );
  XNOR U5091 ( .A(sreg[371]), .B(n4952), .Z(n4954) );
  NANDN U5092 ( .A(sreg[370]), .B(n4911), .Z(n4915) );
  NAND U5093 ( .A(n4913), .B(n4912), .Z(n4914) );
  NAND U5094 ( .A(n4915), .B(n4914), .Z(n4953) );
  XNOR U5095 ( .A(n4954), .B(n4953), .Z(c[371]) );
  NANDN U5096 ( .A(n4917), .B(n4916), .Z(n4921) );
  NANDN U5097 ( .A(n4919), .B(n4918), .Z(n4920) );
  AND U5098 ( .A(n4921), .B(n4920), .Z(n4960) );
  NANDN U5099 ( .A(n4923), .B(n4922), .Z(n4927) );
  NANDN U5100 ( .A(n4925), .B(n4924), .Z(n4926) );
  AND U5101 ( .A(n4927), .B(n4926), .Z(n4958) );
  NAND U5102 ( .A(n26), .B(n4928), .Z(n4930) );
  XOR U5103 ( .A(b[7]), .B(a[118]), .Z(n4969) );
  NAND U5104 ( .A(n10531), .B(n4969), .Z(n4929) );
  AND U5105 ( .A(n4930), .B(n4929), .Z(n4988) );
  NAND U5106 ( .A(n23), .B(n4931), .Z(n4933) );
  XOR U5107 ( .A(b[3]), .B(a[122]), .Z(n4972) );
  NAND U5108 ( .A(n24), .B(n4972), .Z(n4932) );
  NAND U5109 ( .A(n4933), .B(n4932), .Z(n4987) );
  XNOR U5110 ( .A(n4988), .B(n4987), .Z(n4990) );
  NAND U5111 ( .A(n25), .B(n4934), .Z(n4936) );
  XOR U5112 ( .A(b[5]), .B(a[120]), .Z(n4978) );
  NAND U5113 ( .A(n10456), .B(n4978), .Z(n4935) );
  AND U5114 ( .A(n4936), .B(n4935), .Z(n4982) );
  AND U5115 ( .A(b[7]), .B(a[116]), .Z(n4981) );
  XNOR U5116 ( .A(n4982), .B(n4981), .Z(n4983) );
  NAND U5117 ( .A(b[0]), .B(a[124]), .Z(n4937) );
  XNOR U5118 ( .A(b[1]), .B(n4937), .Z(n4939) );
  NANDN U5119 ( .A(b[0]), .B(a[123]), .Z(n4938) );
  NAND U5120 ( .A(n4939), .B(n4938), .Z(n4984) );
  XNOR U5121 ( .A(n4983), .B(n4984), .Z(n4989) );
  XOR U5122 ( .A(n4990), .B(n4989), .Z(n4964) );
  NANDN U5123 ( .A(n4941), .B(n4940), .Z(n4945) );
  NANDN U5124 ( .A(n4943), .B(n4942), .Z(n4944) );
  AND U5125 ( .A(n4945), .B(n4944), .Z(n4963) );
  XNOR U5126 ( .A(n4964), .B(n4963), .Z(n4965) );
  NANDN U5127 ( .A(n4947), .B(n4946), .Z(n4951) );
  NAND U5128 ( .A(n4949), .B(n4948), .Z(n4950) );
  NAND U5129 ( .A(n4951), .B(n4950), .Z(n4966) );
  XNOR U5130 ( .A(n4965), .B(n4966), .Z(n4957) );
  XNOR U5131 ( .A(n4958), .B(n4957), .Z(n4959) );
  XNOR U5132 ( .A(n4960), .B(n4959), .Z(n4993) );
  XNOR U5133 ( .A(sreg[372]), .B(n4993), .Z(n4995) );
  NANDN U5134 ( .A(sreg[371]), .B(n4952), .Z(n4956) );
  NAND U5135 ( .A(n4954), .B(n4953), .Z(n4955) );
  NAND U5136 ( .A(n4956), .B(n4955), .Z(n4994) );
  XNOR U5137 ( .A(n4995), .B(n4994), .Z(c[372]) );
  NANDN U5138 ( .A(n4958), .B(n4957), .Z(n4962) );
  NANDN U5139 ( .A(n4960), .B(n4959), .Z(n4961) );
  AND U5140 ( .A(n4962), .B(n4961), .Z(n5001) );
  NANDN U5141 ( .A(n4964), .B(n4963), .Z(n4968) );
  NANDN U5142 ( .A(n4966), .B(n4965), .Z(n4967) );
  AND U5143 ( .A(n4968), .B(n4967), .Z(n4999) );
  NAND U5144 ( .A(n26), .B(n4969), .Z(n4971) );
  XOR U5145 ( .A(b[7]), .B(a[119]), .Z(n5010) );
  NAND U5146 ( .A(n10531), .B(n5010), .Z(n4970) );
  AND U5147 ( .A(n4971), .B(n4970), .Z(n5029) );
  NAND U5148 ( .A(n23), .B(n4972), .Z(n4974) );
  XOR U5149 ( .A(b[3]), .B(a[123]), .Z(n5013) );
  NAND U5150 ( .A(n24), .B(n5013), .Z(n4973) );
  NAND U5151 ( .A(n4974), .B(n4973), .Z(n5028) );
  XNOR U5152 ( .A(n5029), .B(n5028), .Z(n5031) );
  NAND U5153 ( .A(b[0]), .B(a[125]), .Z(n4975) );
  XNOR U5154 ( .A(b[1]), .B(n4975), .Z(n4977) );
  NANDN U5155 ( .A(b[0]), .B(a[124]), .Z(n4976) );
  NAND U5156 ( .A(n4977), .B(n4976), .Z(n5025) );
  NAND U5157 ( .A(n25), .B(n4978), .Z(n4980) );
  XOR U5158 ( .A(b[5]), .B(a[121]), .Z(n5019) );
  NAND U5159 ( .A(n10456), .B(n5019), .Z(n4979) );
  AND U5160 ( .A(n4980), .B(n4979), .Z(n5023) );
  AND U5161 ( .A(b[7]), .B(a[117]), .Z(n5022) );
  XNOR U5162 ( .A(n5023), .B(n5022), .Z(n5024) );
  XNOR U5163 ( .A(n5025), .B(n5024), .Z(n5030) );
  XOR U5164 ( .A(n5031), .B(n5030), .Z(n5005) );
  NANDN U5165 ( .A(n4982), .B(n4981), .Z(n4986) );
  NANDN U5166 ( .A(n4984), .B(n4983), .Z(n4985) );
  AND U5167 ( .A(n4986), .B(n4985), .Z(n5004) );
  XNOR U5168 ( .A(n5005), .B(n5004), .Z(n5006) );
  NANDN U5169 ( .A(n4988), .B(n4987), .Z(n4992) );
  NAND U5170 ( .A(n4990), .B(n4989), .Z(n4991) );
  NAND U5171 ( .A(n4992), .B(n4991), .Z(n5007) );
  XNOR U5172 ( .A(n5006), .B(n5007), .Z(n4998) );
  XNOR U5173 ( .A(n4999), .B(n4998), .Z(n5000) );
  XNOR U5174 ( .A(n5001), .B(n5000), .Z(n5034) );
  XNOR U5175 ( .A(sreg[373]), .B(n5034), .Z(n5036) );
  NANDN U5176 ( .A(sreg[372]), .B(n4993), .Z(n4997) );
  NAND U5177 ( .A(n4995), .B(n4994), .Z(n4996) );
  NAND U5178 ( .A(n4997), .B(n4996), .Z(n5035) );
  XNOR U5179 ( .A(n5036), .B(n5035), .Z(c[373]) );
  NANDN U5180 ( .A(n4999), .B(n4998), .Z(n5003) );
  NANDN U5181 ( .A(n5001), .B(n5000), .Z(n5002) );
  AND U5182 ( .A(n5003), .B(n5002), .Z(n5042) );
  NANDN U5183 ( .A(n5005), .B(n5004), .Z(n5009) );
  NANDN U5184 ( .A(n5007), .B(n5006), .Z(n5008) );
  AND U5185 ( .A(n5009), .B(n5008), .Z(n5040) );
  NAND U5186 ( .A(n26), .B(n5010), .Z(n5012) );
  XOR U5187 ( .A(b[7]), .B(a[120]), .Z(n5051) );
  NAND U5188 ( .A(n10531), .B(n5051), .Z(n5011) );
  AND U5189 ( .A(n5012), .B(n5011), .Z(n5070) );
  NAND U5190 ( .A(n23), .B(n5013), .Z(n5015) );
  XOR U5191 ( .A(b[3]), .B(a[124]), .Z(n5054) );
  NAND U5192 ( .A(n24), .B(n5054), .Z(n5014) );
  NAND U5193 ( .A(n5015), .B(n5014), .Z(n5069) );
  XNOR U5194 ( .A(n5070), .B(n5069), .Z(n5072) );
  NAND U5195 ( .A(b[0]), .B(a[126]), .Z(n5016) );
  XNOR U5196 ( .A(b[1]), .B(n5016), .Z(n5018) );
  NANDN U5197 ( .A(b[0]), .B(a[125]), .Z(n5017) );
  NAND U5198 ( .A(n5018), .B(n5017), .Z(n5066) );
  NAND U5199 ( .A(n25), .B(n5019), .Z(n5021) );
  XOR U5200 ( .A(b[5]), .B(a[122]), .Z(n5060) );
  NAND U5201 ( .A(n10456), .B(n5060), .Z(n5020) );
  AND U5202 ( .A(n5021), .B(n5020), .Z(n5064) );
  AND U5203 ( .A(b[7]), .B(a[118]), .Z(n5063) );
  XNOR U5204 ( .A(n5064), .B(n5063), .Z(n5065) );
  XNOR U5205 ( .A(n5066), .B(n5065), .Z(n5071) );
  XOR U5206 ( .A(n5072), .B(n5071), .Z(n5046) );
  NANDN U5207 ( .A(n5023), .B(n5022), .Z(n5027) );
  NANDN U5208 ( .A(n5025), .B(n5024), .Z(n5026) );
  AND U5209 ( .A(n5027), .B(n5026), .Z(n5045) );
  XNOR U5210 ( .A(n5046), .B(n5045), .Z(n5047) );
  NANDN U5211 ( .A(n5029), .B(n5028), .Z(n5033) );
  NAND U5212 ( .A(n5031), .B(n5030), .Z(n5032) );
  NAND U5213 ( .A(n5033), .B(n5032), .Z(n5048) );
  XNOR U5214 ( .A(n5047), .B(n5048), .Z(n5039) );
  XNOR U5215 ( .A(n5040), .B(n5039), .Z(n5041) );
  XNOR U5216 ( .A(n5042), .B(n5041), .Z(n5075) );
  XNOR U5217 ( .A(sreg[374]), .B(n5075), .Z(n5077) );
  NANDN U5218 ( .A(sreg[373]), .B(n5034), .Z(n5038) );
  NAND U5219 ( .A(n5036), .B(n5035), .Z(n5037) );
  NAND U5220 ( .A(n5038), .B(n5037), .Z(n5076) );
  XNOR U5221 ( .A(n5077), .B(n5076), .Z(c[374]) );
  NANDN U5222 ( .A(n5040), .B(n5039), .Z(n5044) );
  NANDN U5223 ( .A(n5042), .B(n5041), .Z(n5043) );
  AND U5224 ( .A(n5044), .B(n5043), .Z(n5083) );
  NANDN U5225 ( .A(n5046), .B(n5045), .Z(n5050) );
  NANDN U5226 ( .A(n5048), .B(n5047), .Z(n5049) );
  AND U5227 ( .A(n5050), .B(n5049), .Z(n5081) );
  NAND U5228 ( .A(n26), .B(n5051), .Z(n5053) );
  XOR U5229 ( .A(b[7]), .B(a[121]), .Z(n5092) );
  NAND U5230 ( .A(n10531), .B(n5092), .Z(n5052) );
  AND U5231 ( .A(n5053), .B(n5052), .Z(n5111) );
  NAND U5232 ( .A(n23), .B(n5054), .Z(n5056) );
  XOR U5233 ( .A(b[3]), .B(a[125]), .Z(n5095) );
  NAND U5234 ( .A(n24), .B(n5095), .Z(n5055) );
  NAND U5235 ( .A(n5056), .B(n5055), .Z(n5110) );
  XNOR U5236 ( .A(n5111), .B(n5110), .Z(n5113) );
  NAND U5237 ( .A(b[0]), .B(a[127]), .Z(n5057) );
  XNOR U5238 ( .A(b[1]), .B(n5057), .Z(n5059) );
  NANDN U5239 ( .A(b[0]), .B(a[126]), .Z(n5058) );
  NAND U5240 ( .A(n5059), .B(n5058), .Z(n5107) );
  NAND U5241 ( .A(n25), .B(n5060), .Z(n5062) );
  XOR U5242 ( .A(b[5]), .B(a[123]), .Z(n5101) );
  NAND U5243 ( .A(n10456), .B(n5101), .Z(n5061) );
  AND U5244 ( .A(n5062), .B(n5061), .Z(n5105) );
  AND U5245 ( .A(b[7]), .B(a[119]), .Z(n5104) );
  XNOR U5246 ( .A(n5105), .B(n5104), .Z(n5106) );
  XNOR U5247 ( .A(n5107), .B(n5106), .Z(n5112) );
  XOR U5248 ( .A(n5113), .B(n5112), .Z(n5087) );
  NANDN U5249 ( .A(n5064), .B(n5063), .Z(n5068) );
  NANDN U5250 ( .A(n5066), .B(n5065), .Z(n5067) );
  AND U5251 ( .A(n5068), .B(n5067), .Z(n5086) );
  XNOR U5252 ( .A(n5087), .B(n5086), .Z(n5088) );
  NANDN U5253 ( .A(n5070), .B(n5069), .Z(n5074) );
  NAND U5254 ( .A(n5072), .B(n5071), .Z(n5073) );
  NAND U5255 ( .A(n5074), .B(n5073), .Z(n5089) );
  XNOR U5256 ( .A(n5088), .B(n5089), .Z(n5080) );
  XNOR U5257 ( .A(n5081), .B(n5080), .Z(n5082) );
  XNOR U5258 ( .A(n5083), .B(n5082), .Z(n5116) );
  XNOR U5259 ( .A(sreg[375]), .B(n5116), .Z(n5118) );
  NANDN U5260 ( .A(sreg[374]), .B(n5075), .Z(n5079) );
  NAND U5261 ( .A(n5077), .B(n5076), .Z(n5078) );
  NAND U5262 ( .A(n5079), .B(n5078), .Z(n5117) );
  XNOR U5263 ( .A(n5118), .B(n5117), .Z(c[375]) );
  NANDN U5264 ( .A(n5081), .B(n5080), .Z(n5085) );
  NANDN U5265 ( .A(n5083), .B(n5082), .Z(n5084) );
  AND U5266 ( .A(n5085), .B(n5084), .Z(n5124) );
  NANDN U5267 ( .A(n5087), .B(n5086), .Z(n5091) );
  NANDN U5268 ( .A(n5089), .B(n5088), .Z(n5090) );
  AND U5269 ( .A(n5091), .B(n5090), .Z(n5122) );
  NAND U5270 ( .A(n26), .B(n5092), .Z(n5094) );
  XOR U5271 ( .A(b[7]), .B(a[122]), .Z(n5133) );
  NAND U5272 ( .A(n10531), .B(n5133), .Z(n5093) );
  AND U5273 ( .A(n5094), .B(n5093), .Z(n5152) );
  NAND U5274 ( .A(n23), .B(n5095), .Z(n5097) );
  XOR U5275 ( .A(b[3]), .B(a[126]), .Z(n5136) );
  NAND U5276 ( .A(n24), .B(n5136), .Z(n5096) );
  NAND U5277 ( .A(n5097), .B(n5096), .Z(n5151) );
  XNOR U5278 ( .A(n5152), .B(n5151), .Z(n5154) );
  NAND U5279 ( .A(b[0]), .B(a[128]), .Z(n5098) );
  XNOR U5280 ( .A(b[1]), .B(n5098), .Z(n5100) );
  NANDN U5281 ( .A(b[0]), .B(a[127]), .Z(n5099) );
  NAND U5282 ( .A(n5100), .B(n5099), .Z(n5148) );
  NAND U5283 ( .A(n25), .B(n5101), .Z(n5103) );
  XOR U5284 ( .A(b[5]), .B(a[124]), .Z(n5142) );
  NAND U5285 ( .A(n10456), .B(n5142), .Z(n5102) );
  AND U5286 ( .A(n5103), .B(n5102), .Z(n5146) );
  AND U5287 ( .A(b[7]), .B(a[120]), .Z(n5145) );
  XNOR U5288 ( .A(n5146), .B(n5145), .Z(n5147) );
  XNOR U5289 ( .A(n5148), .B(n5147), .Z(n5153) );
  XOR U5290 ( .A(n5154), .B(n5153), .Z(n5128) );
  NANDN U5291 ( .A(n5105), .B(n5104), .Z(n5109) );
  NANDN U5292 ( .A(n5107), .B(n5106), .Z(n5108) );
  AND U5293 ( .A(n5109), .B(n5108), .Z(n5127) );
  XNOR U5294 ( .A(n5128), .B(n5127), .Z(n5129) );
  NANDN U5295 ( .A(n5111), .B(n5110), .Z(n5115) );
  NAND U5296 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U5297 ( .A(n5115), .B(n5114), .Z(n5130) );
  XNOR U5298 ( .A(n5129), .B(n5130), .Z(n5121) );
  XNOR U5299 ( .A(n5122), .B(n5121), .Z(n5123) );
  XNOR U5300 ( .A(n5124), .B(n5123), .Z(n5157) );
  XNOR U5301 ( .A(sreg[376]), .B(n5157), .Z(n5159) );
  NANDN U5302 ( .A(sreg[375]), .B(n5116), .Z(n5120) );
  NAND U5303 ( .A(n5118), .B(n5117), .Z(n5119) );
  NAND U5304 ( .A(n5120), .B(n5119), .Z(n5158) );
  XNOR U5305 ( .A(n5159), .B(n5158), .Z(c[376]) );
  NANDN U5306 ( .A(n5122), .B(n5121), .Z(n5126) );
  NANDN U5307 ( .A(n5124), .B(n5123), .Z(n5125) );
  AND U5308 ( .A(n5126), .B(n5125), .Z(n5165) );
  NANDN U5309 ( .A(n5128), .B(n5127), .Z(n5132) );
  NANDN U5310 ( .A(n5130), .B(n5129), .Z(n5131) );
  AND U5311 ( .A(n5132), .B(n5131), .Z(n5163) );
  NAND U5312 ( .A(n26), .B(n5133), .Z(n5135) );
  XOR U5313 ( .A(b[7]), .B(a[123]), .Z(n5174) );
  NAND U5314 ( .A(n10531), .B(n5174), .Z(n5134) );
  AND U5315 ( .A(n5135), .B(n5134), .Z(n5193) );
  NAND U5316 ( .A(n23), .B(n5136), .Z(n5138) );
  XOR U5317 ( .A(b[3]), .B(a[127]), .Z(n5177) );
  NAND U5318 ( .A(n24), .B(n5177), .Z(n5137) );
  NAND U5319 ( .A(n5138), .B(n5137), .Z(n5192) );
  XNOR U5320 ( .A(n5193), .B(n5192), .Z(n5195) );
  NAND U5321 ( .A(b[0]), .B(a[129]), .Z(n5139) );
  XNOR U5322 ( .A(b[1]), .B(n5139), .Z(n5141) );
  NANDN U5323 ( .A(b[0]), .B(a[128]), .Z(n5140) );
  NAND U5324 ( .A(n5141), .B(n5140), .Z(n5189) );
  NAND U5325 ( .A(n25), .B(n5142), .Z(n5144) );
  XOR U5326 ( .A(b[5]), .B(a[125]), .Z(n5183) );
  NAND U5327 ( .A(n10456), .B(n5183), .Z(n5143) );
  AND U5328 ( .A(n5144), .B(n5143), .Z(n5187) );
  AND U5329 ( .A(b[7]), .B(a[121]), .Z(n5186) );
  XNOR U5330 ( .A(n5187), .B(n5186), .Z(n5188) );
  XNOR U5331 ( .A(n5189), .B(n5188), .Z(n5194) );
  XOR U5332 ( .A(n5195), .B(n5194), .Z(n5169) );
  NANDN U5333 ( .A(n5146), .B(n5145), .Z(n5150) );
  NANDN U5334 ( .A(n5148), .B(n5147), .Z(n5149) );
  AND U5335 ( .A(n5150), .B(n5149), .Z(n5168) );
  XNOR U5336 ( .A(n5169), .B(n5168), .Z(n5170) );
  NANDN U5337 ( .A(n5152), .B(n5151), .Z(n5156) );
  NAND U5338 ( .A(n5154), .B(n5153), .Z(n5155) );
  NAND U5339 ( .A(n5156), .B(n5155), .Z(n5171) );
  XNOR U5340 ( .A(n5170), .B(n5171), .Z(n5162) );
  XNOR U5341 ( .A(n5163), .B(n5162), .Z(n5164) );
  XNOR U5342 ( .A(n5165), .B(n5164), .Z(n5198) );
  XNOR U5343 ( .A(sreg[377]), .B(n5198), .Z(n5200) );
  NANDN U5344 ( .A(sreg[376]), .B(n5157), .Z(n5161) );
  NAND U5345 ( .A(n5159), .B(n5158), .Z(n5160) );
  NAND U5346 ( .A(n5161), .B(n5160), .Z(n5199) );
  XNOR U5347 ( .A(n5200), .B(n5199), .Z(c[377]) );
  NANDN U5348 ( .A(n5163), .B(n5162), .Z(n5167) );
  NANDN U5349 ( .A(n5165), .B(n5164), .Z(n5166) );
  AND U5350 ( .A(n5167), .B(n5166), .Z(n5206) );
  NANDN U5351 ( .A(n5169), .B(n5168), .Z(n5173) );
  NANDN U5352 ( .A(n5171), .B(n5170), .Z(n5172) );
  AND U5353 ( .A(n5173), .B(n5172), .Z(n5204) );
  NAND U5354 ( .A(n26), .B(n5174), .Z(n5176) );
  XOR U5355 ( .A(b[7]), .B(a[124]), .Z(n5215) );
  NAND U5356 ( .A(n10531), .B(n5215), .Z(n5175) );
  AND U5357 ( .A(n5176), .B(n5175), .Z(n5234) );
  NAND U5358 ( .A(n23), .B(n5177), .Z(n5179) );
  XOR U5359 ( .A(b[3]), .B(a[128]), .Z(n5218) );
  NAND U5360 ( .A(n24), .B(n5218), .Z(n5178) );
  NAND U5361 ( .A(n5179), .B(n5178), .Z(n5233) );
  XNOR U5362 ( .A(n5234), .B(n5233), .Z(n5236) );
  NAND U5363 ( .A(b[0]), .B(a[130]), .Z(n5180) );
  XNOR U5364 ( .A(b[1]), .B(n5180), .Z(n5182) );
  NANDN U5365 ( .A(b[0]), .B(a[129]), .Z(n5181) );
  NAND U5366 ( .A(n5182), .B(n5181), .Z(n5230) );
  NAND U5367 ( .A(n25), .B(n5183), .Z(n5185) );
  XOR U5368 ( .A(b[5]), .B(a[126]), .Z(n5221) );
  NAND U5369 ( .A(n10456), .B(n5221), .Z(n5184) );
  AND U5370 ( .A(n5185), .B(n5184), .Z(n5228) );
  AND U5371 ( .A(b[7]), .B(a[122]), .Z(n5227) );
  XNOR U5372 ( .A(n5228), .B(n5227), .Z(n5229) );
  XNOR U5373 ( .A(n5230), .B(n5229), .Z(n5235) );
  XOR U5374 ( .A(n5236), .B(n5235), .Z(n5210) );
  NANDN U5375 ( .A(n5187), .B(n5186), .Z(n5191) );
  NANDN U5376 ( .A(n5189), .B(n5188), .Z(n5190) );
  AND U5377 ( .A(n5191), .B(n5190), .Z(n5209) );
  XNOR U5378 ( .A(n5210), .B(n5209), .Z(n5211) );
  NANDN U5379 ( .A(n5193), .B(n5192), .Z(n5197) );
  NAND U5380 ( .A(n5195), .B(n5194), .Z(n5196) );
  NAND U5381 ( .A(n5197), .B(n5196), .Z(n5212) );
  XNOR U5382 ( .A(n5211), .B(n5212), .Z(n5203) );
  XNOR U5383 ( .A(n5204), .B(n5203), .Z(n5205) );
  XNOR U5384 ( .A(n5206), .B(n5205), .Z(n5239) );
  XNOR U5385 ( .A(sreg[378]), .B(n5239), .Z(n5241) );
  NANDN U5386 ( .A(sreg[377]), .B(n5198), .Z(n5202) );
  NAND U5387 ( .A(n5200), .B(n5199), .Z(n5201) );
  NAND U5388 ( .A(n5202), .B(n5201), .Z(n5240) );
  XNOR U5389 ( .A(n5241), .B(n5240), .Z(c[378]) );
  NANDN U5390 ( .A(n5204), .B(n5203), .Z(n5208) );
  NANDN U5391 ( .A(n5206), .B(n5205), .Z(n5207) );
  AND U5392 ( .A(n5208), .B(n5207), .Z(n5247) );
  NANDN U5393 ( .A(n5210), .B(n5209), .Z(n5214) );
  NANDN U5394 ( .A(n5212), .B(n5211), .Z(n5213) );
  AND U5395 ( .A(n5214), .B(n5213), .Z(n5245) );
  NAND U5396 ( .A(n26), .B(n5215), .Z(n5217) );
  XOR U5397 ( .A(b[7]), .B(a[125]), .Z(n5256) );
  NAND U5398 ( .A(n10531), .B(n5256), .Z(n5216) );
  AND U5399 ( .A(n5217), .B(n5216), .Z(n5275) );
  NAND U5400 ( .A(n23), .B(n5218), .Z(n5220) );
  XOR U5401 ( .A(b[3]), .B(a[129]), .Z(n5259) );
  NAND U5402 ( .A(n24), .B(n5259), .Z(n5219) );
  NAND U5403 ( .A(n5220), .B(n5219), .Z(n5274) );
  XNOR U5404 ( .A(n5275), .B(n5274), .Z(n5277) );
  NAND U5405 ( .A(n25), .B(n5221), .Z(n5223) );
  XOR U5406 ( .A(b[5]), .B(a[127]), .Z(n5265) );
  NAND U5407 ( .A(n10456), .B(n5265), .Z(n5222) );
  AND U5408 ( .A(n5223), .B(n5222), .Z(n5269) );
  AND U5409 ( .A(b[7]), .B(a[123]), .Z(n5268) );
  XNOR U5410 ( .A(n5269), .B(n5268), .Z(n5270) );
  NAND U5411 ( .A(b[0]), .B(a[131]), .Z(n5224) );
  XNOR U5412 ( .A(b[1]), .B(n5224), .Z(n5226) );
  NANDN U5413 ( .A(b[0]), .B(a[130]), .Z(n5225) );
  NAND U5414 ( .A(n5226), .B(n5225), .Z(n5271) );
  XNOR U5415 ( .A(n5270), .B(n5271), .Z(n5276) );
  XOR U5416 ( .A(n5277), .B(n5276), .Z(n5251) );
  NANDN U5417 ( .A(n5228), .B(n5227), .Z(n5232) );
  NANDN U5418 ( .A(n5230), .B(n5229), .Z(n5231) );
  AND U5419 ( .A(n5232), .B(n5231), .Z(n5250) );
  XNOR U5420 ( .A(n5251), .B(n5250), .Z(n5252) );
  NANDN U5421 ( .A(n5234), .B(n5233), .Z(n5238) );
  NAND U5422 ( .A(n5236), .B(n5235), .Z(n5237) );
  NAND U5423 ( .A(n5238), .B(n5237), .Z(n5253) );
  XNOR U5424 ( .A(n5252), .B(n5253), .Z(n5244) );
  XNOR U5425 ( .A(n5245), .B(n5244), .Z(n5246) );
  XNOR U5426 ( .A(n5247), .B(n5246), .Z(n5280) );
  XNOR U5427 ( .A(sreg[379]), .B(n5280), .Z(n5282) );
  NANDN U5428 ( .A(sreg[378]), .B(n5239), .Z(n5243) );
  NAND U5429 ( .A(n5241), .B(n5240), .Z(n5242) );
  NAND U5430 ( .A(n5243), .B(n5242), .Z(n5281) );
  XNOR U5431 ( .A(n5282), .B(n5281), .Z(c[379]) );
  NANDN U5432 ( .A(n5245), .B(n5244), .Z(n5249) );
  NANDN U5433 ( .A(n5247), .B(n5246), .Z(n5248) );
  AND U5434 ( .A(n5249), .B(n5248), .Z(n5288) );
  NANDN U5435 ( .A(n5251), .B(n5250), .Z(n5255) );
  NANDN U5436 ( .A(n5253), .B(n5252), .Z(n5254) );
  AND U5437 ( .A(n5255), .B(n5254), .Z(n5286) );
  NAND U5438 ( .A(n26), .B(n5256), .Z(n5258) );
  XOR U5439 ( .A(b[7]), .B(a[126]), .Z(n5297) );
  NAND U5440 ( .A(n10531), .B(n5297), .Z(n5257) );
  AND U5441 ( .A(n5258), .B(n5257), .Z(n5316) );
  NAND U5442 ( .A(n23), .B(n5259), .Z(n5261) );
  XOR U5443 ( .A(b[3]), .B(a[130]), .Z(n5300) );
  NAND U5444 ( .A(n24), .B(n5300), .Z(n5260) );
  NAND U5445 ( .A(n5261), .B(n5260), .Z(n5315) );
  XNOR U5446 ( .A(n5316), .B(n5315), .Z(n5318) );
  NAND U5447 ( .A(b[0]), .B(a[132]), .Z(n5262) );
  XNOR U5448 ( .A(b[1]), .B(n5262), .Z(n5264) );
  NANDN U5449 ( .A(b[0]), .B(a[131]), .Z(n5263) );
  NAND U5450 ( .A(n5264), .B(n5263), .Z(n5312) );
  NAND U5451 ( .A(n25), .B(n5265), .Z(n5267) );
  XOR U5452 ( .A(b[5]), .B(a[128]), .Z(n5306) );
  NAND U5453 ( .A(n10456), .B(n5306), .Z(n5266) );
  AND U5454 ( .A(n5267), .B(n5266), .Z(n5310) );
  AND U5455 ( .A(b[7]), .B(a[124]), .Z(n5309) );
  XNOR U5456 ( .A(n5310), .B(n5309), .Z(n5311) );
  XNOR U5457 ( .A(n5312), .B(n5311), .Z(n5317) );
  XOR U5458 ( .A(n5318), .B(n5317), .Z(n5292) );
  NANDN U5459 ( .A(n5269), .B(n5268), .Z(n5273) );
  NANDN U5460 ( .A(n5271), .B(n5270), .Z(n5272) );
  AND U5461 ( .A(n5273), .B(n5272), .Z(n5291) );
  XNOR U5462 ( .A(n5292), .B(n5291), .Z(n5293) );
  NANDN U5463 ( .A(n5275), .B(n5274), .Z(n5279) );
  NAND U5464 ( .A(n5277), .B(n5276), .Z(n5278) );
  NAND U5465 ( .A(n5279), .B(n5278), .Z(n5294) );
  XNOR U5466 ( .A(n5293), .B(n5294), .Z(n5285) );
  XNOR U5467 ( .A(n5286), .B(n5285), .Z(n5287) );
  XNOR U5468 ( .A(n5288), .B(n5287), .Z(n5321) );
  XNOR U5469 ( .A(sreg[380]), .B(n5321), .Z(n5323) );
  NANDN U5470 ( .A(sreg[379]), .B(n5280), .Z(n5284) );
  NAND U5471 ( .A(n5282), .B(n5281), .Z(n5283) );
  NAND U5472 ( .A(n5284), .B(n5283), .Z(n5322) );
  XNOR U5473 ( .A(n5323), .B(n5322), .Z(c[380]) );
  NANDN U5474 ( .A(n5286), .B(n5285), .Z(n5290) );
  NANDN U5475 ( .A(n5288), .B(n5287), .Z(n5289) );
  AND U5476 ( .A(n5290), .B(n5289), .Z(n5329) );
  NANDN U5477 ( .A(n5292), .B(n5291), .Z(n5296) );
  NANDN U5478 ( .A(n5294), .B(n5293), .Z(n5295) );
  AND U5479 ( .A(n5296), .B(n5295), .Z(n5327) );
  NAND U5480 ( .A(n26), .B(n5297), .Z(n5299) );
  XOR U5481 ( .A(b[7]), .B(a[127]), .Z(n5338) );
  NAND U5482 ( .A(n10531), .B(n5338), .Z(n5298) );
  AND U5483 ( .A(n5299), .B(n5298), .Z(n5357) );
  NAND U5484 ( .A(n23), .B(n5300), .Z(n5302) );
  XOR U5485 ( .A(b[3]), .B(a[131]), .Z(n5341) );
  NAND U5486 ( .A(n24), .B(n5341), .Z(n5301) );
  NAND U5487 ( .A(n5302), .B(n5301), .Z(n5356) );
  XNOR U5488 ( .A(n5357), .B(n5356), .Z(n5359) );
  NAND U5489 ( .A(b[0]), .B(a[133]), .Z(n5303) );
  XNOR U5490 ( .A(b[1]), .B(n5303), .Z(n5305) );
  NANDN U5491 ( .A(b[0]), .B(a[132]), .Z(n5304) );
  NAND U5492 ( .A(n5305), .B(n5304), .Z(n5353) );
  NAND U5493 ( .A(n25), .B(n5306), .Z(n5308) );
  XOR U5494 ( .A(b[5]), .B(a[129]), .Z(n5347) );
  NAND U5495 ( .A(n10456), .B(n5347), .Z(n5307) );
  AND U5496 ( .A(n5308), .B(n5307), .Z(n5351) );
  AND U5497 ( .A(b[7]), .B(a[125]), .Z(n5350) );
  XNOR U5498 ( .A(n5351), .B(n5350), .Z(n5352) );
  XNOR U5499 ( .A(n5353), .B(n5352), .Z(n5358) );
  XOR U5500 ( .A(n5359), .B(n5358), .Z(n5333) );
  NANDN U5501 ( .A(n5310), .B(n5309), .Z(n5314) );
  NANDN U5502 ( .A(n5312), .B(n5311), .Z(n5313) );
  AND U5503 ( .A(n5314), .B(n5313), .Z(n5332) );
  XNOR U5504 ( .A(n5333), .B(n5332), .Z(n5334) );
  NANDN U5505 ( .A(n5316), .B(n5315), .Z(n5320) );
  NAND U5506 ( .A(n5318), .B(n5317), .Z(n5319) );
  NAND U5507 ( .A(n5320), .B(n5319), .Z(n5335) );
  XNOR U5508 ( .A(n5334), .B(n5335), .Z(n5326) );
  XNOR U5509 ( .A(n5327), .B(n5326), .Z(n5328) );
  XNOR U5510 ( .A(n5329), .B(n5328), .Z(n5362) );
  XNOR U5511 ( .A(sreg[381]), .B(n5362), .Z(n5364) );
  NANDN U5512 ( .A(sreg[380]), .B(n5321), .Z(n5325) );
  NAND U5513 ( .A(n5323), .B(n5322), .Z(n5324) );
  NAND U5514 ( .A(n5325), .B(n5324), .Z(n5363) );
  XNOR U5515 ( .A(n5364), .B(n5363), .Z(c[381]) );
  NANDN U5516 ( .A(n5327), .B(n5326), .Z(n5331) );
  NANDN U5517 ( .A(n5329), .B(n5328), .Z(n5330) );
  AND U5518 ( .A(n5331), .B(n5330), .Z(n5370) );
  NANDN U5519 ( .A(n5333), .B(n5332), .Z(n5337) );
  NANDN U5520 ( .A(n5335), .B(n5334), .Z(n5336) );
  AND U5521 ( .A(n5337), .B(n5336), .Z(n5368) );
  NAND U5522 ( .A(n26), .B(n5338), .Z(n5340) );
  XOR U5523 ( .A(b[7]), .B(a[128]), .Z(n5379) );
  NAND U5524 ( .A(n10531), .B(n5379), .Z(n5339) );
  AND U5525 ( .A(n5340), .B(n5339), .Z(n5398) );
  NAND U5526 ( .A(n23), .B(n5341), .Z(n5343) );
  XOR U5527 ( .A(b[3]), .B(a[132]), .Z(n5382) );
  NAND U5528 ( .A(n24), .B(n5382), .Z(n5342) );
  NAND U5529 ( .A(n5343), .B(n5342), .Z(n5397) );
  XNOR U5530 ( .A(n5398), .B(n5397), .Z(n5400) );
  NAND U5531 ( .A(b[0]), .B(a[134]), .Z(n5344) );
  XNOR U5532 ( .A(b[1]), .B(n5344), .Z(n5346) );
  NANDN U5533 ( .A(b[0]), .B(a[133]), .Z(n5345) );
  NAND U5534 ( .A(n5346), .B(n5345), .Z(n5394) );
  NAND U5535 ( .A(n25), .B(n5347), .Z(n5349) );
  XOR U5536 ( .A(b[5]), .B(a[130]), .Z(n5385) );
  NAND U5537 ( .A(n10456), .B(n5385), .Z(n5348) );
  AND U5538 ( .A(n5349), .B(n5348), .Z(n5392) );
  AND U5539 ( .A(b[7]), .B(a[126]), .Z(n5391) );
  XNOR U5540 ( .A(n5392), .B(n5391), .Z(n5393) );
  XNOR U5541 ( .A(n5394), .B(n5393), .Z(n5399) );
  XOR U5542 ( .A(n5400), .B(n5399), .Z(n5374) );
  NANDN U5543 ( .A(n5351), .B(n5350), .Z(n5355) );
  NANDN U5544 ( .A(n5353), .B(n5352), .Z(n5354) );
  AND U5545 ( .A(n5355), .B(n5354), .Z(n5373) );
  XNOR U5546 ( .A(n5374), .B(n5373), .Z(n5375) );
  NANDN U5547 ( .A(n5357), .B(n5356), .Z(n5361) );
  NAND U5548 ( .A(n5359), .B(n5358), .Z(n5360) );
  NAND U5549 ( .A(n5361), .B(n5360), .Z(n5376) );
  XNOR U5550 ( .A(n5375), .B(n5376), .Z(n5367) );
  XNOR U5551 ( .A(n5368), .B(n5367), .Z(n5369) );
  XNOR U5552 ( .A(n5370), .B(n5369), .Z(n5403) );
  XNOR U5553 ( .A(sreg[382]), .B(n5403), .Z(n5405) );
  NANDN U5554 ( .A(sreg[381]), .B(n5362), .Z(n5366) );
  NAND U5555 ( .A(n5364), .B(n5363), .Z(n5365) );
  NAND U5556 ( .A(n5366), .B(n5365), .Z(n5404) );
  XNOR U5557 ( .A(n5405), .B(n5404), .Z(c[382]) );
  NANDN U5558 ( .A(n5368), .B(n5367), .Z(n5372) );
  NANDN U5559 ( .A(n5370), .B(n5369), .Z(n5371) );
  AND U5560 ( .A(n5372), .B(n5371), .Z(n5411) );
  NANDN U5561 ( .A(n5374), .B(n5373), .Z(n5378) );
  NANDN U5562 ( .A(n5376), .B(n5375), .Z(n5377) );
  AND U5563 ( .A(n5378), .B(n5377), .Z(n5409) );
  NAND U5564 ( .A(n26), .B(n5379), .Z(n5381) );
  XOR U5565 ( .A(b[7]), .B(a[129]), .Z(n5420) );
  NAND U5566 ( .A(n10531), .B(n5420), .Z(n5380) );
  AND U5567 ( .A(n5381), .B(n5380), .Z(n5439) );
  NAND U5568 ( .A(n23), .B(n5382), .Z(n5384) );
  XOR U5569 ( .A(b[3]), .B(a[133]), .Z(n5423) );
  NAND U5570 ( .A(n24), .B(n5423), .Z(n5383) );
  NAND U5571 ( .A(n5384), .B(n5383), .Z(n5438) );
  XNOR U5572 ( .A(n5439), .B(n5438), .Z(n5441) );
  NAND U5573 ( .A(n25), .B(n5385), .Z(n5387) );
  XOR U5574 ( .A(b[5]), .B(a[131]), .Z(n5429) );
  NAND U5575 ( .A(n10456), .B(n5429), .Z(n5386) );
  AND U5576 ( .A(n5387), .B(n5386), .Z(n5433) );
  AND U5577 ( .A(b[7]), .B(a[127]), .Z(n5432) );
  XNOR U5578 ( .A(n5433), .B(n5432), .Z(n5434) );
  NAND U5579 ( .A(b[0]), .B(a[135]), .Z(n5388) );
  XNOR U5580 ( .A(b[1]), .B(n5388), .Z(n5390) );
  NANDN U5581 ( .A(b[0]), .B(a[134]), .Z(n5389) );
  NAND U5582 ( .A(n5390), .B(n5389), .Z(n5435) );
  XNOR U5583 ( .A(n5434), .B(n5435), .Z(n5440) );
  XOR U5584 ( .A(n5441), .B(n5440), .Z(n5415) );
  NANDN U5585 ( .A(n5392), .B(n5391), .Z(n5396) );
  NANDN U5586 ( .A(n5394), .B(n5393), .Z(n5395) );
  AND U5587 ( .A(n5396), .B(n5395), .Z(n5414) );
  XNOR U5588 ( .A(n5415), .B(n5414), .Z(n5416) );
  NANDN U5589 ( .A(n5398), .B(n5397), .Z(n5402) );
  NAND U5590 ( .A(n5400), .B(n5399), .Z(n5401) );
  NAND U5591 ( .A(n5402), .B(n5401), .Z(n5417) );
  XNOR U5592 ( .A(n5416), .B(n5417), .Z(n5408) );
  XNOR U5593 ( .A(n5409), .B(n5408), .Z(n5410) );
  XNOR U5594 ( .A(n5411), .B(n5410), .Z(n5444) );
  XNOR U5595 ( .A(sreg[383]), .B(n5444), .Z(n5446) );
  NANDN U5596 ( .A(sreg[382]), .B(n5403), .Z(n5407) );
  NAND U5597 ( .A(n5405), .B(n5404), .Z(n5406) );
  NAND U5598 ( .A(n5407), .B(n5406), .Z(n5445) );
  XNOR U5599 ( .A(n5446), .B(n5445), .Z(c[383]) );
  NANDN U5600 ( .A(n5409), .B(n5408), .Z(n5413) );
  NANDN U5601 ( .A(n5411), .B(n5410), .Z(n5412) );
  AND U5602 ( .A(n5413), .B(n5412), .Z(n5452) );
  NANDN U5603 ( .A(n5415), .B(n5414), .Z(n5419) );
  NANDN U5604 ( .A(n5417), .B(n5416), .Z(n5418) );
  AND U5605 ( .A(n5419), .B(n5418), .Z(n5450) );
  NAND U5606 ( .A(n26), .B(n5420), .Z(n5422) );
  XOR U5607 ( .A(b[7]), .B(a[130]), .Z(n5461) );
  NAND U5608 ( .A(n10531), .B(n5461), .Z(n5421) );
  AND U5609 ( .A(n5422), .B(n5421), .Z(n5480) );
  NAND U5610 ( .A(n23), .B(n5423), .Z(n5425) );
  XOR U5611 ( .A(b[3]), .B(a[134]), .Z(n5464) );
  NAND U5612 ( .A(n24), .B(n5464), .Z(n5424) );
  NAND U5613 ( .A(n5425), .B(n5424), .Z(n5479) );
  XNOR U5614 ( .A(n5480), .B(n5479), .Z(n5482) );
  NAND U5615 ( .A(b[0]), .B(a[136]), .Z(n5426) );
  XNOR U5616 ( .A(b[1]), .B(n5426), .Z(n5428) );
  NANDN U5617 ( .A(b[0]), .B(a[135]), .Z(n5427) );
  NAND U5618 ( .A(n5428), .B(n5427), .Z(n5476) );
  NAND U5619 ( .A(n25), .B(n5429), .Z(n5431) );
  XOR U5620 ( .A(b[5]), .B(a[132]), .Z(n5470) );
  NAND U5621 ( .A(n10456), .B(n5470), .Z(n5430) );
  AND U5622 ( .A(n5431), .B(n5430), .Z(n5474) );
  AND U5623 ( .A(b[7]), .B(a[128]), .Z(n5473) );
  XNOR U5624 ( .A(n5474), .B(n5473), .Z(n5475) );
  XNOR U5625 ( .A(n5476), .B(n5475), .Z(n5481) );
  XOR U5626 ( .A(n5482), .B(n5481), .Z(n5456) );
  NANDN U5627 ( .A(n5433), .B(n5432), .Z(n5437) );
  NANDN U5628 ( .A(n5435), .B(n5434), .Z(n5436) );
  AND U5629 ( .A(n5437), .B(n5436), .Z(n5455) );
  XNOR U5630 ( .A(n5456), .B(n5455), .Z(n5457) );
  NANDN U5631 ( .A(n5439), .B(n5438), .Z(n5443) );
  NAND U5632 ( .A(n5441), .B(n5440), .Z(n5442) );
  NAND U5633 ( .A(n5443), .B(n5442), .Z(n5458) );
  XNOR U5634 ( .A(n5457), .B(n5458), .Z(n5449) );
  XNOR U5635 ( .A(n5450), .B(n5449), .Z(n5451) );
  XNOR U5636 ( .A(n5452), .B(n5451), .Z(n5485) );
  XNOR U5637 ( .A(sreg[384]), .B(n5485), .Z(n5487) );
  NANDN U5638 ( .A(sreg[383]), .B(n5444), .Z(n5448) );
  NAND U5639 ( .A(n5446), .B(n5445), .Z(n5447) );
  NAND U5640 ( .A(n5448), .B(n5447), .Z(n5486) );
  XNOR U5641 ( .A(n5487), .B(n5486), .Z(c[384]) );
  NANDN U5642 ( .A(n5450), .B(n5449), .Z(n5454) );
  NANDN U5643 ( .A(n5452), .B(n5451), .Z(n5453) );
  AND U5644 ( .A(n5454), .B(n5453), .Z(n5493) );
  NANDN U5645 ( .A(n5456), .B(n5455), .Z(n5460) );
  NANDN U5646 ( .A(n5458), .B(n5457), .Z(n5459) );
  AND U5647 ( .A(n5460), .B(n5459), .Z(n5491) );
  NAND U5648 ( .A(n26), .B(n5461), .Z(n5463) );
  XOR U5649 ( .A(b[7]), .B(a[131]), .Z(n5502) );
  NAND U5650 ( .A(n10531), .B(n5502), .Z(n5462) );
  AND U5651 ( .A(n5463), .B(n5462), .Z(n5521) );
  NAND U5652 ( .A(n23), .B(n5464), .Z(n5466) );
  XOR U5653 ( .A(b[3]), .B(a[135]), .Z(n5505) );
  NAND U5654 ( .A(n24), .B(n5505), .Z(n5465) );
  NAND U5655 ( .A(n5466), .B(n5465), .Z(n5520) );
  XNOR U5656 ( .A(n5521), .B(n5520), .Z(n5523) );
  NAND U5657 ( .A(b[0]), .B(a[137]), .Z(n5467) );
  XNOR U5658 ( .A(b[1]), .B(n5467), .Z(n5469) );
  NANDN U5659 ( .A(b[0]), .B(a[136]), .Z(n5468) );
  NAND U5660 ( .A(n5469), .B(n5468), .Z(n5517) );
  NAND U5661 ( .A(n25), .B(n5470), .Z(n5472) );
  XOR U5662 ( .A(b[5]), .B(a[133]), .Z(n5508) );
  NAND U5663 ( .A(n10456), .B(n5508), .Z(n5471) );
  AND U5664 ( .A(n5472), .B(n5471), .Z(n5515) );
  AND U5665 ( .A(b[7]), .B(a[129]), .Z(n5514) );
  XNOR U5666 ( .A(n5515), .B(n5514), .Z(n5516) );
  XNOR U5667 ( .A(n5517), .B(n5516), .Z(n5522) );
  XOR U5668 ( .A(n5523), .B(n5522), .Z(n5497) );
  NANDN U5669 ( .A(n5474), .B(n5473), .Z(n5478) );
  NANDN U5670 ( .A(n5476), .B(n5475), .Z(n5477) );
  AND U5671 ( .A(n5478), .B(n5477), .Z(n5496) );
  XNOR U5672 ( .A(n5497), .B(n5496), .Z(n5498) );
  NANDN U5673 ( .A(n5480), .B(n5479), .Z(n5484) );
  NAND U5674 ( .A(n5482), .B(n5481), .Z(n5483) );
  NAND U5675 ( .A(n5484), .B(n5483), .Z(n5499) );
  XNOR U5676 ( .A(n5498), .B(n5499), .Z(n5490) );
  XNOR U5677 ( .A(n5491), .B(n5490), .Z(n5492) );
  XNOR U5678 ( .A(n5493), .B(n5492), .Z(n5526) );
  XNOR U5679 ( .A(sreg[385]), .B(n5526), .Z(n5528) );
  NANDN U5680 ( .A(sreg[384]), .B(n5485), .Z(n5489) );
  NAND U5681 ( .A(n5487), .B(n5486), .Z(n5488) );
  NAND U5682 ( .A(n5489), .B(n5488), .Z(n5527) );
  XNOR U5683 ( .A(n5528), .B(n5527), .Z(c[385]) );
  NANDN U5684 ( .A(n5491), .B(n5490), .Z(n5495) );
  NANDN U5685 ( .A(n5493), .B(n5492), .Z(n5494) );
  AND U5686 ( .A(n5495), .B(n5494), .Z(n5534) );
  NANDN U5687 ( .A(n5497), .B(n5496), .Z(n5501) );
  NANDN U5688 ( .A(n5499), .B(n5498), .Z(n5500) );
  AND U5689 ( .A(n5501), .B(n5500), .Z(n5532) );
  NAND U5690 ( .A(n26), .B(n5502), .Z(n5504) );
  XOR U5691 ( .A(b[7]), .B(a[132]), .Z(n5543) );
  NAND U5692 ( .A(n10531), .B(n5543), .Z(n5503) );
  AND U5693 ( .A(n5504), .B(n5503), .Z(n5562) );
  NAND U5694 ( .A(n23), .B(n5505), .Z(n5507) );
  XOR U5695 ( .A(b[3]), .B(a[136]), .Z(n5546) );
  NAND U5696 ( .A(n24), .B(n5546), .Z(n5506) );
  NAND U5697 ( .A(n5507), .B(n5506), .Z(n5561) );
  XNOR U5698 ( .A(n5562), .B(n5561), .Z(n5564) );
  NAND U5699 ( .A(n25), .B(n5508), .Z(n5510) );
  XOR U5700 ( .A(b[5]), .B(a[134]), .Z(n5552) );
  NAND U5701 ( .A(n10456), .B(n5552), .Z(n5509) );
  AND U5702 ( .A(n5510), .B(n5509), .Z(n5556) );
  AND U5703 ( .A(b[7]), .B(a[130]), .Z(n5555) );
  XNOR U5704 ( .A(n5556), .B(n5555), .Z(n5557) );
  NAND U5705 ( .A(b[0]), .B(a[138]), .Z(n5511) );
  XNOR U5706 ( .A(b[1]), .B(n5511), .Z(n5513) );
  NANDN U5707 ( .A(b[0]), .B(a[137]), .Z(n5512) );
  NAND U5708 ( .A(n5513), .B(n5512), .Z(n5558) );
  XNOR U5709 ( .A(n5557), .B(n5558), .Z(n5563) );
  XOR U5710 ( .A(n5564), .B(n5563), .Z(n5538) );
  NANDN U5711 ( .A(n5515), .B(n5514), .Z(n5519) );
  NANDN U5712 ( .A(n5517), .B(n5516), .Z(n5518) );
  AND U5713 ( .A(n5519), .B(n5518), .Z(n5537) );
  XNOR U5714 ( .A(n5538), .B(n5537), .Z(n5539) );
  NANDN U5715 ( .A(n5521), .B(n5520), .Z(n5525) );
  NAND U5716 ( .A(n5523), .B(n5522), .Z(n5524) );
  NAND U5717 ( .A(n5525), .B(n5524), .Z(n5540) );
  XNOR U5718 ( .A(n5539), .B(n5540), .Z(n5531) );
  XNOR U5719 ( .A(n5532), .B(n5531), .Z(n5533) );
  XNOR U5720 ( .A(n5534), .B(n5533), .Z(n5567) );
  XNOR U5721 ( .A(sreg[386]), .B(n5567), .Z(n5569) );
  NANDN U5722 ( .A(sreg[385]), .B(n5526), .Z(n5530) );
  NAND U5723 ( .A(n5528), .B(n5527), .Z(n5529) );
  NAND U5724 ( .A(n5530), .B(n5529), .Z(n5568) );
  XNOR U5725 ( .A(n5569), .B(n5568), .Z(c[386]) );
  NANDN U5726 ( .A(n5532), .B(n5531), .Z(n5536) );
  NANDN U5727 ( .A(n5534), .B(n5533), .Z(n5535) );
  AND U5728 ( .A(n5536), .B(n5535), .Z(n5575) );
  NANDN U5729 ( .A(n5538), .B(n5537), .Z(n5542) );
  NANDN U5730 ( .A(n5540), .B(n5539), .Z(n5541) );
  AND U5731 ( .A(n5542), .B(n5541), .Z(n5573) );
  NAND U5732 ( .A(n26), .B(n5543), .Z(n5545) );
  XOR U5733 ( .A(b[7]), .B(a[133]), .Z(n5584) );
  NAND U5734 ( .A(n10531), .B(n5584), .Z(n5544) );
  AND U5735 ( .A(n5545), .B(n5544), .Z(n5603) );
  NAND U5736 ( .A(n23), .B(n5546), .Z(n5548) );
  XOR U5737 ( .A(b[3]), .B(a[137]), .Z(n5587) );
  NAND U5738 ( .A(n24), .B(n5587), .Z(n5547) );
  NAND U5739 ( .A(n5548), .B(n5547), .Z(n5602) );
  XNOR U5740 ( .A(n5603), .B(n5602), .Z(n5605) );
  NAND U5741 ( .A(b[0]), .B(a[139]), .Z(n5549) );
  XNOR U5742 ( .A(b[1]), .B(n5549), .Z(n5551) );
  NANDN U5743 ( .A(b[0]), .B(a[138]), .Z(n5550) );
  NAND U5744 ( .A(n5551), .B(n5550), .Z(n5599) );
  NAND U5745 ( .A(n25), .B(n5552), .Z(n5554) );
  XOR U5746 ( .A(b[5]), .B(a[135]), .Z(n5590) );
  NAND U5747 ( .A(n10456), .B(n5590), .Z(n5553) );
  AND U5748 ( .A(n5554), .B(n5553), .Z(n5597) );
  AND U5749 ( .A(b[7]), .B(a[131]), .Z(n5596) );
  XNOR U5750 ( .A(n5597), .B(n5596), .Z(n5598) );
  XNOR U5751 ( .A(n5599), .B(n5598), .Z(n5604) );
  XOR U5752 ( .A(n5605), .B(n5604), .Z(n5579) );
  NANDN U5753 ( .A(n5556), .B(n5555), .Z(n5560) );
  NANDN U5754 ( .A(n5558), .B(n5557), .Z(n5559) );
  AND U5755 ( .A(n5560), .B(n5559), .Z(n5578) );
  XNOR U5756 ( .A(n5579), .B(n5578), .Z(n5580) );
  NANDN U5757 ( .A(n5562), .B(n5561), .Z(n5566) );
  NAND U5758 ( .A(n5564), .B(n5563), .Z(n5565) );
  NAND U5759 ( .A(n5566), .B(n5565), .Z(n5581) );
  XNOR U5760 ( .A(n5580), .B(n5581), .Z(n5572) );
  XNOR U5761 ( .A(n5573), .B(n5572), .Z(n5574) );
  XNOR U5762 ( .A(n5575), .B(n5574), .Z(n5608) );
  XNOR U5763 ( .A(sreg[387]), .B(n5608), .Z(n5610) );
  NANDN U5764 ( .A(sreg[386]), .B(n5567), .Z(n5571) );
  NAND U5765 ( .A(n5569), .B(n5568), .Z(n5570) );
  NAND U5766 ( .A(n5571), .B(n5570), .Z(n5609) );
  XNOR U5767 ( .A(n5610), .B(n5609), .Z(c[387]) );
  NANDN U5768 ( .A(n5573), .B(n5572), .Z(n5577) );
  NANDN U5769 ( .A(n5575), .B(n5574), .Z(n5576) );
  AND U5770 ( .A(n5577), .B(n5576), .Z(n5616) );
  NANDN U5771 ( .A(n5579), .B(n5578), .Z(n5583) );
  NANDN U5772 ( .A(n5581), .B(n5580), .Z(n5582) );
  AND U5773 ( .A(n5583), .B(n5582), .Z(n5614) );
  NAND U5774 ( .A(n26), .B(n5584), .Z(n5586) );
  XOR U5775 ( .A(b[7]), .B(a[134]), .Z(n5625) );
  NAND U5776 ( .A(n10531), .B(n5625), .Z(n5585) );
  AND U5777 ( .A(n5586), .B(n5585), .Z(n5644) );
  NAND U5778 ( .A(n23), .B(n5587), .Z(n5589) );
  XOR U5779 ( .A(b[3]), .B(a[138]), .Z(n5628) );
  NAND U5780 ( .A(n24), .B(n5628), .Z(n5588) );
  NAND U5781 ( .A(n5589), .B(n5588), .Z(n5643) );
  XNOR U5782 ( .A(n5644), .B(n5643), .Z(n5646) );
  NAND U5783 ( .A(n25), .B(n5590), .Z(n5592) );
  XOR U5784 ( .A(b[5]), .B(a[136]), .Z(n5634) );
  NAND U5785 ( .A(n10456), .B(n5634), .Z(n5591) );
  AND U5786 ( .A(n5592), .B(n5591), .Z(n5638) );
  AND U5787 ( .A(b[7]), .B(a[132]), .Z(n5637) );
  XNOR U5788 ( .A(n5638), .B(n5637), .Z(n5639) );
  NAND U5789 ( .A(b[0]), .B(a[140]), .Z(n5593) );
  XNOR U5790 ( .A(b[1]), .B(n5593), .Z(n5595) );
  NANDN U5791 ( .A(b[0]), .B(a[139]), .Z(n5594) );
  NAND U5792 ( .A(n5595), .B(n5594), .Z(n5640) );
  XNOR U5793 ( .A(n5639), .B(n5640), .Z(n5645) );
  XOR U5794 ( .A(n5646), .B(n5645), .Z(n5620) );
  NANDN U5795 ( .A(n5597), .B(n5596), .Z(n5601) );
  NANDN U5796 ( .A(n5599), .B(n5598), .Z(n5600) );
  AND U5797 ( .A(n5601), .B(n5600), .Z(n5619) );
  XNOR U5798 ( .A(n5620), .B(n5619), .Z(n5621) );
  NANDN U5799 ( .A(n5603), .B(n5602), .Z(n5607) );
  NAND U5800 ( .A(n5605), .B(n5604), .Z(n5606) );
  NAND U5801 ( .A(n5607), .B(n5606), .Z(n5622) );
  XNOR U5802 ( .A(n5621), .B(n5622), .Z(n5613) );
  XNOR U5803 ( .A(n5614), .B(n5613), .Z(n5615) );
  XNOR U5804 ( .A(n5616), .B(n5615), .Z(n5649) );
  XNOR U5805 ( .A(sreg[388]), .B(n5649), .Z(n5651) );
  NANDN U5806 ( .A(sreg[387]), .B(n5608), .Z(n5612) );
  NAND U5807 ( .A(n5610), .B(n5609), .Z(n5611) );
  NAND U5808 ( .A(n5612), .B(n5611), .Z(n5650) );
  XNOR U5809 ( .A(n5651), .B(n5650), .Z(c[388]) );
  NANDN U5810 ( .A(n5614), .B(n5613), .Z(n5618) );
  NANDN U5811 ( .A(n5616), .B(n5615), .Z(n5617) );
  AND U5812 ( .A(n5618), .B(n5617), .Z(n5657) );
  NANDN U5813 ( .A(n5620), .B(n5619), .Z(n5624) );
  NANDN U5814 ( .A(n5622), .B(n5621), .Z(n5623) );
  AND U5815 ( .A(n5624), .B(n5623), .Z(n5655) );
  NAND U5816 ( .A(n26), .B(n5625), .Z(n5627) );
  XOR U5817 ( .A(b[7]), .B(a[135]), .Z(n5666) );
  NAND U5818 ( .A(n10531), .B(n5666), .Z(n5626) );
  AND U5819 ( .A(n5627), .B(n5626), .Z(n5685) );
  NAND U5820 ( .A(n23), .B(n5628), .Z(n5630) );
  XOR U5821 ( .A(b[3]), .B(a[139]), .Z(n5669) );
  NAND U5822 ( .A(n24), .B(n5669), .Z(n5629) );
  NAND U5823 ( .A(n5630), .B(n5629), .Z(n5684) );
  XNOR U5824 ( .A(n5685), .B(n5684), .Z(n5687) );
  NAND U5825 ( .A(b[0]), .B(a[141]), .Z(n5631) );
  XNOR U5826 ( .A(b[1]), .B(n5631), .Z(n5633) );
  NANDN U5827 ( .A(b[0]), .B(a[140]), .Z(n5632) );
  NAND U5828 ( .A(n5633), .B(n5632), .Z(n5681) );
  NAND U5829 ( .A(n25), .B(n5634), .Z(n5636) );
  XOR U5830 ( .A(b[5]), .B(a[137]), .Z(n5672) );
  NAND U5831 ( .A(n10456), .B(n5672), .Z(n5635) );
  AND U5832 ( .A(n5636), .B(n5635), .Z(n5679) );
  AND U5833 ( .A(b[7]), .B(a[133]), .Z(n5678) );
  XNOR U5834 ( .A(n5679), .B(n5678), .Z(n5680) );
  XNOR U5835 ( .A(n5681), .B(n5680), .Z(n5686) );
  XOR U5836 ( .A(n5687), .B(n5686), .Z(n5661) );
  NANDN U5837 ( .A(n5638), .B(n5637), .Z(n5642) );
  NANDN U5838 ( .A(n5640), .B(n5639), .Z(n5641) );
  AND U5839 ( .A(n5642), .B(n5641), .Z(n5660) );
  XNOR U5840 ( .A(n5661), .B(n5660), .Z(n5662) );
  NANDN U5841 ( .A(n5644), .B(n5643), .Z(n5648) );
  NAND U5842 ( .A(n5646), .B(n5645), .Z(n5647) );
  NAND U5843 ( .A(n5648), .B(n5647), .Z(n5663) );
  XNOR U5844 ( .A(n5662), .B(n5663), .Z(n5654) );
  XNOR U5845 ( .A(n5655), .B(n5654), .Z(n5656) );
  XNOR U5846 ( .A(n5657), .B(n5656), .Z(n5690) );
  XNOR U5847 ( .A(sreg[389]), .B(n5690), .Z(n5692) );
  NANDN U5848 ( .A(sreg[388]), .B(n5649), .Z(n5653) );
  NAND U5849 ( .A(n5651), .B(n5650), .Z(n5652) );
  NAND U5850 ( .A(n5653), .B(n5652), .Z(n5691) );
  XNOR U5851 ( .A(n5692), .B(n5691), .Z(c[389]) );
  NANDN U5852 ( .A(n5655), .B(n5654), .Z(n5659) );
  NANDN U5853 ( .A(n5657), .B(n5656), .Z(n5658) );
  AND U5854 ( .A(n5659), .B(n5658), .Z(n5698) );
  NANDN U5855 ( .A(n5661), .B(n5660), .Z(n5665) );
  NANDN U5856 ( .A(n5663), .B(n5662), .Z(n5664) );
  AND U5857 ( .A(n5665), .B(n5664), .Z(n5696) );
  NAND U5858 ( .A(n26), .B(n5666), .Z(n5668) );
  XOR U5859 ( .A(b[7]), .B(a[136]), .Z(n5707) );
  NAND U5860 ( .A(n10531), .B(n5707), .Z(n5667) );
  AND U5861 ( .A(n5668), .B(n5667), .Z(n5726) );
  NAND U5862 ( .A(n23), .B(n5669), .Z(n5671) );
  XOR U5863 ( .A(b[3]), .B(a[140]), .Z(n5710) );
  NAND U5864 ( .A(n24), .B(n5710), .Z(n5670) );
  NAND U5865 ( .A(n5671), .B(n5670), .Z(n5725) );
  XNOR U5866 ( .A(n5726), .B(n5725), .Z(n5728) );
  NAND U5867 ( .A(n25), .B(n5672), .Z(n5674) );
  XOR U5868 ( .A(b[5]), .B(a[138]), .Z(n5716) );
  NAND U5869 ( .A(n10456), .B(n5716), .Z(n5673) );
  AND U5870 ( .A(n5674), .B(n5673), .Z(n5720) );
  AND U5871 ( .A(b[7]), .B(a[134]), .Z(n5719) );
  XNOR U5872 ( .A(n5720), .B(n5719), .Z(n5721) );
  NAND U5873 ( .A(b[0]), .B(a[142]), .Z(n5675) );
  XNOR U5874 ( .A(b[1]), .B(n5675), .Z(n5677) );
  NANDN U5875 ( .A(b[0]), .B(a[141]), .Z(n5676) );
  NAND U5876 ( .A(n5677), .B(n5676), .Z(n5722) );
  XNOR U5877 ( .A(n5721), .B(n5722), .Z(n5727) );
  XOR U5878 ( .A(n5728), .B(n5727), .Z(n5702) );
  NANDN U5879 ( .A(n5679), .B(n5678), .Z(n5683) );
  NANDN U5880 ( .A(n5681), .B(n5680), .Z(n5682) );
  AND U5881 ( .A(n5683), .B(n5682), .Z(n5701) );
  XNOR U5882 ( .A(n5702), .B(n5701), .Z(n5703) );
  NANDN U5883 ( .A(n5685), .B(n5684), .Z(n5689) );
  NAND U5884 ( .A(n5687), .B(n5686), .Z(n5688) );
  NAND U5885 ( .A(n5689), .B(n5688), .Z(n5704) );
  XNOR U5886 ( .A(n5703), .B(n5704), .Z(n5695) );
  XNOR U5887 ( .A(n5696), .B(n5695), .Z(n5697) );
  XNOR U5888 ( .A(n5698), .B(n5697), .Z(n5731) );
  XNOR U5889 ( .A(sreg[390]), .B(n5731), .Z(n5733) );
  NANDN U5890 ( .A(sreg[389]), .B(n5690), .Z(n5694) );
  NAND U5891 ( .A(n5692), .B(n5691), .Z(n5693) );
  NAND U5892 ( .A(n5694), .B(n5693), .Z(n5732) );
  XNOR U5893 ( .A(n5733), .B(n5732), .Z(c[390]) );
  NANDN U5894 ( .A(n5696), .B(n5695), .Z(n5700) );
  NANDN U5895 ( .A(n5698), .B(n5697), .Z(n5699) );
  AND U5896 ( .A(n5700), .B(n5699), .Z(n5739) );
  NANDN U5897 ( .A(n5702), .B(n5701), .Z(n5706) );
  NANDN U5898 ( .A(n5704), .B(n5703), .Z(n5705) );
  AND U5899 ( .A(n5706), .B(n5705), .Z(n5737) );
  NAND U5900 ( .A(n26), .B(n5707), .Z(n5709) );
  XOR U5901 ( .A(b[7]), .B(a[137]), .Z(n5748) );
  NAND U5902 ( .A(n10531), .B(n5748), .Z(n5708) );
  AND U5903 ( .A(n5709), .B(n5708), .Z(n5767) );
  NAND U5904 ( .A(n23), .B(n5710), .Z(n5712) );
  XOR U5905 ( .A(b[3]), .B(a[141]), .Z(n5751) );
  NAND U5906 ( .A(n24), .B(n5751), .Z(n5711) );
  NAND U5907 ( .A(n5712), .B(n5711), .Z(n5766) );
  XNOR U5908 ( .A(n5767), .B(n5766), .Z(n5769) );
  NAND U5909 ( .A(b[0]), .B(a[143]), .Z(n5713) );
  XNOR U5910 ( .A(b[1]), .B(n5713), .Z(n5715) );
  NANDN U5911 ( .A(b[0]), .B(a[142]), .Z(n5714) );
  NAND U5912 ( .A(n5715), .B(n5714), .Z(n5763) );
  NAND U5913 ( .A(n25), .B(n5716), .Z(n5718) );
  XOR U5914 ( .A(b[5]), .B(a[139]), .Z(n5757) );
  NAND U5915 ( .A(n10456), .B(n5757), .Z(n5717) );
  AND U5916 ( .A(n5718), .B(n5717), .Z(n5761) );
  AND U5917 ( .A(b[7]), .B(a[135]), .Z(n5760) );
  XNOR U5918 ( .A(n5761), .B(n5760), .Z(n5762) );
  XNOR U5919 ( .A(n5763), .B(n5762), .Z(n5768) );
  XOR U5920 ( .A(n5769), .B(n5768), .Z(n5743) );
  NANDN U5921 ( .A(n5720), .B(n5719), .Z(n5724) );
  NANDN U5922 ( .A(n5722), .B(n5721), .Z(n5723) );
  AND U5923 ( .A(n5724), .B(n5723), .Z(n5742) );
  XNOR U5924 ( .A(n5743), .B(n5742), .Z(n5744) );
  NANDN U5925 ( .A(n5726), .B(n5725), .Z(n5730) );
  NAND U5926 ( .A(n5728), .B(n5727), .Z(n5729) );
  NAND U5927 ( .A(n5730), .B(n5729), .Z(n5745) );
  XNOR U5928 ( .A(n5744), .B(n5745), .Z(n5736) );
  XNOR U5929 ( .A(n5737), .B(n5736), .Z(n5738) );
  XNOR U5930 ( .A(n5739), .B(n5738), .Z(n5772) );
  XNOR U5931 ( .A(sreg[391]), .B(n5772), .Z(n5774) );
  NANDN U5932 ( .A(sreg[390]), .B(n5731), .Z(n5735) );
  NAND U5933 ( .A(n5733), .B(n5732), .Z(n5734) );
  NAND U5934 ( .A(n5735), .B(n5734), .Z(n5773) );
  XNOR U5935 ( .A(n5774), .B(n5773), .Z(c[391]) );
  NANDN U5936 ( .A(n5737), .B(n5736), .Z(n5741) );
  NANDN U5937 ( .A(n5739), .B(n5738), .Z(n5740) );
  AND U5938 ( .A(n5741), .B(n5740), .Z(n5780) );
  NANDN U5939 ( .A(n5743), .B(n5742), .Z(n5747) );
  NANDN U5940 ( .A(n5745), .B(n5744), .Z(n5746) );
  AND U5941 ( .A(n5747), .B(n5746), .Z(n5778) );
  NAND U5942 ( .A(n26), .B(n5748), .Z(n5750) );
  XOR U5943 ( .A(b[7]), .B(a[138]), .Z(n5789) );
  NAND U5944 ( .A(n10531), .B(n5789), .Z(n5749) );
  AND U5945 ( .A(n5750), .B(n5749), .Z(n5808) );
  NAND U5946 ( .A(n23), .B(n5751), .Z(n5753) );
  XOR U5947 ( .A(b[3]), .B(a[142]), .Z(n5792) );
  NAND U5948 ( .A(n24), .B(n5792), .Z(n5752) );
  NAND U5949 ( .A(n5753), .B(n5752), .Z(n5807) );
  XNOR U5950 ( .A(n5808), .B(n5807), .Z(n5810) );
  NAND U5951 ( .A(b[0]), .B(a[144]), .Z(n5754) );
  XNOR U5952 ( .A(b[1]), .B(n5754), .Z(n5756) );
  NANDN U5953 ( .A(b[0]), .B(a[143]), .Z(n5755) );
  NAND U5954 ( .A(n5756), .B(n5755), .Z(n5804) );
  NAND U5955 ( .A(n25), .B(n5757), .Z(n5759) );
  XOR U5956 ( .A(b[5]), .B(a[140]), .Z(n5795) );
  NAND U5957 ( .A(n10456), .B(n5795), .Z(n5758) );
  AND U5958 ( .A(n5759), .B(n5758), .Z(n5802) );
  AND U5959 ( .A(b[7]), .B(a[136]), .Z(n5801) );
  XNOR U5960 ( .A(n5802), .B(n5801), .Z(n5803) );
  XNOR U5961 ( .A(n5804), .B(n5803), .Z(n5809) );
  XOR U5962 ( .A(n5810), .B(n5809), .Z(n5784) );
  NANDN U5963 ( .A(n5761), .B(n5760), .Z(n5765) );
  NANDN U5964 ( .A(n5763), .B(n5762), .Z(n5764) );
  AND U5965 ( .A(n5765), .B(n5764), .Z(n5783) );
  XNOR U5966 ( .A(n5784), .B(n5783), .Z(n5785) );
  NANDN U5967 ( .A(n5767), .B(n5766), .Z(n5771) );
  NAND U5968 ( .A(n5769), .B(n5768), .Z(n5770) );
  NAND U5969 ( .A(n5771), .B(n5770), .Z(n5786) );
  XNOR U5970 ( .A(n5785), .B(n5786), .Z(n5777) );
  XNOR U5971 ( .A(n5778), .B(n5777), .Z(n5779) );
  XNOR U5972 ( .A(n5780), .B(n5779), .Z(n5813) );
  XNOR U5973 ( .A(sreg[392]), .B(n5813), .Z(n5815) );
  NANDN U5974 ( .A(sreg[391]), .B(n5772), .Z(n5776) );
  NAND U5975 ( .A(n5774), .B(n5773), .Z(n5775) );
  NAND U5976 ( .A(n5776), .B(n5775), .Z(n5814) );
  XNOR U5977 ( .A(n5815), .B(n5814), .Z(c[392]) );
  NANDN U5978 ( .A(n5778), .B(n5777), .Z(n5782) );
  NANDN U5979 ( .A(n5780), .B(n5779), .Z(n5781) );
  AND U5980 ( .A(n5782), .B(n5781), .Z(n5821) );
  NANDN U5981 ( .A(n5784), .B(n5783), .Z(n5788) );
  NANDN U5982 ( .A(n5786), .B(n5785), .Z(n5787) );
  AND U5983 ( .A(n5788), .B(n5787), .Z(n5819) );
  NAND U5984 ( .A(n26), .B(n5789), .Z(n5791) );
  XOR U5985 ( .A(b[7]), .B(a[139]), .Z(n5830) );
  NAND U5986 ( .A(n10531), .B(n5830), .Z(n5790) );
  AND U5987 ( .A(n5791), .B(n5790), .Z(n5849) );
  NAND U5988 ( .A(n23), .B(n5792), .Z(n5794) );
  XOR U5989 ( .A(b[3]), .B(a[143]), .Z(n5833) );
  NAND U5990 ( .A(n24), .B(n5833), .Z(n5793) );
  NAND U5991 ( .A(n5794), .B(n5793), .Z(n5848) );
  XNOR U5992 ( .A(n5849), .B(n5848), .Z(n5851) );
  NAND U5993 ( .A(n25), .B(n5795), .Z(n5797) );
  XOR U5994 ( .A(b[5]), .B(a[141]), .Z(n5836) );
  NAND U5995 ( .A(n10456), .B(n5836), .Z(n5796) );
  AND U5996 ( .A(n5797), .B(n5796), .Z(n5843) );
  AND U5997 ( .A(b[7]), .B(a[137]), .Z(n5842) );
  XNOR U5998 ( .A(n5843), .B(n5842), .Z(n5844) );
  NAND U5999 ( .A(b[0]), .B(a[145]), .Z(n5798) );
  XNOR U6000 ( .A(b[1]), .B(n5798), .Z(n5800) );
  NANDN U6001 ( .A(b[0]), .B(a[144]), .Z(n5799) );
  NAND U6002 ( .A(n5800), .B(n5799), .Z(n5845) );
  XNOR U6003 ( .A(n5844), .B(n5845), .Z(n5850) );
  XOR U6004 ( .A(n5851), .B(n5850), .Z(n5825) );
  NANDN U6005 ( .A(n5802), .B(n5801), .Z(n5806) );
  NANDN U6006 ( .A(n5804), .B(n5803), .Z(n5805) );
  AND U6007 ( .A(n5806), .B(n5805), .Z(n5824) );
  XNOR U6008 ( .A(n5825), .B(n5824), .Z(n5826) );
  NANDN U6009 ( .A(n5808), .B(n5807), .Z(n5812) );
  NAND U6010 ( .A(n5810), .B(n5809), .Z(n5811) );
  NAND U6011 ( .A(n5812), .B(n5811), .Z(n5827) );
  XNOR U6012 ( .A(n5826), .B(n5827), .Z(n5818) );
  XNOR U6013 ( .A(n5819), .B(n5818), .Z(n5820) );
  XNOR U6014 ( .A(n5821), .B(n5820), .Z(n5854) );
  XNOR U6015 ( .A(sreg[393]), .B(n5854), .Z(n5856) );
  NANDN U6016 ( .A(sreg[392]), .B(n5813), .Z(n5817) );
  NAND U6017 ( .A(n5815), .B(n5814), .Z(n5816) );
  NAND U6018 ( .A(n5817), .B(n5816), .Z(n5855) );
  XNOR U6019 ( .A(n5856), .B(n5855), .Z(c[393]) );
  NANDN U6020 ( .A(n5819), .B(n5818), .Z(n5823) );
  NANDN U6021 ( .A(n5821), .B(n5820), .Z(n5822) );
  AND U6022 ( .A(n5823), .B(n5822), .Z(n5862) );
  NANDN U6023 ( .A(n5825), .B(n5824), .Z(n5829) );
  NANDN U6024 ( .A(n5827), .B(n5826), .Z(n5828) );
  AND U6025 ( .A(n5829), .B(n5828), .Z(n5860) );
  NAND U6026 ( .A(n26), .B(n5830), .Z(n5832) );
  XOR U6027 ( .A(b[7]), .B(a[140]), .Z(n5871) );
  NAND U6028 ( .A(n10531), .B(n5871), .Z(n5831) );
  AND U6029 ( .A(n5832), .B(n5831), .Z(n5890) );
  NAND U6030 ( .A(n23), .B(n5833), .Z(n5835) );
  XOR U6031 ( .A(b[3]), .B(a[144]), .Z(n5874) );
  NAND U6032 ( .A(n24), .B(n5874), .Z(n5834) );
  NAND U6033 ( .A(n5835), .B(n5834), .Z(n5889) );
  XNOR U6034 ( .A(n5890), .B(n5889), .Z(n5892) );
  NAND U6035 ( .A(n25), .B(n5836), .Z(n5838) );
  XOR U6036 ( .A(b[5]), .B(a[142]), .Z(n5877) );
  NAND U6037 ( .A(n10456), .B(n5877), .Z(n5837) );
  AND U6038 ( .A(n5838), .B(n5837), .Z(n5884) );
  AND U6039 ( .A(b[7]), .B(a[138]), .Z(n5883) );
  XNOR U6040 ( .A(n5884), .B(n5883), .Z(n5885) );
  NAND U6041 ( .A(b[0]), .B(a[146]), .Z(n5839) );
  XNOR U6042 ( .A(b[1]), .B(n5839), .Z(n5841) );
  NANDN U6043 ( .A(b[0]), .B(a[145]), .Z(n5840) );
  NAND U6044 ( .A(n5841), .B(n5840), .Z(n5886) );
  XNOR U6045 ( .A(n5885), .B(n5886), .Z(n5891) );
  XOR U6046 ( .A(n5892), .B(n5891), .Z(n5866) );
  NANDN U6047 ( .A(n5843), .B(n5842), .Z(n5847) );
  NANDN U6048 ( .A(n5845), .B(n5844), .Z(n5846) );
  AND U6049 ( .A(n5847), .B(n5846), .Z(n5865) );
  XNOR U6050 ( .A(n5866), .B(n5865), .Z(n5867) );
  NANDN U6051 ( .A(n5849), .B(n5848), .Z(n5853) );
  NAND U6052 ( .A(n5851), .B(n5850), .Z(n5852) );
  NAND U6053 ( .A(n5853), .B(n5852), .Z(n5868) );
  XNOR U6054 ( .A(n5867), .B(n5868), .Z(n5859) );
  XNOR U6055 ( .A(n5860), .B(n5859), .Z(n5861) );
  XNOR U6056 ( .A(n5862), .B(n5861), .Z(n5895) );
  XNOR U6057 ( .A(sreg[394]), .B(n5895), .Z(n5897) );
  NANDN U6058 ( .A(sreg[393]), .B(n5854), .Z(n5858) );
  NAND U6059 ( .A(n5856), .B(n5855), .Z(n5857) );
  NAND U6060 ( .A(n5858), .B(n5857), .Z(n5896) );
  XNOR U6061 ( .A(n5897), .B(n5896), .Z(c[394]) );
  NANDN U6062 ( .A(n5860), .B(n5859), .Z(n5864) );
  NANDN U6063 ( .A(n5862), .B(n5861), .Z(n5863) );
  AND U6064 ( .A(n5864), .B(n5863), .Z(n5903) );
  NANDN U6065 ( .A(n5866), .B(n5865), .Z(n5870) );
  NANDN U6066 ( .A(n5868), .B(n5867), .Z(n5869) );
  AND U6067 ( .A(n5870), .B(n5869), .Z(n5901) );
  NAND U6068 ( .A(n26), .B(n5871), .Z(n5873) );
  XOR U6069 ( .A(b[7]), .B(a[141]), .Z(n5912) );
  NAND U6070 ( .A(n10531), .B(n5912), .Z(n5872) );
  AND U6071 ( .A(n5873), .B(n5872), .Z(n5931) );
  NAND U6072 ( .A(n23), .B(n5874), .Z(n5876) );
  XOR U6073 ( .A(b[3]), .B(a[145]), .Z(n5915) );
  NAND U6074 ( .A(n24), .B(n5915), .Z(n5875) );
  NAND U6075 ( .A(n5876), .B(n5875), .Z(n5930) );
  XNOR U6076 ( .A(n5931), .B(n5930), .Z(n5933) );
  NAND U6077 ( .A(n25), .B(n5877), .Z(n5879) );
  XOR U6078 ( .A(b[5]), .B(a[143]), .Z(n5921) );
  NAND U6079 ( .A(n10456), .B(n5921), .Z(n5878) );
  AND U6080 ( .A(n5879), .B(n5878), .Z(n5925) );
  AND U6081 ( .A(b[7]), .B(a[139]), .Z(n5924) );
  XNOR U6082 ( .A(n5925), .B(n5924), .Z(n5926) );
  NAND U6083 ( .A(b[0]), .B(a[147]), .Z(n5880) );
  XNOR U6084 ( .A(b[1]), .B(n5880), .Z(n5882) );
  NANDN U6085 ( .A(b[0]), .B(a[146]), .Z(n5881) );
  NAND U6086 ( .A(n5882), .B(n5881), .Z(n5927) );
  XNOR U6087 ( .A(n5926), .B(n5927), .Z(n5932) );
  XOR U6088 ( .A(n5933), .B(n5932), .Z(n5907) );
  NANDN U6089 ( .A(n5884), .B(n5883), .Z(n5888) );
  NANDN U6090 ( .A(n5886), .B(n5885), .Z(n5887) );
  AND U6091 ( .A(n5888), .B(n5887), .Z(n5906) );
  XNOR U6092 ( .A(n5907), .B(n5906), .Z(n5908) );
  NANDN U6093 ( .A(n5890), .B(n5889), .Z(n5894) );
  NAND U6094 ( .A(n5892), .B(n5891), .Z(n5893) );
  NAND U6095 ( .A(n5894), .B(n5893), .Z(n5909) );
  XNOR U6096 ( .A(n5908), .B(n5909), .Z(n5900) );
  XNOR U6097 ( .A(n5901), .B(n5900), .Z(n5902) );
  XNOR U6098 ( .A(n5903), .B(n5902), .Z(n5936) );
  XNOR U6099 ( .A(sreg[395]), .B(n5936), .Z(n5938) );
  NANDN U6100 ( .A(sreg[394]), .B(n5895), .Z(n5899) );
  NAND U6101 ( .A(n5897), .B(n5896), .Z(n5898) );
  NAND U6102 ( .A(n5899), .B(n5898), .Z(n5937) );
  XNOR U6103 ( .A(n5938), .B(n5937), .Z(c[395]) );
  NANDN U6104 ( .A(n5901), .B(n5900), .Z(n5905) );
  NANDN U6105 ( .A(n5903), .B(n5902), .Z(n5904) );
  AND U6106 ( .A(n5905), .B(n5904), .Z(n5944) );
  NANDN U6107 ( .A(n5907), .B(n5906), .Z(n5911) );
  NANDN U6108 ( .A(n5909), .B(n5908), .Z(n5910) );
  AND U6109 ( .A(n5911), .B(n5910), .Z(n5942) );
  NAND U6110 ( .A(n26), .B(n5912), .Z(n5914) );
  XOR U6111 ( .A(b[7]), .B(a[142]), .Z(n5953) );
  NAND U6112 ( .A(n10531), .B(n5953), .Z(n5913) );
  AND U6113 ( .A(n5914), .B(n5913), .Z(n5972) );
  NAND U6114 ( .A(n23), .B(n5915), .Z(n5917) );
  XOR U6115 ( .A(b[3]), .B(a[146]), .Z(n5956) );
  NAND U6116 ( .A(n24), .B(n5956), .Z(n5916) );
  NAND U6117 ( .A(n5917), .B(n5916), .Z(n5971) );
  XNOR U6118 ( .A(n5972), .B(n5971), .Z(n5974) );
  NAND U6119 ( .A(b[0]), .B(a[148]), .Z(n5918) );
  XNOR U6120 ( .A(b[1]), .B(n5918), .Z(n5920) );
  NANDN U6121 ( .A(b[0]), .B(a[147]), .Z(n5919) );
  NAND U6122 ( .A(n5920), .B(n5919), .Z(n5968) );
  NAND U6123 ( .A(n25), .B(n5921), .Z(n5923) );
  XOR U6124 ( .A(b[5]), .B(a[144]), .Z(n5962) );
  NAND U6125 ( .A(n10456), .B(n5962), .Z(n5922) );
  AND U6126 ( .A(n5923), .B(n5922), .Z(n5966) );
  AND U6127 ( .A(b[7]), .B(a[140]), .Z(n5965) );
  XNOR U6128 ( .A(n5966), .B(n5965), .Z(n5967) );
  XNOR U6129 ( .A(n5968), .B(n5967), .Z(n5973) );
  XOR U6130 ( .A(n5974), .B(n5973), .Z(n5948) );
  NANDN U6131 ( .A(n5925), .B(n5924), .Z(n5929) );
  NANDN U6132 ( .A(n5927), .B(n5926), .Z(n5928) );
  AND U6133 ( .A(n5929), .B(n5928), .Z(n5947) );
  XNOR U6134 ( .A(n5948), .B(n5947), .Z(n5949) );
  NANDN U6135 ( .A(n5931), .B(n5930), .Z(n5935) );
  NAND U6136 ( .A(n5933), .B(n5932), .Z(n5934) );
  NAND U6137 ( .A(n5935), .B(n5934), .Z(n5950) );
  XNOR U6138 ( .A(n5949), .B(n5950), .Z(n5941) );
  XNOR U6139 ( .A(n5942), .B(n5941), .Z(n5943) );
  XNOR U6140 ( .A(n5944), .B(n5943), .Z(n5977) );
  XNOR U6141 ( .A(sreg[396]), .B(n5977), .Z(n5979) );
  NANDN U6142 ( .A(sreg[395]), .B(n5936), .Z(n5940) );
  NAND U6143 ( .A(n5938), .B(n5937), .Z(n5939) );
  NAND U6144 ( .A(n5940), .B(n5939), .Z(n5978) );
  XNOR U6145 ( .A(n5979), .B(n5978), .Z(c[396]) );
  NANDN U6146 ( .A(n5942), .B(n5941), .Z(n5946) );
  NANDN U6147 ( .A(n5944), .B(n5943), .Z(n5945) );
  AND U6148 ( .A(n5946), .B(n5945), .Z(n5985) );
  NANDN U6149 ( .A(n5948), .B(n5947), .Z(n5952) );
  NANDN U6150 ( .A(n5950), .B(n5949), .Z(n5951) );
  AND U6151 ( .A(n5952), .B(n5951), .Z(n5983) );
  NAND U6152 ( .A(n26), .B(n5953), .Z(n5955) );
  XOR U6153 ( .A(b[7]), .B(a[143]), .Z(n5994) );
  NAND U6154 ( .A(n10531), .B(n5994), .Z(n5954) );
  AND U6155 ( .A(n5955), .B(n5954), .Z(n6013) );
  NAND U6156 ( .A(n23), .B(n5956), .Z(n5958) );
  XOR U6157 ( .A(b[3]), .B(a[147]), .Z(n5997) );
  NAND U6158 ( .A(n24), .B(n5997), .Z(n5957) );
  NAND U6159 ( .A(n5958), .B(n5957), .Z(n6012) );
  XNOR U6160 ( .A(n6013), .B(n6012), .Z(n6015) );
  NAND U6161 ( .A(b[0]), .B(a[149]), .Z(n5959) );
  XNOR U6162 ( .A(b[1]), .B(n5959), .Z(n5961) );
  NANDN U6163 ( .A(b[0]), .B(a[148]), .Z(n5960) );
  NAND U6164 ( .A(n5961), .B(n5960), .Z(n6009) );
  NAND U6165 ( .A(n25), .B(n5962), .Z(n5964) );
  XOR U6166 ( .A(b[5]), .B(a[145]), .Z(n6000) );
  NAND U6167 ( .A(n10456), .B(n6000), .Z(n5963) );
  AND U6168 ( .A(n5964), .B(n5963), .Z(n6007) );
  AND U6169 ( .A(b[7]), .B(a[141]), .Z(n6006) );
  XNOR U6170 ( .A(n6007), .B(n6006), .Z(n6008) );
  XNOR U6171 ( .A(n6009), .B(n6008), .Z(n6014) );
  XOR U6172 ( .A(n6015), .B(n6014), .Z(n5989) );
  NANDN U6173 ( .A(n5966), .B(n5965), .Z(n5970) );
  NANDN U6174 ( .A(n5968), .B(n5967), .Z(n5969) );
  AND U6175 ( .A(n5970), .B(n5969), .Z(n5988) );
  XNOR U6176 ( .A(n5989), .B(n5988), .Z(n5990) );
  NANDN U6177 ( .A(n5972), .B(n5971), .Z(n5976) );
  NAND U6178 ( .A(n5974), .B(n5973), .Z(n5975) );
  NAND U6179 ( .A(n5976), .B(n5975), .Z(n5991) );
  XNOR U6180 ( .A(n5990), .B(n5991), .Z(n5982) );
  XNOR U6181 ( .A(n5983), .B(n5982), .Z(n5984) );
  XNOR U6182 ( .A(n5985), .B(n5984), .Z(n6018) );
  XNOR U6183 ( .A(sreg[397]), .B(n6018), .Z(n6020) );
  NANDN U6184 ( .A(sreg[396]), .B(n5977), .Z(n5981) );
  NAND U6185 ( .A(n5979), .B(n5978), .Z(n5980) );
  NAND U6186 ( .A(n5981), .B(n5980), .Z(n6019) );
  XNOR U6187 ( .A(n6020), .B(n6019), .Z(c[397]) );
  NANDN U6188 ( .A(n5983), .B(n5982), .Z(n5987) );
  NANDN U6189 ( .A(n5985), .B(n5984), .Z(n5986) );
  AND U6190 ( .A(n5987), .B(n5986), .Z(n6026) );
  NANDN U6191 ( .A(n5989), .B(n5988), .Z(n5993) );
  NANDN U6192 ( .A(n5991), .B(n5990), .Z(n5992) );
  AND U6193 ( .A(n5993), .B(n5992), .Z(n6024) );
  NAND U6194 ( .A(n26), .B(n5994), .Z(n5996) );
  XOR U6195 ( .A(b[7]), .B(a[144]), .Z(n6035) );
  NAND U6196 ( .A(n10531), .B(n6035), .Z(n5995) );
  AND U6197 ( .A(n5996), .B(n5995), .Z(n6054) );
  NAND U6198 ( .A(n23), .B(n5997), .Z(n5999) );
  XOR U6199 ( .A(b[3]), .B(a[148]), .Z(n6038) );
  NAND U6200 ( .A(n24), .B(n6038), .Z(n5998) );
  NAND U6201 ( .A(n5999), .B(n5998), .Z(n6053) );
  XNOR U6202 ( .A(n6054), .B(n6053), .Z(n6056) );
  NAND U6203 ( .A(n25), .B(n6000), .Z(n6002) );
  XOR U6204 ( .A(b[5]), .B(a[146]), .Z(n6044) );
  NAND U6205 ( .A(n10456), .B(n6044), .Z(n6001) );
  AND U6206 ( .A(n6002), .B(n6001), .Z(n6048) );
  AND U6207 ( .A(b[7]), .B(a[142]), .Z(n6047) );
  XNOR U6208 ( .A(n6048), .B(n6047), .Z(n6049) );
  NAND U6209 ( .A(b[0]), .B(a[150]), .Z(n6003) );
  XNOR U6210 ( .A(b[1]), .B(n6003), .Z(n6005) );
  NANDN U6211 ( .A(b[0]), .B(a[149]), .Z(n6004) );
  NAND U6212 ( .A(n6005), .B(n6004), .Z(n6050) );
  XNOR U6213 ( .A(n6049), .B(n6050), .Z(n6055) );
  XOR U6214 ( .A(n6056), .B(n6055), .Z(n6030) );
  NANDN U6215 ( .A(n6007), .B(n6006), .Z(n6011) );
  NANDN U6216 ( .A(n6009), .B(n6008), .Z(n6010) );
  AND U6217 ( .A(n6011), .B(n6010), .Z(n6029) );
  XNOR U6218 ( .A(n6030), .B(n6029), .Z(n6031) );
  NANDN U6219 ( .A(n6013), .B(n6012), .Z(n6017) );
  NAND U6220 ( .A(n6015), .B(n6014), .Z(n6016) );
  NAND U6221 ( .A(n6017), .B(n6016), .Z(n6032) );
  XNOR U6222 ( .A(n6031), .B(n6032), .Z(n6023) );
  XNOR U6223 ( .A(n6024), .B(n6023), .Z(n6025) );
  XNOR U6224 ( .A(n6026), .B(n6025), .Z(n6059) );
  XNOR U6225 ( .A(sreg[398]), .B(n6059), .Z(n6061) );
  NANDN U6226 ( .A(sreg[397]), .B(n6018), .Z(n6022) );
  NAND U6227 ( .A(n6020), .B(n6019), .Z(n6021) );
  NAND U6228 ( .A(n6022), .B(n6021), .Z(n6060) );
  XNOR U6229 ( .A(n6061), .B(n6060), .Z(c[398]) );
  NANDN U6230 ( .A(n6024), .B(n6023), .Z(n6028) );
  NANDN U6231 ( .A(n6026), .B(n6025), .Z(n6027) );
  AND U6232 ( .A(n6028), .B(n6027), .Z(n6067) );
  NANDN U6233 ( .A(n6030), .B(n6029), .Z(n6034) );
  NANDN U6234 ( .A(n6032), .B(n6031), .Z(n6033) );
  AND U6235 ( .A(n6034), .B(n6033), .Z(n6065) );
  NAND U6236 ( .A(n26), .B(n6035), .Z(n6037) );
  XOR U6237 ( .A(b[7]), .B(a[145]), .Z(n6076) );
  NAND U6238 ( .A(n10531), .B(n6076), .Z(n6036) );
  AND U6239 ( .A(n6037), .B(n6036), .Z(n6095) );
  NAND U6240 ( .A(n23), .B(n6038), .Z(n6040) );
  XOR U6241 ( .A(b[3]), .B(a[149]), .Z(n6079) );
  NAND U6242 ( .A(n24), .B(n6079), .Z(n6039) );
  NAND U6243 ( .A(n6040), .B(n6039), .Z(n6094) );
  XNOR U6244 ( .A(n6095), .B(n6094), .Z(n6097) );
  NAND U6245 ( .A(b[0]), .B(a[151]), .Z(n6041) );
  XNOR U6246 ( .A(b[1]), .B(n6041), .Z(n6043) );
  NANDN U6247 ( .A(b[0]), .B(a[150]), .Z(n6042) );
  NAND U6248 ( .A(n6043), .B(n6042), .Z(n6091) );
  NAND U6249 ( .A(n25), .B(n6044), .Z(n6046) );
  XOR U6250 ( .A(b[5]), .B(a[147]), .Z(n6085) );
  NAND U6251 ( .A(n10456), .B(n6085), .Z(n6045) );
  AND U6252 ( .A(n6046), .B(n6045), .Z(n6089) );
  AND U6253 ( .A(b[7]), .B(a[143]), .Z(n6088) );
  XNOR U6254 ( .A(n6089), .B(n6088), .Z(n6090) );
  XNOR U6255 ( .A(n6091), .B(n6090), .Z(n6096) );
  XOR U6256 ( .A(n6097), .B(n6096), .Z(n6071) );
  NANDN U6257 ( .A(n6048), .B(n6047), .Z(n6052) );
  NANDN U6258 ( .A(n6050), .B(n6049), .Z(n6051) );
  AND U6259 ( .A(n6052), .B(n6051), .Z(n6070) );
  XNOR U6260 ( .A(n6071), .B(n6070), .Z(n6072) );
  NANDN U6261 ( .A(n6054), .B(n6053), .Z(n6058) );
  NAND U6262 ( .A(n6056), .B(n6055), .Z(n6057) );
  NAND U6263 ( .A(n6058), .B(n6057), .Z(n6073) );
  XNOR U6264 ( .A(n6072), .B(n6073), .Z(n6064) );
  XNOR U6265 ( .A(n6065), .B(n6064), .Z(n6066) );
  XNOR U6266 ( .A(n6067), .B(n6066), .Z(n6100) );
  XNOR U6267 ( .A(sreg[399]), .B(n6100), .Z(n6102) );
  NANDN U6268 ( .A(sreg[398]), .B(n6059), .Z(n6063) );
  NAND U6269 ( .A(n6061), .B(n6060), .Z(n6062) );
  NAND U6270 ( .A(n6063), .B(n6062), .Z(n6101) );
  XNOR U6271 ( .A(n6102), .B(n6101), .Z(c[399]) );
  NANDN U6272 ( .A(n6065), .B(n6064), .Z(n6069) );
  NANDN U6273 ( .A(n6067), .B(n6066), .Z(n6068) );
  AND U6274 ( .A(n6069), .B(n6068), .Z(n6108) );
  NANDN U6275 ( .A(n6071), .B(n6070), .Z(n6075) );
  NANDN U6276 ( .A(n6073), .B(n6072), .Z(n6074) );
  AND U6277 ( .A(n6075), .B(n6074), .Z(n6106) );
  NAND U6278 ( .A(n26), .B(n6076), .Z(n6078) );
  XOR U6279 ( .A(b[7]), .B(a[146]), .Z(n6117) );
  NAND U6280 ( .A(n10531), .B(n6117), .Z(n6077) );
  AND U6281 ( .A(n6078), .B(n6077), .Z(n6136) );
  NAND U6282 ( .A(n23), .B(n6079), .Z(n6081) );
  XOR U6283 ( .A(b[3]), .B(a[150]), .Z(n6120) );
  NAND U6284 ( .A(n24), .B(n6120), .Z(n6080) );
  NAND U6285 ( .A(n6081), .B(n6080), .Z(n6135) );
  XNOR U6286 ( .A(n6136), .B(n6135), .Z(n6138) );
  NAND U6287 ( .A(b[0]), .B(a[152]), .Z(n6082) );
  XNOR U6288 ( .A(b[1]), .B(n6082), .Z(n6084) );
  NANDN U6289 ( .A(b[0]), .B(a[151]), .Z(n6083) );
  NAND U6290 ( .A(n6084), .B(n6083), .Z(n6132) );
  NAND U6291 ( .A(n25), .B(n6085), .Z(n6087) );
  XOR U6292 ( .A(b[5]), .B(a[148]), .Z(n6123) );
  NAND U6293 ( .A(n10456), .B(n6123), .Z(n6086) );
  AND U6294 ( .A(n6087), .B(n6086), .Z(n6130) );
  AND U6295 ( .A(b[7]), .B(a[144]), .Z(n6129) );
  XNOR U6296 ( .A(n6130), .B(n6129), .Z(n6131) );
  XNOR U6297 ( .A(n6132), .B(n6131), .Z(n6137) );
  XOR U6298 ( .A(n6138), .B(n6137), .Z(n6112) );
  NANDN U6299 ( .A(n6089), .B(n6088), .Z(n6093) );
  NANDN U6300 ( .A(n6091), .B(n6090), .Z(n6092) );
  AND U6301 ( .A(n6093), .B(n6092), .Z(n6111) );
  XNOR U6302 ( .A(n6112), .B(n6111), .Z(n6113) );
  NANDN U6303 ( .A(n6095), .B(n6094), .Z(n6099) );
  NAND U6304 ( .A(n6097), .B(n6096), .Z(n6098) );
  NAND U6305 ( .A(n6099), .B(n6098), .Z(n6114) );
  XNOR U6306 ( .A(n6113), .B(n6114), .Z(n6105) );
  XNOR U6307 ( .A(n6106), .B(n6105), .Z(n6107) );
  XNOR U6308 ( .A(n6108), .B(n6107), .Z(n6141) );
  XNOR U6309 ( .A(sreg[400]), .B(n6141), .Z(n6143) );
  NANDN U6310 ( .A(sreg[399]), .B(n6100), .Z(n6104) );
  NAND U6311 ( .A(n6102), .B(n6101), .Z(n6103) );
  NAND U6312 ( .A(n6104), .B(n6103), .Z(n6142) );
  XNOR U6313 ( .A(n6143), .B(n6142), .Z(c[400]) );
  NANDN U6314 ( .A(n6106), .B(n6105), .Z(n6110) );
  NANDN U6315 ( .A(n6108), .B(n6107), .Z(n6109) );
  AND U6316 ( .A(n6110), .B(n6109), .Z(n6149) );
  NANDN U6317 ( .A(n6112), .B(n6111), .Z(n6116) );
  NANDN U6318 ( .A(n6114), .B(n6113), .Z(n6115) );
  AND U6319 ( .A(n6116), .B(n6115), .Z(n6147) );
  NAND U6320 ( .A(n26), .B(n6117), .Z(n6119) );
  XOR U6321 ( .A(b[7]), .B(a[147]), .Z(n6158) );
  NAND U6322 ( .A(n10531), .B(n6158), .Z(n6118) );
  AND U6323 ( .A(n6119), .B(n6118), .Z(n6177) );
  NAND U6324 ( .A(n23), .B(n6120), .Z(n6122) );
  XOR U6325 ( .A(b[3]), .B(a[151]), .Z(n6161) );
  NAND U6326 ( .A(n24), .B(n6161), .Z(n6121) );
  NAND U6327 ( .A(n6122), .B(n6121), .Z(n6176) );
  XNOR U6328 ( .A(n6177), .B(n6176), .Z(n6179) );
  NAND U6329 ( .A(n25), .B(n6123), .Z(n6125) );
  XOR U6330 ( .A(b[5]), .B(a[149]), .Z(n6167) );
  NAND U6331 ( .A(n10456), .B(n6167), .Z(n6124) );
  AND U6332 ( .A(n6125), .B(n6124), .Z(n6171) );
  AND U6333 ( .A(b[7]), .B(a[145]), .Z(n6170) );
  XNOR U6334 ( .A(n6171), .B(n6170), .Z(n6172) );
  NAND U6335 ( .A(b[0]), .B(a[153]), .Z(n6126) );
  XNOR U6336 ( .A(b[1]), .B(n6126), .Z(n6128) );
  NANDN U6337 ( .A(b[0]), .B(a[152]), .Z(n6127) );
  NAND U6338 ( .A(n6128), .B(n6127), .Z(n6173) );
  XNOR U6339 ( .A(n6172), .B(n6173), .Z(n6178) );
  XOR U6340 ( .A(n6179), .B(n6178), .Z(n6153) );
  NANDN U6341 ( .A(n6130), .B(n6129), .Z(n6134) );
  NANDN U6342 ( .A(n6132), .B(n6131), .Z(n6133) );
  AND U6343 ( .A(n6134), .B(n6133), .Z(n6152) );
  XNOR U6344 ( .A(n6153), .B(n6152), .Z(n6154) );
  NANDN U6345 ( .A(n6136), .B(n6135), .Z(n6140) );
  NAND U6346 ( .A(n6138), .B(n6137), .Z(n6139) );
  NAND U6347 ( .A(n6140), .B(n6139), .Z(n6155) );
  XNOR U6348 ( .A(n6154), .B(n6155), .Z(n6146) );
  XNOR U6349 ( .A(n6147), .B(n6146), .Z(n6148) );
  XNOR U6350 ( .A(n6149), .B(n6148), .Z(n6182) );
  XNOR U6351 ( .A(sreg[401]), .B(n6182), .Z(n6184) );
  NANDN U6352 ( .A(sreg[400]), .B(n6141), .Z(n6145) );
  NAND U6353 ( .A(n6143), .B(n6142), .Z(n6144) );
  NAND U6354 ( .A(n6145), .B(n6144), .Z(n6183) );
  XNOR U6355 ( .A(n6184), .B(n6183), .Z(c[401]) );
  NANDN U6356 ( .A(n6147), .B(n6146), .Z(n6151) );
  NANDN U6357 ( .A(n6149), .B(n6148), .Z(n6150) );
  AND U6358 ( .A(n6151), .B(n6150), .Z(n6190) );
  NANDN U6359 ( .A(n6153), .B(n6152), .Z(n6157) );
  NANDN U6360 ( .A(n6155), .B(n6154), .Z(n6156) );
  AND U6361 ( .A(n6157), .B(n6156), .Z(n6188) );
  NAND U6362 ( .A(n26), .B(n6158), .Z(n6160) );
  XOR U6363 ( .A(b[7]), .B(a[148]), .Z(n6199) );
  NAND U6364 ( .A(n10531), .B(n6199), .Z(n6159) );
  AND U6365 ( .A(n6160), .B(n6159), .Z(n6218) );
  NAND U6366 ( .A(n23), .B(n6161), .Z(n6163) );
  XOR U6367 ( .A(b[3]), .B(a[152]), .Z(n6202) );
  NAND U6368 ( .A(n24), .B(n6202), .Z(n6162) );
  NAND U6369 ( .A(n6163), .B(n6162), .Z(n6217) );
  XNOR U6370 ( .A(n6218), .B(n6217), .Z(n6220) );
  NAND U6371 ( .A(b[0]), .B(a[154]), .Z(n6164) );
  XNOR U6372 ( .A(b[1]), .B(n6164), .Z(n6166) );
  NANDN U6373 ( .A(b[0]), .B(a[153]), .Z(n6165) );
  NAND U6374 ( .A(n6166), .B(n6165), .Z(n6214) );
  NAND U6375 ( .A(n25), .B(n6167), .Z(n6169) );
  XOR U6376 ( .A(b[5]), .B(a[150]), .Z(n6208) );
  NAND U6377 ( .A(n10456), .B(n6208), .Z(n6168) );
  AND U6378 ( .A(n6169), .B(n6168), .Z(n6212) );
  AND U6379 ( .A(b[7]), .B(a[146]), .Z(n6211) );
  XNOR U6380 ( .A(n6212), .B(n6211), .Z(n6213) );
  XNOR U6381 ( .A(n6214), .B(n6213), .Z(n6219) );
  XOR U6382 ( .A(n6220), .B(n6219), .Z(n6194) );
  NANDN U6383 ( .A(n6171), .B(n6170), .Z(n6175) );
  NANDN U6384 ( .A(n6173), .B(n6172), .Z(n6174) );
  AND U6385 ( .A(n6175), .B(n6174), .Z(n6193) );
  XNOR U6386 ( .A(n6194), .B(n6193), .Z(n6195) );
  NANDN U6387 ( .A(n6177), .B(n6176), .Z(n6181) );
  NAND U6388 ( .A(n6179), .B(n6178), .Z(n6180) );
  NAND U6389 ( .A(n6181), .B(n6180), .Z(n6196) );
  XNOR U6390 ( .A(n6195), .B(n6196), .Z(n6187) );
  XNOR U6391 ( .A(n6188), .B(n6187), .Z(n6189) );
  XNOR U6392 ( .A(n6190), .B(n6189), .Z(n6223) );
  XNOR U6393 ( .A(sreg[402]), .B(n6223), .Z(n6225) );
  NANDN U6394 ( .A(sreg[401]), .B(n6182), .Z(n6186) );
  NAND U6395 ( .A(n6184), .B(n6183), .Z(n6185) );
  NAND U6396 ( .A(n6186), .B(n6185), .Z(n6224) );
  XNOR U6397 ( .A(n6225), .B(n6224), .Z(c[402]) );
  NANDN U6398 ( .A(n6188), .B(n6187), .Z(n6192) );
  NANDN U6399 ( .A(n6190), .B(n6189), .Z(n6191) );
  AND U6400 ( .A(n6192), .B(n6191), .Z(n6231) );
  NANDN U6401 ( .A(n6194), .B(n6193), .Z(n6198) );
  NANDN U6402 ( .A(n6196), .B(n6195), .Z(n6197) );
  AND U6403 ( .A(n6198), .B(n6197), .Z(n6229) );
  NAND U6404 ( .A(n26), .B(n6199), .Z(n6201) );
  XOR U6405 ( .A(b[7]), .B(a[149]), .Z(n6240) );
  NAND U6406 ( .A(n10531), .B(n6240), .Z(n6200) );
  AND U6407 ( .A(n6201), .B(n6200), .Z(n6259) );
  NAND U6408 ( .A(n23), .B(n6202), .Z(n6204) );
  XOR U6409 ( .A(b[3]), .B(a[153]), .Z(n6243) );
  NAND U6410 ( .A(n24), .B(n6243), .Z(n6203) );
  NAND U6411 ( .A(n6204), .B(n6203), .Z(n6258) );
  XNOR U6412 ( .A(n6259), .B(n6258), .Z(n6261) );
  NAND U6413 ( .A(b[0]), .B(a[155]), .Z(n6205) );
  XNOR U6414 ( .A(b[1]), .B(n6205), .Z(n6207) );
  NANDN U6415 ( .A(b[0]), .B(a[154]), .Z(n6206) );
  NAND U6416 ( .A(n6207), .B(n6206), .Z(n6255) );
  NAND U6417 ( .A(n25), .B(n6208), .Z(n6210) );
  XOR U6418 ( .A(b[5]), .B(a[151]), .Z(n6249) );
  NAND U6419 ( .A(n10456), .B(n6249), .Z(n6209) );
  AND U6420 ( .A(n6210), .B(n6209), .Z(n6253) );
  AND U6421 ( .A(b[7]), .B(a[147]), .Z(n6252) );
  XNOR U6422 ( .A(n6253), .B(n6252), .Z(n6254) );
  XNOR U6423 ( .A(n6255), .B(n6254), .Z(n6260) );
  XOR U6424 ( .A(n6261), .B(n6260), .Z(n6235) );
  NANDN U6425 ( .A(n6212), .B(n6211), .Z(n6216) );
  NANDN U6426 ( .A(n6214), .B(n6213), .Z(n6215) );
  AND U6427 ( .A(n6216), .B(n6215), .Z(n6234) );
  XNOR U6428 ( .A(n6235), .B(n6234), .Z(n6236) );
  NANDN U6429 ( .A(n6218), .B(n6217), .Z(n6222) );
  NAND U6430 ( .A(n6220), .B(n6219), .Z(n6221) );
  NAND U6431 ( .A(n6222), .B(n6221), .Z(n6237) );
  XNOR U6432 ( .A(n6236), .B(n6237), .Z(n6228) );
  XNOR U6433 ( .A(n6229), .B(n6228), .Z(n6230) );
  XNOR U6434 ( .A(n6231), .B(n6230), .Z(n6264) );
  XNOR U6435 ( .A(sreg[403]), .B(n6264), .Z(n6266) );
  NANDN U6436 ( .A(sreg[402]), .B(n6223), .Z(n6227) );
  NAND U6437 ( .A(n6225), .B(n6224), .Z(n6226) );
  NAND U6438 ( .A(n6227), .B(n6226), .Z(n6265) );
  XNOR U6439 ( .A(n6266), .B(n6265), .Z(c[403]) );
  NANDN U6440 ( .A(n6229), .B(n6228), .Z(n6233) );
  NANDN U6441 ( .A(n6231), .B(n6230), .Z(n6232) );
  AND U6442 ( .A(n6233), .B(n6232), .Z(n6272) );
  NANDN U6443 ( .A(n6235), .B(n6234), .Z(n6239) );
  NANDN U6444 ( .A(n6237), .B(n6236), .Z(n6238) );
  AND U6445 ( .A(n6239), .B(n6238), .Z(n6270) );
  NAND U6446 ( .A(n26), .B(n6240), .Z(n6242) );
  XOR U6447 ( .A(b[7]), .B(a[150]), .Z(n6281) );
  NAND U6448 ( .A(n10531), .B(n6281), .Z(n6241) );
  AND U6449 ( .A(n6242), .B(n6241), .Z(n6300) );
  NAND U6450 ( .A(n23), .B(n6243), .Z(n6245) );
  XOR U6451 ( .A(b[3]), .B(a[154]), .Z(n6284) );
  NAND U6452 ( .A(n24), .B(n6284), .Z(n6244) );
  NAND U6453 ( .A(n6245), .B(n6244), .Z(n6299) );
  XNOR U6454 ( .A(n6300), .B(n6299), .Z(n6302) );
  NAND U6455 ( .A(b[0]), .B(a[156]), .Z(n6246) );
  XNOR U6456 ( .A(b[1]), .B(n6246), .Z(n6248) );
  NANDN U6457 ( .A(b[0]), .B(a[155]), .Z(n6247) );
  NAND U6458 ( .A(n6248), .B(n6247), .Z(n6296) );
  NAND U6459 ( .A(n25), .B(n6249), .Z(n6251) );
  XOR U6460 ( .A(b[5]), .B(a[152]), .Z(n6290) );
  NAND U6461 ( .A(n10456), .B(n6290), .Z(n6250) );
  AND U6462 ( .A(n6251), .B(n6250), .Z(n6294) );
  AND U6463 ( .A(b[7]), .B(a[148]), .Z(n6293) );
  XNOR U6464 ( .A(n6294), .B(n6293), .Z(n6295) );
  XNOR U6465 ( .A(n6296), .B(n6295), .Z(n6301) );
  XOR U6466 ( .A(n6302), .B(n6301), .Z(n6276) );
  NANDN U6467 ( .A(n6253), .B(n6252), .Z(n6257) );
  NANDN U6468 ( .A(n6255), .B(n6254), .Z(n6256) );
  AND U6469 ( .A(n6257), .B(n6256), .Z(n6275) );
  XNOR U6470 ( .A(n6276), .B(n6275), .Z(n6277) );
  NANDN U6471 ( .A(n6259), .B(n6258), .Z(n6263) );
  NAND U6472 ( .A(n6261), .B(n6260), .Z(n6262) );
  NAND U6473 ( .A(n6263), .B(n6262), .Z(n6278) );
  XNOR U6474 ( .A(n6277), .B(n6278), .Z(n6269) );
  XNOR U6475 ( .A(n6270), .B(n6269), .Z(n6271) );
  XNOR U6476 ( .A(n6272), .B(n6271), .Z(n6305) );
  XNOR U6477 ( .A(sreg[404]), .B(n6305), .Z(n6307) );
  NANDN U6478 ( .A(sreg[403]), .B(n6264), .Z(n6268) );
  NAND U6479 ( .A(n6266), .B(n6265), .Z(n6267) );
  NAND U6480 ( .A(n6268), .B(n6267), .Z(n6306) );
  XNOR U6481 ( .A(n6307), .B(n6306), .Z(c[404]) );
  NANDN U6482 ( .A(n6270), .B(n6269), .Z(n6274) );
  NANDN U6483 ( .A(n6272), .B(n6271), .Z(n6273) );
  AND U6484 ( .A(n6274), .B(n6273), .Z(n6313) );
  NANDN U6485 ( .A(n6276), .B(n6275), .Z(n6280) );
  NANDN U6486 ( .A(n6278), .B(n6277), .Z(n6279) );
  AND U6487 ( .A(n6280), .B(n6279), .Z(n6311) );
  NAND U6488 ( .A(n26), .B(n6281), .Z(n6283) );
  XOR U6489 ( .A(b[7]), .B(a[151]), .Z(n6322) );
  NAND U6490 ( .A(n10531), .B(n6322), .Z(n6282) );
  AND U6491 ( .A(n6283), .B(n6282), .Z(n6341) );
  NAND U6492 ( .A(n23), .B(n6284), .Z(n6286) );
  XOR U6493 ( .A(b[3]), .B(a[155]), .Z(n6325) );
  NAND U6494 ( .A(n24), .B(n6325), .Z(n6285) );
  NAND U6495 ( .A(n6286), .B(n6285), .Z(n6340) );
  XNOR U6496 ( .A(n6341), .B(n6340), .Z(n6343) );
  NAND U6497 ( .A(b[0]), .B(a[157]), .Z(n6287) );
  XNOR U6498 ( .A(b[1]), .B(n6287), .Z(n6289) );
  NANDN U6499 ( .A(b[0]), .B(a[156]), .Z(n6288) );
  NAND U6500 ( .A(n6289), .B(n6288), .Z(n6337) );
  NAND U6501 ( .A(n25), .B(n6290), .Z(n6292) );
  XOR U6502 ( .A(b[5]), .B(a[153]), .Z(n6331) );
  NAND U6503 ( .A(n10456), .B(n6331), .Z(n6291) );
  AND U6504 ( .A(n6292), .B(n6291), .Z(n6335) );
  AND U6505 ( .A(b[7]), .B(a[149]), .Z(n6334) );
  XNOR U6506 ( .A(n6335), .B(n6334), .Z(n6336) );
  XNOR U6507 ( .A(n6337), .B(n6336), .Z(n6342) );
  XOR U6508 ( .A(n6343), .B(n6342), .Z(n6317) );
  NANDN U6509 ( .A(n6294), .B(n6293), .Z(n6298) );
  NANDN U6510 ( .A(n6296), .B(n6295), .Z(n6297) );
  AND U6511 ( .A(n6298), .B(n6297), .Z(n6316) );
  XNOR U6512 ( .A(n6317), .B(n6316), .Z(n6318) );
  NANDN U6513 ( .A(n6300), .B(n6299), .Z(n6304) );
  NAND U6514 ( .A(n6302), .B(n6301), .Z(n6303) );
  NAND U6515 ( .A(n6304), .B(n6303), .Z(n6319) );
  XNOR U6516 ( .A(n6318), .B(n6319), .Z(n6310) );
  XNOR U6517 ( .A(n6311), .B(n6310), .Z(n6312) );
  XNOR U6518 ( .A(n6313), .B(n6312), .Z(n6346) );
  XNOR U6519 ( .A(sreg[405]), .B(n6346), .Z(n6348) );
  NANDN U6520 ( .A(sreg[404]), .B(n6305), .Z(n6309) );
  NAND U6521 ( .A(n6307), .B(n6306), .Z(n6308) );
  NAND U6522 ( .A(n6309), .B(n6308), .Z(n6347) );
  XNOR U6523 ( .A(n6348), .B(n6347), .Z(c[405]) );
  NANDN U6524 ( .A(n6311), .B(n6310), .Z(n6315) );
  NANDN U6525 ( .A(n6313), .B(n6312), .Z(n6314) );
  AND U6526 ( .A(n6315), .B(n6314), .Z(n6354) );
  NANDN U6527 ( .A(n6317), .B(n6316), .Z(n6321) );
  NANDN U6528 ( .A(n6319), .B(n6318), .Z(n6320) );
  AND U6529 ( .A(n6321), .B(n6320), .Z(n6352) );
  NAND U6530 ( .A(n26), .B(n6322), .Z(n6324) );
  XOR U6531 ( .A(b[7]), .B(a[152]), .Z(n6363) );
  NAND U6532 ( .A(n10531), .B(n6363), .Z(n6323) );
  AND U6533 ( .A(n6324), .B(n6323), .Z(n6382) );
  NAND U6534 ( .A(n23), .B(n6325), .Z(n6327) );
  XOR U6535 ( .A(b[3]), .B(a[156]), .Z(n6366) );
  NAND U6536 ( .A(n24), .B(n6366), .Z(n6326) );
  NAND U6537 ( .A(n6327), .B(n6326), .Z(n6381) );
  XNOR U6538 ( .A(n6382), .B(n6381), .Z(n6384) );
  NAND U6539 ( .A(b[0]), .B(a[158]), .Z(n6328) );
  XNOR U6540 ( .A(b[1]), .B(n6328), .Z(n6330) );
  NANDN U6541 ( .A(b[0]), .B(a[157]), .Z(n6329) );
  NAND U6542 ( .A(n6330), .B(n6329), .Z(n6378) );
  NAND U6543 ( .A(n25), .B(n6331), .Z(n6333) );
  XOR U6544 ( .A(b[5]), .B(a[154]), .Z(n6372) );
  NAND U6545 ( .A(n10456), .B(n6372), .Z(n6332) );
  AND U6546 ( .A(n6333), .B(n6332), .Z(n6376) );
  AND U6547 ( .A(b[7]), .B(a[150]), .Z(n6375) );
  XNOR U6548 ( .A(n6376), .B(n6375), .Z(n6377) );
  XNOR U6549 ( .A(n6378), .B(n6377), .Z(n6383) );
  XOR U6550 ( .A(n6384), .B(n6383), .Z(n6358) );
  NANDN U6551 ( .A(n6335), .B(n6334), .Z(n6339) );
  NANDN U6552 ( .A(n6337), .B(n6336), .Z(n6338) );
  AND U6553 ( .A(n6339), .B(n6338), .Z(n6357) );
  XNOR U6554 ( .A(n6358), .B(n6357), .Z(n6359) );
  NANDN U6555 ( .A(n6341), .B(n6340), .Z(n6345) );
  NAND U6556 ( .A(n6343), .B(n6342), .Z(n6344) );
  NAND U6557 ( .A(n6345), .B(n6344), .Z(n6360) );
  XNOR U6558 ( .A(n6359), .B(n6360), .Z(n6351) );
  XNOR U6559 ( .A(n6352), .B(n6351), .Z(n6353) );
  XNOR U6560 ( .A(n6354), .B(n6353), .Z(n6387) );
  XNOR U6561 ( .A(sreg[406]), .B(n6387), .Z(n6389) );
  NANDN U6562 ( .A(sreg[405]), .B(n6346), .Z(n6350) );
  NAND U6563 ( .A(n6348), .B(n6347), .Z(n6349) );
  NAND U6564 ( .A(n6350), .B(n6349), .Z(n6388) );
  XNOR U6565 ( .A(n6389), .B(n6388), .Z(c[406]) );
  NANDN U6566 ( .A(n6352), .B(n6351), .Z(n6356) );
  NANDN U6567 ( .A(n6354), .B(n6353), .Z(n6355) );
  AND U6568 ( .A(n6356), .B(n6355), .Z(n6395) );
  NANDN U6569 ( .A(n6358), .B(n6357), .Z(n6362) );
  NANDN U6570 ( .A(n6360), .B(n6359), .Z(n6361) );
  AND U6571 ( .A(n6362), .B(n6361), .Z(n6393) );
  NAND U6572 ( .A(n26), .B(n6363), .Z(n6365) );
  XOR U6573 ( .A(b[7]), .B(a[153]), .Z(n6404) );
  NAND U6574 ( .A(n10531), .B(n6404), .Z(n6364) );
  AND U6575 ( .A(n6365), .B(n6364), .Z(n6423) );
  NAND U6576 ( .A(n23), .B(n6366), .Z(n6368) );
  XOR U6577 ( .A(b[3]), .B(a[157]), .Z(n6407) );
  NAND U6578 ( .A(n24), .B(n6407), .Z(n6367) );
  NAND U6579 ( .A(n6368), .B(n6367), .Z(n6422) );
  XNOR U6580 ( .A(n6423), .B(n6422), .Z(n6425) );
  NAND U6581 ( .A(b[0]), .B(a[159]), .Z(n6369) );
  XNOR U6582 ( .A(b[1]), .B(n6369), .Z(n6371) );
  NANDN U6583 ( .A(b[0]), .B(a[158]), .Z(n6370) );
  NAND U6584 ( .A(n6371), .B(n6370), .Z(n6419) );
  NAND U6585 ( .A(n25), .B(n6372), .Z(n6374) );
  XOR U6586 ( .A(b[5]), .B(a[155]), .Z(n6413) );
  NAND U6587 ( .A(n10456), .B(n6413), .Z(n6373) );
  AND U6588 ( .A(n6374), .B(n6373), .Z(n6417) );
  AND U6589 ( .A(b[7]), .B(a[151]), .Z(n6416) );
  XNOR U6590 ( .A(n6417), .B(n6416), .Z(n6418) );
  XNOR U6591 ( .A(n6419), .B(n6418), .Z(n6424) );
  XOR U6592 ( .A(n6425), .B(n6424), .Z(n6399) );
  NANDN U6593 ( .A(n6376), .B(n6375), .Z(n6380) );
  NANDN U6594 ( .A(n6378), .B(n6377), .Z(n6379) );
  AND U6595 ( .A(n6380), .B(n6379), .Z(n6398) );
  XNOR U6596 ( .A(n6399), .B(n6398), .Z(n6400) );
  NANDN U6597 ( .A(n6382), .B(n6381), .Z(n6386) );
  NAND U6598 ( .A(n6384), .B(n6383), .Z(n6385) );
  NAND U6599 ( .A(n6386), .B(n6385), .Z(n6401) );
  XNOR U6600 ( .A(n6400), .B(n6401), .Z(n6392) );
  XNOR U6601 ( .A(n6393), .B(n6392), .Z(n6394) );
  XNOR U6602 ( .A(n6395), .B(n6394), .Z(n6428) );
  XNOR U6603 ( .A(sreg[407]), .B(n6428), .Z(n6430) );
  NANDN U6604 ( .A(sreg[406]), .B(n6387), .Z(n6391) );
  NAND U6605 ( .A(n6389), .B(n6388), .Z(n6390) );
  NAND U6606 ( .A(n6391), .B(n6390), .Z(n6429) );
  XNOR U6607 ( .A(n6430), .B(n6429), .Z(c[407]) );
  NANDN U6608 ( .A(n6393), .B(n6392), .Z(n6397) );
  NANDN U6609 ( .A(n6395), .B(n6394), .Z(n6396) );
  AND U6610 ( .A(n6397), .B(n6396), .Z(n6436) );
  NANDN U6611 ( .A(n6399), .B(n6398), .Z(n6403) );
  NANDN U6612 ( .A(n6401), .B(n6400), .Z(n6402) );
  AND U6613 ( .A(n6403), .B(n6402), .Z(n6434) );
  NAND U6614 ( .A(n26), .B(n6404), .Z(n6406) );
  XOR U6615 ( .A(b[7]), .B(a[154]), .Z(n6445) );
  NAND U6616 ( .A(n10531), .B(n6445), .Z(n6405) );
  AND U6617 ( .A(n6406), .B(n6405), .Z(n6464) );
  NAND U6618 ( .A(n23), .B(n6407), .Z(n6409) );
  XOR U6619 ( .A(b[3]), .B(a[158]), .Z(n6448) );
  NAND U6620 ( .A(n24), .B(n6448), .Z(n6408) );
  NAND U6621 ( .A(n6409), .B(n6408), .Z(n6463) );
  XNOR U6622 ( .A(n6464), .B(n6463), .Z(n6466) );
  NAND U6623 ( .A(b[0]), .B(a[160]), .Z(n6410) );
  XNOR U6624 ( .A(b[1]), .B(n6410), .Z(n6412) );
  NANDN U6625 ( .A(b[0]), .B(a[159]), .Z(n6411) );
  NAND U6626 ( .A(n6412), .B(n6411), .Z(n6460) );
  NAND U6627 ( .A(n25), .B(n6413), .Z(n6415) );
  XOR U6628 ( .A(b[5]), .B(a[156]), .Z(n6454) );
  NAND U6629 ( .A(n10456), .B(n6454), .Z(n6414) );
  AND U6630 ( .A(n6415), .B(n6414), .Z(n6458) );
  AND U6631 ( .A(b[7]), .B(a[152]), .Z(n6457) );
  XNOR U6632 ( .A(n6458), .B(n6457), .Z(n6459) );
  XNOR U6633 ( .A(n6460), .B(n6459), .Z(n6465) );
  XOR U6634 ( .A(n6466), .B(n6465), .Z(n6440) );
  NANDN U6635 ( .A(n6417), .B(n6416), .Z(n6421) );
  NANDN U6636 ( .A(n6419), .B(n6418), .Z(n6420) );
  AND U6637 ( .A(n6421), .B(n6420), .Z(n6439) );
  XNOR U6638 ( .A(n6440), .B(n6439), .Z(n6441) );
  NANDN U6639 ( .A(n6423), .B(n6422), .Z(n6427) );
  NAND U6640 ( .A(n6425), .B(n6424), .Z(n6426) );
  NAND U6641 ( .A(n6427), .B(n6426), .Z(n6442) );
  XNOR U6642 ( .A(n6441), .B(n6442), .Z(n6433) );
  XNOR U6643 ( .A(n6434), .B(n6433), .Z(n6435) );
  XNOR U6644 ( .A(n6436), .B(n6435), .Z(n6469) );
  XNOR U6645 ( .A(sreg[408]), .B(n6469), .Z(n6471) );
  NANDN U6646 ( .A(sreg[407]), .B(n6428), .Z(n6432) );
  NAND U6647 ( .A(n6430), .B(n6429), .Z(n6431) );
  NAND U6648 ( .A(n6432), .B(n6431), .Z(n6470) );
  XNOR U6649 ( .A(n6471), .B(n6470), .Z(c[408]) );
  NANDN U6650 ( .A(n6434), .B(n6433), .Z(n6438) );
  NANDN U6651 ( .A(n6436), .B(n6435), .Z(n6437) );
  AND U6652 ( .A(n6438), .B(n6437), .Z(n6477) );
  NANDN U6653 ( .A(n6440), .B(n6439), .Z(n6444) );
  NANDN U6654 ( .A(n6442), .B(n6441), .Z(n6443) );
  AND U6655 ( .A(n6444), .B(n6443), .Z(n6475) );
  NAND U6656 ( .A(n26), .B(n6445), .Z(n6447) );
  XOR U6657 ( .A(b[7]), .B(a[155]), .Z(n6486) );
  NAND U6658 ( .A(n10531), .B(n6486), .Z(n6446) );
  AND U6659 ( .A(n6447), .B(n6446), .Z(n6505) );
  NAND U6660 ( .A(n23), .B(n6448), .Z(n6450) );
  XOR U6661 ( .A(b[3]), .B(a[159]), .Z(n6489) );
  NAND U6662 ( .A(n24), .B(n6489), .Z(n6449) );
  NAND U6663 ( .A(n6450), .B(n6449), .Z(n6504) );
  XNOR U6664 ( .A(n6505), .B(n6504), .Z(n6507) );
  NAND U6665 ( .A(b[0]), .B(a[161]), .Z(n6451) );
  XNOR U6666 ( .A(b[1]), .B(n6451), .Z(n6453) );
  NANDN U6667 ( .A(b[0]), .B(a[160]), .Z(n6452) );
  NAND U6668 ( .A(n6453), .B(n6452), .Z(n6501) );
  NAND U6669 ( .A(n25), .B(n6454), .Z(n6456) );
  XOR U6670 ( .A(b[5]), .B(a[157]), .Z(n6495) );
  NAND U6671 ( .A(n10456), .B(n6495), .Z(n6455) );
  AND U6672 ( .A(n6456), .B(n6455), .Z(n6499) );
  AND U6673 ( .A(b[7]), .B(a[153]), .Z(n6498) );
  XNOR U6674 ( .A(n6499), .B(n6498), .Z(n6500) );
  XNOR U6675 ( .A(n6501), .B(n6500), .Z(n6506) );
  XOR U6676 ( .A(n6507), .B(n6506), .Z(n6481) );
  NANDN U6677 ( .A(n6458), .B(n6457), .Z(n6462) );
  NANDN U6678 ( .A(n6460), .B(n6459), .Z(n6461) );
  AND U6679 ( .A(n6462), .B(n6461), .Z(n6480) );
  XNOR U6680 ( .A(n6481), .B(n6480), .Z(n6482) );
  NANDN U6681 ( .A(n6464), .B(n6463), .Z(n6468) );
  NAND U6682 ( .A(n6466), .B(n6465), .Z(n6467) );
  NAND U6683 ( .A(n6468), .B(n6467), .Z(n6483) );
  XNOR U6684 ( .A(n6482), .B(n6483), .Z(n6474) );
  XNOR U6685 ( .A(n6475), .B(n6474), .Z(n6476) );
  XNOR U6686 ( .A(n6477), .B(n6476), .Z(n6510) );
  XNOR U6687 ( .A(sreg[409]), .B(n6510), .Z(n6512) );
  NANDN U6688 ( .A(sreg[408]), .B(n6469), .Z(n6473) );
  NAND U6689 ( .A(n6471), .B(n6470), .Z(n6472) );
  NAND U6690 ( .A(n6473), .B(n6472), .Z(n6511) );
  XNOR U6691 ( .A(n6512), .B(n6511), .Z(c[409]) );
  NANDN U6692 ( .A(n6475), .B(n6474), .Z(n6479) );
  NANDN U6693 ( .A(n6477), .B(n6476), .Z(n6478) );
  AND U6694 ( .A(n6479), .B(n6478), .Z(n6518) );
  NANDN U6695 ( .A(n6481), .B(n6480), .Z(n6485) );
  NANDN U6696 ( .A(n6483), .B(n6482), .Z(n6484) );
  AND U6697 ( .A(n6485), .B(n6484), .Z(n6516) );
  NAND U6698 ( .A(n26), .B(n6486), .Z(n6488) );
  XOR U6699 ( .A(b[7]), .B(a[156]), .Z(n6527) );
  NAND U6700 ( .A(n10531), .B(n6527), .Z(n6487) );
  AND U6701 ( .A(n6488), .B(n6487), .Z(n6546) );
  NAND U6702 ( .A(n23), .B(n6489), .Z(n6491) );
  XOR U6703 ( .A(b[3]), .B(a[160]), .Z(n6530) );
  NAND U6704 ( .A(n24), .B(n6530), .Z(n6490) );
  NAND U6705 ( .A(n6491), .B(n6490), .Z(n6545) );
  XNOR U6706 ( .A(n6546), .B(n6545), .Z(n6548) );
  NAND U6707 ( .A(b[0]), .B(a[162]), .Z(n6492) );
  XNOR U6708 ( .A(b[1]), .B(n6492), .Z(n6494) );
  NANDN U6709 ( .A(b[0]), .B(a[161]), .Z(n6493) );
  NAND U6710 ( .A(n6494), .B(n6493), .Z(n6542) );
  NAND U6711 ( .A(n25), .B(n6495), .Z(n6497) );
  XOR U6712 ( .A(b[5]), .B(a[158]), .Z(n6536) );
  NAND U6713 ( .A(n10456), .B(n6536), .Z(n6496) );
  AND U6714 ( .A(n6497), .B(n6496), .Z(n6540) );
  AND U6715 ( .A(b[7]), .B(a[154]), .Z(n6539) );
  XNOR U6716 ( .A(n6540), .B(n6539), .Z(n6541) );
  XNOR U6717 ( .A(n6542), .B(n6541), .Z(n6547) );
  XOR U6718 ( .A(n6548), .B(n6547), .Z(n6522) );
  NANDN U6719 ( .A(n6499), .B(n6498), .Z(n6503) );
  NANDN U6720 ( .A(n6501), .B(n6500), .Z(n6502) );
  AND U6721 ( .A(n6503), .B(n6502), .Z(n6521) );
  XNOR U6722 ( .A(n6522), .B(n6521), .Z(n6523) );
  NANDN U6723 ( .A(n6505), .B(n6504), .Z(n6509) );
  NAND U6724 ( .A(n6507), .B(n6506), .Z(n6508) );
  NAND U6725 ( .A(n6509), .B(n6508), .Z(n6524) );
  XNOR U6726 ( .A(n6523), .B(n6524), .Z(n6515) );
  XNOR U6727 ( .A(n6516), .B(n6515), .Z(n6517) );
  XNOR U6728 ( .A(n6518), .B(n6517), .Z(n6551) );
  XNOR U6729 ( .A(sreg[410]), .B(n6551), .Z(n6553) );
  NANDN U6730 ( .A(sreg[409]), .B(n6510), .Z(n6514) );
  NAND U6731 ( .A(n6512), .B(n6511), .Z(n6513) );
  NAND U6732 ( .A(n6514), .B(n6513), .Z(n6552) );
  XNOR U6733 ( .A(n6553), .B(n6552), .Z(c[410]) );
  NANDN U6734 ( .A(n6516), .B(n6515), .Z(n6520) );
  NANDN U6735 ( .A(n6518), .B(n6517), .Z(n6519) );
  AND U6736 ( .A(n6520), .B(n6519), .Z(n6559) );
  NANDN U6737 ( .A(n6522), .B(n6521), .Z(n6526) );
  NANDN U6738 ( .A(n6524), .B(n6523), .Z(n6525) );
  AND U6739 ( .A(n6526), .B(n6525), .Z(n6557) );
  NAND U6740 ( .A(n26), .B(n6527), .Z(n6529) );
  XOR U6741 ( .A(b[7]), .B(a[157]), .Z(n6568) );
  NAND U6742 ( .A(n10531), .B(n6568), .Z(n6528) );
  AND U6743 ( .A(n6529), .B(n6528), .Z(n6587) );
  NAND U6744 ( .A(n23), .B(n6530), .Z(n6532) );
  XOR U6745 ( .A(b[3]), .B(a[161]), .Z(n6571) );
  NAND U6746 ( .A(n24), .B(n6571), .Z(n6531) );
  NAND U6747 ( .A(n6532), .B(n6531), .Z(n6586) );
  XNOR U6748 ( .A(n6587), .B(n6586), .Z(n6589) );
  NAND U6749 ( .A(b[0]), .B(a[163]), .Z(n6533) );
  XNOR U6750 ( .A(b[1]), .B(n6533), .Z(n6535) );
  NANDN U6751 ( .A(b[0]), .B(a[162]), .Z(n6534) );
  NAND U6752 ( .A(n6535), .B(n6534), .Z(n6583) );
  NAND U6753 ( .A(n25), .B(n6536), .Z(n6538) );
  XOR U6754 ( .A(b[5]), .B(a[159]), .Z(n6577) );
  NAND U6755 ( .A(n10456), .B(n6577), .Z(n6537) );
  AND U6756 ( .A(n6538), .B(n6537), .Z(n6581) );
  AND U6757 ( .A(b[7]), .B(a[155]), .Z(n6580) );
  XNOR U6758 ( .A(n6581), .B(n6580), .Z(n6582) );
  XNOR U6759 ( .A(n6583), .B(n6582), .Z(n6588) );
  XOR U6760 ( .A(n6589), .B(n6588), .Z(n6563) );
  NANDN U6761 ( .A(n6540), .B(n6539), .Z(n6544) );
  NANDN U6762 ( .A(n6542), .B(n6541), .Z(n6543) );
  AND U6763 ( .A(n6544), .B(n6543), .Z(n6562) );
  XNOR U6764 ( .A(n6563), .B(n6562), .Z(n6564) );
  NANDN U6765 ( .A(n6546), .B(n6545), .Z(n6550) );
  NAND U6766 ( .A(n6548), .B(n6547), .Z(n6549) );
  NAND U6767 ( .A(n6550), .B(n6549), .Z(n6565) );
  XNOR U6768 ( .A(n6564), .B(n6565), .Z(n6556) );
  XNOR U6769 ( .A(n6557), .B(n6556), .Z(n6558) );
  XNOR U6770 ( .A(n6559), .B(n6558), .Z(n6592) );
  XNOR U6771 ( .A(sreg[411]), .B(n6592), .Z(n6594) );
  NANDN U6772 ( .A(sreg[410]), .B(n6551), .Z(n6555) );
  NAND U6773 ( .A(n6553), .B(n6552), .Z(n6554) );
  NAND U6774 ( .A(n6555), .B(n6554), .Z(n6593) );
  XNOR U6775 ( .A(n6594), .B(n6593), .Z(c[411]) );
  NANDN U6776 ( .A(n6557), .B(n6556), .Z(n6561) );
  NANDN U6777 ( .A(n6559), .B(n6558), .Z(n6560) );
  AND U6778 ( .A(n6561), .B(n6560), .Z(n6600) );
  NANDN U6779 ( .A(n6563), .B(n6562), .Z(n6567) );
  NANDN U6780 ( .A(n6565), .B(n6564), .Z(n6566) );
  AND U6781 ( .A(n6567), .B(n6566), .Z(n6598) );
  NAND U6782 ( .A(n26), .B(n6568), .Z(n6570) );
  XOR U6783 ( .A(b[7]), .B(a[158]), .Z(n6609) );
  NAND U6784 ( .A(n10531), .B(n6609), .Z(n6569) );
  AND U6785 ( .A(n6570), .B(n6569), .Z(n6628) );
  NAND U6786 ( .A(n23), .B(n6571), .Z(n6573) );
  XOR U6787 ( .A(b[3]), .B(a[162]), .Z(n6612) );
  NAND U6788 ( .A(n24), .B(n6612), .Z(n6572) );
  NAND U6789 ( .A(n6573), .B(n6572), .Z(n6627) );
  XNOR U6790 ( .A(n6628), .B(n6627), .Z(n6630) );
  NAND U6791 ( .A(b[0]), .B(a[164]), .Z(n6574) );
  XNOR U6792 ( .A(b[1]), .B(n6574), .Z(n6576) );
  NANDN U6793 ( .A(b[0]), .B(a[163]), .Z(n6575) );
  NAND U6794 ( .A(n6576), .B(n6575), .Z(n6624) );
  NAND U6795 ( .A(n25), .B(n6577), .Z(n6579) );
  XOR U6796 ( .A(b[5]), .B(a[160]), .Z(n6618) );
  NAND U6797 ( .A(n10456), .B(n6618), .Z(n6578) );
  AND U6798 ( .A(n6579), .B(n6578), .Z(n6622) );
  AND U6799 ( .A(b[7]), .B(a[156]), .Z(n6621) );
  XNOR U6800 ( .A(n6622), .B(n6621), .Z(n6623) );
  XNOR U6801 ( .A(n6624), .B(n6623), .Z(n6629) );
  XOR U6802 ( .A(n6630), .B(n6629), .Z(n6604) );
  NANDN U6803 ( .A(n6581), .B(n6580), .Z(n6585) );
  NANDN U6804 ( .A(n6583), .B(n6582), .Z(n6584) );
  AND U6805 ( .A(n6585), .B(n6584), .Z(n6603) );
  XNOR U6806 ( .A(n6604), .B(n6603), .Z(n6605) );
  NANDN U6807 ( .A(n6587), .B(n6586), .Z(n6591) );
  NAND U6808 ( .A(n6589), .B(n6588), .Z(n6590) );
  NAND U6809 ( .A(n6591), .B(n6590), .Z(n6606) );
  XNOR U6810 ( .A(n6605), .B(n6606), .Z(n6597) );
  XNOR U6811 ( .A(n6598), .B(n6597), .Z(n6599) );
  XNOR U6812 ( .A(n6600), .B(n6599), .Z(n6633) );
  XNOR U6813 ( .A(sreg[412]), .B(n6633), .Z(n6635) );
  NANDN U6814 ( .A(sreg[411]), .B(n6592), .Z(n6596) );
  NAND U6815 ( .A(n6594), .B(n6593), .Z(n6595) );
  NAND U6816 ( .A(n6596), .B(n6595), .Z(n6634) );
  XNOR U6817 ( .A(n6635), .B(n6634), .Z(c[412]) );
  NANDN U6818 ( .A(n6598), .B(n6597), .Z(n6602) );
  NANDN U6819 ( .A(n6600), .B(n6599), .Z(n6601) );
  AND U6820 ( .A(n6602), .B(n6601), .Z(n6641) );
  NANDN U6821 ( .A(n6604), .B(n6603), .Z(n6608) );
  NANDN U6822 ( .A(n6606), .B(n6605), .Z(n6607) );
  AND U6823 ( .A(n6608), .B(n6607), .Z(n6639) );
  NAND U6824 ( .A(n26), .B(n6609), .Z(n6611) );
  XOR U6825 ( .A(b[7]), .B(a[159]), .Z(n6650) );
  NAND U6826 ( .A(n10531), .B(n6650), .Z(n6610) );
  AND U6827 ( .A(n6611), .B(n6610), .Z(n6669) );
  NAND U6828 ( .A(n23), .B(n6612), .Z(n6614) );
  XOR U6829 ( .A(b[3]), .B(a[163]), .Z(n6653) );
  NAND U6830 ( .A(n24), .B(n6653), .Z(n6613) );
  NAND U6831 ( .A(n6614), .B(n6613), .Z(n6668) );
  XNOR U6832 ( .A(n6669), .B(n6668), .Z(n6671) );
  NAND U6833 ( .A(b[0]), .B(a[165]), .Z(n6615) );
  XNOR U6834 ( .A(b[1]), .B(n6615), .Z(n6617) );
  NANDN U6835 ( .A(b[0]), .B(a[164]), .Z(n6616) );
  NAND U6836 ( .A(n6617), .B(n6616), .Z(n6665) );
  NAND U6837 ( .A(n25), .B(n6618), .Z(n6620) );
  XOR U6838 ( .A(b[5]), .B(a[161]), .Z(n6659) );
  NAND U6839 ( .A(n10456), .B(n6659), .Z(n6619) );
  AND U6840 ( .A(n6620), .B(n6619), .Z(n6663) );
  AND U6841 ( .A(b[7]), .B(a[157]), .Z(n6662) );
  XNOR U6842 ( .A(n6663), .B(n6662), .Z(n6664) );
  XNOR U6843 ( .A(n6665), .B(n6664), .Z(n6670) );
  XOR U6844 ( .A(n6671), .B(n6670), .Z(n6645) );
  NANDN U6845 ( .A(n6622), .B(n6621), .Z(n6626) );
  NANDN U6846 ( .A(n6624), .B(n6623), .Z(n6625) );
  AND U6847 ( .A(n6626), .B(n6625), .Z(n6644) );
  XNOR U6848 ( .A(n6645), .B(n6644), .Z(n6646) );
  NANDN U6849 ( .A(n6628), .B(n6627), .Z(n6632) );
  NAND U6850 ( .A(n6630), .B(n6629), .Z(n6631) );
  NAND U6851 ( .A(n6632), .B(n6631), .Z(n6647) );
  XNOR U6852 ( .A(n6646), .B(n6647), .Z(n6638) );
  XNOR U6853 ( .A(n6639), .B(n6638), .Z(n6640) );
  XNOR U6854 ( .A(n6641), .B(n6640), .Z(n6674) );
  XNOR U6855 ( .A(sreg[413]), .B(n6674), .Z(n6676) );
  NANDN U6856 ( .A(sreg[412]), .B(n6633), .Z(n6637) );
  NAND U6857 ( .A(n6635), .B(n6634), .Z(n6636) );
  NAND U6858 ( .A(n6637), .B(n6636), .Z(n6675) );
  XNOR U6859 ( .A(n6676), .B(n6675), .Z(c[413]) );
  NANDN U6860 ( .A(n6639), .B(n6638), .Z(n6643) );
  NANDN U6861 ( .A(n6641), .B(n6640), .Z(n6642) );
  AND U6862 ( .A(n6643), .B(n6642), .Z(n6682) );
  NANDN U6863 ( .A(n6645), .B(n6644), .Z(n6649) );
  NANDN U6864 ( .A(n6647), .B(n6646), .Z(n6648) );
  AND U6865 ( .A(n6649), .B(n6648), .Z(n6680) );
  NAND U6866 ( .A(n26), .B(n6650), .Z(n6652) );
  XOR U6867 ( .A(b[7]), .B(a[160]), .Z(n6691) );
  NAND U6868 ( .A(n10531), .B(n6691), .Z(n6651) );
  AND U6869 ( .A(n6652), .B(n6651), .Z(n6710) );
  NAND U6870 ( .A(n23), .B(n6653), .Z(n6655) );
  XOR U6871 ( .A(b[3]), .B(a[164]), .Z(n6694) );
  NAND U6872 ( .A(n24), .B(n6694), .Z(n6654) );
  NAND U6873 ( .A(n6655), .B(n6654), .Z(n6709) );
  XNOR U6874 ( .A(n6710), .B(n6709), .Z(n6712) );
  AND U6875 ( .A(b[0]), .B(a[166]), .Z(n6656) );
  XOR U6876 ( .A(b[1]), .B(n6656), .Z(n6658) );
  NANDN U6877 ( .A(b[0]), .B(a[165]), .Z(n6657) );
  AND U6878 ( .A(n6658), .B(n6657), .Z(n6705) );
  NAND U6879 ( .A(n25), .B(n6659), .Z(n6661) );
  XOR U6880 ( .A(b[5]), .B(a[162]), .Z(n6700) );
  NAND U6881 ( .A(n10456), .B(n6700), .Z(n6660) );
  AND U6882 ( .A(n6661), .B(n6660), .Z(n6704) );
  AND U6883 ( .A(b[7]), .B(a[158]), .Z(n6703) );
  XOR U6884 ( .A(n6704), .B(n6703), .Z(n6706) );
  XNOR U6885 ( .A(n6705), .B(n6706), .Z(n6711) );
  XOR U6886 ( .A(n6712), .B(n6711), .Z(n6686) );
  NANDN U6887 ( .A(n6663), .B(n6662), .Z(n6667) );
  NANDN U6888 ( .A(n6665), .B(n6664), .Z(n6666) );
  AND U6889 ( .A(n6667), .B(n6666), .Z(n6685) );
  XNOR U6890 ( .A(n6686), .B(n6685), .Z(n6687) );
  NANDN U6891 ( .A(n6669), .B(n6668), .Z(n6673) );
  NAND U6892 ( .A(n6671), .B(n6670), .Z(n6672) );
  NAND U6893 ( .A(n6673), .B(n6672), .Z(n6688) );
  XNOR U6894 ( .A(n6687), .B(n6688), .Z(n6679) );
  XNOR U6895 ( .A(n6680), .B(n6679), .Z(n6681) );
  XNOR U6896 ( .A(n6682), .B(n6681), .Z(n6715) );
  XNOR U6897 ( .A(sreg[414]), .B(n6715), .Z(n6717) );
  NANDN U6898 ( .A(sreg[413]), .B(n6674), .Z(n6678) );
  NAND U6899 ( .A(n6676), .B(n6675), .Z(n6677) );
  NAND U6900 ( .A(n6678), .B(n6677), .Z(n6716) );
  XNOR U6901 ( .A(n6717), .B(n6716), .Z(c[414]) );
  NANDN U6902 ( .A(n6680), .B(n6679), .Z(n6684) );
  NANDN U6903 ( .A(n6682), .B(n6681), .Z(n6683) );
  AND U6904 ( .A(n6684), .B(n6683), .Z(n6723) );
  NANDN U6905 ( .A(n6686), .B(n6685), .Z(n6690) );
  NANDN U6906 ( .A(n6688), .B(n6687), .Z(n6689) );
  AND U6907 ( .A(n6690), .B(n6689), .Z(n6721) );
  NAND U6908 ( .A(n26), .B(n6691), .Z(n6693) );
  XOR U6909 ( .A(b[7]), .B(a[161]), .Z(n6732) );
  NAND U6910 ( .A(n10531), .B(n6732), .Z(n6692) );
  AND U6911 ( .A(n6693), .B(n6692), .Z(n6751) );
  NAND U6912 ( .A(n23), .B(n6694), .Z(n6696) );
  XOR U6913 ( .A(b[3]), .B(a[165]), .Z(n6735) );
  NAND U6914 ( .A(n24), .B(n6735), .Z(n6695) );
  NAND U6915 ( .A(n6696), .B(n6695), .Z(n6750) );
  XNOR U6916 ( .A(n6751), .B(n6750), .Z(n6753) );
  NAND U6917 ( .A(b[0]), .B(a[167]), .Z(n6697) );
  XNOR U6918 ( .A(b[1]), .B(n6697), .Z(n6699) );
  NANDN U6919 ( .A(b[0]), .B(a[166]), .Z(n6698) );
  NAND U6920 ( .A(n6699), .B(n6698), .Z(n6747) );
  NAND U6921 ( .A(n25), .B(n6700), .Z(n6702) );
  XOR U6922 ( .A(b[5]), .B(a[163]), .Z(n6738) );
  NAND U6923 ( .A(n10456), .B(n6738), .Z(n6701) );
  AND U6924 ( .A(n6702), .B(n6701), .Z(n6745) );
  AND U6925 ( .A(b[7]), .B(a[159]), .Z(n6744) );
  XNOR U6926 ( .A(n6745), .B(n6744), .Z(n6746) );
  XNOR U6927 ( .A(n6747), .B(n6746), .Z(n6752) );
  XOR U6928 ( .A(n6753), .B(n6752), .Z(n6727) );
  NANDN U6929 ( .A(n6704), .B(n6703), .Z(n6708) );
  NANDN U6930 ( .A(n6706), .B(n6705), .Z(n6707) );
  AND U6931 ( .A(n6708), .B(n6707), .Z(n6726) );
  XNOR U6932 ( .A(n6727), .B(n6726), .Z(n6728) );
  NANDN U6933 ( .A(n6710), .B(n6709), .Z(n6714) );
  NAND U6934 ( .A(n6712), .B(n6711), .Z(n6713) );
  NAND U6935 ( .A(n6714), .B(n6713), .Z(n6729) );
  XNOR U6936 ( .A(n6728), .B(n6729), .Z(n6720) );
  XNOR U6937 ( .A(n6721), .B(n6720), .Z(n6722) );
  XNOR U6938 ( .A(n6723), .B(n6722), .Z(n6756) );
  XNOR U6939 ( .A(sreg[415]), .B(n6756), .Z(n6758) );
  NANDN U6940 ( .A(sreg[414]), .B(n6715), .Z(n6719) );
  NAND U6941 ( .A(n6717), .B(n6716), .Z(n6718) );
  NAND U6942 ( .A(n6719), .B(n6718), .Z(n6757) );
  XNOR U6943 ( .A(n6758), .B(n6757), .Z(c[415]) );
  NANDN U6944 ( .A(n6721), .B(n6720), .Z(n6725) );
  NANDN U6945 ( .A(n6723), .B(n6722), .Z(n6724) );
  AND U6946 ( .A(n6725), .B(n6724), .Z(n6764) );
  NANDN U6947 ( .A(n6727), .B(n6726), .Z(n6731) );
  NANDN U6948 ( .A(n6729), .B(n6728), .Z(n6730) );
  AND U6949 ( .A(n6731), .B(n6730), .Z(n6762) );
  NAND U6950 ( .A(n26), .B(n6732), .Z(n6734) );
  XOR U6951 ( .A(b[7]), .B(a[162]), .Z(n6773) );
  NAND U6952 ( .A(n10531), .B(n6773), .Z(n6733) );
  AND U6953 ( .A(n6734), .B(n6733), .Z(n6792) );
  NAND U6954 ( .A(n23), .B(n6735), .Z(n6737) );
  XOR U6955 ( .A(b[3]), .B(a[166]), .Z(n6776) );
  NAND U6956 ( .A(n24), .B(n6776), .Z(n6736) );
  NAND U6957 ( .A(n6737), .B(n6736), .Z(n6791) );
  XNOR U6958 ( .A(n6792), .B(n6791), .Z(n6794) );
  NAND U6959 ( .A(n25), .B(n6738), .Z(n6740) );
  XOR U6960 ( .A(b[5]), .B(a[164]), .Z(n6782) );
  NAND U6961 ( .A(n10456), .B(n6782), .Z(n6739) );
  AND U6962 ( .A(n6740), .B(n6739), .Z(n6786) );
  AND U6963 ( .A(b[7]), .B(a[160]), .Z(n6785) );
  XNOR U6964 ( .A(n6786), .B(n6785), .Z(n6787) );
  NAND U6965 ( .A(b[0]), .B(a[168]), .Z(n6741) );
  XNOR U6966 ( .A(b[1]), .B(n6741), .Z(n6743) );
  NANDN U6967 ( .A(b[0]), .B(a[167]), .Z(n6742) );
  NAND U6968 ( .A(n6743), .B(n6742), .Z(n6788) );
  XNOR U6969 ( .A(n6787), .B(n6788), .Z(n6793) );
  XOR U6970 ( .A(n6794), .B(n6793), .Z(n6768) );
  NANDN U6971 ( .A(n6745), .B(n6744), .Z(n6749) );
  NANDN U6972 ( .A(n6747), .B(n6746), .Z(n6748) );
  AND U6973 ( .A(n6749), .B(n6748), .Z(n6767) );
  XNOR U6974 ( .A(n6768), .B(n6767), .Z(n6769) );
  NANDN U6975 ( .A(n6751), .B(n6750), .Z(n6755) );
  NAND U6976 ( .A(n6753), .B(n6752), .Z(n6754) );
  NAND U6977 ( .A(n6755), .B(n6754), .Z(n6770) );
  XNOR U6978 ( .A(n6769), .B(n6770), .Z(n6761) );
  XNOR U6979 ( .A(n6762), .B(n6761), .Z(n6763) );
  XNOR U6980 ( .A(n6764), .B(n6763), .Z(n6797) );
  XNOR U6981 ( .A(sreg[416]), .B(n6797), .Z(n6799) );
  NANDN U6982 ( .A(sreg[415]), .B(n6756), .Z(n6760) );
  NAND U6983 ( .A(n6758), .B(n6757), .Z(n6759) );
  NAND U6984 ( .A(n6760), .B(n6759), .Z(n6798) );
  XNOR U6985 ( .A(n6799), .B(n6798), .Z(c[416]) );
  NANDN U6986 ( .A(n6762), .B(n6761), .Z(n6766) );
  NANDN U6987 ( .A(n6764), .B(n6763), .Z(n6765) );
  AND U6988 ( .A(n6766), .B(n6765), .Z(n6805) );
  NANDN U6989 ( .A(n6768), .B(n6767), .Z(n6772) );
  NANDN U6990 ( .A(n6770), .B(n6769), .Z(n6771) );
  AND U6991 ( .A(n6772), .B(n6771), .Z(n6803) );
  NAND U6992 ( .A(n26), .B(n6773), .Z(n6775) );
  XOR U6993 ( .A(b[7]), .B(a[163]), .Z(n6814) );
  NAND U6994 ( .A(n10531), .B(n6814), .Z(n6774) );
  AND U6995 ( .A(n6775), .B(n6774), .Z(n6833) );
  NAND U6996 ( .A(n23), .B(n6776), .Z(n6778) );
  XOR U6997 ( .A(b[3]), .B(a[167]), .Z(n6817) );
  NAND U6998 ( .A(n24), .B(n6817), .Z(n6777) );
  NAND U6999 ( .A(n6778), .B(n6777), .Z(n6832) );
  XNOR U7000 ( .A(n6833), .B(n6832), .Z(n6835) );
  NAND U7001 ( .A(b[0]), .B(a[169]), .Z(n6779) );
  XNOR U7002 ( .A(b[1]), .B(n6779), .Z(n6781) );
  NANDN U7003 ( .A(b[0]), .B(a[168]), .Z(n6780) );
  NAND U7004 ( .A(n6781), .B(n6780), .Z(n6829) );
  NAND U7005 ( .A(n25), .B(n6782), .Z(n6784) );
  XOR U7006 ( .A(b[5]), .B(a[165]), .Z(n6820) );
  NAND U7007 ( .A(n10456), .B(n6820), .Z(n6783) );
  AND U7008 ( .A(n6784), .B(n6783), .Z(n6827) );
  AND U7009 ( .A(b[7]), .B(a[161]), .Z(n6826) );
  XNOR U7010 ( .A(n6827), .B(n6826), .Z(n6828) );
  XNOR U7011 ( .A(n6829), .B(n6828), .Z(n6834) );
  XOR U7012 ( .A(n6835), .B(n6834), .Z(n6809) );
  NANDN U7013 ( .A(n6786), .B(n6785), .Z(n6790) );
  NANDN U7014 ( .A(n6788), .B(n6787), .Z(n6789) );
  AND U7015 ( .A(n6790), .B(n6789), .Z(n6808) );
  XNOR U7016 ( .A(n6809), .B(n6808), .Z(n6810) );
  NANDN U7017 ( .A(n6792), .B(n6791), .Z(n6796) );
  NAND U7018 ( .A(n6794), .B(n6793), .Z(n6795) );
  NAND U7019 ( .A(n6796), .B(n6795), .Z(n6811) );
  XNOR U7020 ( .A(n6810), .B(n6811), .Z(n6802) );
  XNOR U7021 ( .A(n6803), .B(n6802), .Z(n6804) );
  XNOR U7022 ( .A(n6805), .B(n6804), .Z(n6838) );
  XNOR U7023 ( .A(sreg[417]), .B(n6838), .Z(n6840) );
  NANDN U7024 ( .A(sreg[416]), .B(n6797), .Z(n6801) );
  NAND U7025 ( .A(n6799), .B(n6798), .Z(n6800) );
  NAND U7026 ( .A(n6801), .B(n6800), .Z(n6839) );
  XNOR U7027 ( .A(n6840), .B(n6839), .Z(c[417]) );
  NANDN U7028 ( .A(n6803), .B(n6802), .Z(n6807) );
  NANDN U7029 ( .A(n6805), .B(n6804), .Z(n6806) );
  AND U7030 ( .A(n6807), .B(n6806), .Z(n6846) );
  NANDN U7031 ( .A(n6809), .B(n6808), .Z(n6813) );
  NANDN U7032 ( .A(n6811), .B(n6810), .Z(n6812) );
  AND U7033 ( .A(n6813), .B(n6812), .Z(n6844) );
  NAND U7034 ( .A(n26), .B(n6814), .Z(n6816) );
  XOR U7035 ( .A(b[7]), .B(a[164]), .Z(n6855) );
  NAND U7036 ( .A(n10531), .B(n6855), .Z(n6815) );
  AND U7037 ( .A(n6816), .B(n6815), .Z(n6874) );
  NAND U7038 ( .A(n23), .B(n6817), .Z(n6819) );
  XOR U7039 ( .A(b[3]), .B(a[168]), .Z(n6858) );
  NAND U7040 ( .A(n24), .B(n6858), .Z(n6818) );
  NAND U7041 ( .A(n6819), .B(n6818), .Z(n6873) );
  XNOR U7042 ( .A(n6874), .B(n6873), .Z(n6876) );
  NAND U7043 ( .A(n25), .B(n6820), .Z(n6822) );
  XOR U7044 ( .A(b[5]), .B(a[166]), .Z(n6864) );
  NAND U7045 ( .A(n10456), .B(n6864), .Z(n6821) );
  AND U7046 ( .A(n6822), .B(n6821), .Z(n6868) );
  AND U7047 ( .A(b[7]), .B(a[162]), .Z(n6867) );
  XNOR U7048 ( .A(n6868), .B(n6867), .Z(n6869) );
  NAND U7049 ( .A(b[0]), .B(a[170]), .Z(n6823) );
  XNOR U7050 ( .A(b[1]), .B(n6823), .Z(n6825) );
  NANDN U7051 ( .A(b[0]), .B(a[169]), .Z(n6824) );
  NAND U7052 ( .A(n6825), .B(n6824), .Z(n6870) );
  XNOR U7053 ( .A(n6869), .B(n6870), .Z(n6875) );
  XOR U7054 ( .A(n6876), .B(n6875), .Z(n6850) );
  NANDN U7055 ( .A(n6827), .B(n6826), .Z(n6831) );
  NANDN U7056 ( .A(n6829), .B(n6828), .Z(n6830) );
  AND U7057 ( .A(n6831), .B(n6830), .Z(n6849) );
  XNOR U7058 ( .A(n6850), .B(n6849), .Z(n6851) );
  NANDN U7059 ( .A(n6833), .B(n6832), .Z(n6837) );
  NAND U7060 ( .A(n6835), .B(n6834), .Z(n6836) );
  NAND U7061 ( .A(n6837), .B(n6836), .Z(n6852) );
  XNOR U7062 ( .A(n6851), .B(n6852), .Z(n6843) );
  XNOR U7063 ( .A(n6844), .B(n6843), .Z(n6845) );
  XNOR U7064 ( .A(n6846), .B(n6845), .Z(n6879) );
  XNOR U7065 ( .A(sreg[418]), .B(n6879), .Z(n6881) );
  NANDN U7066 ( .A(sreg[417]), .B(n6838), .Z(n6842) );
  NAND U7067 ( .A(n6840), .B(n6839), .Z(n6841) );
  NAND U7068 ( .A(n6842), .B(n6841), .Z(n6880) );
  XNOR U7069 ( .A(n6881), .B(n6880), .Z(c[418]) );
  NANDN U7070 ( .A(n6844), .B(n6843), .Z(n6848) );
  NANDN U7071 ( .A(n6846), .B(n6845), .Z(n6847) );
  AND U7072 ( .A(n6848), .B(n6847), .Z(n6887) );
  NANDN U7073 ( .A(n6850), .B(n6849), .Z(n6854) );
  NANDN U7074 ( .A(n6852), .B(n6851), .Z(n6853) );
  AND U7075 ( .A(n6854), .B(n6853), .Z(n6885) );
  NAND U7076 ( .A(n26), .B(n6855), .Z(n6857) );
  XOR U7077 ( .A(b[7]), .B(a[165]), .Z(n6896) );
  NAND U7078 ( .A(n10531), .B(n6896), .Z(n6856) );
  AND U7079 ( .A(n6857), .B(n6856), .Z(n6915) );
  NAND U7080 ( .A(n23), .B(n6858), .Z(n6860) );
  XOR U7081 ( .A(b[3]), .B(a[169]), .Z(n6899) );
  NAND U7082 ( .A(n24), .B(n6899), .Z(n6859) );
  NAND U7083 ( .A(n6860), .B(n6859), .Z(n6914) );
  XNOR U7084 ( .A(n6915), .B(n6914), .Z(n6917) );
  NAND U7085 ( .A(b[0]), .B(a[171]), .Z(n6861) );
  XNOR U7086 ( .A(b[1]), .B(n6861), .Z(n6863) );
  NANDN U7087 ( .A(b[0]), .B(a[170]), .Z(n6862) );
  NAND U7088 ( .A(n6863), .B(n6862), .Z(n6911) );
  NAND U7089 ( .A(n25), .B(n6864), .Z(n6866) );
  XOR U7090 ( .A(b[5]), .B(a[167]), .Z(n6905) );
  NAND U7091 ( .A(n10456), .B(n6905), .Z(n6865) );
  AND U7092 ( .A(n6866), .B(n6865), .Z(n6909) );
  AND U7093 ( .A(b[7]), .B(a[163]), .Z(n6908) );
  XNOR U7094 ( .A(n6909), .B(n6908), .Z(n6910) );
  XNOR U7095 ( .A(n6911), .B(n6910), .Z(n6916) );
  XOR U7096 ( .A(n6917), .B(n6916), .Z(n6891) );
  NANDN U7097 ( .A(n6868), .B(n6867), .Z(n6872) );
  NANDN U7098 ( .A(n6870), .B(n6869), .Z(n6871) );
  AND U7099 ( .A(n6872), .B(n6871), .Z(n6890) );
  XNOR U7100 ( .A(n6891), .B(n6890), .Z(n6892) );
  NANDN U7101 ( .A(n6874), .B(n6873), .Z(n6878) );
  NAND U7102 ( .A(n6876), .B(n6875), .Z(n6877) );
  NAND U7103 ( .A(n6878), .B(n6877), .Z(n6893) );
  XNOR U7104 ( .A(n6892), .B(n6893), .Z(n6884) );
  XNOR U7105 ( .A(n6885), .B(n6884), .Z(n6886) );
  XNOR U7106 ( .A(n6887), .B(n6886), .Z(n6920) );
  XNOR U7107 ( .A(sreg[419]), .B(n6920), .Z(n6922) );
  NANDN U7108 ( .A(sreg[418]), .B(n6879), .Z(n6883) );
  NAND U7109 ( .A(n6881), .B(n6880), .Z(n6882) );
  NAND U7110 ( .A(n6883), .B(n6882), .Z(n6921) );
  XNOR U7111 ( .A(n6922), .B(n6921), .Z(c[419]) );
  NANDN U7112 ( .A(n6885), .B(n6884), .Z(n6889) );
  NANDN U7113 ( .A(n6887), .B(n6886), .Z(n6888) );
  AND U7114 ( .A(n6889), .B(n6888), .Z(n6928) );
  NANDN U7115 ( .A(n6891), .B(n6890), .Z(n6895) );
  NANDN U7116 ( .A(n6893), .B(n6892), .Z(n6894) );
  AND U7117 ( .A(n6895), .B(n6894), .Z(n6926) );
  NAND U7118 ( .A(n26), .B(n6896), .Z(n6898) );
  XOR U7119 ( .A(b[7]), .B(a[166]), .Z(n6937) );
  NAND U7120 ( .A(n10531), .B(n6937), .Z(n6897) );
  AND U7121 ( .A(n6898), .B(n6897), .Z(n6956) );
  NAND U7122 ( .A(n23), .B(n6899), .Z(n6901) );
  XOR U7123 ( .A(b[3]), .B(a[170]), .Z(n6940) );
  NAND U7124 ( .A(n24), .B(n6940), .Z(n6900) );
  NAND U7125 ( .A(n6901), .B(n6900), .Z(n6955) );
  XNOR U7126 ( .A(n6956), .B(n6955), .Z(n6958) );
  NAND U7127 ( .A(b[0]), .B(a[172]), .Z(n6902) );
  XNOR U7128 ( .A(b[1]), .B(n6902), .Z(n6904) );
  NANDN U7129 ( .A(b[0]), .B(a[171]), .Z(n6903) );
  NAND U7130 ( .A(n6904), .B(n6903), .Z(n6952) );
  NAND U7131 ( .A(n25), .B(n6905), .Z(n6907) );
  XOR U7132 ( .A(b[5]), .B(a[168]), .Z(n6946) );
  NAND U7133 ( .A(n10456), .B(n6946), .Z(n6906) );
  AND U7134 ( .A(n6907), .B(n6906), .Z(n6950) );
  AND U7135 ( .A(b[7]), .B(a[164]), .Z(n6949) );
  XNOR U7136 ( .A(n6950), .B(n6949), .Z(n6951) );
  XNOR U7137 ( .A(n6952), .B(n6951), .Z(n6957) );
  XOR U7138 ( .A(n6958), .B(n6957), .Z(n6932) );
  NANDN U7139 ( .A(n6909), .B(n6908), .Z(n6913) );
  NANDN U7140 ( .A(n6911), .B(n6910), .Z(n6912) );
  AND U7141 ( .A(n6913), .B(n6912), .Z(n6931) );
  XNOR U7142 ( .A(n6932), .B(n6931), .Z(n6933) );
  NANDN U7143 ( .A(n6915), .B(n6914), .Z(n6919) );
  NAND U7144 ( .A(n6917), .B(n6916), .Z(n6918) );
  NAND U7145 ( .A(n6919), .B(n6918), .Z(n6934) );
  XNOR U7146 ( .A(n6933), .B(n6934), .Z(n6925) );
  XNOR U7147 ( .A(n6926), .B(n6925), .Z(n6927) );
  XNOR U7148 ( .A(n6928), .B(n6927), .Z(n6961) );
  XNOR U7149 ( .A(sreg[420]), .B(n6961), .Z(n6963) );
  NANDN U7150 ( .A(sreg[419]), .B(n6920), .Z(n6924) );
  NAND U7151 ( .A(n6922), .B(n6921), .Z(n6923) );
  NAND U7152 ( .A(n6924), .B(n6923), .Z(n6962) );
  XNOR U7153 ( .A(n6963), .B(n6962), .Z(c[420]) );
  NANDN U7154 ( .A(n6926), .B(n6925), .Z(n6930) );
  NANDN U7155 ( .A(n6928), .B(n6927), .Z(n6929) );
  AND U7156 ( .A(n6930), .B(n6929), .Z(n6969) );
  NANDN U7157 ( .A(n6932), .B(n6931), .Z(n6936) );
  NANDN U7158 ( .A(n6934), .B(n6933), .Z(n6935) );
  AND U7159 ( .A(n6936), .B(n6935), .Z(n6967) );
  NAND U7160 ( .A(n26), .B(n6937), .Z(n6939) );
  XOR U7161 ( .A(b[7]), .B(a[167]), .Z(n6978) );
  NAND U7162 ( .A(n10531), .B(n6978), .Z(n6938) );
  AND U7163 ( .A(n6939), .B(n6938), .Z(n6997) );
  NAND U7164 ( .A(n23), .B(n6940), .Z(n6942) );
  XOR U7165 ( .A(b[3]), .B(a[171]), .Z(n6981) );
  NAND U7166 ( .A(n24), .B(n6981), .Z(n6941) );
  NAND U7167 ( .A(n6942), .B(n6941), .Z(n6996) );
  XNOR U7168 ( .A(n6997), .B(n6996), .Z(n6999) );
  NAND U7169 ( .A(b[0]), .B(a[173]), .Z(n6943) );
  XNOR U7170 ( .A(b[1]), .B(n6943), .Z(n6945) );
  NANDN U7171 ( .A(b[0]), .B(a[172]), .Z(n6944) );
  NAND U7172 ( .A(n6945), .B(n6944), .Z(n6993) );
  NAND U7173 ( .A(n25), .B(n6946), .Z(n6948) );
  XOR U7174 ( .A(b[5]), .B(a[169]), .Z(n6987) );
  NAND U7175 ( .A(n10456), .B(n6987), .Z(n6947) );
  AND U7176 ( .A(n6948), .B(n6947), .Z(n6991) );
  AND U7177 ( .A(b[7]), .B(a[165]), .Z(n6990) );
  XNOR U7178 ( .A(n6991), .B(n6990), .Z(n6992) );
  XNOR U7179 ( .A(n6993), .B(n6992), .Z(n6998) );
  XOR U7180 ( .A(n6999), .B(n6998), .Z(n6973) );
  NANDN U7181 ( .A(n6950), .B(n6949), .Z(n6954) );
  NANDN U7182 ( .A(n6952), .B(n6951), .Z(n6953) );
  AND U7183 ( .A(n6954), .B(n6953), .Z(n6972) );
  XNOR U7184 ( .A(n6973), .B(n6972), .Z(n6974) );
  NANDN U7185 ( .A(n6956), .B(n6955), .Z(n6960) );
  NAND U7186 ( .A(n6958), .B(n6957), .Z(n6959) );
  NAND U7187 ( .A(n6960), .B(n6959), .Z(n6975) );
  XNOR U7188 ( .A(n6974), .B(n6975), .Z(n6966) );
  XNOR U7189 ( .A(n6967), .B(n6966), .Z(n6968) );
  XNOR U7190 ( .A(n6969), .B(n6968), .Z(n7002) );
  XNOR U7191 ( .A(sreg[421]), .B(n7002), .Z(n7004) );
  NANDN U7192 ( .A(sreg[420]), .B(n6961), .Z(n6965) );
  NAND U7193 ( .A(n6963), .B(n6962), .Z(n6964) );
  NAND U7194 ( .A(n6965), .B(n6964), .Z(n7003) );
  XNOR U7195 ( .A(n7004), .B(n7003), .Z(c[421]) );
  NANDN U7196 ( .A(n6967), .B(n6966), .Z(n6971) );
  NANDN U7197 ( .A(n6969), .B(n6968), .Z(n6970) );
  AND U7198 ( .A(n6971), .B(n6970), .Z(n7010) );
  NANDN U7199 ( .A(n6973), .B(n6972), .Z(n6977) );
  NANDN U7200 ( .A(n6975), .B(n6974), .Z(n6976) );
  AND U7201 ( .A(n6977), .B(n6976), .Z(n7008) );
  NAND U7202 ( .A(n26), .B(n6978), .Z(n6980) );
  XOR U7203 ( .A(b[7]), .B(a[168]), .Z(n7019) );
  NAND U7204 ( .A(n10531), .B(n7019), .Z(n6979) );
  AND U7205 ( .A(n6980), .B(n6979), .Z(n7038) );
  NAND U7206 ( .A(n23), .B(n6981), .Z(n6983) );
  XOR U7207 ( .A(b[3]), .B(a[172]), .Z(n7022) );
  NAND U7208 ( .A(n24), .B(n7022), .Z(n6982) );
  NAND U7209 ( .A(n6983), .B(n6982), .Z(n7037) );
  XNOR U7210 ( .A(n7038), .B(n7037), .Z(n7040) );
  NAND U7211 ( .A(b[0]), .B(a[174]), .Z(n6984) );
  XNOR U7212 ( .A(b[1]), .B(n6984), .Z(n6986) );
  NANDN U7213 ( .A(b[0]), .B(a[173]), .Z(n6985) );
  NAND U7214 ( .A(n6986), .B(n6985), .Z(n7034) );
  NAND U7215 ( .A(n25), .B(n6987), .Z(n6989) );
  XOR U7216 ( .A(b[5]), .B(a[170]), .Z(n7028) );
  NAND U7217 ( .A(n10456), .B(n7028), .Z(n6988) );
  AND U7218 ( .A(n6989), .B(n6988), .Z(n7032) );
  AND U7219 ( .A(b[7]), .B(a[166]), .Z(n7031) );
  XNOR U7220 ( .A(n7032), .B(n7031), .Z(n7033) );
  XNOR U7221 ( .A(n7034), .B(n7033), .Z(n7039) );
  XOR U7222 ( .A(n7040), .B(n7039), .Z(n7014) );
  NANDN U7223 ( .A(n6991), .B(n6990), .Z(n6995) );
  NANDN U7224 ( .A(n6993), .B(n6992), .Z(n6994) );
  AND U7225 ( .A(n6995), .B(n6994), .Z(n7013) );
  XNOR U7226 ( .A(n7014), .B(n7013), .Z(n7015) );
  NANDN U7227 ( .A(n6997), .B(n6996), .Z(n7001) );
  NAND U7228 ( .A(n6999), .B(n6998), .Z(n7000) );
  NAND U7229 ( .A(n7001), .B(n7000), .Z(n7016) );
  XNOR U7230 ( .A(n7015), .B(n7016), .Z(n7007) );
  XNOR U7231 ( .A(n7008), .B(n7007), .Z(n7009) );
  XNOR U7232 ( .A(n7010), .B(n7009), .Z(n7043) );
  XNOR U7233 ( .A(sreg[422]), .B(n7043), .Z(n7045) );
  NANDN U7234 ( .A(sreg[421]), .B(n7002), .Z(n7006) );
  NAND U7235 ( .A(n7004), .B(n7003), .Z(n7005) );
  NAND U7236 ( .A(n7006), .B(n7005), .Z(n7044) );
  XNOR U7237 ( .A(n7045), .B(n7044), .Z(c[422]) );
  NANDN U7238 ( .A(n7008), .B(n7007), .Z(n7012) );
  NANDN U7239 ( .A(n7010), .B(n7009), .Z(n7011) );
  AND U7240 ( .A(n7012), .B(n7011), .Z(n7051) );
  NANDN U7241 ( .A(n7014), .B(n7013), .Z(n7018) );
  NANDN U7242 ( .A(n7016), .B(n7015), .Z(n7017) );
  AND U7243 ( .A(n7018), .B(n7017), .Z(n7049) );
  NAND U7244 ( .A(n26), .B(n7019), .Z(n7021) );
  XOR U7245 ( .A(b[7]), .B(a[169]), .Z(n7060) );
  NAND U7246 ( .A(n10531), .B(n7060), .Z(n7020) );
  AND U7247 ( .A(n7021), .B(n7020), .Z(n7079) );
  NAND U7248 ( .A(n23), .B(n7022), .Z(n7024) );
  XOR U7249 ( .A(b[3]), .B(a[173]), .Z(n7063) );
  NAND U7250 ( .A(n24), .B(n7063), .Z(n7023) );
  NAND U7251 ( .A(n7024), .B(n7023), .Z(n7078) );
  XNOR U7252 ( .A(n7079), .B(n7078), .Z(n7081) );
  NAND U7253 ( .A(b[0]), .B(a[175]), .Z(n7025) );
  XNOR U7254 ( .A(b[1]), .B(n7025), .Z(n7027) );
  NANDN U7255 ( .A(b[0]), .B(a[174]), .Z(n7026) );
  NAND U7256 ( .A(n7027), .B(n7026), .Z(n7075) );
  NAND U7257 ( .A(n25), .B(n7028), .Z(n7030) );
  XOR U7258 ( .A(b[5]), .B(a[171]), .Z(n7069) );
  NAND U7259 ( .A(n10456), .B(n7069), .Z(n7029) );
  AND U7260 ( .A(n7030), .B(n7029), .Z(n7073) );
  AND U7261 ( .A(b[7]), .B(a[167]), .Z(n7072) );
  XNOR U7262 ( .A(n7073), .B(n7072), .Z(n7074) );
  XNOR U7263 ( .A(n7075), .B(n7074), .Z(n7080) );
  XOR U7264 ( .A(n7081), .B(n7080), .Z(n7055) );
  NANDN U7265 ( .A(n7032), .B(n7031), .Z(n7036) );
  NANDN U7266 ( .A(n7034), .B(n7033), .Z(n7035) );
  AND U7267 ( .A(n7036), .B(n7035), .Z(n7054) );
  XNOR U7268 ( .A(n7055), .B(n7054), .Z(n7056) );
  NANDN U7269 ( .A(n7038), .B(n7037), .Z(n7042) );
  NAND U7270 ( .A(n7040), .B(n7039), .Z(n7041) );
  NAND U7271 ( .A(n7042), .B(n7041), .Z(n7057) );
  XNOR U7272 ( .A(n7056), .B(n7057), .Z(n7048) );
  XNOR U7273 ( .A(n7049), .B(n7048), .Z(n7050) );
  XNOR U7274 ( .A(n7051), .B(n7050), .Z(n7084) );
  XNOR U7275 ( .A(sreg[423]), .B(n7084), .Z(n7086) );
  NANDN U7276 ( .A(sreg[422]), .B(n7043), .Z(n7047) );
  NAND U7277 ( .A(n7045), .B(n7044), .Z(n7046) );
  NAND U7278 ( .A(n7047), .B(n7046), .Z(n7085) );
  XNOR U7279 ( .A(n7086), .B(n7085), .Z(c[423]) );
  NANDN U7280 ( .A(n7049), .B(n7048), .Z(n7053) );
  NANDN U7281 ( .A(n7051), .B(n7050), .Z(n7052) );
  AND U7282 ( .A(n7053), .B(n7052), .Z(n7092) );
  NANDN U7283 ( .A(n7055), .B(n7054), .Z(n7059) );
  NANDN U7284 ( .A(n7057), .B(n7056), .Z(n7058) );
  AND U7285 ( .A(n7059), .B(n7058), .Z(n7090) );
  NAND U7286 ( .A(n26), .B(n7060), .Z(n7062) );
  XOR U7287 ( .A(b[7]), .B(a[170]), .Z(n7101) );
  NAND U7288 ( .A(n10531), .B(n7101), .Z(n7061) );
  AND U7289 ( .A(n7062), .B(n7061), .Z(n7120) );
  NAND U7290 ( .A(n23), .B(n7063), .Z(n7065) );
  XOR U7291 ( .A(b[3]), .B(a[174]), .Z(n7104) );
  NAND U7292 ( .A(n24), .B(n7104), .Z(n7064) );
  NAND U7293 ( .A(n7065), .B(n7064), .Z(n7119) );
  XNOR U7294 ( .A(n7120), .B(n7119), .Z(n7122) );
  NAND U7295 ( .A(b[0]), .B(a[176]), .Z(n7066) );
  XNOR U7296 ( .A(b[1]), .B(n7066), .Z(n7068) );
  NANDN U7297 ( .A(b[0]), .B(a[175]), .Z(n7067) );
  NAND U7298 ( .A(n7068), .B(n7067), .Z(n7116) );
  NAND U7299 ( .A(n25), .B(n7069), .Z(n7071) );
  XOR U7300 ( .A(b[5]), .B(a[172]), .Z(n7110) );
  NAND U7301 ( .A(n10456), .B(n7110), .Z(n7070) );
  AND U7302 ( .A(n7071), .B(n7070), .Z(n7114) );
  AND U7303 ( .A(b[7]), .B(a[168]), .Z(n7113) );
  XNOR U7304 ( .A(n7114), .B(n7113), .Z(n7115) );
  XNOR U7305 ( .A(n7116), .B(n7115), .Z(n7121) );
  XOR U7306 ( .A(n7122), .B(n7121), .Z(n7096) );
  NANDN U7307 ( .A(n7073), .B(n7072), .Z(n7077) );
  NANDN U7308 ( .A(n7075), .B(n7074), .Z(n7076) );
  AND U7309 ( .A(n7077), .B(n7076), .Z(n7095) );
  XNOR U7310 ( .A(n7096), .B(n7095), .Z(n7097) );
  NANDN U7311 ( .A(n7079), .B(n7078), .Z(n7083) );
  NAND U7312 ( .A(n7081), .B(n7080), .Z(n7082) );
  NAND U7313 ( .A(n7083), .B(n7082), .Z(n7098) );
  XNOR U7314 ( .A(n7097), .B(n7098), .Z(n7089) );
  XNOR U7315 ( .A(n7090), .B(n7089), .Z(n7091) );
  XNOR U7316 ( .A(n7092), .B(n7091), .Z(n7125) );
  XNOR U7317 ( .A(sreg[424]), .B(n7125), .Z(n7127) );
  NANDN U7318 ( .A(sreg[423]), .B(n7084), .Z(n7088) );
  NAND U7319 ( .A(n7086), .B(n7085), .Z(n7087) );
  NAND U7320 ( .A(n7088), .B(n7087), .Z(n7126) );
  XNOR U7321 ( .A(n7127), .B(n7126), .Z(c[424]) );
  NANDN U7322 ( .A(n7090), .B(n7089), .Z(n7094) );
  NANDN U7323 ( .A(n7092), .B(n7091), .Z(n7093) );
  AND U7324 ( .A(n7094), .B(n7093), .Z(n7133) );
  NANDN U7325 ( .A(n7096), .B(n7095), .Z(n7100) );
  NANDN U7326 ( .A(n7098), .B(n7097), .Z(n7099) );
  AND U7327 ( .A(n7100), .B(n7099), .Z(n7131) );
  NAND U7328 ( .A(n26), .B(n7101), .Z(n7103) );
  XOR U7329 ( .A(b[7]), .B(a[171]), .Z(n7142) );
  NAND U7330 ( .A(n10531), .B(n7142), .Z(n7102) );
  AND U7331 ( .A(n7103), .B(n7102), .Z(n7161) );
  NAND U7332 ( .A(n23), .B(n7104), .Z(n7106) );
  XOR U7333 ( .A(b[3]), .B(a[175]), .Z(n7145) );
  NAND U7334 ( .A(n24), .B(n7145), .Z(n7105) );
  NAND U7335 ( .A(n7106), .B(n7105), .Z(n7160) );
  XNOR U7336 ( .A(n7161), .B(n7160), .Z(n7163) );
  NAND U7337 ( .A(b[0]), .B(a[177]), .Z(n7107) );
  XNOR U7338 ( .A(b[1]), .B(n7107), .Z(n7109) );
  NANDN U7339 ( .A(b[0]), .B(a[176]), .Z(n7108) );
  NAND U7340 ( .A(n7109), .B(n7108), .Z(n7157) );
  NAND U7341 ( .A(n25), .B(n7110), .Z(n7112) );
  XOR U7342 ( .A(b[5]), .B(a[173]), .Z(n7148) );
  NAND U7343 ( .A(n10456), .B(n7148), .Z(n7111) );
  AND U7344 ( .A(n7112), .B(n7111), .Z(n7155) );
  AND U7345 ( .A(b[7]), .B(a[169]), .Z(n7154) );
  XNOR U7346 ( .A(n7155), .B(n7154), .Z(n7156) );
  XNOR U7347 ( .A(n7157), .B(n7156), .Z(n7162) );
  XOR U7348 ( .A(n7163), .B(n7162), .Z(n7137) );
  NANDN U7349 ( .A(n7114), .B(n7113), .Z(n7118) );
  NANDN U7350 ( .A(n7116), .B(n7115), .Z(n7117) );
  AND U7351 ( .A(n7118), .B(n7117), .Z(n7136) );
  XNOR U7352 ( .A(n7137), .B(n7136), .Z(n7138) );
  NANDN U7353 ( .A(n7120), .B(n7119), .Z(n7124) );
  NAND U7354 ( .A(n7122), .B(n7121), .Z(n7123) );
  NAND U7355 ( .A(n7124), .B(n7123), .Z(n7139) );
  XNOR U7356 ( .A(n7138), .B(n7139), .Z(n7130) );
  XNOR U7357 ( .A(n7131), .B(n7130), .Z(n7132) );
  XNOR U7358 ( .A(n7133), .B(n7132), .Z(n7166) );
  XNOR U7359 ( .A(sreg[425]), .B(n7166), .Z(n7168) );
  NANDN U7360 ( .A(sreg[424]), .B(n7125), .Z(n7129) );
  NAND U7361 ( .A(n7127), .B(n7126), .Z(n7128) );
  NAND U7362 ( .A(n7129), .B(n7128), .Z(n7167) );
  XNOR U7363 ( .A(n7168), .B(n7167), .Z(c[425]) );
  NANDN U7364 ( .A(n7131), .B(n7130), .Z(n7135) );
  NANDN U7365 ( .A(n7133), .B(n7132), .Z(n7134) );
  AND U7366 ( .A(n7135), .B(n7134), .Z(n7174) );
  NANDN U7367 ( .A(n7137), .B(n7136), .Z(n7141) );
  NANDN U7368 ( .A(n7139), .B(n7138), .Z(n7140) );
  AND U7369 ( .A(n7141), .B(n7140), .Z(n7172) );
  NAND U7370 ( .A(n26), .B(n7142), .Z(n7144) );
  XOR U7371 ( .A(b[7]), .B(a[172]), .Z(n7183) );
  NAND U7372 ( .A(n10531), .B(n7183), .Z(n7143) );
  AND U7373 ( .A(n7144), .B(n7143), .Z(n7202) );
  NAND U7374 ( .A(n23), .B(n7145), .Z(n7147) );
  XOR U7375 ( .A(b[3]), .B(a[176]), .Z(n7186) );
  NAND U7376 ( .A(n24), .B(n7186), .Z(n7146) );
  NAND U7377 ( .A(n7147), .B(n7146), .Z(n7201) );
  XNOR U7378 ( .A(n7202), .B(n7201), .Z(n7204) );
  NAND U7379 ( .A(n25), .B(n7148), .Z(n7150) );
  XOR U7380 ( .A(b[5]), .B(a[174]), .Z(n7192) );
  NAND U7381 ( .A(n10456), .B(n7192), .Z(n7149) );
  AND U7382 ( .A(n7150), .B(n7149), .Z(n7196) );
  AND U7383 ( .A(b[7]), .B(a[170]), .Z(n7195) );
  XNOR U7384 ( .A(n7196), .B(n7195), .Z(n7197) );
  NAND U7385 ( .A(b[0]), .B(a[178]), .Z(n7151) );
  XNOR U7386 ( .A(b[1]), .B(n7151), .Z(n7153) );
  NANDN U7387 ( .A(b[0]), .B(a[177]), .Z(n7152) );
  NAND U7388 ( .A(n7153), .B(n7152), .Z(n7198) );
  XNOR U7389 ( .A(n7197), .B(n7198), .Z(n7203) );
  XOR U7390 ( .A(n7204), .B(n7203), .Z(n7178) );
  NANDN U7391 ( .A(n7155), .B(n7154), .Z(n7159) );
  NANDN U7392 ( .A(n7157), .B(n7156), .Z(n7158) );
  AND U7393 ( .A(n7159), .B(n7158), .Z(n7177) );
  XNOR U7394 ( .A(n7178), .B(n7177), .Z(n7179) );
  NANDN U7395 ( .A(n7161), .B(n7160), .Z(n7165) );
  NAND U7396 ( .A(n7163), .B(n7162), .Z(n7164) );
  NAND U7397 ( .A(n7165), .B(n7164), .Z(n7180) );
  XNOR U7398 ( .A(n7179), .B(n7180), .Z(n7171) );
  XNOR U7399 ( .A(n7172), .B(n7171), .Z(n7173) );
  XNOR U7400 ( .A(n7174), .B(n7173), .Z(n7207) );
  XNOR U7401 ( .A(sreg[426]), .B(n7207), .Z(n7209) );
  NANDN U7402 ( .A(sreg[425]), .B(n7166), .Z(n7170) );
  NAND U7403 ( .A(n7168), .B(n7167), .Z(n7169) );
  NAND U7404 ( .A(n7170), .B(n7169), .Z(n7208) );
  XNOR U7405 ( .A(n7209), .B(n7208), .Z(c[426]) );
  NANDN U7406 ( .A(n7172), .B(n7171), .Z(n7176) );
  NANDN U7407 ( .A(n7174), .B(n7173), .Z(n7175) );
  AND U7408 ( .A(n7176), .B(n7175), .Z(n7215) );
  NANDN U7409 ( .A(n7178), .B(n7177), .Z(n7182) );
  NANDN U7410 ( .A(n7180), .B(n7179), .Z(n7181) );
  AND U7411 ( .A(n7182), .B(n7181), .Z(n7213) );
  NAND U7412 ( .A(n26), .B(n7183), .Z(n7185) );
  XOR U7413 ( .A(b[7]), .B(a[173]), .Z(n7224) );
  NAND U7414 ( .A(n10531), .B(n7224), .Z(n7184) );
  AND U7415 ( .A(n7185), .B(n7184), .Z(n7243) );
  NAND U7416 ( .A(n23), .B(n7186), .Z(n7188) );
  XOR U7417 ( .A(b[3]), .B(a[177]), .Z(n7227) );
  NAND U7418 ( .A(n24), .B(n7227), .Z(n7187) );
  NAND U7419 ( .A(n7188), .B(n7187), .Z(n7242) );
  XNOR U7420 ( .A(n7243), .B(n7242), .Z(n7245) );
  NAND U7421 ( .A(b[0]), .B(a[179]), .Z(n7189) );
  XNOR U7422 ( .A(b[1]), .B(n7189), .Z(n7191) );
  NANDN U7423 ( .A(b[0]), .B(a[178]), .Z(n7190) );
  NAND U7424 ( .A(n7191), .B(n7190), .Z(n7239) );
  NAND U7425 ( .A(n25), .B(n7192), .Z(n7194) );
  XOR U7426 ( .A(b[5]), .B(a[175]), .Z(n7233) );
  NAND U7427 ( .A(n10456), .B(n7233), .Z(n7193) );
  AND U7428 ( .A(n7194), .B(n7193), .Z(n7237) );
  AND U7429 ( .A(b[7]), .B(a[171]), .Z(n7236) );
  XNOR U7430 ( .A(n7237), .B(n7236), .Z(n7238) );
  XNOR U7431 ( .A(n7239), .B(n7238), .Z(n7244) );
  XOR U7432 ( .A(n7245), .B(n7244), .Z(n7219) );
  NANDN U7433 ( .A(n7196), .B(n7195), .Z(n7200) );
  NANDN U7434 ( .A(n7198), .B(n7197), .Z(n7199) );
  AND U7435 ( .A(n7200), .B(n7199), .Z(n7218) );
  XNOR U7436 ( .A(n7219), .B(n7218), .Z(n7220) );
  NANDN U7437 ( .A(n7202), .B(n7201), .Z(n7206) );
  NAND U7438 ( .A(n7204), .B(n7203), .Z(n7205) );
  NAND U7439 ( .A(n7206), .B(n7205), .Z(n7221) );
  XNOR U7440 ( .A(n7220), .B(n7221), .Z(n7212) );
  XNOR U7441 ( .A(n7213), .B(n7212), .Z(n7214) );
  XNOR U7442 ( .A(n7215), .B(n7214), .Z(n7248) );
  XNOR U7443 ( .A(sreg[427]), .B(n7248), .Z(n7250) );
  NANDN U7444 ( .A(sreg[426]), .B(n7207), .Z(n7211) );
  NAND U7445 ( .A(n7209), .B(n7208), .Z(n7210) );
  NAND U7446 ( .A(n7211), .B(n7210), .Z(n7249) );
  XNOR U7447 ( .A(n7250), .B(n7249), .Z(c[427]) );
  NANDN U7448 ( .A(n7213), .B(n7212), .Z(n7217) );
  NANDN U7449 ( .A(n7215), .B(n7214), .Z(n7216) );
  AND U7450 ( .A(n7217), .B(n7216), .Z(n7256) );
  NANDN U7451 ( .A(n7219), .B(n7218), .Z(n7223) );
  NANDN U7452 ( .A(n7221), .B(n7220), .Z(n7222) );
  AND U7453 ( .A(n7223), .B(n7222), .Z(n7254) );
  NAND U7454 ( .A(n26), .B(n7224), .Z(n7226) );
  XOR U7455 ( .A(b[7]), .B(a[174]), .Z(n7265) );
  NAND U7456 ( .A(n10531), .B(n7265), .Z(n7225) );
  AND U7457 ( .A(n7226), .B(n7225), .Z(n7284) );
  NAND U7458 ( .A(n23), .B(n7227), .Z(n7229) );
  XOR U7459 ( .A(b[3]), .B(a[178]), .Z(n7268) );
  NAND U7460 ( .A(n24), .B(n7268), .Z(n7228) );
  NAND U7461 ( .A(n7229), .B(n7228), .Z(n7283) );
  XNOR U7462 ( .A(n7284), .B(n7283), .Z(n7286) );
  NAND U7463 ( .A(b[0]), .B(a[180]), .Z(n7230) );
  XNOR U7464 ( .A(b[1]), .B(n7230), .Z(n7232) );
  NANDN U7465 ( .A(b[0]), .B(a[179]), .Z(n7231) );
  NAND U7466 ( .A(n7232), .B(n7231), .Z(n7280) );
  NAND U7467 ( .A(n25), .B(n7233), .Z(n7235) );
  XOR U7468 ( .A(b[5]), .B(a[176]), .Z(n7274) );
  NAND U7469 ( .A(n10456), .B(n7274), .Z(n7234) );
  AND U7470 ( .A(n7235), .B(n7234), .Z(n7278) );
  AND U7471 ( .A(b[7]), .B(a[172]), .Z(n7277) );
  XNOR U7472 ( .A(n7278), .B(n7277), .Z(n7279) );
  XNOR U7473 ( .A(n7280), .B(n7279), .Z(n7285) );
  XOR U7474 ( .A(n7286), .B(n7285), .Z(n7260) );
  NANDN U7475 ( .A(n7237), .B(n7236), .Z(n7241) );
  NANDN U7476 ( .A(n7239), .B(n7238), .Z(n7240) );
  AND U7477 ( .A(n7241), .B(n7240), .Z(n7259) );
  XNOR U7478 ( .A(n7260), .B(n7259), .Z(n7261) );
  NANDN U7479 ( .A(n7243), .B(n7242), .Z(n7247) );
  NAND U7480 ( .A(n7245), .B(n7244), .Z(n7246) );
  NAND U7481 ( .A(n7247), .B(n7246), .Z(n7262) );
  XNOR U7482 ( .A(n7261), .B(n7262), .Z(n7253) );
  XNOR U7483 ( .A(n7254), .B(n7253), .Z(n7255) );
  XNOR U7484 ( .A(n7256), .B(n7255), .Z(n7289) );
  XNOR U7485 ( .A(sreg[428]), .B(n7289), .Z(n7291) );
  NANDN U7486 ( .A(sreg[427]), .B(n7248), .Z(n7252) );
  NAND U7487 ( .A(n7250), .B(n7249), .Z(n7251) );
  NAND U7488 ( .A(n7252), .B(n7251), .Z(n7290) );
  XNOR U7489 ( .A(n7291), .B(n7290), .Z(c[428]) );
  NANDN U7490 ( .A(n7254), .B(n7253), .Z(n7258) );
  NANDN U7491 ( .A(n7256), .B(n7255), .Z(n7257) );
  AND U7492 ( .A(n7258), .B(n7257), .Z(n7297) );
  NANDN U7493 ( .A(n7260), .B(n7259), .Z(n7264) );
  NANDN U7494 ( .A(n7262), .B(n7261), .Z(n7263) );
  AND U7495 ( .A(n7264), .B(n7263), .Z(n7295) );
  NAND U7496 ( .A(n26), .B(n7265), .Z(n7267) );
  XOR U7497 ( .A(b[7]), .B(a[175]), .Z(n7306) );
  NAND U7498 ( .A(n10531), .B(n7306), .Z(n7266) );
  AND U7499 ( .A(n7267), .B(n7266), .Z(n7325) );
  NAND U7500 ( .A(n23), .B(n7268), .Z(n7270) );
  XOR U7501 ( .A(b[3]), .B(a[179]), .Z(n7309) );
  NAND U7502 ( .A(n24), .B(n7309), .Z(n7269) );
  NAND U7503 ( .A(n7270), .B(n7269), .Z(n7324) );
  XNOR U7504 ( .A(n7325), .B(n7324), .Z(n7327) );
  NAND U7505 ( .A(b[0]), .B(a[181]), .Z(n7271) );
  XNOR U7506 ( .A(b[1]), .B(n7271), .Z(n7273) );
  NANDN U7507 ( .A(b[0]), .B(a[180]), .Z(n7272) );
  NAND U7508 ( .A(n7273), .B(n7272), .Z(n7321) );
  NAND U7509 ( .A(n25), .B(n7274), .Z(n7276) );
  XOR U7510 ( .A(b[5]), .B(a[177]), .Z(n7315) );
  NAND U7511 ( .A(n10456), .B(n7315), .Z(n7275) );
  AND U7512 ( .A(n7276), .B(n7275), .Z(n7319) );
  AND U7513 ( .A(b[7]), .B(a[173]), .Z(n7318) );
  XNOR U7514 ( .A(n7319), .B(n7318), .Z(n7320) );
  XNOR U7515 ( .A(n7321), .B(n7320), .Z(n7326) );
  XOR U7516 ( .A(n7327), .B(n7326), .Z(n7301) );
  NANDN U7517 ( .A(n7278), .B(n7277), .Z(n7282) );
  NANDN U7518 ( .A(n7280), .B(n7279), .Z(n7281) );
  AND U7519 ( .A(n7282), .B(n7281), .Z(n7300) );
  XNOR U7520 ( .A(n7301), .B(n7300), .Z(n7302) );
  NANDN U7521 ( .A(n7284), .B(n7283), .Z(n7288) );
  NAND U7522 ( .A(n7286), .B(n7285), .Z(n7287) );
  NAND U7523 ( .A(n7288), .B(n7287), .Z(n7303) );
  XNOR U7524 ( .A(n7302), .B(n7303), .Z(n7294) );
  XNOR U7525 ( .A(n7295), .B(n7294), .Z(n7296) );
  XNOR U7526 ( .A(n7297), .B(n7296), .Z(n7330) );
  XNOR U7527 ( .A(sreg[429]), .B(n7330), .Z(n7332) );
  NANDN U7528 ( .A(sreg[428]), .B(n7289), .Z(n7293) );
  NAND U7529 ( .A(n7291), .B(n7290), .Z(n7292) );
  NAND U7530 ( .A(n7293), .B(n7292), .Z(n7331) );
  XNOR U7531 ( .A(n7332), .B(n7331), .Z(c[429]) );
  NANDN U7532 ( .A(n7295), .B(n7294), .Z(n7299) );
  NANDN U7533 ( .A(n7297), .B(n7296), .Z(n7298) );
  AND U7534 ( .A(n7299), .B(n7298), .Z(n7338) );
  NANDN U7535 ( .A(n7301), .B(n7300), .Z(n7305) );
  NANDN U7536 ( .A(n7303), .B(n7302), .Z(n7304) );
  AND U7537 ( .A(n7305), .B(n7304), .Z(n7336) );
  NAND U7538 ( .A(n26), .B(n7306), .Z(n7308) );
  XOR U7539 ( .A(b[7]), .B(a[176]), .Z(n7347) );
  NAND U7540 ( .A(n10531), .B(n7347), .Z(n7307) );
  AND U7541 ( .A(n7308), .B(n7307), .Z(n7366) );
  NAND U7542 ( .A(n23), .B(n7309), .Z(n7311) );
  XOR U7543 ( .A(b[3]), .B(a[180]), .Z(n7350) );
  NAND U7544 ( .A(n24), .B(n7350), .Z(n7310) );
  NAND U7545 ( .A(n7311), .B(n7310), .Z(n7365) );
  XNOR U7546 ( .A(n7366), .B(n7365), .Z(n7368) );
  NAND U7547 ( .A(b[0]), .B(a[182]), .Z(n7312) );
  XNOR U7548 ( .A(b[1]), .B(n7312), .Z(n7314) );
  NANDN U7549 ( .A(b[0]), .B(a[181]), .Z(n7313) );
  NAND U7550 ( .A(n7314), .B(n7313), .Z(n7362) );
  NAND U7551 ( .A(n25), .B(n7315), .Z(n7317) );
  XOR U7552 ( .A(b[5]), .B(a[178]), .Z(n7356) );
  NAND U7553 ( .A(n10456), .B(n7356), .Z(n7316) );
  AND U7554 ( .A(n7317), .B(n7316), .Z(n7360) );
  AND U7555 ( .A(b[7]), .B(a[174]), .Z(n7359) );
  XNOR U7556 ( .A(n7360), .B(n7359), .Z(n7361) );
  XNOR U7557 ( .A(n7362), .B(n7361), .Z(n7367) );
  XOR U7558 ( .A(n7368), .B(n7367), .Z(n7342) );
  NANDN U7559 ( .A(n7319), .B(n7318), .Z(n7323) );
  NANDN U7560 ( .A(n7321), .B(n7320), .Z(n7322) );
  AND U7561 ( .A(n7323), .B(n7322), .Z(n7341) );
  XNOR U7562 ( .A(n7342), .B(n7341), .Z(n7343) );
  NANDN U7563 ( .A(n7325), .B(n7324), .Z(n7329) );
  NAND U7564 ( .A(n7327), .B(n7326), .Z(n7328) );
  NAND U7565 ( .A(n7329), .B(n7328), .Z(n7344) );
  XNOR U7566 ( .A(n7343), .B(n7344), .Z(n7335) );
  XNOR U7567 ( .A(n7336), .B(n7335), .Z(n7337) );
  XNOR U7568 ( .A(n7338), .B(n7337), .Z(n7371) );
  XNOR U7569 ( .A(sreg[430]), .B(n7371), .Z(n7373) );
  NANDN U7570 ( .A(sreg[429]), .B(n7330), .Z(n7334) );
  NAND U7571 ( .A(n7332), .B(n7331), .Z(n7333) );
  NAND U7572 ( .A(n7334), .B(n7333), .Z(n7372) );
  XNOR U7573 ( .A(n7373), .B(n7372), .Z(c[430]) );
  NANDN U7574 ( .A(n7336), .B(n7335), .Z(n7340) );
  NANDN U7575 ( .A(n7338), .B(n7337), .Z(n7339) );
  AND U7576 ( .A(n7340), .B(n7339), .Z(n7379) );
  NANDN U7577 ( .A(n7342), .B(n7341), .Z(n7346) );
  NANDN U7578 ( .A(n7344), .B(n7343), .Z(n7345) );
  AND U7579 ( .A(n7346), .B(n7345), .Z(n7377) );
  NAND U7580 ( .A(n26), .B(n7347), .Z(n7349) );
  XOR U7581 ( .A(b[7]), .B(a[177]), .Z(n7388) );
  NAND U7582 ( .A(n10531), .B(n7388), .Z(n7348) );
  AND U7583 ( .A(n7349), .B(n7348), .Z(n7407) );
  NAND U7584 ( .A(n23), .B(n7350), .Z(n7352) );
  XOR U7585 ( .A(b[3]), .B(a[181]), .Z(n7391) );
  NAND U7586 ( .A(n24), .B(n7391), .Z(n7351) );
  NAND U7587 ( .A(n7352), .B(n7351), .Z(n7406) );
  XNOR U7588 ( .A(n7407), .B(n7406), .Z(n7409) );
  NAND U7589 ( .A(b[0]), .B(a[183]), .Z(n7353) );
  XNOR U7590 ( .A(b[1]), .B(n7353), .Z(n7355) );
  NANDN U7591 ( .A(b[0]), .B(a[182]), .Z(n7354) );
  NAND U7592 ( .A(n7355), .B(n7354), .Z(n7403) );
  NAND U7593 ( .A(n25), .B(n7356), .Z(n7358) );
  XOR U7594 ( .A(b[5]), .B(a[179]), .Z(n7397) );
  NAND U7595 ( .A(n10456), .B(n7397), .Z(n7357) );
  AND U7596 ( .A(n7358), .B(n7357), .Z(n7401) );
  AND U7597 ( .A(b[7]), .B(a[175]), .Z(n7400) );
  XNOR U7598 ( .A(n7401), .B(n7400), .Z(n7402) );
  XNOR U7599 ( .A(n7403), .B(n7402), .Z(n7408) );
  XOR U7600 ( .A(n7409), .B(n7408), .Z(n7383) );
  NANDN U7601 ( .A(n7360), .B(n7359), .Z(n7364) );
  NANDN U7602 ( .A(n7362), .B(n7361), .Z(n7363) );
  AND U7603 ( .A(n7364), .B(n7363), .Z(n7382) );
  XNOR U7604 ( .A(n7383), .B(n7382), .Z(n7384) );
  NANDN U7605 ( .A(n7366), .B(n7365), .Z(n7370) );
  NAND U7606 ( .A(n7368), .B(n7367), .Z(n7369) );
  NAND U7607 ( .A(n7370), .B(n7369), .Z(n7385) );
  XNOR U7608 ( .A(n7384), .B(n7385), .Z(n7376) );
  XNOR U7609 ( .A(n7377), .B(n7376), .Z(n7378) );
  XNOR U7610 ( .A(n7379), .B(n7378), .Z(n7412) );
  XNOR U7611 ( .A(sreg[431]), .B(n7412), .Z(n7414) );
  NANDN U7612 ( .A(sreg[430]), .B(n7371), .Z(n7375) );
  NAND U7613 ( .A(n7373), .B(n7372), .Z(n7374) );
  NAND U7614 ( .A(n7375), .B(n7374), .Z(n7413) );
  XNOR U7615 ( .A(n7414), .B(n7413), .Z(c[431]) );
  NANDN U7616 ( .A(n7377), .B(n7376), .Z(n7381) );
  NANDN U7617 ( .A(n7379), .B(n7378), .Z(n7380) );
  AND U7618 ( .A(n7381), .B(n7380), .Z(n7420) );
  NANDN U7619 ( .A(n7383), .B(n7382), .Z(n7387) );
  NANDN U7620 ( .A(n7385), .B(n7384), .Z(n7386) );
  AND U7621 ( .A(n7387), .B(n7386), .Z(n7418) );
  NAND U7622 ( .A(n26), .B(n7388), .Z(n7390) );
  XOR U7623 ( .A(b[7]), .B(a[178]), .Z(n7429) );
  NAND U7624 ( .A(n10531), .B(n7429), .Z(n7389) );
  AND U7625 ( .A(n7390), .B(n7389), .Z(n7448) );
  NAND U7626 ( .A(n23), .B(n7391), .Z(n7393) );
  XOR U7627 ( .A(b[3]), .B(a[182]), .Z(n7432) );
  NAND U7628 ( .A(n24), .B(n7432), .Z(n7392) );
  NAND U7629 ( .A(n7393), .B(n7392), .Z(n7447) );
  XNOR U7630 ( .A(n7448), .B(n7447), .Z(n7450) );
  NAND U7631 ( .A(b[0]), .B(a[184]), .Z(n7394) );
  XNOR U7632 ( .A(b[1]), .B(n7394), .Z(n7396) );
  NANDN U7633 ( .A(b[0]), .B(a[183]), .Z(n7395) );
  NAND U7634 ( .A(n7396), .B(n7395), .Z(n7444) );
  NAND U7635 ( .A(n25), .B(n7397), .Z(n7399) );
  XOR U7636 ( .A(b[5]), .B(a[180]), .Z(n7435) );
  NAND U7637 ( .A(n10456), .B(n7435), .Z(n7398) );
  AND U7638 ( .A(n7399), .B(n7398), .Z(n7442) );
  AND U7639 ( .A(b[7]), .B(a[176]), .Z(n7441) );
  XNOR U7640 ( .A(n7442), .B(n7441), .Z(n7443) );
  XNOR U7641 ( .A(n7444), .B(n7443), .Z(n7449) );
  XOR U7642 ( .A(n7450), .B(n7449), .Z(n7424) );
  NANDN U7643 ( .A(n7401), .B(n7400), .Z(n7405) );
  NANDN U7644 ( .A(n7403), .B(n7402), .Z(n7404) );
  AND U7645 ( .A(n7405), .B(n7404), .Z(n7423) );
  XNOR U7646 ( .A(n7424), .B(n7423), .Z(n7425) );
  NANDN U7647 ( .A(n7407), .B(n7406), .Z(n7411) );
  NAND U7648 ( .A(n7409), .B(n7408), .Z(n7410) );
  NAND U7649 ( .A(n7411), .B(n7410), .Z(n7426) );
  XNOR U7650 ( .A(n7425), .B(n7426), .Z(n7417) );
  XNOR U7651 ( .A(n7418), .B(n7417), .Z(n7419) );
  XNOR U7652 ( .A(n7420), .B(n7419), .Z(n7453) );
  XNOR U7653 ( .A(sreg[432]), .B(n7453), .Z(n7455) );
  NANDN U7654 ( .A(sreg[431]), .B(n7412), .Z(n7416) );
  NAND U7655 ( .A(n7414), .B(n7413), .Z(n7415) );
  NAND U7656 ( .A(n7416), .B(n7415), .Z(n7454) );
  XNOR U7657 ( .A(n7455), .B(n7454), .Z(c[432]) );
  NANDN U7658 ( .A(n7418), .B(n7417), .Z(n7422) );
  NANDN U7659 ( .A(n7420), .B(n7419), .Z(n7421) );
  AND U7660 ( .A(n7422), .B(n7421), .Z(n7461) );
  NANDN U7661 ( .A(n7424), .B(n7423), .Z(n7428) );
  NANDN U7662 ( .A(n7426), .B(n7425), .Z(n7427) );
  AND U7663 ( .A(n7428), .B(n7427), .Z(n7459) );
  NAND U7664 ( .A(n26), .B(n7429), .Z(n7431) );
  XOR U7665 ( .A(b[7]), .B(a[179]), .Z(n7470) );
  NAND U7666 ( .A(n10531), .B(n7470), .Z(n7430) );
  AND U7667 ( .A(n7431), .B(n7430), .Z(n7489) );
  NAND U7668 ( .A(n23), .B(n7432), .Z(n7434) );
  XOR U7669 ( .A(b[3]), .B(a[183]), .Z(n7473) );
  NAND U7670 ( .A(n24), .B(n7473), .Z(n7433) );
  NAND U7671 ( .A(n7434), .B(n7433), .Z(n7488) );
  XNOR U7672 ( .A(n7489), .B(n7488), .Z(n7491) );
  NAND U7673 ( .A(n25), .B(n7435), .Z(n7437) );
  XOR U7674 ( .A(b[5]), .B(a[181]), .Z(n7479) );
  NAND U7675 ( .A(n10456), .B(n7479), .Z(n7436) );
  AND U7676 ( .A(n7437), .B(n7436), .Z(n7483) );
  AND U7677 ( .A(b[7]), .B(a[177]), .Z(n7482) );
  XNOR U7678 ( .A(n7483), .B(n7482), .Z(n7484) );
  NAND U7679 ( .A(b[0]), .B(a[185]), .Z(n7438) );
  XNOR U7680 ( .A(b[1]), .B(n7438), .Z(n7440) );
  NANDN U7681 ( .A(b[0]), .B(a[184]), .Z(n7439) );
  NAND U7682 ( .A(n7440), .B(n7439), .Z(n7485) );
  XNOR U7683 ( .A(n7484), .B(n7485), .Z(n7490) );
  XOR U7684 ( .A(n7491), .B(n7490), .Z(n7465) );
  NANDN U7685 ( .A(n7442), .B(n7441), .Z(n7446) );
  NANDN U7686 ( .A(n7444), .B(n7443), .Z(n7445) );
  AND U7687 ( .A(n7446), .B(n7445), .Z(n7464) );
  XNOR U7688 ( .A(n7465), .B(n7464), .Z(n7466) );
  NANDN U7689 ( .A(n7448), .B(n7447), .Z(n7452) );
  NAND U7690 ( .A(n7450), .B(n7449), .Z(n7451) );
  NAND U7691 ( .A(n7452), .B(n7451), .Z(n7467) );
  XNOR U7692 ( .A(n7466), .B(n7467), .Z(n7458) );
  XNOR U7693 ( .A(n7459), .B(n7458), .Z(n7460) );
  XNOR U7694 ( .A(n7461), .B(n7460), .Z(n7494) );
  XNOR U7695 ( .A(sreg[433]), .B(n7494), .Z(n7496) );
  NANDN U7696 ( .A(sreg[432]), .B(n7453), .Z(n7457) );
  NAND U7697 ( .A(n7455), .B(n7454), .Z(n7456) );
  NAND U7698 ( .A(n7457), .B(n7456), .Z(n7495) );
  XNOR U7699 ( .A(n7496), .B(n7495), .Z(c[433]) );
  NANDN U7700 ( .A(n7459), .B(n7458), .Z(n7463) );
  NANDN U7701 ( .A(n7461), .B(n7460), .Z(n7462) );
  AND U7702 ( .A(n7463), .B(n7462), .Z(n7502) );
  NANDN U7703 ( .A(n7465), .B(n7464), .Z(n7469) );
  NANDN U7704 ( .A(n7467), .B(n7466), .Z(n7468) );
  AND U7705 ( .A(n7469), .B(n7468), .Z(n7500) );
  NAND U7706 ( .A(n26), .B(n7470), .Z(n7472) );
  XOR U7707 ( .A(b[7]), .B(a[180]), .Z(n7511) );
  NAND U7708 ( .A(n10531), .B(n7511), .Z(n7471) );
  AND U7709 ( .A(n7472), .B(n7471), .Z(n7530) );
  NAND U7710 ( .A(n23), .B(n7473), .Z(n7475) );
  XOR U7711 ( .A(b[3]), .B(a[184]), .Z(n7514) );
  NAND U7712 ( .A(n24), .B(n7514), .Z(n7474) );
  NAND U7713 ( .A(n7475), .B(n7474), .Z(n7529) );
  XNOR U7714 ( .A(n7530), .B(n7529), .Z(n7532) );
  NAND U7715 ( .A(b[0]), .B(a[186]), .Z(n7476) );
  XNOR U7716 ( .A(b[1]), .B(n7476), .Z(n7478) );
  NANDN U7717 ( .A(b[0]), .B(a[185]), .Z(n7477) );
  NAND U7718 ( .A(n7478), .B(n7477), .Z(n7526) );
  NAND U7719 ( .A(n25), .B(n7479), .Z(n7481) );
  XOR U7720 ( .A(b[5]), .B(a[182]), .Z(n7520) );
  NAND U7721 ( .A(n10456), .B(n7520), .Z(n7480) );
  AND U7722 ( .A(n7481), .B(n7480), .Z(n7524) );
  AND U7723 ( .A(b[7]), .B(a[178]), .Z(n7523) );
  XNOR U7724 ( .A(n7524), .B(n7523), .Z(n7525) );
  XNOR U7725 ( .A(n7526), .B(n7525), .Z(n7531) );
  XOR U7726 ( .A(n7532), .B(n7531), .Z(n7506) );
  NANDN U7727 ( .A(n7483), .B(n7482), .Z(n7487) );
  NANDN U7728 ( .A(n7485), .B(n7484), .Z(n7486) );
  AND U7729 ( .A(n7487), .B(n7486), .Z(n7505) );
  XNOR U7730 ( .A(n7506), .B(n7505), .Z(n7507) );
  NANDN U7731 ( .A(n7489), .B(n7488), .Z(n7493) );
  NAND U7732 ( .A(n7491), .B(n7490), .Z(n7492) );
  NAND U7733 ( .A(n7493), .B(n7492), .Z(n7508) );
  XNOR U7734 ( .A(n7507), .B(n7508), .Z(n7499) );
  XNOR U7735 ( .A(n7500), .B(n7499), .Z(n7501) );
  XNOR U7736 ( .A(n7502), .B(n7501), .Z(n7535) );
  XNOR U7737 ( .A(sreg[434]), .B(n7535), .Z(n7537) );
  NANDN U7738 ( .A(sreg[433]), .B(n7494), .Z(n7498) );
  NAND U7739 ( .A(n7496), .B(n7495), .Z(n7497) );
  NAND U7740 ( .A(n7498), .B(n7497), .Z(n7536) );
  XNOR U7741 ( .A(n7537), .B(n7536), .Z(c[434]) );
  NANDN U7742 ( .A(n7500), .B(n7499), .Z(n7504) );
  NANDN U7743 ( .A(n7502), .B(n7501), .Z(n7503) );
  AND U7744 ( .A(n7504), .B(n7503), .Z(n7543) );
  NANDN U7745 ( .A(n7506), .B(n7505), .Z(n7510) );
  NANDN U7746 ( .A(n7508), .B(n7507), .Z(n7509) );
  AND U7747 ( .A(n7510), .B(n7509), .Z(n7541) );
  NAND U7748 ( .A(n26), .B(n7511), .Z(n7513) );
  XOR U7749 ( .A(b[7]), .B(a[181]), .Z(n7552) );
  NAND U7750 ( .A(n10531), .B(n7552), .Z(n7512) );
  AND U7751 ( .A(n7513), .B(n7512), .Z(n7571) );
  NAND U7752 ( .A(n23), .B(n7514), .Z(n7516) );
  XOR U7753 ( .A(b[3]), .B(a[185]), .Z(n7555) );
  NAND U7754 ( .A(n24), .B(n7555), .Z(n7515) );
  NAND U7755 ( .A(n7516), .B(n7515), .Z(n7570) );
  XNOR U7756 ( .A(n7571), .B(n7570), .Z(n7573) );
  NAND U7757 ( .A(b[0]), .B(a[187]), .Z(n7517) );
  XNOR U7758 ( .A(b[1]), .B(n7517), .Z(n7519) );
  NANDN U7759 ( .A(b[0]), .B(a[186]), .Z(n7518) );
  NAND U7760 ( .A(n7519), .B(n7518), .Z(n7567) );
  NAND U7761 ( .A(n25), .B(n7520), .Z(n7522) );
  XOR U7762 ( .A(b[5]), .B(a[183]), .Z(n7561) );
  NAND U7763 ( .A(n10456), .B(n7561), .Z(n7521) );
  AND U7764 ( .A(n7522), .B(n7521), .Z(n7565) );
  AND U7765 ( .A(b[7]), .B(a[179]), .Z(n7564) );
  XNOR U7766 ( .A(n7565), .B(n7564), .Z(n7566) );
  XNOR U7767 ( .A(n7567), .B(n7566), .Z(n7572) );
  XOR U7768 ( .A(n7573), .B(n7572), .Z(n7547) );
  NANDN U7769 ( .A(n7524), .B(n7523), .Z(n7528) );
  NANDN U7770 ( .A(n7526), .B(n7525), .Z(n7527) );
  AND U7771 ( .A(n7528), .B(n7527), .Z(n7546) );
  XNOR U7772 ( .A(n7547), .B(n7546), .Z(n7548) );
  NANDN U7773 ( .A(n7530), .B(n7529), .Z(n7534) );
  NAND U7774 ( .A(n7532), .B(n7531), .Z(n7533) );
  NAND U7775 ( .A(n7534), .B(n7533), .Z(n7549) );
  XNOR U7776 ( .A(n7548), .B(n7549), .Z(n7540) );
  XNOR U7777 ( .A(n7541), .B(n7540), .Z(n7542) );
  XNOR U7778 ( .A(n7543), .B(n7542), .Z(n7576) );
  XNOR U7779 ( .A(sreg[435]), .B(n7576), .Z(n7578) );
  NANDN U7780 ( .A(sreg[434]), .B(n7535), .Z(n7539) );
  NAND U7781 ( .A(n7537), .B(n7536), .Z(n7538) );
  NAND U7782 ( .A(n7539), .B(n7538), .Z(n7577) );
  XNOR U7783 ( .A(n7578), .B(n7577), .Z(c[435]) );
  NANDN U7784 ( .A(n7541), .B(n7540), .Z(n7545) );
  NANDN U7785 ( .A(n7543), .B(n7542), .Z(n7544) );
  AND U7786 ( .A(n7545), .B(n7544), .Z(n7584) );
  NANDN U7787 ( .A(n7547), .B(n7546), .Z(n7551) );
  NANDN U7788 ( .A(n7549), .B(n7548), .Z(n7550) );
  AND U7789 ( .A(n7551), .B(n7550), .Z(n7582) );
  NAND U7790 ( .A(n26), .B(n7552), .Z(n7554) );
  XOR U7791 ( .A(b[7]), .B(a[182]), .Z(n7593) );
  NAND U7792 ( .A(n10531), .B(n7593), .Z(n7553) );
  AND U7793 ( .A(n7554), .B(n7553), .Z(n7612) );
  NAND U7794 ( .A(n23), .B(n7555), .Z(n7557) );
  XOR U7795 ( .A(b[3]), .B(a[186]), .Z(n7596) );
  NAND U7796 ( .A(n24), .B(n7596), .Z(n7556) );
  NAND U7797 ( .A(n7557), .B(n7556), .Z(n7611) );
  XNOR U7798 ( .A(n7612), .B(n7611), .Z(n7614) );
  NAND U7799 ( .A(b[0]), .B(a[188]), .Z(n7558) );
  XNOR U7800 ( .A(b[1]), .B(n7558), .Z(n7560) );
  NANDN U7801 ( .A(b[0]), .B(a[187]), .Z(n7559) );
  NAND U7802 ( .A(n7560), .B(n7559), .Z(n7608) );
  NAND U7803 ( .A(n25), .B(n7561), .Z(n7563) );
  XOR U7804 ( .A(b[5]), .B(a[184]), .Z(n7599) );
  NAND U7805 ( .A(n10456), .B(n7599), .Z(n7562) );
  AND U7806 ( .A(n7563), .B(n7562), .Z(n7606) );
  AND U7807 ( .A(b[7]), .B(a[180]), .Z(n7605) );
  XNOR U7808 ( .A(n7606), .B(n7605), .Z(n7607) );
  XNOR U7809 ( .A(n7608), .B(n7607), .Z(n7613) );
  XOR U7810 ( .A(n7614), .B(n7613), .Z(n7588) );
  NANDN U7811 ( .A(n7565), .B(n7564), .Z(n7569) );
  NANDN U7812 ( .A(n7567), .B(n7566), .Z(n7568) );
  AND U7813 ( .A(n7569), .B(n7568), .Z(n7587) );
  XNOR U7814 ( .A(n7588), .B(n7587), .Z(n7589) );
  NANDN U7815 ( .A(n7571), .B(n7570), .Z(n7575) );
  NAND U7816 ( .A(n7573), .B(n7572), .Z(n7574) );
  NAND U7817 ( .A(n7575), .B(n7574), .Z(n7590) );
  XNOR U7818 ( .A(n7589), .B(n7590), .Z(n7581) );
  XNOR U7819 ( .A(n7582), .B(n7581), .Z(n7583) );
  XNOR U7820 ( .A(n7584), .B(n7583), .Z(n7617) );
  XNOR U7821 ( .A(sreg[436]), .B(n7617), .Z(n7619) );
  NANDN U7822 ( .A(sreg[435]), .B(n7576), .Z(n7580) );
  NAND U7823 ( .A(n7578), .B(n7577), .Z(n7579) );
  NAND U7824 ( .A(n7580), .B(n7579), .Z(n7618) );
  XNOR U7825 ( .A(n7619), .B(n7618), .Z(c[436]) );
  NANDN U7826 ( .A(n7582), .B(n7581), .Z(n7586) );
  NANDN U7827 ( .A(n7584), .B(n7583), .Z(n7585) );
  AND U7828 ( .A(n7586), .B(n7585), .Z(n7625) );
  NANDN U7829 ( .A(n7588), .B(n7587), .Z(n7592) );
  NANDN U7830 ( .A(n7590), .B(n7589), .Z(n7591) );
  AND U7831 ( .A(n7592), .B(n7591), .Z(n7623) );
  NAND U7832 ( .A(n26), .B(n7593), .Z(n7595) );
  XOR U7833 ( .A(b[7]), .B(a[183]), .Z(n7634) );
  NAND U7834 ( .A(n10531), .B(n7634), .Z(n7594) );
  AND U7835 ( .A(n7595), .B(n7594), .Z(n7653) );
  NAND U7836 ( .A(n23), .B(n7596), .Z(n7598) );
  XOR U7837 ( .A(b[3]), .B(a[187]), .Z(n7637) );
  NAND U7838 ( .A(n24), .B(n7637), .Z(n7597) );
  NAND U7839 ( .A(n7598), .B(n7597), .Z(n7652) );
  XNOR U7840 ( .A(n7653), .B(n7652), .Z(n7655) );
  NAND U7841 ( .A(n25), .B(n7599), .Z(n7601) );
  XOR U7842 ( .A(b[5]), .B(a[185]), .Z(n7643) );
  NAND U7843 ( .A(n10456), .B(n7643), .Z(n7600) );
  AND U7844 ( .A(n7601), .B(n7600), .Z(n7647) );
  AND U7845 ( .A(b[7]), .B(a[181]), .Z(n7646) );
  XNOR U7846 ( .A(n7647), .B(n7646), .Z(n7648) );
  NAND U7847 ( .A(b[0]), .B(a[189]), .Z(n7602) );
  XNOR U7848 ( .A(b[1]), .B(n7602), .Z(n7604) );
  NANDN U7849 ( .A(b[0]), .B(a[188]), .Z(n7603) );
  NAND U7850 ( .A(n7604), .B(n7603), .Z(n7649) );
  XNOR U7851 ( .A(n7648), .B(n7649), .Z(n7654) );
  XOR U7852 ( .A(n7655), .B(n7654), .Z(n7629) );
  NANDN U7853 ( .A(n7606), .B(n7605), .Z(n7610) );
  NANDN U7854 ( .A(n7608), .B(n7607), .Z(n7609) );
  AND U7855 ( .A(n7610), .B(n7609), .Z(n7628) );
  XNOR U7856 ( .A(n7629), .B(n7628), .Z(n7630) );
  NANDN U7857 ( .A(n7612), .B(n7611), .Z(n7616) );
  NAND U7858 ( .A(n7614), .B(n7613), .Z(n7615) );
  NAND U7859 ( .A(n7616), .B(n7615), .Z(n7631) );
  XNOR U7860 ( .A(n7630), .B(n7631), .Z(n7622) );
  XNOR U7861 ( .A(n7623), .B(n7622), .Z(n7624) );
  XNOR U7862 ( .A(n7625), .B(n7624), .Z(n7658) );
  XNOR U7863 ( .A(sreg[437]), .B(n7658), .Z(n7660) );
  NANDN U7864 ( .A(sreg[436]), .B(n7617), .Z(n7621) );
  NAND U7865 ( .A(n7619), .B(n7618), .Z(n7620) );
  NAND U7866 ( .A(n7621), .B(n7620), .Z(n7659) );
  XNOR U7867 ( .A(n7660), .B(n7659), .Z(c[437]) );
  NANDN U7868 ( .A(n7623), .B(n7622), .Z(n7627) );
  NANDN U7869 ( .A(n7625), .B(n7624), .Z(n7626) );
  AND U7870 ( .A(n7627), .B(n7626), .Z(n7666) );
  NANDN U7871 ( .A(n7629), .B(n7628), .Z(n7633) );
  NANDN U7872 ( .A(n7631), .B(n7630), .Z(n7632) );
  AND U7873 ( .A(n7633), .B(n7632), .Z(n7664) );
  NAND U7874 ( .A(n26), .B(n7634), .Z(n7636) );
  XOR U7875 ( .A(b[7]), .B(a[184]), .Z(n7675) );
  NAND U7876 ( .A(n10531), .B(n7675), .Z(n7635) );
  AND U7877 ( .A(n7636), .B(n7635), .Z(n7694) );
  NAND U7878 ( .A(n23), .B(n7637), .Z(n7639) );
  XOR U7879 ( .A(b[3]), .B(a[188]), .Z(n7678) );
  NAND U7880 ( .A(n24), .B(n7678), .Z(n7638) );
  NAND U7881 ( .A(n7639), .B(n7638), .Z(n7693) );
  XNOR U7882 ( .A(n7694), .B(n7693), .Z(n7696) );
  NAND U7883 ( .A(b[0]), .B(a[190]), .Z(n7640) );
  XNOR U7884 ( .A(b[1]), .B(n7640), .Z(n7642) );
  NANDN U7885 ( .A(b[0]), .B(a[189]), .Z(n7641) );
  NAND U7886 ( .A(n7642), .B(n7641), .Z(n7690) );
  NAND U7887 ( .A(n25), .B(n7643), .Z(n7645) );
  XOR U7888 ( .A(b[5]), .B(a[186]), .Z(n7684) );
  NAND U7889 ( .A(n10456), .B(n7684), .Z(n7644) );
  AND U7890 ( .A(n7645), .B(n7644), .Z(n7688) );
  AND U7891 ( .A(b[7]), .B(a[182]), .Z(n7687) );
  XNOR U7892 ( .A(n7688), .B(n7687), .Z(n7689) );
  XNOR U7893 ( .A(n7690), .B(n7689), .Z(n7695) );
  XOR U7894 ( .A(n7696), .B(n7695), .Z(n7670) );
  NANDN U7895 ( .A(n7647), .B(n7646), .Z(n7651) );
  NANDN U7896 ( .A(n7649), .B(n7648), .Z(n7650) );
  AND U7897 ( .A(n7651), .B(n7650), .Z(n7669) );
  XNOR U7898 ( .A(n7670), .B(n7669), .Z(n7671) );
  NANDN U7899 ( .A(n7653), .B(n7652), .Z(n7657) );
  NAND U7900 ( .A(n7655), .B(n7654), .Z(n7656) );
  NAND U7901 ( .A(n7657), .B(n7656), .Z(n7672) );
  XNOR U7902 ( .A(n7671), .B(n7672), .Z(n7663) );
  XNOR U7903 ( .A(n7664), .B(n7663), .Z(n7665) );
  XNOR U7904 ( .A(n7666), .B(n7665), .Z(n7699) );
  XNOR U7905 ( .A(sreg[438]), .B(n7699), .Z(n7701) );
  NANDN U7906 ( .A(sreg[437]), .B(n7658), .Z(n7662) );
  NAND U7907 ( .A(n7660), .B(n7659), .Z(n7661) );
  NAND U7908 ( .A(n7662), .B(n7661), .Z(n7700) );
  XNOR U7909 ( .A(n7701), .B(n7700), .Z(c[438]) );
  NANDN U7910 ( .A(n7664), .B(n7663), .Z(n7668) );
  NANDN U7911 ( .A(n7666), .B(n7665), .Z(n7667) );
  AND U7912 ( .A(n7668), .B(n7667), .Z(n7707) );
  NANDN U7913 ( .A(n7670), .B(n7669), .Z(n7674) );
  NANDN U7914 ( .A(n7672), .B(n7671), .Z(n7673) );
  AND U7915 ( .A(n7674), .B(n7673), .Z(n7705) );
  NAND U7916 ( .A(n26), .B(n7675), .Z(n7677) );
  XOR U7917 ( .A(b[7]), .B(a[185]), .Z(n7716) );
  NAND U7918 ( .A(n10531), .B(n7716), .Z(n7676) );
  AND U7919 ( .A(n7677), .B(n7676), .Z(n7735) );
  NAND U7920 ( .A(n23), .B(n7678), .Z(n7680) );
  XOR U7921 ( .A(b[3]), .B(a[189]), .Z(n7719) );
  NAND U7922 ( .A(n24), .B(n7719), .Z(n7679) );
  NAND U7923 ( .A(n7680), .B(n7679), .Z(n7734) );
  XNOR U7924 ( .A(n7735), .B(n7734), .Z(n7737) );
  NAND U7925 ( .A(b[0]), .B(a[191]), .Z(n7681) );
  XNOR U7926 ( .A(b[1]), .B(n7681), .Z(n7683) );
  NANDN U7927 ( .A(b[0]), .B(a[190]), .Z(n7682) );
  NAND U7928 ( .A(n7683), .B(n7682), .Z(n7731) );
  NAND U7929 ( .A(n25), .B(n7684), .Z(n7686) );
  XOR U7930 ( .A(b[5]), .B(a[187]), .Z(n7725) );
  NAND U7931 ( .A(n10456), .B(n7725), .Z(n7685) );
  AND U7932 ( .A(n7686), .B(n7685), .Z(n7729) );
  AND U7933 ( .A(b[7]), .B(a[183]), .Z(n7728) );
  XNOR U7934 ( .A(n7729), .B(n7728), .Z(n7730) );
  XNOR U7935 ( .A(n7731), .B(n7730), .Z(n7736) );
  XOR U7936 ( .A(n7737), .B(n7736), .Z(n7711) );
  NANDN U7937 ( .A(n7688), .B(n7687), .Z(n7692) );
  NANDN U7938 ( .A(n7690), .B(n7689), .Z(n7691) );
  AND U7939 ( .A(n7692), .B(n7691), .Z(n7710) );
  XNOR U7940 ( .A(n7711), .B(n7710), .Z(n7712) );
  NANDN U7941 ( .A(n7694), .B(n7693), .Z(n7698) );
  NAND U7942 ( .A(n7696), .B(n7695), .Z(n7697) );
  NAND U7943 ( .A(n7698), .B(n7697), .Z(n7713) );
  XNOR U7944 ( .A(n7712), .B(n7713), .Z(n7704) );
  XNOR U7945 ( .A(n7705), .B(n7704), .Z(n7706) );
  XNOR U7946 ( .A(n7707), .B(n7706), .Z(n7740) );
  XNOR U7947 ( .A(sreg[439]), .B(n7740), .Z(n7742) );
  NANDN U7948 ( .A(sreg[438]), .B(n7699), .Z(n7703) );
  NAND U7949 ( .A(n7701), .B(n7700), .Z(n7702) );
  NAND U7950 ( .A(n7703), .B(n7702), .Z(n7741) );
  XNOR U7951 ( .A(n7742), .B(n7741), .Z(c[439]) );
  NANDN U7952 ( .A(n7705), .B(n7704), .Z(n7709) );
  NANDN U7953 ( .A(n7707), .B(n7706), .Z(n7708) );
  AND U7954 ( .A(n7709), .B(n7708), .Z(n7748) );
  NANDN U7955 ( .A(n7711), .B(n7710), .Z(n7715) );
  NANDN U7956 ( .A(n7713), .B(n7712), .Z(n7714) );
  AND U7957 ( .A(n7715), .B(n7714), .Z(n7746) );
  NAND U7958 ( .A(n26), .B(n7716), .Z(n7718) );
  XOR U7959 ( .A(b[7]), .B(a[186]), .Z(n7757) );
  NAND U7960 ( .A(n10531), .B(n7757), .Z(n7717) );
  AND U7961 ( .A(n7718), .B(n7717), .Z(n7776) );
  NAND U7962 ( .A(n23), .B(n7719), .Z(n7721) );
  XOR U7963 ( .A(b[3]), .B(a[190]), .Z(n7760) );
  NAND U7964 ( .A(n24), .B(n7760), .Z(n7720) );
  NAND U7965 ( .A(n7721), .B(n7720), .Z(n7775) );
  XNOR U7966 ( .A(n7776), .B(n7775), .Z(n7778) );
  NAND U7967 ( .A(b[0]), .B(a[192]), .Z(n7722) );
  XNOR U7968 ( .A(b[1]), .B(n7722), .Z(n7724) );
  NANDN U7969 ( .A(b[0]), .B(a[191]), .Z(n7723) );
  NAND U7970 ( .A(n7724), .B(n7723), .Z(n7772) );
  NAND U7971 ( .A(n25), .B(n7725), .Z(n7727) );
  XOR U7972 ( .A(b[5]), .B(a[188]), .Z(n7763) );
  NAND U7973 ( .A(n10456), .B(n7763), .Z(n7726) );
  AND U7974 ( .A(n7727), .B(n7726), .Z(n7770) );
  AND U7975 ( .A(b[7]), .B(a[184]), .Z(n7769) );
  XNOR U7976 ( .A(n7770), .B(n7769), .Z(n7771) );
  XNOR U7977 ( .A(n7772), .B(n7771), .Z(n7777) );
  XOR U7978 ( .A(n7778), .B(n7777), .Z(n7752) );
  NANDN U7979 ( .A(n7729), .B(n7728), .Z(n7733) );
  NANDN U7980 ( .A(n7731), .B(n7730), .Z(n7732) );
  AND U7981 ( .A(n7733), .B(n7732), .Z(n7751) );
  XNOR U7982 ( .A(n7752), .B(n7751), .Z(n7753) );
  NANDN U7983 ( .A(n7735), .B(n7734), .Z(n7739) );
  NAND U7984 ( .A(n7737), .B(n7736), .Z(n7738) );
  NAND U7985 ( .A(n7739), .B(n7738), .Z(n7754) );
  XNOR U7986 ( .A(n7753), .B(n7754), .Z(n7745) );
  XNOR U7987 ( .A(n7746), .B(n7745), .Z(n7747) );
  XNOR U7988 ( .A(n7748), .B(n7747), .Z(n7781) );
  XNOR U7989 ( .A(sreg[440]), .B(n7781), .Z(n7783) );
  NANDN U7990 ( .A(sreg[439]), .B(n7740), .Z(n7744) );
  NAND U7991 ( .A(n7742), .B(n7741), .Z(n7743) );
  NAND U7992 ( .A(n7744), .B(n7743), .Z(n7782) );
  XNOR U7993 ( .A(n7783), .B(n7782), .Z(c[440]) );
  NANDN U7994 ( .A(n7746), .B(n7745), .Z(n7750) );
  NANDN U7995 ( .A(n7748), .B(n7747), .Z(n7749) );
  AND U7996 ( .A(n7750), .B(n7749), .Z(n7789) );
  NANDN U7997 ( .A(n7752), .B(n7751), .Z(n7756) );
  NANDN U7998 ( .A(n7754), .B(n7753), .Z(n7755) );
  AND U7999 ( .A(n7756), .B(n7755), .Z(n7787) );
  NAND U8000 ( .A(n26), .B(n7757), .Z(n7759) );
  XOR U8001 ( .A(b[7]), .B(a[187]), .Z(n7798) );
  NAND U8002 ( .A(n10531), .B(n7798), .Z(n7758) );
  AND U8003 ( .A(n7759), .B(n7758), .Z(n7817) );
  NAND U8004 ( .A(n23), .B(n7760), .Z(n7762) );
  XOR U8005 ( .A(b[3]), .B(a[191]), .Z(n7801) );
  NAND U8006 ( .A(n24), .B(n7801), .Z(n7761) );
  NAND U8007 ( .A(n7762), .B(n7761), .Z(n7816) );
  XNOR U8008 ( .A(n7817), .B(n7816), .Z(n7819) );
  NAND U8009 ( .A(n25), .B(n7763), .Z(n7765) );
  XOR U8010 ( .A(b[5]), .B(a[189]), .Z(n7807) );
  NAND U8011 ( .A(n10456), .B(n7807), .Z(n7764) );
  AND U8012 ( .A(n7765), .B(n7764), .Z(n7811) );
  AND U8013 ( .A(b[7]), .B(a[185]), .Z(n7810) );
  XNOR U8014 ( .A(n7811), .B(n7810), .Z(n7812) );
  NAND U8015 ( .A(b[0]), .B(a[193]), .Z(n7766) );
  XNOR U8016 ( .A(b[1]), .B(n7766), .Z(n7768) );
  NANDN U8017 ( .A(b[0]), .B(a[192]), .Z(n7767) );
  NAND U8018 ( .A(n7768), .B(n7767), .Z(n7813) );
  XNOR U8019 ( .A(n7812), .B(n7813), .Z(n7818) );
  XOR U8020 ( .A(n7819), .B(n7818), .Z(n7793) );
  NANDN U8021 ( .A(n7770), .B(n7769), .Z(n7774) );
  NANDN U8022 ( .A(n7772), .B(n7771), .Z(n7773) );
  AND U8023 ( .A(n7774), .B(n7773), .Z(n7792) );
  XNOR U8024 ( .A(n7793), .B(n7792), .Z(n7794) );
  NANDN U8025 ( .A(n7776), .B(n7775), .Z(n7780) );
  NAND U8026 ( .A(n7778), .B(n7777), .Z(n7779) );
  NAND U8027 ( .A(n7780), .B(n7779), .Z(n7795) );
  XNOR U8028 ( .A(n7794), .B(n7795), .Z(n7786) );
  XNOR U8029 ( .A(n7787), .B(n7786), .Z(n7788) );
  XNOR U8030 ( .A(n7789), .B(n7788), .Z(n7822) );
  XNOR U8031 ( .A(sreg[441]), .B(n7822), .Z(n7824) );
  NANDN U8032 ( .A(sreg[440]), .B(n7781), .Z(n7785) );
  NAND U8033 ( .A(n7783), .B(n7782), .Z(n7784) );
  NAND U8034 ( .A(n7785), .B(n7784), .Z(n7823) );
  XNOR U8035 ( .A(n7824), .B(n7823), .Z(c[441]) );
  NANDN U8036 ( .A(n7787), .B(n7786), .Z(n7791) );
  NANDN U8037 ( .A(n7789), .B(n7788), .Z(n7790) );
  AND U8038 ( .A(n7791), .B(n7790), .Z(n7830) );
  NANDN U8039 ( .A(n7793), .B(n7792), .Z(n7797) );
  NANDN U8040 ( .A(n7795), .B(n7794), .Z(n7796) );
  AND U8041 ( .A(n7797), .B(n7796), .Z(n7828) );
  NAND U8042 ( .A(n26), .B(n7798), .Z(n7800) );
  XOR U8043 ( .A(b[7]), .B(a[188]), .Z(n7839) );
  NAND U8044 ( .A(n10531), .B(n7839), .Z(n7799) );
  AND U8045 ( .A(n7800), .B(n7799), .Z(n7858) );
  NAND U8046 ( .A(n23), .B(n7801), .Z(n7803) );
  XOR U8047 ( .A(b[3]), .B(a[192]), .Z(n7842) );
  NAND U8048 ( .A(n24), .B(n7842), .Z(n7802) );
  NAND U8049 ( .A(n7803), .B(n7802), .Z(n7857) );
  XNOR U8050 ( .A(n7858), .B(n7857), .Z(n7860) );
  NAND U8051 ( .A(b[0]), .B(a[194]), .Z(n7804) );
  XNOR U8052 ( .A(b[1]), .B(n7804), .Z(n7806) );
  NANDN U8053 ( .A(b[0]), .B(a[193]), .Z(n7805) );
  NAND U8054 ( .A(n7806), .B(n7805), .Z(n7854) );
  NAND U8055 ( .A(n25), .B(n7807), .Z(n7809) );
  XOR U8056 ( .A(b[5]), .B(a[190]), .Z(n7848) );
  NAND U8057 ( .A(n10456), .B(n7848), .Z(n7808) );
  AND U8058 ( .A(n7809), .B(n7808), .Z(n7852) );
  AND U8059 ( .A(b[7]), .B(a[186]), .Z(n7851) );
  XNOR U8060 ( .A(n7852), .B(n7851), .Z(n7853) );
  XNOR U8061 ( .A(n7854), .B(n7853), .Z(n7859) );
  XOR U8062 ( .A(n7860), .B(n7859), .Z(n7834) );
  NANDN U8063 ( .A(n7811), .B(n7810), .Z(n7815) );
  NANDN U8064 ( .A(n7813), .B(n7812), .Z(n7814) );
  AND U8065 ( .A(n7815), .B(n7814), .Z(n7833) );
  XNOR U8066 ( .A(n7834), .B(n7833), .Z(n7835) );
  NANDN U8067 ( .A(n7817), .B(n7816), .Z(n7821) );
  NAND U8068 ( .A(n7819), .B(n7818), .Z(n7820) );
  NAND U8069 ( .A(n7821), .B(n7820), .Z(n7836) );
  XNOR U8070 ( .A(n7835), .B(n7836), .Z(n7827) );
  XNOR U8071 ( .A(n7828), .B(n7827), .Z(n7829) );
  XNOR U8072 ( .A(n7830), .B(n7829), .Z(n7863) );
  XNOR U8073 ( .A(sreg[442]), .B(n7863), .Z(n7865) );
  NANDN U8074 ( .A(sreg[441]), .B(n7822), .Z(n7826) );
  NAND U8075 ( .A(n7824), .B(n7823), .Z(n7825) );
  NAND U8076 ( .A(n7826), .B(n7825), .Z(n7864) );
  XNOR U8077 ( .A(n7865), .B(n7864), .Z(c[442]) );
  NANDN U8078 ( .A(n7828), .B(n7827), .Z(n7832) );
  NANDN U8079 ( .A(n7830), .B(n7829), .Z(n7831) );
  AND U8080 ( .A(n7832), .B(n7831), .Z(n7871) );
  NANDN U8081 ( .A(n7834), .B(n7833), .Z(n7838) );
  NANDN U8082 ( .A(n7836), .B(n7835), .Z(n7837) );
  AND U8083 ( .A(n7838), .B(n7837), .Z(n7869) );
  NAND U8084 ( .A(n26), .B(n7839), .Z(n7841) );
  XOR U8085 ( .A(b[7]), .B(a[189]), .Z(n7880) );
  NAND U8086 ( .A(n10531), .B(n7880), .Z(n7840) );
  AND U8087 ( .A(n7841), .B(n7840), .Z(n7899) );
  NAND U8088 ( .A(n23), .B(n7842), .Z(n7844) );
  XOR U8089 ( .A(b[3]), .B(a[193]), .Z(n7883) );
  NAND U8090 ( .A(n24), .B(n7883), .Z(n7843) );
  NAND U8091 ( .A(n7844), .B(n7843), .Z(n7898) );
  XNOR U8092 ( .A(n7899), .B(n7898), .Z(n7901) );
  NAND U8093 ( .A(b[0]), .B(a[195]), .Z(n7845) );
  XNOR U8094 ( .A(b[1]), .B(n7845), .Z(n7847) );
  NANDN U8095 ( .A(b[0]), .B(a[194]), .Z(n7846) );
  NAND U8096 ( .A(n7847), .B(n7846), .Z(n7895) );
  NAND U8097 ( .A(n25), .B(n7848), .Z(n7850) );
  XOR U8098 ( .A(b[5]), .B(a[191]), .Z(n7889) );
  NAND U8099 ( .A(n10456), .B(n7889), .Z(n7849) );
  AND U8100 ( .A(n7850), .B(n7849), .Z(n7893) );
  AND U8101 ( .A(b[7]), .B(a[187]), .Z(n7892) );
  XNOR U8102 ( .A(n7893), .B(n7892), .Z(n7894) );
  XNOR U8103 ( .A(n7895), .B(n7894), .Z(n7900) );
  XOR U8104 ( .A(n7901), .B(n7900), .Z(n7875) );
  NANDN U8105 ( .A(n7852), .B(n7851), .Z(n7856) );
  NANDN U8106 ( .A(n7854), .B(n7853), .Z(n7855) );
  AND U8107 ( .A(n7856), .B(n7855), .Z(n7874) );
  XNOR U8108 ( .A(n7875), .B(n7874), .Z(n7876) );
  NANDN U8109 ( .A(n7858), .B(n7857), .Z(n7862) );
  NAND U8110 ( .A(n7860), .B(n7859), .Z(n7861) );
  NAND U8111 ( .A(n7862), .B(n7861), .Z(n7877) );
  XNOR U8112 ( .A(n7876), .B(n7877), .Z(n7868) );
  XNOR U8113 ( .A(n7869), .B(n7868), .Z(n7870) );
  XNOR U8114 ( .A(n7871), .B(n7870), .Z(n7904) );
  XNOR U8115 ( .A(sreg[443]), .B(n7904), .Z(n7906) );
  NANDN U8116 ( .A(sreg[442]), .B(n7863), .Z(n7867) );
  NAND U8117 ( .A(n7865), .B(n7864), .Z(n7866) );
  NAND U8118 ( .A(n7867), .B(n7866), .Z(n7905) );
  XNOR U8119 ( .A(n7906), .B(n7905), .Z(c[443]) );
  NANDN U8120 ( .A(n7869), .B(n7868), .Z(n7873) );
  NANDN U8121 ( .A(n7871), .B(n7870), .Z(n7872) );
  AND U8122 ( .A(n7873), .B(n7872), .Z(n7912) );
  NANDN U8123 ( .A(n7875), .B(n7874), .Z(n7879) );
  NANDN U8124 ( .A(n7877), .B(n7876), .Z(n7878) );
  AND U8125 ( .A(n7879), .B(n7878), .Z(n7910) );
  NAND U8126 ( .A(n26), .B(n7880), .Z(n7882) );
  XOR U8127 ( .A(b[7]), .B(a[190]), .Z(n7921) );
  NAND U8128 ( .A(n10531), .B(n7921), .Z(n7881) );
  AND U8129 ( .A(n7882), .B(n7881), .Z(n7940) );
  NAND U8130 ( .A(n23), .B(n7883), .Z(n7885) );
  XOR U8131 ( .A(b[3]), .B(a[194]), .Z(n7924) );
  NAND U8132 ( .A(n24), .B(n7924), .Z(n7884) );
  NAND U8133 ( .A(n7885), .B(n7884), .Z(n7939) );
  XNOR U8134 ( .A(n7940), .B(n7939), .Z(n7942) );
  NAND U8135 ( .A(b[0]), .B(a[196]), .Z(n7886) );
  XNOR U8136 ( .A(b[1]), .B(n7886), .Z(n7888) );
  NANDN U8137 ( .A(b[0]), .B(a[195]), .Z(n7887) );
  NAND U8138 ( .A(n7888), .B(n7887), .Z(n7936) );
  NAND U8139 ( .A(n25), .B(n7889), .Z(n7891) );
  XOR U8140 ( .A(b[5]), .B(a[192]), .Z(n7930) );
  NAND U8141 ( .A(n10456), .B(n7930), .Z(n7890) );
  AND U8142 ( .A(n7891), .B(n7890), .Z(n7934) );
  AND U8143 ( .A(b[7]), .B(a[188]), .Z(n7933) );
  XNOR U8144 ( .A(n7934), .B(n7933), .Z(n7935) );
  XNOR U8145 ( .A(n7936), .B(n7935), .Z(n7941) );
  XOR U8146 ( .A(n7942), .B(n7941), .Z(n7916) );
  NANDN U8147 ( .A(n7893), .B(n7892), .Z(n7897) );
  NANDN U8148 ( .A(n7895), .B(n7894), .Z(n7896) );
  AND U8149 ( .A(n7897), .B(n7896), .Z(n7915) );
  XNOR U8150 ( .A(n7916), .B(n7915), .Z(n7917) );
  NANDN U8151 ( .A(n7899), .B(n7898), .Z(n7903) );
  NAND U8152 ( .A(n7901), .B(n7900), .Z(n7902) );
  NAND U8153 ( .A(n7903), .B(n7902), .Z(n7918) );
  XNOR U8154 ( .A(n7917), .B(n7918), .Z(n7909) );
  XNOR U8155 ( .A(n7910), .B(n7909), .Z(n7911) );
  XNOR U8156 ( .A(n7912), .B(n7911), .Z(n7945) );
  XNOR U8157 ( .A(sreg[444]), .B(n7945), .Z(n7947) );
  NANDN U8158 ( .A(sreg[443]), .B(n7904), .Z(n7908) );
  NAND U8159 ( .A(n7906), .B(n7905), .Z(n7907) );
  NAND U8160 ( .A(n7908), .B(n7907), .Z(n7946) );
  XNOR U8161 ( .A(n7947), .B(n7946), .Z(c[444]) );
  NANDN U8162 ( .A(n7910), .B(n7909), .Z(n7914) );
  NANDN U8163 ( .A(n7912), .B(n7911), .Z(n7913) );
  AND U8164 ( .A(n7914), .B(n7913), .Z(n7953) );
  NANDN U8165 ( .A(n7916), .B(n7915), .Z(n7920) );
  NANDN U8166 ( .A(n7918), .B(n7917), .Z(n7919) );
  AND U8167 ( .A(n7920), .B(n7919), .Z(n7951) );
  NAND U8168 ( .A(n26), .B(n7921), .Z(n7923) );
  XOR U8169 ( .A(b[7]), .B(a[191]), .Z(n7962) );
  NAND U8170 ( .A(n10531), .B(n7962), .Z(n7922) );
  AND U8171 ( .A(n7923), .B(n7922), .Z(n7981) );
  NAND U8172 ( .A(n23), .B(n7924), .Z(n7926) );
  XOR U8173 ( .A(b[3]), .B(a[195]), .Z(n7965) );
  NAND U8174 ( .A(n24), .B(n7965), .Z(n7925) );
  NAND U8175 ( .A(n7926), .B(n7925), .Z(n7980) );
  XNOR U8176 ( .A(n7981), .B(n7980), .Z(n7983) );
  NAND U8177 ( .A(b[0]), .B(a[197]), .Z(n7927) );
  XNOR U8178 ( .A(b[1]), .B(n7927), .Z(n7929) );
  NANDN U8179 ( .A(b[0]), .B(a[196]), .Z(n7928) );
  NAND U8180 ( .A(n7929), .B(n7928), .Z(n7977) );
  NAND U8181 ( .A(n25), .B(n7930), .Z(n7932) );
  XOR U8182 ( .A(b[5]), .B(a[193]), .Z(n7971) );
  NAND U8183 ( .A(n10456), .B(n7971), .Z(n7931) );
  AND U8184 ( .A(n7932), .B(n7931), .Z(n7975) );
  AND U8185 ( .A(b[7]), .B(a[189]), .Z(n7974) );
  XNOR U8186 ( .A(n7975), .B(n7974), .Z(n7976) );
  XNOR U8187 ( .A(n7977), .B(n7976), .Z(n7982) );
  XOR U8188 ( .A(n7983), .B(n7982), .Z(n7957) );
  NANDN U8189 ( .A(n7934), .B(n7933), .Z(n7938) );
  NANDN U8190 ( .A(n7936), .B(n7935), .Z(n7937) );
  AND U8191 ( .A(n7938), .B(n7937), .Z(n7956) );
  XNOR U8192 ( .A(n7957), .B(n7956), .Z(n7958) );
  NANDN U8193 ( .A(n7940), .B(n7939), .Z(n7944) );
  NAND U8194 ( .A(n7942), .B(n7941), .Z(n7943) );
  NAND U8195 ( .A(n7944), .B(n7943), .Z(n7959) );
  XNOR U8196 ( .A(n7958), .B(n7959), .Z(n7950) );
  XNOR U8197 ( .A(n7951), .B(n7950), .Z(n7952) );
  XNOR U8198 ( .A(n7953), .B(n7952), .Z(n7986) );
  XNOR U8199 ( .A(sreg[445]), .B(n7986), .Z(n7988) );
  NANDN U8200 ( .A(sreg[444]), .B(n7945), .Z(n7949) );
  NAND U8201 ( .A(n7947), .B(n7946), .Z(n7948) );
  NAND U8202 ( .A(n7949), .B(n7948), .Z(n7987) );
  XNOR U8203 ( .A(n7988), .B(n7987), .Z(c[445]) );
  NANDN U8204 ( .A(n7951), .B(n7950), .Z(n7955) );
  NANDN U8205 ( .A(n7953), .B(n7952), .Z(n7954) );
  AND U8206 ( .A(n7955), .B(n7954), .Z(n7994) );
  NANDN U8207 ( .A(n7957), .B(n7956), .Z(n7961) );
  NANDN U8208 ( .A(n7959), .B(n7958), .Z(n7960) );
  AND U8209 ( .A(n7961), .B(n7960), .Z(n7992) );
  NAND U8210 ( .A(n26), .B(n7962), .Z(n7964) );
  XOR U8211 ( .A(b[7]), .B(a[192]), .Z(n8003) );
  NAND U8212 ( .A(n10531), .B(n8003), .Z(n7963) );
  AND U8213 ( .A(n7964), .B(n7963), .Z(n8022) );
  NAND U8214 ( .A(n23), .B(n7965), .Z(n7967) );
  XOR U8215 ( .A(b[3]), .B(a[196]), .Z(n8006) );
  NAND U8216 ( .A(n24), .B(n8006), .Z(n7966) );
  NAND U8217 ( .A(n7967), .B(n7966), .Z(n8021) );
  XNOR U8218 ( .A(n8022), .B(n8021), .Z(n8024) );
  NAND U8219 ( .A(b[0]), .B(a[198]), .Z(n7968) );
  XNOR U8220 ( .A(b[1]), .B(n7968), .Z(n7970) );
  NANDN U8221 ( .A(b[0]), .B(a[197]), .Z(n7969) );
  NAND U8222 ( .A(n7970), .B(n7969), .Z(n8018) );
  NAND U8223 ( .A(n25), .B(n7971), .Z(n7973) );
  XOR U8224 ( .A(b[5]), .B(a[194]), .Z(n8012) );
  NAND U8225 ( .A(n10456), .B(n8012), .Z(n7972) );
  AND U8226 ( .A(n7973), .B(n7972), .Z(n8016) );
  AND U8227 ( .A(b[7]), .B(a[190]), .Z(n8015) );
  XNOR U8228 ( .A(n8016), .B(n8015), .Z(n8017) );
  XNOR U8229 ( .A(n8018), .B(n8017), .Z(n8023) );
  XOR U8230 ( .A(n8024), .B(n8023), .Z(n7998) );
  NANDN U8231 ( .A(n7975), .B(n7974), .Z(n7979) );
  NANDN U8232 ( .A(n7977), .B(n7976), .Z(n7978) );
  AND U8233 ( .A(n7979), .B(n7978), .Z(n7997) );
  XNOR U8234 ( .A(n7998), .B(n7997), .Z(n7999) );
  NANDN U8235 ( .A(n7981), .B(n7980), .Z(n7985) );
  NAND U8236 ( .A(n7983), .B(n7982), .Z(n7984) );
  NAND U8237 ( .A(n7985), .B(n7984), .Z(n8000) );
  XNOR U8238 ( .A(n7999), .B(n8000), .Z(n7991) );
  XNOR U8239 ( .A(n7992), .B(n7991), .Z(n7993) );
  XNOR U8240 ( .A(n7994), .B(n7993), .Z(n8027) );
  XNOR U8241 ( .A(sreg[446]), .B(n8027), .Z(n8029) );
  NANDN U8242 ( .A(sreg[445]), .B(n7986), .Z(n7990) );
  NAND U8243 ( .A(n7988), .B(n7987), .Z(n7989) );
  NAND U8244 ( .A(n7990), .B(n7989), .Z(n8028) );
  XNOR U8245 ( .A(n8029), .B(n8028), .Z(c[446]) );
  NANDN U8246 ( .A(n7992), .B(n7991), .Z(n7996) );
  NANDN U8247 ( .A(n7994), .B(n7993), .Z(n7995) );
  AND U8248 ( .A(n7996), .B(n7995), .Z(n8035) );
  NANDN U8249 ( .A(n7998), .B(n7997), .Z(n8002) );
  NANDN U8250 ( .A(n8000), .B(n7999), .Z(n8001) );
  AND U8251 ( .A(n8002), .B(n8001), .Z(n8033) );
  NAND U8252 ( .A(n26), .B(n8003), .Z(n8005) );
  XOR U8253 ( .A(b[7]), .B(a[193]), .Z(n8044) );
  NAND U8254 ( .A(n10531), .B(n8044), .Z(n8004) );
  AND U8255 ( .A(n8005), .B(n8004), .Z(n8063) );
  NAND U8256 ( .A(n23), .B(n8006), .Z(n8008) );
  XOR U8257 ( .A(b[3]), .B(a[197]), .Z(n8047) );
  NAND U8258 ( .A(n24), .B(n8047), .Z(n8007) );
  NAND U8259 ( .A(n8008), .B(n8007), .Z(n8062) );
  XNOR U8260 ( .A(n8063), .B(n8062), .Z(n8065) );
  NAND U8261 ( .A(b[0]), .B(a[199]), .Z(n8009) );
  XNOR U8262 ( .A(b[1]), .B(n8009), .Z(n8011) );
  NANDN U8263 ( .A(b[0]), .B(a[198]), .Z(n8010) );
  NAND U8264 ( .A(n8011), .B(n8010), .Z(n8059) );
  NAND U8265 ( .A(n25), .B(n8012), .Z(n8014) );
  XOR U8266 ( .A(b[5]), .B(a[195]), .Z(n8050) );
  NAND U8267 ( .A(n10456), .B(n8050), .Z(n8013) );
  AND U8268 ( .A(n8014), .B(n8013), .Z(n8057) );
  AND U8269 ( .A(b[7]), .B(a[191]), .Z(n8056) );
  XNOR U8270 ( .A(n8057), .B(n8056), .Z(n8058) );
  XNOR U8271 ( .A(n8059), .B(n8058), .Z(n8064) );
  XOR U8272 ( .A(n8065), .B(n8064), .Z(n8039) );
  NANDN U8273 ( .A(n8016), .B(n8015), .Z(n8020) );
  NANDN U8274 ( .A(n8018), .B(n8017), .Z(n8019) );
  AND U8275 ( .A(n8020), .B(n8019), .Z(n8038) );
  XNOR U8276 ( .A(n8039), .B(n8038), .Z(n8040) );
  NANDN U8277 ( .A(n8022), .B(n8021), .Z(n8026) );
  NAND U8278 ( .A(n8024), .B(n8023), .Z(n8025) );
  NAND U8279 ( .A(n8026), .B(n8025), .Z(n8041) );
  XNOR U8280 ( .A(n8040), .B(n8041), .Z(n8032) );
  XNOR U8281 ( .A(n8033), .B(n8032), .Z(n8034) );
  XNOR U8282 ( .A(n8035), .B(n8034), .Z(n8068) );
  XNOR U8283 ( .A(sreg[447]), .B(n8068), .Z(n8070) );
  NANDN U8284 ( .A(sreg[446]), .B(n8027), .Z(n8031) );
  NAND U8285 ( .A(n8029), .B(n8028), .Z(n8030) );
  NAND U8286 ( .A(n8031), .B(n8030), .Z(n8069) );
  XNOR U8287 ( .A(n8070), .B(n8069), .Z(c[447]) );
  NANDN U8288 ( .A(n8033), .B(n8032), .Z(n8037) );
  NANDN U8289 ( .A(n8035), .B(n8034), .Z(n8036) );
  AND U8290 ( .A(n8037), .B(n8036), .Z(n8076) );
  NANDN U8291 ( .A(n8039), .B(n8038), .Z(n8043) );
  NANDN U8292 ( .A(n8041), .B(n8040), .Z(n8042) );
  AND U8293 ( .A(n8043), .B(n8042), .Z(n8074) );
  NAND U8294 ( .A(n26), .B(n8044), .Z(n8046) );
  XOR U8295 ( .A(b[7]), .B(a[194]), .Z(n8085) );
  NAND U8296 ( .A(n10531), .B(n8085), .Z(n8045) );
  AND U8297 ( .A(n8046), .B(n8045), .Z(n8104) );
  NAND U8298 ( .A(n23), .B(n8047), .Z(n8049) );
  XOR U8299 ( .A(b[3]), .B(a[198]), .Z(n8088) );
  NAND U8300 ( .A(n24), .B(n8088), .Z(n8048) );
  NAND U8301 ( .A(n8049), .B(n8048), .Z(n8103) );
  XNOR U8302 ( .A(n8104), .B(n8103), .Z(n8106) );
  NAND U8303 ( .A(n25), .B(n8050), .Z(n8052) );
  XOR U8304 ( .A(b[5]), .B(a[196]), .Z(n8094) );
  NAND U8305 ( .A(n10456), .B(n8094), .Z(n8051) );
  AND U8306 ( .A(n8052), .B(n8051), .Z(n8098) );
  AND U8307 ( .A(b[7]), .B(a[192]), .Z(n8097) );
  XNOR U8308 ( .A(n8098), .B(n8097), .Z(n8099) );
  NAND U8309 ( .A(b[0]), .B(a[200]), .Z(n8053) );
  XNOR U8310 ( .A(b[1]), .B(n8053), .Z(n8055) );
  NANDN U8311 ( .A(b[0]), .B(a[199]), .Z(n8054) );
  NAND U8312 ( .A(n8055), .B(n8054), .Z(n8100) );
  XNOR U8313 ( .A(n8099), .B(n8100), .Z(n8105) );
  XOR U8314 ( .A(n8106), .B(n8105), .Z(n8080) );
  NANDN U8315 ( .A(n8057), .B(n8056), .Z(n8061) );
  NANDN U8316 ( .A(n8059), .B(n8058), .Z(n8060) );
  AND U8317 ( .A(n8061), .B(n8060), .Z(n8079) );
  XNOR U8318 ( .A(n8080), .B(n8079), .Z(n8081) );
  NANDN U8319 ( .A(n8063), .B(n8062), .Z(n8067) );
  NAND U8320 ( .A(n8065), .B(n8064), .Z(n8066) );
  NAND U8321 ( .A(n8067), .B(n8066), .Z(n8082) );
  XNOR U8322 ( .A(n8081), .B(n8082), .Z(n8073) );
  XNOR U8323 ( .A(n8074), .B(n8073), .Z(n8075) );
  XNOR U8324 ( .A(n8076), .B(n8075), .Z(n8109) );
  XNOR U8325 ( .A(sreg[448]), .B(n8109), .Z(n8111) );
  NANDN U8326 ( .A(sreg[447]), .B(n8068), .Z(n8072) );
  NAND U8327 ( .A(n8070), .B(n8069), .Z(n8071) );
  NAND U8328 ( .A(n8072), .B(n8071), .Z(n8110) );
  XNOR U8329 ( .A(n8111), .B(n8110), .Z(c[448]) );
  NANDN U8330 ( .A(n8074), .B(n8073), .Z(n8078) );
  NANDN U8331 ( .A(n8076), .B(n8075), .Z(n8077) );
  AND U8332 ( .A(n8078), .B(n8077), .Z(n8117) );
  NANDN U8333 ( .A(n8080), .B(n8079), .Z(n8084) );
  NANDN U8334 ( .A(n8082), .B(n8081), .Z(n8083) );
  AND U8335 ( .A(n8084), .B(n8083), .Z(n8115) );
  NAND U8336 ( .A(n26), .B(n8085), .Z(n8087) );
  XOR U8337 ( .A(b[7]), .B(a[195]), .Z(n8126) );
  NAND U8338 ( .A(n10531), .B(n8126), .Z(n8086) );
  AND U8339 ( .A(n8087), .B(n8086), .Z(n8145) );
  NAND U8340 ( .A(n23), .B(n8088), .Z(n8090) );
  XOR U8341 ( .A(b[3]), .B(a[199]), .Z(n8129) );
  NAND U8342 ( .A(n24), .B(n8129), .Z(n8089) );
  NAND U8343 ( .A(n8090), .B(n8089), .Z(n8144) );
  XNOR U8344 ( .A(n8145), .B(n8144), .Z(n8147) );
  NAND U8345 ( .A(b[0]), .B(a[201]), .Z(n8091) );
  XNOR U8346 ( .A(b[1]), .B(n8091), .Z(n8093) );
  NANDN U8347 ( .A(b[0]), .B(a[200]), .Z(n8092) );
  NAND U8348 ( .A(n8093), .B(n8092), .Z(n8141) );
  NAND U8349 ( .A(n25), .B(n8094), .Z(n8096) );
  XOR U8350 ( .A(b[5]), .B(a[197]), .Z(n8135) );
  NAND U8351 ( .A(n10456), .B(n8135), .Z(n8095) );
  AND U8352 ( .A(n8096), .B(n8095), .Z(n8139) );
  AND U8353 ( .A(b[7]), .B(a[193]), .Z(n8138) );
  XNOR U8354 ( .A(n8139), .B(n8138), .Z(n8140) );
  XNOR U8355 ( .A(n8141), .B(n8140), .Z(n8146) );
  XOR U8356 ( .A(n8147), .B(n8146), .Z(n8121) );
  NANDN U8357 ( .A(n8098), .B(n8097), .Z(n8102) );
  NANDN U8358 ( .A(n8100), .B(n8099), .Z(n8101) );
  AND U8359 ( .A(n8102), .B(n8101), .Z(n8120) );
  XNOR U8360 ( .A(n8121), .B(n8120), .Z(n8122) );
  NANDN U8361 ( .A(n8104), .B(n8103), .Z(n8108) );
  NAND U8362 ( .A(n8106), .B(n8105), .Z(n8107) );
  NAND U8363 ( .A(n8108), .B(n8107), .Z(n8123) );
  XNOR U8364 ( .A(n8122), .B(n8123), .Z(n8114) );
  XNOR U8365 ( .A(n8115), .B(n8114), .Z(n8116) );
  XNOR U8366 ( .A(n8117), .B(n8116), .Z(n8150) );
  XNOR U8367 ( .A(sreg[449]), .B(n8150), .Z(n8152) );
  NANDN U8368 ( .A(sreg[448]), .B(n8109), .Z(n8113) );
  NAND U8369 ( .A(n8111), .B(n8110), .Z(n8112) );
  NAND U8370 ( .A(n8113), .B(n8112), .Z(n8151) );
  XNOR U8371 ( .A(n8152), .B(n8151), .Z(c[449]) );
  NANDN U8372 ( .A(n8115), .B(n8114), .Z(n8119) );
  NANDN U8373 ( .A(n8117), .B(n8116), .Z(n8118) );
  AND U8374 ( .A(n8119), .B(n8118), .Z(n8158) );
  NANDN U8375 ( .A(n8121), .B(n8120), .Z(n8125) );
  NANDN U8376 ( .A(n8123), .B(n8122), .Z(n8124) );
  AND U8377 ( .A(n8125), .B(n8124), .Z(n8156) );
  NAND U8378 ( .A(n26), .B(n8126), .Z(n8128) );
  XOR U8379 ( .A(b[7]), .B(a[196]), .Z(n8167) );
  NAND U8380 ( .A(n10531), .B(n8167), .Z(n8127) );
  AND U8381 ( .A(n8128), .B(n8127), .Z(n8186) );
  NAND U8382 ( .A(n23), .B(n8129), .Z(n8131) );
  XOR U8383 ( .A(b[3]), .B(a[200]), .Z(n8170) );
  NAND U8384 ( .A(n24), .B(n8170), .Z(n8130) );
  NAND U8385 ( .A(n8131), .B(n8130), .Z(n8185) );
  XNOR U8386 ( .A(n8186), .B(n8185), .Z(n8188) );
  NAND U8387 ( .A(b[0]), .B(a[202]), .Z(n8132) );
  XNOR U8388 ( .A(b[1]), .B(n8132), .Z(n8134) );
  NANDN U8389 ( .A(b[0]), .B(a[201]), .Z(n8133) );
  NAND U8390 ( .A(n8134), .B(n8133), .Z(n8182) );
  NAND U8391 ( .A(n25), .B(n8135), .Z(n8137) );
  XOR U8392 ( .A(b[5]), .B(a[198]), .Z(n8176) );
  NAND U8393 ( .A(n10456), .B(n8176), .Z(n8136) );
  AND U8394 ( .A(n8137), .B(n8136), .Z(n8180) );
  AND U8395 ( .A(b[7]), .B(a[194]), .Z(n8179) );
  XNOR U8396 ( .A(n8180), .B(n8179), .Z(n8181) );
  XNOR U8397 ( .A(n8182), .B(n8181), .Z(n8187) );
  XOR U8398 ( .A(n8188), .B(n8187), .Z(n8162) );
  NANDN U8399 ( .A(n8139), .B(n8138), .Z(n8143) );
  NANDN U8400 ( .A(n8141), .B(n8140), .Z(n8142) );
  AND U8401 ( .A(n8143), .B(n8142), .Z(n8161) );
  XNOR U8402 ( .A(n8162), .B(n8161), .Z(n8163) );
  NANDN U8403 ( .A(n8145), .B(n8144), .Z(n8149) );
  NAND U8404 ( .A(n8147), .B(n8146), .Z(n8148) );
  NAND U8405 ( .A(n8149), .B(n8148), .Z(n8164) );
  XNOR U8406 ( .A(n8163), .B(n8164), .Z(n8155) );
  XNOR U8407 ( .A(n8156), .B(n8155), .Z(n8157) );
  XNOR U8408 ( .A(n8158), .B(n8157), .Z(n8191) );
  XNOR U8409 ( .A(sreg[450]), .B(n8191), .Z(n8193) );
  NANDN U8410 ( .A(sreg[449]), .B(n8150), .Z(n8154) );
  NAND U8411 ( .A(n8152), .B(n8151), .Z(n8153) );
  NAND U8412 ( .A(n8154), .B(n8153), .Z(n8192) );
  XNOR U8413 ( .A(n8193), .B(n8192), .Z(c[450]) );
  NANDN U8414 ( .A(n8156), .B(n8155), .Z(n8160) );
  NANDN U8415 ( .A(n8158), .B(n8157), .Z(n8159) );
  AND U8416 ( .A(n8160), .B(n8159), .Z(n8199) );
  NANDN U8417 ( .A(n8162), .B(n8161), .Z(n8166) );
  NANDN U8418 ( .A(n8164), .B(n8163), .Z(n8165) );
  AND U8419 ( .A(n8166), .B(n8165), .Z(n8197) );
  NAND U8420 ( .A(n26), .B(n8167), .Z(n8169) );
  XOR U8421 ( .A(b[7]), .B(a[197]), .Z(n8208) );
  NAND U8422 ( .A(n10531), .B(n8208), .Z(n8168) );
  AND U8423 ( .A(n8169), .B(n8168), .Z(n8227) );
  NAND U8424 ( .A(n23), .B(n8170), .Z(n8172) );
  XOR U8425 ( .A(b[3]), .B(a[201]), .Z(n8211) );
  NAND U8426 ( .A(n24), .B(n8211), .Z(n8171) );
  NAND U8427 ( .A(n8172), .B(n8171), .Z(n8226) );
  XNOR U8428 ( .A(n8227), .B(n8226), .Z(n8229) );
  NAND U8429 ( .A(b[0]), .B(a[203]), .Z(n8173) );
  XNOR U8430 ( .A(b[1]), .B(n8173), .Z(n8175) );
  NANDN U8431 ( .A(b[0]), .B(a[202]), .Z(n8174) );
  NAND U8432 ( .A(n8175), .B(n8174), .Z(n8223) );
  NAND U8433 ( .A(n25), .B(n8176), .Z(n8178) );
  XOR U8434 ( .A(b[5]), .B(a[199]), .Z(n8217) );
  NAND U8435 ( .A(n10456), .B(n8217), .Z(n8177) );
  AND U8436 ( .A(n8178), .B(n8177), .Z(n8221) );
  AND U8437 ( .A(b[7]), .B(a[195]), .Z(n8220) );
  XNOR U8438 ( .A(n8221), .B(n8220), .Z(n8222) );
  XNOR U8439 ( .A(n8223), .B(n8222), .Z(n8228) );
  XOR U8440 ( .A(n8229), .B(n8228), .Z(n8203) );
  NANDN U8441 ( .A(n8180), .B(n8179), .Z(n8184) );
  NANDN U8442 ( .A(n8182), .B(n8181), .Z(n8183) );
  AND U8443 ( .A(n8184), .B(n8183), .Z(n8202) );
  XNOR U8444 ( .A(n8203), .B(n8202), .Z(n8204) );
  NANDN U8445 ( .A(n8186), .B(n8185), .Z(n8190) );
  NAND U8446 ( .A(n8188), .B(n8187), .Z(n8189) );
  NAND U8447 ( .A(n8190), .B(n8189), .Z(n8205) );
  XNOR U8448 ( .A(n8204), .B(n8205), .Z(n8196) );
  XNOR U8449 ( .A(n8197), .B(n8196), .Z(n8198) );
  XNOR U8450 ( .A(n8199), .B(n8198), .Z(n8232) );
  XNOR U8451 ( .A(sreg[451]), .B(n8232), .Z(n8234) );
  NANDN U8452 ( .A(sreg[450]), .B(n8191), .Z(n8195) );
  NAND U8453 ( .A(n8193), .B(n8192), .Z(n8194) );
  NAND U8454 ( .A(n8195), .B(n8194), .Z(n8233) );
  XNOR U8455 ( .A(n8234), .B(n8233), .Z(c[451]) );
  NANDN U8456 ( .A(n8197), .B(n8196), .Z(n8201) );
  NANDN U8457 ( .A(n8199), .B(n8198), .Z(n8200) );
  AND U8458 ( .A(n8201), .B(n8200), .Z(n8240) );
  NANDN U8459 ( .A(n8203), .B(n8202), .Z(n8207) );
  NANDN U8460 ( .A(n8205), .B(n8204), .Z(n8206) );
  AND U8461 ( .A(n8207), .B(n8206), .Z(n8238) );
  NAND U8462 ( .A(n26), .B(n8208), .Z(n8210) );
  XOR U8463 ( .A(b[7]), .B(a[198]), .Z(n8249) );
  NAND U8464 ( .A(n10531), .B(n8249), .Z(n8209) );
  AND U8465 ( .A(n8210), .B(n8209), .Z(n8268) );
  NAND U8466 ( .A(n23), .B(n8211), .Z(n8213) );
  XOR U8467 ( .A(b[3]), .B(a[202]), .Z(n8252) );
  NAND U8468 ( .A(n24), .B(n8252), .Z(n8212) );
  NAND U8469 ( .A(n8213), .B(n8212), .Z(n8267) );
  XNOR U8470 ( .A(n8268), .B(n8267), .Z(n8270) );
  NAND U8471 ( .A(b[0]), .B(a[204]), .Z(n8214) );
  XNOR U8472 ( .A(b[1]), .B(n8214), .Z(n8216) );
  NANDN U8473 ( .A(b[0]), .B(a[203]), .Z(n8215) );
  NAND U8474 ( .A(n8216), .B(n8215), .Z(n8264) );
  NAND U8475 ( .A(n25), .B(n8217), .Z(n8219) );
  XOR U8476 ( .A(b[5]), .B(a[200]), .Z(n8258) );
  NAND U8477 ( .A(n10456), .B(n8258), .Z(n8218) );
  AND U8478 ( .A(n8219), .B(n8218), .Z(n8262) );
  AND U8479 ( .A(b[7]), .B(a[196]), .Z(n8261) );
  XNOR U8480 ( .A(n8262), .B(n8261), .Z(n8263) );
  XNOR U8481 ( .A(n8264), .B(n8263), .Z(n8269) );
  XOR U8482 ( .A(n8270), .B(n8269), .Z(n8244) );
  NANDN U8483 ( .A(n8221), .B(n8220), .Z(n8225) );
  NANDN U8484 ( .A(n8223), .B(n8222), .Z(n8224) );
  AND U8485 ( .A(n8225), .B(n8224), .Z(n8243) );
  XNOR U8486 ( .A(n8244), .B(n8243), .Z(n8245) );
  NANDN U8487 ( .A(n8227), .B(n8226), .Z(n8231) );
  NAND U8488 ( .A(n8229), .B(n8228), .Z(n8230) );
  NAND U8489 ( .A(n8231), .B(n8230), .Z(n8246) );
  XNOR U8490 ( .A(n8245), .B(n8246), .Z(n8237) );
  XNOR U8491 ( .A(n8238), .B(n8237), .Z(n8239) );
  XNOR U8492 ( .A(n8240), .B(n8239), .Z(n8273) );
  XNOR U8493 ( .A(sreg[452]), .B(n8273), .Z(n8275) );
  NANDN U8494 ( .A(sreg[451]), .B(n8232), .Z(n8236) );
  NAND U8495 ( .A(n8234), .B(n8233), .Z(n8235) );
  NAND U8496 ( .A(n8236), .B(n8235), .Z(n8274) );
  XNOR U8497 ( .A(n8275), .B(n8274), .Z(c[452]) );
  NANDN U8498 ( .A(n8238), .B(n8237), .Z(n8242) );
  NANDN U8499 ( .A(n8240), .B(n8239), .Z(n8241) );
  AND U8500 ( .A(n8242), .B(n8241), .Z(n8281) );
  NANDN U8501 ( .A(n8244), .B(n8243), .Z(n8248) );
  NANDN U8502 ( .A(n8246), .B(n8245), .Z(n8247) );
  AND U8503 ( .A(n8248), .B(n8247), .Z(n8279) );
  NAND U8504 ( .A(n26), .B(n8249), .Z(n8251) );
  XOR U8505 ( .A(b[7]), .B(a[199]), .Z(n8290) );
  NAND U8506 ( .A(n10531), .B(n8290), .Z(n8250) );
  AND U8507 ( .A(n8251), .B(n8250), .Z(n8306) );
  NAND U8508 ( .A(n23), .B(n8252), .Z(n8254) );
  XOR U8509 ( .A(b[3]), .B(a[203]), .Z(n8293) );
  NAND U8510 ( .A(n24), .B(n8293), .Z(n8253) );
  NAND U8511 ( .A(n8254), .B(n8253), .Z(n8305) );
  XNOR U8512 ( .A(n8306), .B(n8305), .Z(n8308) );
  NAND U8513 ( .A(b[0]), .B(a[205]), .Z(n8255) );
  XNOR U8514 ( .A(b[1]), .B(n8255), .Z(n8257) );
  NANDN U8515 ( .A(b[0]), .B(a[204]), .Z(n8256) );
  NAND U8516 ( .A(n8257), .B(n8256), .Z(n8302) );
  NAND U8517 ( .A(n25), .B(n8258), .Z(n8260) );
  XOR U8518 ( .A(b[5]), .B(a[201]), .Z(n8296) );
  NAND U8519 ( .A(n10456), .B(n8296), .Z(n8259) );
  AND U8520 ( .A(n8260), .B(n8259), .Z(n8300) );
  AND U8521 ( .A(b[7]), .B(a[197]), .Z(n8299) );
  XNOR U8522 ( .A(n8300), .B(n8299), .Z(n8301) );
  XNOR U8523 ( .A(n8302), .B(n8301), .Z(n8307) );
  XOR U8524 ( .A(n8308), .B(n8307), .Z(n8285) );
  NANDN U8525 ( .A(n8262), .B(n8261), .Z(n8266) );
  NANDN U8526 ( .A(n8264), .B(n8263), .Z(n8265) );
  AND U8527 ( .A(n8266), .B(n8265), .Z(n8284) );
  XNOR U8528 ( .A(n8285), .B(n8284), .Z(n8286) );
  NANDN U8529 ( .A(n8268), .B(n8267), .Z(n8272) );
  NAND U8530 ( .A(n8270), .B(n8269), .Z(n8271) );
  NAND U8531 ( .A(n8272), .B(n8271), .Z(n8287) );
  XNOR U8532 ( .A(n8286), .B(n8287), .Z(n8278) );
  XNOR U8533 ( .A(n8279), .B(n8278), .Z(n8280) );
  XNOR U8534 ( .A(n8281), .B(n8280), .Z(n8311) );
  XNOR U8535 ( .A(sreg[453]), .B(n8311), .Z(n8313) );
  NANDN U8536 ( .A(sreg[452]), .B(n8273), .Z(n8277) );
  NAND U8537 ( .A(n8275), .B(n8274), .Z(n8276) );
  NAND U8538 ( .A(n8277), .B(n8276), .Z(n8312) );
  XNOR U8539 ( .A(n8313), .B(n8312), .Z(c[453]) );
  NANDN U8540 ( .A(n8279), .B(n8278), .Z(n8283) );
  NANDN U8541 ( .A(n8281), .B(n8280), .Z(n8282) );
  AND U8542 ( .A(n8283), .B(n8282), .Z(n8319) );
  NANDN U8543 ( .A(n8285), .B(n8284), .Z(n8289) );
  NANDN U8544 ( .A(n8287), .B(n8286), .Z(n8288) );
  AND U8545 ( .A(n8289), .B(n8288), .Z(n8317) );
  NAND U8546 ( .A(n26), .B(n8290), .Z(n8292) );
  XOR U8547 ( .A(b[7]), .B(a[200]), .Z(n8328) );
  NAND U8548 ( .A(n10531), .B(n8328), .Z(n8291) );
  AND U8549 ( .A(n8292), .B(n8291), .Z(n8347) );
  NAND U8550 ( .A(n23), .B(n8293), .Z(n8295) );
  XOR U8551 ( .A(b[3]), .B(a[204]), .Z(n8331) );
  NAND U8552 ( .A(n24), .B(n8331), .Z(n8294) );
  NAND U8553 ( .A(n8295), .B(n8294), .Z(n8346) );
  XNOR U8554 ( .A(n8347), .B(n8346), .Z(n8349) );
  NAND U8555 ( .A(n25), .B(n8296), .Z(n8298) );
  XOR U8556 ( .A(b[5]), .B(a[202]), .Z(n8337) );
  NAND U8557 ( .A(n10456), .B(n8337), .Z(n8297) );
  AND U8558 ( .A(n8298), .B(n8297), .Z(n8341) );
  AND U8559 ( .A(b[7]), .B(a[198]), .Z(n8340) );
  XOR U8560 ( .A(n8341), .B(n8340), .Z(n8343) );
  XNOR U8561 ( .A(n8342), .B(n8343), .Z(n8348) );
  XOR U8562 ( .A(n8349), .B(n8348), .Z(n8323) );
  NANDN U8563 ( .A(n8300), .B(n8299), .Z(n8304) );
  NANDN U8564 ( .A(n8302), .B(n8301), .Z(n8303) );
  AND U8565 ( .A(n8304), .B(n8303), .Z(n8322) );
  XNOR U8566 ( .A(n8323), .B(n8322), .Z(n8324) );
  NANDN U8567 ( .A(n8306), .B(n8305), .Z(n8310) );
  NAND U8568 ( .A(n8308), .B(n8307), .Z(n8309) );
  NAND U8569 ( .A(n8310), .B(n8309), .Z(n8325) );
  XNOR U8570 ( .A(n8324), .B(n8325), .Z(n8316) );
  XNOR U8571 ( .A(n8317), .B(n8316), .Z(n8318) );
  XNOR U8572 ( .A(n8319), .B(n8318), .Z(n8352) );
  XNOR U8573 ( .A(sreg[454]), .B(n8352), .Z(n8354) );
  NANDN U8574 ( .A(sreg[453]), .B(n8311), .Z(n8315) );
  NAND U8575 ( .A(n8313), .B(n8312), .Z(n8314) );
  NAND U8576 ( .A(n8315), .B(n8314), .Z(n8353) );
  XNOR U8577 ( .A(n8354), .B(n8353), .Z(c[454]) );
  NANDN U8578 ( .A(n8317), .B(n8316), .Z(n8321) );
  NANDN U8579 ( .A(n8319), .B(n8318), .Z(n8320) );
  AND U8580 ( .A(n8321), .B(n8320), .Z(n8360) );
  NANDN U8581 ( .A(n8323), .B(n8322), .Z(n8327) );
  NANDN U8582 ( .A(n8325), .B(n8324), .Z(n8326) );
  AND U8583 ( .A(n8327), .B(n8326), .Z(n8358) );
  NAND U8584 ( .A(n26), .B(n8328), .Z(n8330) );
  XOR U8585 ( .A(b[7]), .B(a[201]), .Z(n8369) );
  NAND U8586 ( .A(n10531), .B(n8369), .Z(n8329) );
  AND U8587 ( .A(n8330), .B(n8329), .Z(n8388) );
  NAND U8588 ( .A(n23), .B(n8331), .Z(n8333) );
  XOR U8589 ( .A(b[3]), .B(a[205]), .Z(n8372) );
  NAND U8590 ( .A(n24), .B(n8372), .Z(n8332) );
  NAND U8591 ( .A(n8333), .B(n8332), .Z(n8387) );
  XNOR U8592 ( .A(n8388), .B(n8387), .Z(n8390) );
  NAND U8593 ( .A(b[0]), .B(a[207]), .Z(n8334) );
  XNOR U8594 ( .A(b[1]), .B(n8334), .Z(n8336) );
  NANDN U8595 ( .A(b[0]), .B(a[206]), .Z(n8335) );
  NAND U8596 ( .A(n8336), .B(n8335), .Z(n8384) );
  NAND U8597 ( .A(n25), .B(n8337), .Z(n8339) );
  XOR U8598 ( .A(b[5]), .B(a[203]), .Z(n8378) );
  NAND U8599 ( .A(n10456), .B(n8378), .Z(n8338) );
  AND U8600 ( .A(n8339), .B(n8338), .Z(n8382) );
  AND U8601 ( .A(b[7]), .B(a[199]), .Z(n8381) );
  XNOR U8602 ( .A(n8382), .B(n8381), .Z(n8383) );
  XNOR U8603 ( .A(n8384), .B(n8383), .Z(n8389) );
  XOR U8604 ( .A(n8390), .B(n8389), .Z(n8364) );
  NANDN U8605 ( .A(n8341), .B(n8340), .Z(n8345) );
  NANDN U8606 ( .A(n8343), .B(n8342), .Z(n8344) );
  AND U8607 ( .A(n8345), .B(n8344), .Z(n8363) );
  XNOR U8608 ( .A(n8364), .B(n8363), .Z(n8365) );
  NANDN U8609 ( .A(n8347), .B(n8346), .Z(n8351) );
  NAND U8610 ( .A(n8349), .B(n8348), .Z(n8350) );
  NAND U8611 ( .A(n8351), .B(n8350), .Z(n8366) );
  XNOR U8612 ( .A(n8365), .B(n8366), .Z(n8357) );
  XNOR U8613 ( .A(n8358), .B(n8357), .Z(n8359) );
  XNOR U8614 ( .A(n8360), .B(n8359), .Z(n8393) );
  XNOR U8615 ( .A(sreg[455]), .B(n8393), .Z(n8395) );
  NANDN U8616 ( .A(sreg[454]), .B(n8352), .Z(n8356) );
  NAND U8617 ( .A(n8354), .B(n8353), .Z(n8355) );
  NAND U8618 ( .A(n8356), .B(n8355), .Z(n8394) );
  XNOR U8619 ( .A(n8395), .B(n8394), .Z(c[455]) );
  NANDN U8620 ( .A(n8358), .B(n8357), .Z(n8362) );
  NANDN U8621 ( .A(n8360), .B(n8359), .Z(n8361) );
  AND U8622 ( .A(n8362), .B(n8361), .Z(n8401) );
  NANDN U8623 ( .A(n8364), .B(n8363), .Z(n8368) );
  NANDN U8624 ( .A(n8366), .B(n8365), .Z(n8367) );
  AND U8625 ( .A(n8368), .B(n8367), .Z(n8399) );
  NAND U8626 ( .A(n26), .B(n8369), .Z(n8371) );
  XOR U8627 ( .A(b[7]), .B(a[202]), .Z(n8410) );
  NAND U8628 ( .A(n10531), .B(n8410), .Z(n8370) );
  AND U8629 ( .A(n8371), .B(n8370), .Z(n8429) );
  NAND U8630 ( .A(n23), .B(n8372), .Z(n8374) );
  XOR U8631 ( .A(b[3]), .B(a[206]), .Z(n8413) );
  NAND U8632 ( .A(n24), .B(n8413), .Z(n8373) );
  NAND U8633 ( .A(n8374), .B(n8373), .Z(n8428) );
  XNOR U8634 ( .A(n8429), .B(n8428), .Z(n8431) );
  NAND U8635 ( .A(b[0]), .B(a[208]), .Z(n8375) );
  XNOR U8636 ( .A(b[1]), .B(n8375), .Z(n8377) );
  NANDN U8637 ( .A(b[0]), .B(a[207]), .Z(n8376) );
  NAND U8638 ( .A(n8377), .B(n8376), .Z(n8425) );
  NAND U8639 ( .A(n25), .B(n8378), .Z(n8380) );
  XOR U8640 ( .A(b[5]), .B(a[204]), .Z(n8419) );
  NAND U8641 ( .A(n10456), .B(n8419), .Z(n8379) );
  AND U8642 ( .A(n8380), .B(n8379), .Z(n8423) );
  AND U8643 ( .A(b[7]), .B(a[200]), .Z(n8422) );
  XNOR U8644 ( .A(n8423), .B(n8422), .Z(n8424) );
  XNOR U8645 ( .A(n8425), .B(n8424), .Z(n8430) );
  XOR U8646 ( .A(n8431), .B(n8430), .Z(n8405) );
  NANDN U8647 ( .A(n8382), .B(n8381), .Z(n8386) );
  NANDN U8648 ( .A(n8384), .B(n8383), .Z(n8385) );
  AND U8649 ( .A(n8386), .B(n8385), .Z(n8404) );
  XNOR U8650 ( .A(n8405), .B(n8404), .Z(n8406) );
  NANDN U8651 ( .A(n8388), .B(n8387), .Z(n8392) );
  NAND U8652 ( .A(n8390), .B(n8389), .Z(n8391) );
  NAND U8653 ( .A(n8392), .B(n8391), .Z(n8407) );
  XNOR U8654 ( .A(n8406), .B(n8407), .Z(n8398) );
  XNOR U8655 ( .A(n8399), .B(n8398), .Z(n8400) );
  XNOR U8656 ( .A(n8401), .B(n8400), .Z(n8434) );
  XNOR U8657 ( .A(sreg[456]), .B(n8434), .Z(n8436) );
  NANDN U8658 ( .A(sreg[455]), .B(n8393), .Z(n8397) );
  NAND U8659 ( .A(n8395), .B(n8394), .Z(n8396) );
  NAND U8660 ( .A(n8397), .B(n8396), .Z(n8435) );
  XNOR U8661 ( .A(n8436), .B(n8435), .Z(c[456]) );
  NANDN U8662 ( .A(n8399), .B(n8398), .Z(n8403) );
  NANDN U8663 ( .A(n8401), .B(n8400), .Z(n8402) );
  AND U8664 ( .A(n8403), .B(n8402), .Z(n8442) );
  NANDN U8665 ( .A(n8405), .B(n8404), .Z(n8409) );
  NANDN U8666 ( .A(n8407), .B(n8406), .Z(n8408) );
  AND U8667 ( .A(n8409), .B(n8408), .Z(n8440) );
  NAND U8668 ( .A(n26), .B(n8410), .Z(n8412) );
  XOR U8669 ( .A(b[7]), .B(a[203]), .Z(n8451) );
  NAND U8670 ( .A(n10531), .B(n8451), .Z(n8411) );
  AND U8671 ( .A(n8412), .B(n8411), .Z(n8470) );
  NAND U8672 ( .A(n23), .B(n8413), .Z(n8415) );
  XOR U8673 ( .A(b[3]), .B(a[207]), .Z(n8454) );
  NAND U8674 ( .A(n24), .B(n8454), .Z(n8414) );
  NAND U8675 ( .A(n8415), .B(n8414), .Z(n8469) );
  XNOR U8676 ( .A(n8470), .B(n8469), .Z(n8472) );
  NAND U8677 ( .A(b[0]), .B(a[209]), .Z(n8416) );
  XNOR U8678 ( .A(b[1]), .B(n8416), .Z(n8418) );
  NANDN U8679 ( .A(b[0]), .B(a[208]), .Z(n8417) );
  NAND U8680 ( .A(n8418), .B(n8417), .Z(n8466) );
  NAND U8681 ( .A(n25), .B(n8419), .Z(n8421) );
  XOR U8682 ( .A(b[5]), .B(a[205]), .Z(n8457) );
  NAND U8683 ( .A(n10456), .B(n8457), .Z(n8420) );
  AND U8684 ( .A(n8421), .B(n8420), .Z(n8464) );
  AND U8685 ( .A(b[7]), .B(a[201]), .Z(n8463) );
  XNOR U8686 ( .A(n8464), .B(n8463), .Z(n8465) );
  XNOR U8687 ( .A(n8466), .B(n8465), .Z(n8471) );
  XOR U8688 ( .A(n8472), .B(n8471), .Z(n8446) );
  NANDN U8689 ( .A(n8423), .B(n8422), .Z(n8427) );
  NANDN U8690 ( .A(n8425), .B(n8424), .Z(n8426) );
  AND U8691 ( .A(n8427), .B(n8426), .Z(n8445) );
  XNOR U8692 ( .A(n8446), .B(n8445), .Z(n8447) );
  NANDN U8693 ( .A(n8429), .B(n8428), .Z(n8433) );
  NAND U8694 ( .A(n8431), .B(n8430), .Z(n8432) );
  NAND U8695 ( .A(n8433), .B(n8432), .Z(n8448) );
  XNOR U8696 ( .A(n8447), .B(n8448), .Z(n8439) );
  XNOR U8697 ( .A(n8440), .B(n8439), .Z(n8441) );
  XNOR U8698 ( .A(n8442), .B(n8441), .Z(n8475) );
  XNOR U8699 ( .A(sreg[457]), .B(n8475), .Z(n8477) );
  NANDN U8700 ( .A(sreg[456]), .B(n8434), .Z(n8438) );
  NAND U8701 ( .A(n8436), .B(n8435), .Z(n8437) );
  NAND U8702 ( .A(n8438), .B(n8437), .Z(n8476) );
  XNOR U8703 ( .A(n8477), .B(n8476), .Z(c[457]) );
  NANDN U8704 ( .A(n8440), .B(n8439), .Z(n8444) );
  NANDN U8705 ( .A(n8442), .B(n8441), .Z(n8443) );
  AND U8706 ( .A(n8444), .B(n8443), .Z(n8483) );
  NANDN U8707 ( .A(n8446), .B(n8445), .Z(n8450) );
  NANDN U8708 ( .A(n8448), .B(n8447), .Z(n8449) );
  AND U8709 ( .A(n8450), .B(n8449), .Z(n8481) );
  NAND U8710 ( .A(n26), .B(n8451), .Z(n8453) );
  XOR U8711 ( .A(b[7]), .B(a[204]), .Z(n8492) );
  NAND U8712 ( .A(n10531), .B(n8492), .Z(n8452) );
  AND U8713 ( .A(n8453), .B(n8452), .Z(n8511) );
  NAND U8714 ( .A(n23), .B(n8454), .Z(n8456) );
  XOR U8715 ( .A(b[3]), .B(a[208]), .Z(n8495) );
  NAND U8716 ( .A(n24), .B(n8495), .Z(n8455) );
  NAND U8717 ( .A(n8456), .B(n8455), .Z(n8510) );
  XNOR U8718 ( .A(n8511), .B(n8510), .Z(n8513) );
  NAND U8719 ( .A(n25), .B(n8457), .Z(n8459) );
  XOR U8720 ( .A(b[5]), .B(a[206]), .Z(n8501) );
  NAND U8721 ( .A(n10456), .B(n8501), .Z(n8458) );
  AND U8722 ( .A(n8459), .B(n8458), .Z(n8505) );
  AND U8723 ( .A(b[7]), .B(a[202]), .Z(n8504) );
  XNOR U8724 ( .A(n8505), .B(n8504), .Z(n8506) );
  NAND U8725 ( .A(b[0]), .B(a[210]), .Z(n8460) );
  XNOR U8726 ( .A(b[1]), .B(n8460), .Z(n8462) );
  NANDN U8727 ( .A(b[0]), .B(a[209]), .Z(n8461) );
  NAND U8728 ( .A(n8462), .B(n8461), .Z(n8507) );
  XNOR U8729 ( .A(n8506), .B(n8507), .Z(n8512) );
  XOR U8730 ( .A(n8513), .B(n8512), .Z(n8487) );
  NANDN U8731 ( .A(n8464), .B(n8463), .Z(n8468) );
  NANDN U8732 ( .A(n8466), .B(n8465), .Z(n8467) );
  AND U8733 ( .A(n8468), .B(n8467), .Z(n8486) );
  XNOR U8734 ( .A(n8487), .B(n8486), .Z(n8488) );
  NANDN U8735 ( .A(n8470), .B(n8469), .Z(n8474) );
  NAND U8736 ( .A(n8472), .B(n8471), .Z(n8473) );
  NAND U8737 ( .A(n8474), .B(n8473), .Z(n8489) );
  XNOR U8738 ( .A(n8488), .B(n8489), .Z(n8480) );
  XNOR U8739 ( .A(n8481), .B(n8480), .Z(n8482) );
  XNOR U8740 ( .A(n8483), .B(n8482), .Z(n8516) );
  XNOR U8741 ( .A(sreg[458]), .B(n8516), .Z(n8518) );
  NANDN U8742 ( .A(sreg[457]), .B(n8475), .Z(n8479) );
  NAND U8743 ( .A(n8477), .B(n8476), .Z(n8478) );
  NAND U8744 ( .A(n8479), .B(n8478), .Z(n8517) );
  XNOR U8745 ( .A(n8518), .B(n8517), .Z(c[458]) );
  NANDN U8746 ( .A(n8481), .B(n8480), .Z(n8485) );
  NANDN U8747 ( .A(n8483), .B(n8482), .Z(n8484) );
  AND U8748 ( .A(n8485), .B(n8484), .Z(n8528) );
  NANDN U8749 ( .A(n8487), .B(n8486), .Z(n8491) );
  NANDN U8750 ( .A(n8489), .B(n8488), .Z(n8490) );
  AND U8751 ( .A(n8491), .B(n8490), .Z(n8527) );
  NAND U8752 ( .A(n26), .B(n8492), .Z(n8494) );
  XOR U8753 ( .A(b[7]), .B(a[205]), .Z(n8538) );
  NAND U8754 ( .A(n10531), .B(n8538), .Z(n8493) );
  AND U8755 ( .A(n8494), .B(n8493), .Z(n8557) );
  NAND U8756 ( .A(n23), .B(n8495), .Z(n8497) );
  XOR U8757 ( .A(b[3]), .B(a[209]), .Z(n8541) );
  NAND U8758 ( .A(n24), .B(n8541), .Z(n8496) );
  NAND U8759 ( .A(n8497), .B(n8496), .Z(n8556) );
  XNOR U8760 ( .A(n8557), .B(n8556), .Z(n8559) );
  NAND U8761 ( .A(b[0]), .B(a[211]), .Z(n8498) );
  XNOR U8762 ( .A(b[1]), .B(n8498), .Z(n8500) );
  NANDN U8763 ( .A(b[0]), .B(a[210]), .Z(n8499) );
  NAND U8764 ( .A(n8500), .B(n8499), .Z(n8553) );
  NAND U8765 ( .A(n25), .B(n8501), .Z(n8503) );
  XOR U8766 ( .A(b[5]), .B(a[207]), .Z(n8547) );
  NAND U8767 ( .A(n10456), .B(n8547), .Z(n8502) );
  AND U8768 ( .A(n8503), .B(n8502), .Z(n8551) );
  AND U8769 ( .A(b[7]), .B(a[203]), .Z(n8550) );
  XNOR U8770 ( .A(n8551), .B(n8550), .Z(n8552) );
  XNOR U8771 ( .A(n8553), .B(n8552), .Z(n8558) );
  XOR U8772 ( .A(n8559), .B(n8558), .Z(n8533) );
  NANDN U8773 ( .A(n8505), .B(n8504), .Z(n8509) );
  NANDN U8774 ( .A(n8507), .B(n8506), .Z(n8508) );
  AND U8775 ( .A(n8509), .B(n8508), .Z(n8532) );
  XNOR U8776 ( .A(n8533), .B(n8532), .Z(n8534) );
  NANDN U8777 ( .A(n8511), .B(n8510), .Z(n8515) );
  NAND U8778 ( .A(n8513), .B(n8512), .Z(n8514) );
  NAND U8779 ( .A(n8515), .B(n8514), .Z(n8535) );
  XNOR U8780 ( .A(n8534), .B(n8535), .Z(n8526) );
  XOR U8781 ( .A(n8527), .B(n8526), .Z(n8529) );
  XOR U8782 ( .A(n8528), .B(n8529), .Z(n8521) );
  XNOR U8783 ( .A(n8521), .B(sreg[459]), .Z(n8523) );
  NANDN U8784 ( .A(sreg[458]), .B(n8516), .Z(n8520) );
  NAND U8785 ( .A(n8518), .B(n8517), .Z(n8519) );
  AND U8786 ( .A(n8520), .B(n8519), .Z(n8522) );
  XOR U8787 ( .A(n8523), .B(n8522), .Z(c[459]) );
  NANDN U8788 ( .A(n8521), .B(sreg[459]), .Z(n8525) );
  NAND U8789 ( .A(n8523), .B(n8522), .Z(n8524) );
  AND U8790 ( .A(n8525), .B(n8524), .Z(n8600) );
  NANDN U8791 ( .A(n8527), .B(n8526), .Z(n8531) );
  OR U8792 ( .A(n8529), .B(n8528), .Z(n8530) );
  AND U8793 ( .A(n8531), .B(n8530), .Z(n8565) );
  NANDN U8794 ( .A(n8533), .B(n8532), .Z(n8537) );
  NANDN U8795 ( .A(n8535), .B(n8534), .Z(n8536) );
  AND U8796 ( .A(n8537), .B(n8536), .Z(n8563) );
  NAND U8797 ( .A(n26), .B(n8538), .Z(n8540) );
  XOR U8798 ( .A(b[7]), .B(a[206]), .Z(n8574) );
  NAND U8799 ( .A(n10531), .B(n8574), .Z(n8539) );
  AND U8800 ( .A(n8540), .B(n8539), .Z(n8593) );
  NAND U8801 ( .A(n23), .B(n8541), .Z(n8543) );
  XOR U8802 ( .A(b[3]), .B(a[210]), .Z(n8577) );
  NAND U8803 ( .A(n24), .B(n8577), .Z(n8542) );
  NAND U8804 ( .A(n8543), .B(n8542), .Z(n8592) );
  XNOR U8805 ( .A(n8593), .B(n8592), .Z(n8595) );
  NAND U8806 ( .A(b[0]), .B(a[212]), .Z(n8544) );
  XNOR U8807 ( .A(b[1]), .B(n8544), .Z(n8546) );
  NANDN U8808 ( .A(b[0]), .B(a[211]), .Z(n8545) );
  NAND U8809 ( .A(n8546), .B(n8545), .Z(n8589) );
  NAND U8810 ( .A(n25), .B(n8547), .Z(n8549) );
  XOR U8811 ( .A(b[5]), .B(a[208]), .Z(n8583) );
  NAND U8812 ( .A(n10456), .B(n8583), .Z(n8548) );
  AND U8813 ( .A(n8549), .B(n8548), .Z(n8587) );
  AND U8814 ( .A(b[7]), .B(a[204]), .Z(n8586) );
  XNOR U8815 ( .A(n8587), .B(n8586), .Z(n8588) );
  XNOR U8816 ( .A(n8589), .B(n8588), .Z(n8594) );
  XOR U8817 ( .A(n8595), .B(n8594), .Z(n8569) );
  NANDN U8818 ( .A(n8551), .B(n8550), .Z(n8555) );
  NANDN U8819 ( .A(n8553), .B(n8552), .Z(n8554) );
  AND U8820 ( .A(n8555), .B(n8554), .Z(n8568) );
  XNOR U8821 ( .A(n8569), .B(n8568), .Z(n8570) );
  NANDN U8822 ( .A(n8557), .B(n8556), .Z(n8561) );
  NAND U8823 ( .A(n8559), .B(n8558), .Z(n8560) );
  NAND U8824 ( .A(n8561), .B(n8560), .Z(n8571) );
  XNOR U8825 ( .A(n8570), .B(n8571), .Z(n8562) );
  XNOR U8826 ( .A(n8563), .B(n8562), .Z(n8564) );
  XNOR U8827 ( .A(n8565), .B(n8564), .Z(n8598) );
  XNOR U8828 ( .A(sreg[460]), .B(n8598), .Z(n8599) );
  XNOR U8829 ( .A(n8600), .B(n8599), .Z(c[460]) );
  NANDN U8830 ( .A(n8563), .B(n8562), .Z(n8567) );
  NANDN U8831 ( .A(n8565), .B(n8564), .Z(n8566) );
  AND U8832 ( .A(n8567), .B(n8566), .Z(n8606) );
  NANDN U8833 ( .A(n8569), .B(n8568), .Z(n8573) );
  NANDN U8834 ( .A(n8571), .B(n8570), .Z(n8572) );
  AND U8835 ( .A(n8573), .B(n8572), .Z(n8604) );
  NAND U8836 ( .A(n26), .B(n8574), .Z(n8576) );
  XOR U8837 ( .A(b[7]), .B(a[207]), .Z(n8615) );
  NAND U8838 ( .A(n10531), .B(n8615), .Z(n8575) );
  AND U8839 ( .A(n8576), .B(n8575), .Z(n8634) );
  NAND U8840 ( .A(n23), .B(n8577), .Z(n8579) );
  XOR U8841 ( .A(b[3]), .B(a[211]), .Z(n8618) );
  NAND U8842 ( .A(n24), .B(n8618), .Z(n8578) );
  NAND U8843 ( .A(n8579), .B(n8578), .Z(n8633) );
  XNOR U8844 ( .A(n8634), .B(n8633), .Z(n8636) );
  NAND U8845 ( .A(b[0]), .B(a[213]), .Z(n8580) );
  XNOR U8846 ( .A(b[1]), .B(n8580), .Z(n8582) );
  NANDN U8847 ( .A(b[0]), .B(a[212]), .Z(n8581) );
  NAND U8848 ( .A(n8582), .B(n8581), .Z(n8630) );
  NAND U8849 ( .A(n25), .B(n8583), .Z(n8585) );
  XOR U8850 ( .A(b[5]), .B(a[209]), .Z(n8624) );
  NAND U8851 ( .A(n10456), .B(n8624), .Z(n8584) );
  AND U8852 ( .A(n8585), .B(n8584), .Z(n8628) );
  AND U8853 ( .A(b[7]), .B(a[205]), .Z(n8627) );
  XNOR U8854 ( .A(n8628), .B(n8627), .Z(n8629) );
  XNOR U8855 ( .A(n8630), .B(n8629), .Z(n8635) );
  XOR U8856 ( .A(n8636), .B(n8635), .Z(n8610) );
  NANDN U8857 ( .A(n8587), .B(n8586), .Z(n8591) );
  NANDN U8858 ( .A(n8589), .B(n8588), .Z(n8590) );
  AND U8859 ( .A(n8591), .B(n8590), .Z(n8609) );
  XNOR U8860 ( .A(n8610), .B(n8609), .Z(n8611) );
  NANDN U8861 ( .A(n8593), .B(n8592), .Z(n8597) );
  NAND U8862 ( .A(n8595), .B(n8594), .Z(n8596) );
  NAND U8863 ( .A(n8597), .B(n8596), .Z(n8612) );
  XNOR U8864 ( .A(n8611), .B(n8612), .Z(n8603) );
  XNOR U8865 ( .A(n8604), .B(n8603), .Z(n8605) );
  XNOR U8866 ( .A(n8606), .B(n8605), .Z(n8639) );
  XNOR U8867 ( .A(sreg[461]), .B(n8639), .Z(n8641) );
  NANDN U8868 ( .A(sreg[460]), .B(n8598), .Z(n8602) );
  NAND U8869 ( .A(n8600), .B(n8599), .Z(n8601) );
  NAND U8870 ( .A(n8602), .B(n8601), .Z(n8640) );
  XNOR U8871 ( .A(n8641), .B(n8640), .Z(c[461]) );
  NANDN U8872 ( .A(n8604), .B(n8603), .Z(n8608) );
  NANDN U8873 ( .A(n8606), .B(n8605), .Z(n8607) );
  AND U8874 ( .A(n8608), .B(n8607), .Z(n8647) );
  NANDN U8875 ( .A(n8610), .B(n8609), .Z(n8614) );
  NANDN U8876 ( .A(n8612), .B(n8611), .Z(n8613) );
  AND U8877 ( .A(n8614), .B(n8613), .Z(n8645) );
  NAND U8878 ( .A(n26), .B(n8615), .Z(n8617) );
  XOR U8879 ( .A(b[7]), .B(a[208]), .Z(n8656) );
  NAND U8880 ( .A(n10531), .B(n8656), .Z(n8616) );
  AND U8881 ( .A(n8617), .B(n8616), .Z(n8675) );
  NAND U8882 ( .A(n23), .B(n8618), .Z(n8620) );
  XOR U8883 ( .A(b[3]), .B(a[212]), .Z(n8659) );
  NAND U8884 ( .A(n24), .B(n8659), .Z(n8619) );
  NAND U8885 ( .A(n8620), .B(n8619), .Z(n8674) );
  XNOR U8886 ( .A(n8675), .B(n8674), .Z(n8677) );
  NAND U8887 ( .A(b[0]), .B(a[214]), .Z(n8621) );
  XNOR U8888 ( .A(b[1]), .B(n8621), .Z(n8623) );
  NANDN U8889 ( .A(b[0]), .B(a[213]), .Z(n8622) );
  NAND U8890 ( .A(n8623), .B(n8622), .Z(n8671) );
  NAND U8891 ( .A(n25), .B(n8624), .Z(n8626) );
  XOR U8892 ( .A(b[5]), .B(a[210]), .Z(n8665) );
  NAND U8893 ( .A(n10456), .B(n8665), .Z(n8625) );
  AND U8894 ( .A(n8626), .B(n8625), .Z(n8669) );
  AND U8895 ( .A(b[7]), .B(a[206]), .Z(n8668) );
  XNOR U8896 ( .A(n8669), .B(n8668), .Z(n8670) );
  XNOR U8897 ( .A(n8671), .B(n8670), .Z(n8676) );
  XOR U8898 ( .A(n8677), .B(n8676), .Z(n8651) );
  NANDN U8899 ( .A(n8628), .B(n8627), .Z(n8632) );
  NANDN U8900 ( .A(n8630), .B(n8629), .Z(n8631) );
  AND U8901 ( .A(n8632), .B(n8631), .Z(n8650) );
  XNOR U8902 ( .A(n8651), .B(n8650), .Z(n8652) );
  NANDN U8903 ( .A(n8634), .B(n8633), .Z(n8638) );
  NAND U8904 ( .A(n8636), .B(n8635), .Z(n8637) );
  NAND U8905 ( .A(n8638), .B(n8637), .Z(n8653) );
  XNOR U8906 ( .A(n8652), .B(n8653), .Z(n8644) );
  XNOR U8907 ( .A(n8645), .B(n8644), .Z(n8646) );
  XNOR U8908 ( .A(n8647), .B(n8646), .Z(n8680) );
  XNOR U8909 ( .A(sreg[462]), .B(n8680), .Z(n8682) );
  NANDN U8910 ( .A(sreg[461]), .B(n8639), .Z(n8643) );
  NAND U8911 ( .A(n8641), .B(n8640), .Z(n8642) );
  NAND U8912 ( .A(n8643), .B(n8642), .Z(n8681) );
  XNOR U8913 ( .A(n8682), .B(n8681), .Z(c[462]) );
  NANDN U8914 ( .A(n8645), .B(n8644), .Z(n8649) );
  NANDN U8915 ( .A(n8647), .B(n8646), .Z(n8648) );
  AND U8916 ( .A(n8649), .B(n8648), .Z(n8688) );
  NANDN U8917 ( .A(n8651), .B(n8650), .Z(n8655) );
  NANDN U8918 ( .A(n8653), .B(n8652), .Z(n8654) );
  AND U8919 ( .A(n8655), .B(n8654), .Z(n8686) );
  NAND U8920 ( .A(n26), .B(n8656), .Z(n8658) );
  XOR U8921 ( .A(b[7]), .B(a[209]), .Z(n8697) );
  NAND U8922 ( .A(n10531), .B(n8697), .Z(n8657) );
  AND U8923 ( .A(n8658), .B(n8657), .Z(n8716) );
  NAND U8924 ( .A(n23), .B(n8659), .Z(n8661) );
  XOR U8925 ( .A(b[3]), .B(a[213]), .Z(n8700) );
  NAND U8926 ( .A(n24), .B(n8700), .Z(n8660) );
  NAND U8927 ( .A(n8661), .B(n8660), .Z(n8715) );
  XNOR U8928 ( .A(n8716), .B(n8715), .Z(n8718) );
  NAND U8929 ( .A(b[0]), .B(a[215]), .Z(n8662) );
  XNOR U8930 ( .A(b[1]), .B(n8662), .Z(n8664) );
  NANDN U8931 ( .A(b[0]), .B(a[214]), .Z(n8663) );
  NAND U8932 ( .A(n8664), .B(n8663), .Z(n8712) );
  NAND U8933 ( .A(n25), .B(n8665), .Z(n8667) );
  XOR U8934 ( .A(b[5]), .B(a[211]), .Z(n8706) );
  NAND U8935 ( .A(n10456), .B(n8706), .Z(n8666) );
  AND U8936 ( .A(n8667), .B(n8666), .Z(n8710) );
  AND U8937 ( .A(b[7]), .B(a[207]), .Z(n8709) );
  XNOR U8938 ( .A(n8710), .B(n8709), .Z(n8711) );
  XNOR U8939 ( .A(n8712), .B(n8711), .Z(n8717) );
  XOR U8940 ( .A(n8718), .B(n8717), .Z(n8692) );
  NANDN U8941 ( .A(n8669), .B(n8668), .Z(n8673) );
  NANDN U8942 ( .A(n8671), .B(n8670), .Z(n8672) );
  AND U8943 ( .A(n8673), .B(n8672), .Z(n8691) );
  XNOR U8944 ( .A(n8692), .B(n8691), .Z(n8693) );
  NANDN U8945 ( .A(n8675), .B(n8674), .Z(n8679) );
  NAND U8946 ( .A(n8677), .B(n8676), .Z(n8678) );
  NAND U8947 ( .A(n8679), .B(n8678), .Z(n8694) );
  XNOR U8948 ( .A(n8693), .B(n8694), .Z(n8685) );
  XNOR U8949 ( .A(n8686), .B(n8685), .Z(n8687) );
  XNOR U8950 ( .A(n8688), .B(n8687), .Z(n8721) );
  XNOR U8951 ( .A(sreg[463]), .B(n8721), .Z(n8723) );
  NANDN U8952 ( .A(sreg[462]), .B(n8680), .Z(n8684) );
  NAND U8953 ( .A(n8682), .B(n8681), .Z(n8683) );
  NAND U8954 ( .A(n8684), .B(n8683), .Z(n8722) );
  XNOR U8955 ( .A(n8723), .B(n8722), .Z(c[463]) );
  NANDN U8956 ( .A(n8686), .B(n8685), .Z(n8690) );
  NANDN U8957 ( .A(n8688), .B(n8687), .Z(n8689) );
  AND U8958 ( .A(n8690), .B(n8689), .Z(n8729) );
  NANDN U8959 ( .A(n8692), .B(n8691), .Z(n8696) );
  NANDN U8960 ( .A(n8694), .B(n8693), .Z(n8695) );
  AND U8961 ( .A(n8696), .B(n8695), .Z(n8727) );
  NAND U8962 ( .A(n26), .B(n8697), .Z(n8699) );
  XOR U8963 ( .A(b[7]), .B(a[210]), .Z(n8738) );
  NAND U8964 ( .A(n10531), .B(n8738), .Z(n8698) );
  AND U8965 ( .A(n8699), .B(n8698), .Z(n8757) );
  NAND U8966 ( .A(n23), .B(n8700), .Z(n8702) );
  XOR U8967 ( .A(b[3]), .B(a[214]), .Z(n8741) );
  NAND U8968 ( .A(n24), .B(n8741), .Z(n8701) );
  NAND U8969 ( .A(n8702), .B(n8701), .Z(n8756) );
  XNOR U8970 ( .A(n8757), .B(n8756), .Z(n8759) );
  NAND U8971 ( .A(b[0]), .B(a[216]), .Z(n8703) );
  XNOR U8972 ( .A(b[1]), .B(n8703), .Z(n8705) );
  NANDN U8973 ( .A(b[0]), .B(a[215]), .Z(n8704) );
  NAND U8974 ( .A(n8705), .B(n8704), .Z(n8753) );
  NAND U8975 ( .A(n25), .B(n8706), .Z(n8708) );
  XOR U8976 ( .A(b[5]), .B(a[212]), .Z(n8744) );
  NAND U8977 ( .A(n10456), .B(n8744), .Z(n8707) );
  AND U8978 ( .A(n8708), .B(n8707), .Z(n8751) );
  AND U8979 ( .A(b[7]), .B(a[208]), .Z(n8750) );
  XNOR U8980 ( .A(n8751), .B(n8750), .Z(n8752) );
  XNOR U8981 ( .A(n8753), .B(n8752), .Z(n8758) );
  XOR U8982 ( .A(n8759), .B(n8758), .Z(n8733) );
  NANDN U8983 ( .A(n8710), .B(n8709), .Z(n8714) );
  NANDN U8984 ( .A(n8712), .B(n8711), .Z(n8713) );
  AND U8985 ( .A(n8714), .B(n8713), .Z(n8732) );
  XNOR U8986 ( .A(n8733), .B(n8732), .Z(n8734) );
  NANDN U8987 ( .A(n8716), .B(n8715), .Z(n8720) );
  NAND U8988 ( .A(n8718), .B(n8717), .Z(n8719) );
  NAND U8989 ( .A(n8720), .B(n8719), .Z(n8735) );
  XNOR U8990 ( .A(n8734), .B(n8735), .Z(n8726) );
  XNOR U8991 ( .A(n8727), .B(n8726), .Z(n8728) );
  XNOR U8992 ( .A(n8729), .B(n8728), .Z(n8762) );
  XNOR U8993 ( .A(sreg[464]), .B(n8762), .Z(n8764) );
  NANDN U8994 ( .A(sreg[463]), .B(n8721), .Z(n8725) );
  NAND U8995 ( .A(n8723), .B(n8722), .Z(n8724) );
  NAND U8996 ( .A(n8725), .B(n8724), .Z(n8763) );
  XNOR U8997 ( .A(n8764), .B(n8763), .Z(c[464]) );
  NANDN U8998 ( .A(n8727), .B(n8726), .Z(n8731) );
  NANDN U8999 ( .A(n8729), .B(n8728), .Z(n8730) );
  AND U9000 ( .A(n8731), .B(n8730), .Z(n8770) );
  NANDN U9001 ( .A(n8733), .B(n8732), .Z(n8737) );
  NANDN U9002 ( .A(n8735), .B(n8734), .Z(n8736) );
  AND U9003 ( .A(n8737), .B(n8736), .Z(n8768) );
  NAND U9004 ( .A(n26), .B(n8738), .Z(n8740) );
  XOR U9005 ( .A(b[7]), .B(a[211]), .Z(n8779) );
  NAND U9006 ( .A(n10531), .B(n8779), .Z(n8739) );
  AND U9007 ( .A(n8740), .B(n8739), .Z(n8798) );
  NAND U9008 ( .A(n23), .B(n8741), .Z(n8743) );
  XOR U9009 ( .A(b[3]), .B(a[215]), .Z(n8782) );
  NAND U9010 ( .A(n24), .B(n8782), .Z(n8742) );
  NAND U9011 ( .A(n8743), .B(n8742), .Z(n8797) );
  XNOR U9012 ( .A(n8798), .B(n8797), .Z(n8800) );
  NAND U9013 ( .A(n25), .B(n8744), .Z(n8746) );
  XOR U9014 ( .A(b[5]), .B(a[213]), .Z(n8788) );
  NAND U9015 ( .A(n10456), .B(n8788), .Z(n8745) );
  AND U9016 ( .A(n8746), .B(n8745), .Z(n8792) );
  AND U9017 ( .A(b[7]), .B(a[209]), .Z(n8791) );
  XNOR U9018 ( .A(n8792), .B(n8791), .Z(n8793) );
  NAND U9019 ( .A(b[0]), .B(a[217]), .Z(n8747) );
  XNOR U9020 ( .A(b[1]), .B(n8747), .Z(n8749) );
  NANDN U9021 ( .A(b[0]), .B(a[216]), .Z(n8748) );
  NAND U9022 ( .A(n8749), .B(n8748), .Z(n8794) );
  XNOR U9023 ( .A(n8793), .B(n8794), .Z(n8799) );
  XOR U9024 ( .A(n8800), .B(n8799), .Z(n8774) );
  NANDN U9025 ( .A(n8751), .B(n8750), .Z(n8755) );
  NANDN U9026 ( .A(n8753), .B(n8752), .Z(n8754) );
  AND U9027 ( .A(n8755), .B(n8754), .Z(n8773) );
  XNOR U9028 ( .A(n8774), .B(n8773), .Z(n8775) );
  NANDN U9029 ( .A(n8757), .B(n8756), .Z(n8761) );
  NAND U9030 ( .A(n8759), .B(n8758), .Z(n8760) );
  NAND U9031 ( .A(n8761), .B(n8760), .Z(n8776) );
  XNOR U9032 ( .A(n8775), .B(n8776), .Z(n8767) );
  XNOR U9033 ( .A(n8768), .B(n8767), .Z(n8769) );
  XNOR U9034 ( .A(n8770), .B(n8769), .Z(n8803) );
  XNOR U9035 ( .A(sreg[465]), .B(n8803), .Z(n8805) );
  NANDN U9036 ( .A(sreg[464]), .B(n8762), .Z(n8766) );
  NAND U9037 ( .A(n8764), .B(n8763), .Z(n8765) );
  NAND U9038 ( .A(n8766), .B(n8765), .Z(n8804) );
  XNOR U9039 ( .A(n8805), .B(n8804), .Z(c[465]) );
  NANDN U9040 ( .A(n8768), .B(n8767), .Z(n8772) );
  NANDN U9041 ( .A(n8770), .B(n8769), .Z(n8771) );
  AND U9042 ( .A(n8772), .B(n8771), .Z(n8811) );
  NANDN U9043 ( .A(n8774), .B(n8773), .Z(n8778) );
  NANDN U9044 ( .A(n8776), .B(n8775), .Z(n8777) );
  AND U9045 ( .A(n8778), .B(n8777), .Z(n8809) );
  NAND U9046 ( .A(n26), .B(n8779), .Z(n8781) );
  XOR U9047 ( .A(b[7]), .B(a[212]), .Z(n8820) );
  NAND U9048 ( .A(n10531), .B(n8820), .Z(n8780) );
  AND U9049 ( .A(n8781), .B(n8780), .Z(n8839) );
  NAND U9050 ( .A(n23), .B(n8782), .Z(n8784) );
  XOR U9051 ( .A(b[3]), .B(a[216]), .Z(n8823) );
  NAND U9052 ( .A(n24), .B(n8823), .Z(n8783) );
  NAND U9053 ( .A(n8784), .B(n8783), .Z(n8838) );
  XNOR U9054 ( .A(n8839), .B(n8838), .Z(n8841) );
  NAND U9055 ( .A(b[0]), .B(a[218]), .Z(n8785) );
  XNOR U9056 ( .A(b[1]), .B(n8785), .Z(n8787) );
  NANDN U9057 ( .A(b[0]), .B(a[217]), .Z(n8786) );
  NAND U9058 ( .A(n8787), .B(n8786), .Z(n8835) );
  NAND U9059 ( .A(n25), .B(n8788), .Z(n8790) );
  XOR U9060 ( .A(b[5]), .B(a[214]), .Z(n8826) );
  NAND U9061 ( .A(n10456), .B(n8826), .Z(n8789) );
  AND U9062 ( .A(n8790), .B(n8789), .Z(n8833) );
  AND U9063 ( .A(b[7]), .B(a[210]), .Z(n8832) );
  XNOR U9064 ( .A(n8833), .B(n8832), .Z(n8834) );
  XNOR U9065 ( .A(n8835), .B(n8834), .Z(n8840) );
  XOR U9066 ( .A(n8841), .B(n8840), .Z(n8815) );
  NANDN U9067 ( .A(n8792), .B(n8791), .Z(n8796) );
  NANDN U9068 ( .A(n8794), .B(n8793), .Z(n8795) );
  AND U9069 ( .A(n8796), .B(n8795), .Z(n8814) );
  XNOR U9070 ( .A(n8815), .B(n8814), .Z(n8816) );
  NANDN U9071 ( .A(n8798), .B(n8797), .Z(n8802) );
  NAND U9072 ( .A(n8800), .B(n8799), .Z(n8801) );
  NAND U9073 ( .A(n8802), .B(n8801), .Z(n8817) );
  XNOR U9074 ( .A(n8816), .B(n8817), .Z(n8808) );
  XNOR U9075 ( .A(n8809), .B(n8808), .Z(n8810) );
  XNOR U9076 ( .A(n8811), .B(n8810), .Z(n8844) );
  XNOR U9077 ( .A(sreg[466]), .B(n8844), .Z(n8846) );
  NANDN U9078 ( .A(sreg[465]), .B(n8803), .Z(n8807) );
  NAND U9079 ( .A(n8805), .B(n8804), .Z(n8806) );
  NAND U9080 ( .A(n8807), .B(n8806), .Z(n8845) );
  XNOR U9081 ( .A(n8846), .B(n8845), .Z(c[466]) );
  NANDN U9082 ( .A(n8809), .B(n8808), .Z(n8813) );
  NANDN U9083 ( .A(n8811), .B(n8810), .Z(n8812) );
  AND U9084 ( .A(n8813), .B(n8812), .Z(n8852) );
  NANDN U9085 ( .A(n8815), .B(n8814), .Z(n8819) );
  NANDN U9086 ( .A(n8817), .B(n8816), .Z(n8818) );
  AND U9087 ( .A(n8819), .B(n8818), .Z(n8850) );
  NAND U9088 ( .A(n26), .B(n8820), .Z(n8822) );
  XOR U9089 ( .A(b[7]), .B(a[213]), .Z(n8861) );
  NAND U9090 ( .A(n10531), .B(n8861), .Z(n8821) );
  AND U9091 ( .A(n8822), .B(n8821), .Z(n8880) );
  NAND U9092 ( .A(n23), .B(n8823), .Z(n8825) );
  XOR U9093 ( .A(b[3]), .B(a[217]), .Z(n8864) );
  NAND U9094 ( .A(n24), .B(n8864), .Z(n8824) );
  NAND U9095 ( .A(n8825), .B(n8824), .Z(n8879) );
  XNOR U9096 ( .A(n8880), .B(n8879), .Z(n8882) );
  NAND U9097 ( .A(n25), .B(n8826), .Z(n8828) );
  XOR U9098 ( .A(b[5]), .B(a[215]), .Z(n8867) );
  NAND U9099 ( .A(n10456), .B(n8867), .Z(n8827) );
  AND U9100 ( .A(n8828), .B(n8827), .Z(n8874) );
  AND U9101 ( .A(b[7]), .B(a[211]), .Z(n8873) );
  XNOR U9102 ( .A(n8874), .B(n8873), .Z(n8875) );
  NAND U9103 ( .A(b[0]), .B(a[219]), .Z(n8829) );
  XNOR U9104 ( .A(b[1]), .B(n8829), .Z(n8831) );
  NANDN U9105 ( .A(b[0]), .B(a[218]), .Z(n8830) );
  NAND U9106 ( .A(n8831), .B(n8830), .Z(n8876) );
  XNOR U9107 ( .A(n8875), .B(n8876), .Z(n8881) );
  XOR U9108 ( .A(n8882), .B(n8881), .Z(n8856) );
  NANDN U9109 ( .A(n8833), .B(n8832), .Z(n8837) );
  NANDN U9110 ( .A(n8835), .B(n8834), .Z(n8836) );
  AND U9111 ( .A(n8837), .B(n8836), .Z(n8855) );
  XNOR U9112 ( .A(n8856), .B(n8855), .Z(n8857) );
  NANDN U9113 ( .A(n8839), .B(n8838), .Z(n8843) );
  NAND U9114 ( .A(n8841), .B(n8840), .Z(n8842) );
  NAND U9115 ( .A(n8843), .B(n8842), .Z(n8858) );
  XNOR U9116 ( .A(n8857), .B(n8858), .Z(n8849) );
  XNOR U9117 ( .A(n8850), .B(n8849), .Z(n8851) );
  XNOR U9118 ( .A(n8852), .B(n8851), .Z(n8885) );
  XNOR U9119 ( .A(sreg[467]), .B(n8885), .Z(n8887) );
  NANDN U9120 ( .A(sreg[466]), .B(n8844), .Z(n8848) );
  NAND U9121 ( .A(n8846), .B(n8845), .Z(n8847) );
  NAND U9122 ( .A(n8848), .B(n8847), .Z(n8886) );
  XNOR U9123 ( .A(n8887), .B(n8886), .Z(c[467]) );
  NANDN U9124 ( .A(n8850), .B(n8849), .Z(n8854) );
  NANDN U9125 ( .A(n8852), .B(n8851), .Z(n8853) );
  AND U9126 ( .A(n8854), .B(n8853), .Z(n8893) );
  NANDN U9127 ( .A(n8856), .B(n8855), .Z(n8860) );
  NANDN U9128 ( .A(n8858), .B(n8857), .Z(n8859) );
  AND U9129 ( .A(n8860), .B(n8859), .Z(n8891) );
  NAND U9130 ( .A(n26), .B(n8861), .Z(n8863) );
  XOR U9131 ( .A(b[7]), .B(a[214]), .Z(n8902) );
  NAND U9132 ( .A(n10531), .B(n8902), .Z(n8862) );
  AND U9133 ( .A(n8863), .B(n8862), .Z(n8921) );
  NAND U9134 ( .A(n23), .B(n8864), .Z(n8866) );
  XOR U9135 ( .A(b[3]), .B(a[218]), .Z(n8905) );
  NAND U9136 ( .A(n24), .B(n8905), .Z(n8865) );
  NAND U9137 ( .A(n8866), .B(n8865), .Z(n8920) );
  XNOR U9138 ( .A(n8921), .B(n8920), .Z(n8923) );
  NAND U9139 ( .A(n25), .B(n8867), .Z(n8869) );
  XOR U9140 ( .A(b[5]), .B(a[216]), .Z(n8908) );
  NAND U9141 ( .A(n10456), .B(n8908), .Z(n8868) );
  AND U9142 ( .A(n8869), .B(n8868), .Z(n8915) );
  AND U9143 ( .A(b[7]), .B(a[212]), .Z(n8914) );
  XNOR U9144 ( .A(n8915), .B(n8914), .Z(n8916) );
  NAND U9145 ( .A(b[0]), .B(a[220]), .Z(n8870) );
  XNOR U9146 ( .A(b[1]), .B(n8870), .Z(n8872) );
  NANDN U9147 ( .A(b[0]), .B(a[219]), .Z(n8871) );
  NAND U9148 ( .A(n8872), .B(n8871), .Z(n8917) );
  XNOR U9149 ( .A(n8916), .B(n8917), .Z(n8922) );
  XOR U9150 ( .A(n8923), .B(n8922), .Z(n8897) );
  NANDN U9151 ( .A(n8874), .B(n8873), .Z(n8878) );
  NANDN U9152 ( .A(n8876), .B(n8875), .Z(n8877) );
  AND U9153 ( .A(n8878), .B(n8877), .Z(n8896) );
  XNOR U9154 ( .A(n8897), .B(n8896), .Z(n8898) );
  NANDN U9155 ( .A(n8880), .B(n8879), .Z(n8884) );
  NAND U9156 ( .A(n8882), .B(n8881), .Z(n8883) );
  NAND U9157 ( .A(n8884), .B(n8883), .Z(n8899) );
  XNOR U9158 ( .A(n8898), .B(n8899), .Z(n8890) );
  XNOR U9159 ( .A(n8891), .B(n8890), .Z(n8892) );
  XNOR U9160 ( .A(n8893), .B(n8892), .Z(n8926) );
  XNOR U9161 ( .A(sreg[468]), .B(n8926), .Z(n8928) );
  NANDN U9162 ( .A(sreg[467]), .B(n8885), .Z(n8889) );
  NAND U9163 ( .A(n8887), .B(n8886), .Z(n8888) );
  NAND U9164 ( .A(n8889), .B(n8888), .Z(n8927) );
  XNOR U9165 ( .A(n8928), .B(n8927), .Z(c[468]) );
  NANDN U9166 ( .A(n8891), .B(n8890), .Z(n8895) );
  NANDN U9167 ( .A(n8893), .B(n8892), .Z(n8894) );
  AND U9168 ( .A(n8895), .B(n8894), .Z(n8934) );
  NANDN U9169 ( .A(n8897), .B(n8896), .Z(n8901) );
  NANDN U9170 ( .A(n8899), .B(n8898), .Z(n8900) );
  AND U9171 ( .A(n8901), .B(n8900), .Z(n8932) );
  NAND U9172 ( .A(n26), .B(n8902), .Z(n8904) );
  XOR U9173 ( .A(b[7]), .B(a[215]), .Z(n8943) );
  NAND U9174 ( .A(n10531), .B(n8943), .Z(n8903) );
  AND U9175 ( .A(n8904), .B(n8903), .Z(n8962) );
  NAND U9176 ( .A(n23), .B(n8905), .Z(n8907) );
  XOR U9177 ( .A(b[3]), .B(a[219]), .Z(n8946) );
  NAND U9178 ( .A(n24), .B(n8946), .Z(n8906) );
  NAND U9179 ( .A(n8907), .B(n8906), .Z(n8961) );
  XNOR U9180 ( .A(n8962), .B(n8961), .Z(n8964) );
  NAND U9181 ( .A(n25), .B(n8908), .Z(n8910) );
  XOR U9182 ( .A(b[5]), .B(a[217]), .Z(n8952) );
  NAND U9183 ( .A(n10456), .B(n8952), .Z(n8909) );
  AND U9184 ( .A(n8910), .B(n8909), .Z(n8956) );
  AND U9185 ( .A(b[7]), .B(a[213]), .Z(n8955) );
  XNOR U9186 ( .A(n8956), .B(n8955), .Z(n8957) );
  NAND U9187 ( .A(b[0]), .B(a[221]), .Z(n8911) );
  XNOR U9188 ( .A(b[1]), .B(n8911), .Z(n8913) );
  NANDN U9189 ( .A(b[0]), .B(a[220]), .Z(n8912) );
  NAND U9190 ( .A(n8913), .B(n8912), .Z(n8958) );
  XNOR U9191 ( .A(n8957), .B(n8958), .Z(n8963) );
  XOR U9192 ( .A(n8964), .B(n8963), .Z(n8938) );
  NANDN U9193 ( .A(n8915), .B(n8914), .Z(n8919) );
  NANDN U9194 ( .A(n8917), .B(n8916), .Z(n8918) );
  AND U9195 ( .A(n8919), .B(n8918), .Z(n8937) );
  XNOR U9196 ( .A(n8938), .B(n8937), .Z(n8939) );
  NANDN U9197 ( .A(n8921), .B(n8920), .Z(n8925) );
  NAND U9198 ( .A(n8923), .B(n8922), .Z(n8924) );
  NAND U9199 ( .A(n8925), .B(n8924), .Z(n8940) );
  XNOR U9200 ( .A(n8939), .B(n8940), .Z(n8931) );
  XNOR U9201 ( .A(n8932), .B(n8931), .Z(n8933) );
  XNOR U9202 ( .A(n8934), .B(n8933), .Z(n8967) );
  XNOR U9203 ( .A(sreg[469]), .B(n8967), .Z(n8969) );
  NANDN U9204 ( .A(sreg[468]), .B(n8926), .Z(n8930) );
  NAND U9205 ( .A(n8928), .B(n8927), .Z(n8929) );
  NAND U9206 ( .A(n8930), .B(n8929), .Z(n8968) );
  XNOR U9207 ( .A(n8969), .B(n8968), .Z(c[469]) );
  NANDN U9208 ( .A(n8932), .B(n8931), .Z(n8936) );
  NANDN U9209 ( .A(n8934), .B(n8933), .Z(n8935) );
  AND U9210 ( .A(n8936), .B(n8935), .Z(n8975) );
  NANDN U9211 ( .A(n8938), .B(n8937), .Z(n8942) );
  NANDN U9212 ( .A(n8940), .B(n8939), .Z(n8941) );
  AND U9213 ( .A(n8942), .B(n8941), .Z(n8973) );
  NAND U9214 ( .A(n26), .B(n8943), .Z(n8945) );
  XOR U9215 ( .A(b[7]), .B(a[216]), .Z(n8984) );
  NAND U9216 ( .A(n10531), .B(n8984), .Z(n8944) );
  AND U9217 ( .A(n8945), .B(n8944), .Z(n9003) );
  NAND U9218 ( .A(n23), .B(n8946), .Z(n8948) );
  XOR U9219 ( .A(b[3]), .B(a[220]), .Z(n8987) );
  NAND U9220 ( .A(n24), .B(n8987), .Z(n8947) );
  NAND U9221 ( .A(n8948), .B(n8947), .Z(n9002) );
  XNOR U9222 ( .A(n9003), .B(n9002), .Z(n9005) );
  NAND U9223 ( .A(b[0]), .B(a[222]), .Z(n8949) );
  XNOR U9224 ( .A(b[1]), .B(n8949), .Z(n8951) );
  NANDN U9225 ( .A(b[0]), .B(a[221]), .Z(n8950) );
  NAND U9226 ( .A(n8951), .B(n8950), .Z(n8999) );
  NAND U9227 ( .A(n25), .B(n8952), .Z(n8954) );
  XOR U9228 ( .A(b[5]), .B(a[218]), .Z(n8993) );
  NAND U9229 ( .A(n10456), .B(n8993), .Z(n8953) );
  AND U9230 ( .A(n8954), .B(n8953), .Z(n8997) );
  AND U9231 ( .A(b[7]), .B(a[214]), .Z(n8996) );
  XNOR U9232 ( .A(n8997), .B(n8996), .Z(n8998) );
  XNOR U9233 ( .A(n8999), .B(n8998), .Z(n9004) );
  XOR U9234 ( .A(n9005), .B(n9004), .Z(n8979) );
  NANDN U9235 ( .A(n8956), .B(n8955), .Z(n8960) );
  NANDN U9236 ( .A(n8958), .B(n8957), .Z(n8959) );
  AND U9237 ( .A(n8960), .B(n8959), .Z(n8978) );
  XNOR U9238 ( .A(n8979), .B(n8978), .Z(n8980) );
  NANDN U9239 ( .A(n8962), .B(n8961), .Z(n8966) );
  NAND U9240 ( .A(n8964), .B(n8963), .Z(n8965) );
  NAND U9241 ( .A(n8966), .B(n8965), .Z(n8981) );
  XNOR U9242 ( .A(n8980), .B(n8981), .Z(n8972) );
  XNOR U9243 ( .A(n8973), .B(n8972), .Z(n8974) );
  XNOR U9244 ( .A(n8975), .B(n8974), .Z(n9008) );
  XNOR U9245 ( .A(sreg[470]), .B(n9008), .Z(n9010) );
  NANDN U9246 ( .A(sreg[469]), .B(n8967), .Z(n8971) );
  NAND U9247 ( .A(n8969), .B(n8968), .Z(n8970) );
  NAND U9248 ( .A(n8971), .B(n8970), .Z(n9009) );
  XNOR U9249 ( .A(n9010), .B(n9009), .Z(c[470]) );
  NANDN U9250 ( .A(n8973), .B(n8972), .Z(n8977) );
  NANDN U9251 ( .A(n8975), .B(n8974), .Z(n8976) );
  AND U9252 ( .A(n8977), .B(n8976), .Z(n9016) );
  NANDN U9253 ( .A(n8979), .B(n8978), .Z(n8983) );
  NANDN U9254 ( .A(n8981), .B(n8980), .Z(n8982) );
  AND U9255 ( .A(n8983), .B(n8982), .Z(n9014) );
  NAND U9256 ( .A(n26), .B(n8984), .Z(n8986) );
  XOR U9257 ( .A(b[7]), .B(a[217]), .Z(n9025) );
  NAND U9258 ( .A(n10531), .B(n9025), .Z(n8985) );
  AND U9259 ( .A(n8986), .B(n8985), .Z(n9044) );
  NAND U9260 ( .A(n23), .B(n8987), .Z(n8989) );
  XOR U9261 ( .A(b[3]), .B(a[221]), .Z(n9028) );
  NAND U9262 ( .A(n24), .B(n9028), .Z(n8988) );
  NAND U9263 ( .A(n8989), .B(n8988), .Z(n9043) );
  XNOR U9264 ( .A(n9044), .B(n9043), .Z(n9046) );
  NAND U9265 ( .A(b[0]), .B(a[223]), .Z(n8990) );
  XNOR U9266 ( .A(b[1]), .B(n8990), .Z(n8992) );
  NANDN U9267 ( .A(b[0]), .B(a[222]), .Z(n8991) );
  NAND U9268 ( .A(n8992), .B(n8991), .Z(n9040) );
  NAND U9269 ( .A(n25), .B(n8993), .Z(n8995) );
  XOR U9270 ( .A(b[5]), .B(a[219]), .Z(n9034) );
  NAND U9271 ( .A(n10456), .B(n9034), .Z(n8994) );
  AND U9272 ( .A(n8995), .B(n8994), .Z(n9038) );
  AND U9273 ( .A(b[7]), .B(a[215]), .Z(n9037) );
  XNOR U9274 ( .A(n9038), .B(n9037), .Z(n9039) );
  XNOR U9275 ( .A(n9040), .B(n9039), .Z(n9045) );
  XOR U9276 ( .A(n9046), .B(n9045), .Z(n9020) );
  NANDN U9277 ( .A(n8997), .B(n8996), .Z(n9001) );
  NANDN U9278 ( .A(n8999), .B(n8998), .Z(n9000) );
  AND U9279 ( .A(n9001), .B(n9000), .Z(n9019) );
  XNOR U9280 ( .A(n9020), .B(n9019), .Z(n9021) );
  NANDN U9281 ( .A(n9003), .B(n9002), .Z(n9007) );
  NAND U9282 ( .A(n9005), .B(n9004), .Z(n9006) );
  NAND U9283 ( .A(n9007), .B(n9006), .Z(n9022) );
  XNOR U9284 ( .A(n9021), .B(n9022), .Z(n9013) );
  XNOR U9285 ( .A(n9014), .B(n9013), .Z(n9015) );
  XNOR U9286 ( .A(n9016), .B(n9015), .Z(n9049) );
  XNOR U9287 ( .A(sreg[471]), .B(n9049), .Z(n9051) );
  NANDN U9288 ( .A(sreg[470]), .B(n9008), .Z(n9012) );
  NAND U9289 ( .A(n9010), .B(n9009), .Z(n9011) );
  NAND U9290 ( .A(n9012), .B(n9011), .Z(n9050) );
  XNOR U9291 ( .A(n9051), .B(n9050), .Z(c[471]) );
  NANDN U9292 ( .A(n9014), .B(n9013), .Z(n9018) );
  NANDN U9293 ( .A(n9016), .B(n9015), .Z(n9017) );
  AND U9294 ( .A(n9018), .B(n9017), .Z(n9057) );
  NANDN U9295 ( .A(n9020), .B(n9019), .Z(n9024) );
  NANDN U9296 ( .A(n9022), .B(n9021), .Z(n9023) );
  AND U9297 ( .A(n9024), .B(n9023), .Z(n9055) );
  NAND U9298 ( .A(n26), .B(n9025), .Z(n9027) );
  XOR U9299 ( .A(b[7]), .B(a[218]), .Z(n9066) );
  NAND U9300 ( .A(n10531), .B(n9066), .Z(n9026) );
  AND U9301 ( .A(n9027), .B(n9026), .Z(n9085) );
  NAND U9302 ( .A(n23), .B(n9028), .Z(n9030) );
  XOR U9303 ( .A(b[3]), .B(a[222]), .Z(n9069) );
  NAND U9304 ( .A(n24), .B(n9069), .Z(n9029) );
  NAND U9305 ( .A(n9030), .B(n9029), .Z(n9084) );
  XNOR U9306 ( .A(n9085), .B(n9084), .Z(n9087) );
  NAND U9307 ( .A(b[0]), .B(a[224]), .Z(n9031) );
  XNOR U9308 ( .A(b[1]), .B(n9031), .Z(n9033) );
  NANDN U9309 ( .A(b[0]), .B(a[223]), .Z(n9032) );
  NAND U9310 ( .A(n9033), .B(n9032), .Z(n9081) );
  NAND U9311 ( .A(n25), .B(n9034), .Z(n9036) );
  XOR U9312 ( .A(b[5]), .B(a[220]), .Z(n9075) );
  NAND U9313 ( .A(n10456), .B(n9075), .Z(n9035) );
  AND U9314 ( .A(n9036), .B(n9035), .Z(n9079) );
  AND U9315 ( .A(b[7]), .B(a[216]), .Z(n9078) );
  XNOR U9316 ( .A(n9079), .B(n9078), .Z(n9080) );
  XNOR U9317 ( .A(n9081), .B(n9080), .Z(n9086) );
  XOR U9318 ( .A(n9087), .B(n9086), .Z(n9061) );
  NANDN U9319 ( .A(n9038), .B(n9037), .Z(n9042) );
  NANDN U9320 ( .A(n9040), .B(n9039), .Z(n9041) );
  AND U9321 ( .A(n9042), .B(n9041), .Z(n9060) );
  XNOR U9322 ( .A(n9061), .B(n9060), .Z(n9062) );
  NANDN U9323 ( .A(n9044), .B(n9043), .Z(n9048) );
  NAND U9324 ( .A(n9046), .B(n9045), .Z(n9047) );
  NAND U9325 ( .A(n9048), .B(n9047), .Z(n9063) );
  XNOR U9326 ( .A(n9062), .B(n9063), .Z(n9054) );
  XNOR U9327 ( .A(n9055), .B(n9054), .Z(n9056) );
  XNOR U9328 ( .A(n9057), .B(n9056), .Z(n9090) );
  XNOR U9329 ( .A(sreg[472]), .B(n9090), .Z(n9092) );
  NANDN U9330 ( .A(sreg[471]), .B(n9049), .Z(n9053) );
  NAND U9331 ( .A(n9051), .B(n9050), .Z(n9052) );
  NAND U9332 ( .A(n9053), .B(n9052), .Z(n9091) );
  XNOR U9333 ( .A(n9092), .B(n9091), .Z(c[472]) );
  NANDN U9334 ( .A(n9055), .B(n9054), .Z(n9059) );
  NANDN U9335 ( .A(n9057), .B(n9056), .Z(n9058) );
  AND U9336 ( .A(n9059), .B(n9058), .Z(n9098) );
  NANDN U9337 ( .A(n9061), .B(n9060), .Z(n9065) );
  NANDN U9338 ( .A(n9063), .B(n9062), .Z(n9064) );
  AND U9339 ( .A(n9065), .B(n9064), .Z(n9096) );
  NAND U9340 ( .A(n26), .B(n9066), .Z(n9068) );
  XOR U9341 ( .A(b[7]), .B(a[219]), .Z(n9107) );
  NAND U9342 ( .A(n10531), .B(n9107), .Z(n9067) );
  AND U9343 ( .A(n9068), .B(n9067), .Z(n9126) );
  NAND U9344 ( .A(n23), .B(n9069), .Z(n9071) );
  XOR U9345 ( .A(b[3]), .B(a[223]), .Z(n9110) );
  NAND U9346 ( .A(n24), .B(n9110), .Z(n9070) );
  NAND U9347 ( .A(n9071), .B(n9070), .Z(n9125) );
  XNOR U9348 ( .A(n9126), .B(n9125), .Z(n9128) );
  NAND U9349 ( .A(b[0]), .B(a[225]), .Z(n9072) );
  XNOR U9350 ( .A(b[1]), .B(n9072), .Z(n9074) );
  NANDN U9351 ( .A(b[0]), .B(a[224]), .Z(n9073) );
  NAND U9352 ( .A(n9074), .B(n9073), .Z(n9122) );
  NAND U9353 ( .A(n25), .B(n9075), .Z(n9077) );
  XOR U9354 ( .A(b[5]), .B(a[221]), .Z(n9116) );
  NAND U9355 ( .A(n10456), .B(n9116), .Z(n9076) );
  AND U9356 ( .A(n9077), .B(n9076), .Z(n9120) );
  AND U9357 ( .A(b[7]), .B(a[217]), .Z(n9119) );
  XNOR U9358 ( .A(n9120), .B(n9119), .Z(n9121) );
  XNOR U9359 ( .A(n9122), .B(n9121), .Z(n9127) );
  XOR U9360 ( .A(n9128), .B(n9127), .Z(n9102) );
  NANDN U9361 ( .A(n9079), .B(n9078), .Z(n9083) );
  NANDN U9362 ( .A(n9081), .B(n9080), .Z(n9082) );
  AND U9363 ( .A(n9083), .B(n9082), .Z(n9101) );
  XNOR U9364 ( .A(n9102), .B(n9101), .Z(n9103) );
  NANDN U9365 ( .A(n9085), .B(n9084), .Z(n9089) );
  NAND U9366 ( .A(n9087), .B(n9086), .Z(n9088) );
  NAND U9367 ( .A(n9089), .B(n9088), .Z(n9104) );
  XNOR U9368 ( .A(n9103), .B(n9104), .Z(n9095) );
  XNOR U9369 ( .A(n9096), .B(n9095), .Z(n9097) );
  XNOR U9370 ( .A(n9098), .B(n9097), .Z(n9131) );
  XNOR U9371 ( .A(sreg[473]), .B(n9131), .Z(n9133) );
  NANDN U9372 ( .A(sreg[472]), .B(n9090), .Z(n9094) );
  NAND U9373 ( .A(n9092), .B(n9091), .Z(n9093) );
  NAND U9374 ( .A(n9094), .B(n9093), .Z(n9132) );
  XNOR U9375 ( .A(n9133), .B(n9132), .Z(c[473]) );
  NANDN U9376 ( .A(n9096), .B(n9095), .Z(n9100) );
  NANDN U9377 ( .A(n9098), .B(n9097), .Z(n9099) );
  AND U9378 ( .A(n9100), .B(n9099), .Z(n9139) );
  NANDN U9379 ( .A(n9102), .B(n9101), .Z(n9106) );
  NANDN U9380 ( .A(n9104), .B(n9103), .Z(n9105) );
  AND U9381 ( .A(n9106), .B(n9105), .Z(n9137) );
  NAND U9382 ( .A(n26), .B(n9107), .Z(n9109) );
  XOR U9383 ( .A(b[7]), .B(a[220]), .Z(n9148) );
  NAND U9384 ( .A(n10531), .B(n9148), .Z(n9108) );
  AND U9385 ( .A(n9109), .B(n9108), .Z(n9167) );
  NAND U9386 ( .A(n23), .B(n9110), .Z(n9112) );
  XOR U9387 ( .A(b[3]), .B(a[224]), .Z(n9151) );
  NAND U9388 ( .A(n24), .B(n9151), .Z(n9111) );
  NAND U9389 ( .A(n9112), .B(n9111), .Z(n9166) );
  XNOR U9390 ( .A(n9167), .B(n9166), .Z(n9169) );
  NAND U9391 ( .A(b[0]), .B(a[226]), .Z(n9113) );
  XNOR U9392 ( .A(b[1]), .B(n9113), .Z(n9115) );
  NANDN U9393 ( .A(b[0]), .B(a[225]), .Z(n9114) );
  NAND U9394 ( .A(n9115), .B(n9114), .Z(n9163) );
  NAND U9395 ( .A(n25), .B(n9116), .Z(n9118) );
  XOR U9396 ( .A(b[5]), .B(a[222]), .Z(n9154) );
  NAND U9397 ( .A(n10456), .B(n9154), .Z(n9117) );
  AND U9398 ( .A(n9118), .B(n9117), .Z(n9161) );
  AND U9399 ( .A(b[7]), .B(a[218]), .Z(n9160) );
  XNOR U9400 ( .A(n9161), .B(n9160), .Z(n9162) );
  XNOR U9401 ( .A(n9163), .B(n9162), .Z(n9168) );
  XOR U9402 ( .A(n9169), .B(n9168), .Z(n9143) );
  NANDN U9403 ( .A(n9120), .B(n9119), .Z(n9124) );
  NANDN U9404 ( .A(n9122), .B(n9121), .Z(n9123) );
  AND U9405 ( .A(n9124), .B(n9123), .Z(n9142) );
  XNOR U9406 ( .A(n9143), .B(n9142), .Z(n9144) );
  NANDN U9407 ( .A(n9126), .B(n9125), .Z(n9130) );
  NAND U9408 ( .A(n9128), .B(n9127), .Z(n9129) );
  NAND U9409 ( .A(n9130), .B(n9129), .Z(n9145) );
  XNOR U9410 ( .A(n9144), .B(n9145), .Z(n9136) );
  XNOR U9411 ( .A(n9137), .B(n9136), .Z(n9138) );
  XNOR U9412 ( .A(n9139), .B(n9138), .Z(n9172) );
  XNOR U9413 ( .A(sreg[474]), .B(n9172), .Z(n9174) );
  NANDN U9414 ( .A(sreg[473]), .B(n9131), .Z(n9135) );
  NAND U9415 ( .A(n9133), .B(n9132), .Z(n9134) );
  NAND U9416 ( .A(n9135), .B(n9134), .Z(n9173) );
  XNOR U9417 ( .A(n9174), .B(n9173), .Z(c[474]) );
  NANDN U9418 ( .A(n9137), .B(n9136), .Z(n9141) );
  NANDN U9419 ( .A(n9139), .B(n9138), .Z(n9140) );
  AND U9420 ( .A(n9141), .B(n9140), .Z(n9180) );
  NANDN U9421 ( .A(n9143), .B(n9142), .Z(n9147) );
  NANDN U9422 ( .A(n9145), .B(n9144), .Z(n9146) );
  AND U9423 ( .A(n9147), .B(n9146), .Z(n9178) );
  NAND U9424 ( .A(n26), .B(n9148), .Z(n9150) );
  XOR U9425 ( .A(b[7]), .B(a[221]), .Z(n9189) );
  NAND U9426 ( .A(n10531), .B(n9189), .Z(n9149) );
  AND U9427 ( .A(n9150), .B(n9149), .Z(n9208) );
  NAND U9428 ( .A(n23), .B(n9151), .Z(n9153) );
  XOR U9429 ( .A(b[3]), .B(a[225]), .Z(n9192) );
  NAND U9430 ( .A(n24), .B(n9192), .Z(n9152) );
  NAND U9431 ( .A(n9153), .B(n9152), .Z(n9207) );
  XNOR U9432 ( .A(n9208), .B(n9207), .Z(n9210) );
  NAND U9433 ( .A(n25), .B(n9154), .Z(n9156) );
  XOR U9434 ( .A(b[5]), .B(a[223]), .Z(n9198) );
  NAND U9435 ( .A(n10456), .B(n9198), .Z(n9155) );
  AND U9436 ( .A(n9156), .B(n9155), .Z(n9202) );
  AND U9437 ( .A(b[7]), .B(a[219]), .Z(n9201) );
  XNOR U9438 ( .A(n9202), .B(n9201), .Z(n9203) );
  NAND U9439 ( .A(b[0]), .B(a[227]), .Z(n9157) );
  XNOR U9440 ( .A(b[1]), .B(n9157), .Z(n9159) );
  NANDN U9441 ( .A(b[0]), .B(a[226]), .Z(n9158) );
  NAND U9442 ( .A(n9159), .B(n9158), .Z(n9204) );
  XNOR U9443 ( .A(n9203), .B(n9204), .Z(n9209) );
  XOR U9444 ( .A(n9210), .B(n9209), .Z(n9184) );
  NANDN U9445 ( .A(n9161), .B(n9160), .Z(n9165) );
  NANDN U9446 ( .A(n9163), .B(n9162), .Z(n9164) );
  AND U9447 ( .A(n9165), .B(n9164), .Z(n9183) );
  XNOR U9448 ( .A(n9184), .B(n9183), .Z(n9185) );
  NANDN U9449 ( .A(n9167), .B(n9166), .Z(n9171) );
  NAND U9450 ( .A(n9169), .B(n9168), .Z(n9170) );
  NAND U9451 ( .A(n9171), .B(n9170), .Z(n9186) );
  XNOR U9452 ( .A(n9185), .B(n9186), .Z(n9177) );
  XNOR U9453 ( .A(n9178), .B(n9177), .Z(n9179) );
  XNOR U9454 ( .A(n9180), .B(n9179), .Z(n9213) );
  XNOR U9455 ( .A(sreg[475]), .B(n9213), .Z(n9215) );
  NANDN U9456 ( .A(sreg[474]), .B(n9172), .Z(n9176) );
  NAND U9457 ( .A(n9174), .B(n9173), .Z(n9175) );
  NAND U9458 ( .A(n9176), .B(n9175), .Z(n9214) );
  XNOR U9459 ( .A(n9215), .B(n9214), .Z(c[475]) );
  NANDN U9460 ( .A(n9178), .B(n9177), .Z(n9182) );
  NANDN U9461 ( .A(n9180), .B(n9179), .Z(n9181) );
  AND U9462 ( .A(n9182), .B(n9181), .Z(n9221) );
  NANDN U9463 ( .A(n9184), .B(n9183), .Z(n9188) );
  NANDN U9464 ( .A(n9186), .B(n9185), .Z(n9187) );
  AND U9465 ( .A(n9188), .B(n9187), .Z(n9219) );
  NAND U9466 ( .A(n26), .B(n9189), .Z(n9191) );
  XOR U9467 ( .A(b[7]), .B(a[222]), .Z(n9230) );
  NAND U9468 ( .A(n10531), .B(n9230), .Z(n9190) );
  AND U9469 ( .A(n9191), .B(n9190), .Z(n9249) );
  NAND U9470 ( .A(n23), .B(n9192), .Z(n9194) );
  XOR U9471 ( .A(b[3]), .B(a[226]), .Z(n9233) );
  NAND U9472 ( .A(n24), .B(n9233), .Z(n9193) );
  NAND U9473 ( .A(n9194), .B(n9193), .Z(n9248) );
  XNOR U9474 ( .A(n9249), .B(n9248), .Z(n9251) );
  NAND U9475 ( .A(b[0]), .B(a[228]), .Z(n9195) );
  XNOR U9476 ( .A(b[1]), .B(n9195), .Z(n9197) );
  NANDN U9477 ( .A(b[0]), .B(a[227]), .Z(n9196) );
  NAND U9478 ( .A(n9197), .B(n9196), .Z(n9245) );
  NAND U9479 ( .A(n25), .B(n9198), .Z(n9200) );
  XOR U9480 ( .A(b[5]), .B(a[224]), .Z(n9239) );
  NAND U9481 ( .A(n10456), .B(n9239), .Z(n9199) );
  AND U9482 ( .A(n9200), .B(n9199), .Z(n9243) );
  AND U9483 ( .A(b[7]), .B(a[220]), .Z(n9242) );
  XNOR U9484 ( .A(n9243), .B(n9242), .Z(n9244) );
  XNOR U9485 ( .A(n9245), .B(n9244), .Z(n9250) );
  XOR U9486 ( .A(n9251), .B(n9250), .Z(n9225) );
  NANDN U9487 ( .A(n9202), .B(n9201), .Z(n9206) );
  NANDN U9488 ( .A(n9204), .B(n9203), .Z(n9205) );
  AND U9489 ( .A(n9206), .B(n9205), .Z(n9224) );
  XNOR U9490 ( .A(n9225), .B(n9224), .Z(n9226) );
  NANDN U9491 ( .A(n9208), .B(n9207), .Z(n9212) );
  NAND U9492 ( .A(n9210), .B(n9209), .Z(n9211) );
  NAND U9493 ( .A(n9212), .B(n9211), .Z(n9227) );
  XNOR U9494 ( .A(n9226), .B(n9227), .Z(n9218) );
  XNOR U9495 ( .A(n9219), .B(n9218), .Z(n9220) );
  XNOR U9496 ( .A(n9221), .B(n9220), .Z(n9254) );
  XNOR U9497 ( .A(sreg[476]), .B(n9254), .Z(n9256) );
  NANDN U9498 ( .A(sreg[475]), .B(n9213), .Z(n9217) );
  NAND U9499 ( .A(n9215), .B(n9214), .Z(n9216) );
  NAND U9500 ( .A(n9217), .B(n9216), .Z(n9255) );
  XNOR U9501 ( .A(n9256), .B(n9255), .Z(c[476]) );
  NANDN U9502 ( .A(n9219), .B(n9218), .Z(n9223) );
  NANDN U9503 ( .A(n9221), .B(n9220), .Z(n9222) );
  AND U9504 ( .A(n9223), .B(n9222), .Z(n9262) );
  NANDN U9505 ( .A(n9225), .B(n9224), .Z(n9229) );
  NANDN U9506 ( .A(n9227), .B(n9226), .Z(n9228) );
  AND U9507 ( .A(n9229), .B(n9228), .Z(n9260) );
  NAND U9508 ( .A(n26), .B(n9230), .Z(n9232) );
  XOR U9509 ( .A(b[7]), .B(a[223]), .Z(n9271) );
  NAND U9510 ( .A(n10531), .B(n9271), .Z(n9231) );
  AND U9511 ( .A(n9232), .B(n9231), .Z(n9290) );
  NAND U9512 ( .A(n23), .B(n9233), .Z(n9235) );
  XOR U9513 ( .A(b[3]), .B(a[227]), .Z(n9274) );
  NAND U9514 ( .A(n24), .B(n9274), .Z(n9234) );
  NAND U9515 ( .A(n9235), .B(n9234), .Z(n9289) );
  XNOR U9516 ( .A(n9290), .B(n9289), .Z(n9292) );
  NAND U9517 ( .A(b[0]), .B(a[229]), .Z(n9236) );
  XNOR U9518 ( .A(b[1]), .B(n9236), .Z(n9238) );
  NANDN U9519 ( .A(b[0]), .B(a[228]), .Z(n9237) );
  NAND U9520 ( .A(n9238), .B(n9237), .Z(n9286) );
  NAND U9521 ( .A(n25), .B(n9239), .Z(n9241) );
  XOR U9522 ( .A(b[5]), .B(a[225]), .Z(n9280) );
  NAND U9523 ( .A(n10456), .B(n9280), .Z(n9240) );
  AND U9524 ( .A(n9241), .B(n9240), .Z(n9284) );
  AND U9525 ( .A(b[7]), .B(a[221]), .Z(n9283) );
  XNOR U9526 ( .A(n9284), .B(n9283), .Z(n9285) );
  XNOR U9527 ( .A(n9286), .B(n9285), .Z(n9291) );
  XOR U9528 ( .A(n9292), .B(n9291), .Z(n9266) );
  NANDN U9529 ( .A(n9243), .B(n9242), .Z(n9247) );
  NANDN U9530 ( .A(n9245), .B(n9244), .Z(n9246) );
  AND U9531 ( .A(n9247), .B(n9246), .Z(n9265) );
  XNOR U9532 ( .A(n9266), .B(n9265), .Z(n9267) );
  NANDN U9533 ( .A(n9249), .B(n9248), .Z(n9253) );
  NAND U9534 ( .A(n9251), .B(n9250), .Z(n9252) );
  NAND U9535 ( .A(n9253), .B(n9252), .Z(n9268) );
  XNOR U9536 ( .A(n9267), .B(n9268), .Z(n9259) );
  XNOR U9537 ( .A(n9260), .B(n9259), .Z(n9261) );
  XNOR U9538 ( .A(n9262), .B(n9261), .Z(n9295) );
  XNOR U9539 ( .A(sreg[477]), .B(n9295), .Z(n9297) );
  NANDN U9540 ( .A(sreg[476]), .B(n9254), .Z(n9258) );
  NAND U9541 ( .A(n9256), .B(n9255), .Z(n9257) );
  NAND U9542 ( .A(n9258), .B(n9257), .Z(n9296) );
  XNOR U9543 ( .A(n9297), .B(n9296), .Z(c[477]) );
  NANDN U9544 ( .A(n9260), .B(n9259), .Z(n9264) );
  NANDN U9545 ( .A(n9262), .B(n9261), .Z(n9263) );
  AND U9546 ( .A(n9264), .B(n9263), .Z(n9303) );
  NANDN U9547 ( .A(n9266), .B(n9265), .Z(n9270) );
  NANDN U9548 ( .A(n9268), .B(n9267), .Z(n9269) );
  AND U9549 ( .A(n9270), .B(n9269), .Z(n9301) );
  NAND U9550 ( .A(n26), .B(n9271), .Z(n9273) );
  XOR U9551 ( .A(b[7]), .B(a[224]), .Z(n9312) );
  NAND U9552 ( .A(n10531), .B(n9312), .Z(n9272) );
  AND U9553 ( .A(n9273), .B(n9272), .Z(n9331) );
  NAND U9554 ( .A(n23), .B(n9274), .Z(n9276) );
  XOR U9555 ( .A(b[3]), .B(a[228]), .Z(n9315) );
  NAND U9556 ( .A(n24), .B(n9315), .Z(n9275) );
  NAND U9557 ( .A(n9276), .B(n9275), .Z(n9330) );
  XNOR U9558 ( .A(n9331), .B(n9330), .Z(n9333) );
  NAND U9559 ( .A(b[0]), .B(a[230]), .Z(n9277) );
  XNOR U9560 ( .A(b[1]), .B(n9277), .Z(n9279) );
  NANDN U9561 ( .A(b[0]), .B(a[229]), .Z(n9278) );
  NAND U9562 ( .A(n9279), .B(n9278), .Z(n9327) );
  NAND U9563 ( .A(n25), .B(n9280), .Z(n9282) );
  XOR U9564 ( .A(b[5]), .B(a[226]), .Z(n9321) );
  NAND U9565 ( .A(n10456), .B(n9321), .Z(n9281) );
  AND U9566 ( .A(n9282), .B(n9281), .Z(n9325) );
  AND U9567 ( .A(b[7]), .B(a[222]), .Z(n9324) );
  XNOR U9568 ( .A(n9325), .B(n9324), .Z(n9326) );
  XNOR U9569 ( .A(n9327), .B(n9326), .Z(n9332) );
  XOR U9570 ( .A(n9333), .B(n9332), .Z(n9307) );
  NANDN U9571 ( .A(n9284), .B(n9283), .Z(n9288) );
  NANDN U9572 ( .A(n9286), .B(n9285), .Z(n9287) );
  AND U9573 ( .A(n9288), .B(n9287), .Z(n9306) );
  XNOR U9574 ( .A(n9307), .B(n9306), .Z(n9308) );
  NANDN U9575 ( .A(n9290), .B(n9289), .Z(n9294) );
  NAND U9576 ( .A(n9292), .B(n9291), .Z(n9293) );
  NAND U9577 ( .A(n9294), .B(n9293), .Z(n9309) );
  XNOR U9578 ( .A(n9308), .B(n9309), .Z(n9300) );
  XNOR U9579 ( .A(n9301), .B(n9300), .Z(n9302) );
  XNOR U9580 ( .A(n9303), .B(n9302), .Z(n9336) );
  XNOR U9581 ( .A(sreg[478]), .B(n9336), .Z(n9338) );
  NANDN U9582 ( .A(sreg[477]), .B(n9295), .Z(n9299) );
  NAND U9583 ( .A(n9297), .B(n9296), .Z(n9298) );
  NAND U9584 ( .A(n9299), .B(n9298), .Z(n9337) );
  XNOR U9585 ( .A(n9338), .B(n9337), .Z(c[478]) );
  NANDN U9586 ( .A(n9301), .B(n9300), .Z(n9305) );
  NANDN U9587 ( .A(n9303), .B(n9302), .Z(n9304) );
  AND U9588 ( .A(n9305), .B(n9304), .Z(n9344) );
  NANDN U9589 ( .A(n9307), .B(n9306), .Z(n9311) );
  NANDN U9590 ( .A(n9309), .B(n9308), .Z(n9310) );
  AND U9591 ( .A(n9311), .B(n9310), .Z(n9342) );
  NAND U9592 ( .A(n26), .B(n9312), .Z(n9314) );
  XOR U9593 ( .A(b[7]), .B(a[225]), .Z(n9353) );
  NAND U9594 ( .A(n10531), .B(n9353), .Z(n9313) );
  AND U9595 ( .A(n9314), .B(n9313), .Z(n9372) );
  NAND U9596 ( .A(n23), .B(n9315), .Z(n9317) );
  XOR U9597 ( .A(b[3]), .B(a[229]), .Z(n9356) );
  NAND U9598 ( .A(n24), .B(n9356), .Z(n9316) );
  NAND U9599 ( .A(n9317), .B(n9316), .Z(n9371) );
  XNOR U9600 ( .A(n9372), .B(n9371), .Z(n9374) );
  NAND U9601 ( .A(b[0]), .B(a[231]), .Z(n9318) );
  XNOR U9602 ( .A(b[1]), .B(n9318), .Z(n9320) );
  NANDN U9603 ( .A(b[0]), .B(a[230]), .Z(n9319) );
  NAND U9604 ( .A(n9320), .B(n9319), .Z(n9368) );
  NAND U9605 ( .A(n25), .B(n9321), .Z(n9323) );
  XOR U9606 ( .A(b[5]), .B(a[227]), .Z(n9362) );
  NAND U9607 ( .A(n10456), .B(n9362), .Z(n9322) );
  AND U9608 ( .A(n9323), .B(n9322), .Z(n9366) );
  AND U9609 ( .A(b[7]), .B(a[223]), .Z(n9365) );
  XNOR U9610 ( .A(n9366), .B(n9365), .Z(n9367) );
  XNOR U9611 ( .A(n9368), .B(n9367), .Z(n9373) );
  XOR U9612 ( .A(n9374), .B(n9373), .Z(n9348) );
  NANDN U9613 ( .A(n9325), .B(n9324), .Z(n9329) );
  NANDN U9614 ( .A(n9327), .B(n9326), .Z(n9328) );
  AND U9615 ( .A(n9329), .B(n9328), .Z(n9347) );
  XNOR U9616 ( .A(n9348), .B(n9347), .Z(n9349) );
  NANDN U9617 ( .A(n9331), .B(n9330), .Z(n9335) );
  NAND U9618 ( .A(n9333), .B(n9332), .Z(n9334) );
  NAND U9619 ( .A(n9335), .B(n9334), .Z(n9350) );
  XNOR U9620 ( .A(n9349), .B(n9350), .Z(n9341) );
  XNOR U9621 ( .A(n9342), .B(n9341), .Z(n9343) );
  XNOR U9622 ( .A(n9344), .B(n9343), .Z(n9377) );
  XNOR U9623 ( .A(sreg[479]), .B(n9377), .Z(n9379) );
  NANDN U9624 ( .A(sreg[478]), .B(n9336), .Z(n9340) );
  NAND U9625 ( .A(n9338), .B(n9337), .Z(n9339) );
  NAND U9626 ( .A(n9340), .B(n9339), .Z(n9378) );
  XNOR U9627 ( .A(n9379), .B(n9378), .Z(c[479]) );
  NANDN U9628 ( .A(n9342), .B(n9341), .Z(n9346) );
  NANDN U9629 ( .A(n9344), .B(n9343), .Z(n9345) );
  AND U9630 ( .A(n9346), .B(n9345), .Z(n9385) );
  NANDN U9631 ( .A(n9348), .B(n9347), .Z(n9352) );
  NANDN U9632 ( .A(n9350), .B(n9349), .Z(n9351) );
  AND U9633 ( .A(n9352), .B(n9351), .Z(n9383) );
  NAND U9634 ( .A(n26), .B(n9353), .Z(n9355) );
  XOR U9635 ( .A(b[7]), .B(a[226]), .Z(n9394) );
  NAND U9636 ( .A(n10531), .B(n9394), .Z(n9354) );
  AND U9637 ( .A(n9355), .B(n9354), .Z(n9413) );
  NAND U9638 ( .A(n23), .B(n9356), .Z(n9358) );
  XOR U9639 ( .A(b[3]), .B(a[230]), .Z(n9397) );
  NAND U9640 ( .A(n24), .B(n9397), .Z(n9357) );
  NAND U9641 ( .A(n9358), .B(n9357), .Z(n9412) );
  XNOR U9642 ( .A(n9413), .B(n9412), .Z(n9415) );
  NAND U9643 ( .A(b[0]), .B(a[232]), .Z(n9359) );
  XNOR U9644 ( .A(b[1]), .B(n9359), .Z(n9361) );
  NANDN U9645 ( .A(b[0]), .B(a[231]), .Z(n9360) );
  NAND U9646 ( .A(n9361), .B(n9360), .Z(n9409) );
  NAND U9647 ( .A(n25), .B(n9362), .Z(n9364) );
  XOR U9648 ( .A(b[5]), .B(a[228]), .Z(n9400) );
  NAND U9649 ( .A(n10456), .B(n9400), .Z(n9363) );
  AND U9650 ( .A(n9364), .B(n9363), .Z(n9407) );
  AND U9651 ( .A(b[7]), .B(a[224]), .Z(n9406) );
  XNOR U9652 ( .A(n9407), .B(n9406), .Z(n9408) );
  XNOR U9653 ( .A(n9409), .B(n9408), .Z(n9414) );
  XOR U9654 ( .A(n9415), .B(n9414), .Z(n9389) );
  NANDN U9655 ( .A(n9366), .B(n9365), .Z(n9370) );
  NANDN U9656 ( .A(n9368), .B(n9367), .Z(n9369) );
  AND U9657 ( .A(n9370), .B(n9369), .Z(n9388) );
  XNOR U9658 ( .A(n9389), .B(n9388), .Z(n9390) );
  NANDN U9659 ( .A(n9372), .B(n9371), .Z(n9376) );
  NAND U9660 ( .A(n9374), .B(n9373), .Z(n9375) );
  NAND U9661 ( .A(n9376), .B(n9375), .Z(n9391) );
  XNOR U9662 ( .A(n9390), .B(n9391), .Z(n9382) );
  XNOR U9663 ( .A(n9383), .B(n9382), .Z(n9384) );
  XNOR U9664 ( .A(n9385), .B(n9384), .Z(n9418) );
  XNOR U9665 ( .A(sreg[480]), .B(n9418), .Z(n9420) );
  NANDN U9666 ( .A(sreg[479]), .B(n9377), .Z(n9381) );
  NAND U9667 ( .A(n9379), .B(n9378), .Z(n9380) );
  NAND U9668 ( .A(n9381), .B(n9380), .Z(n9419) );
  XNOR U9669 ( .A(n9420), .B(n9419), .Z(c[480]) );
  NANDN U9670 ( .A(n9383), .B(n9382), .Z(n9387) );
  NANDN U9671 ( .A(n9385), .B(n9384), .Z(n9386) );
  AND U9672 ( .A(n9387), .B(n9386), .Z(n9426) );
  NANDN U9673 ( .A(n9389), .B(n9388), .Z(n9393) );
  NANDN U9674 ( .A(n9391), .B(n9390), .Z(n9392) );
  AND U9675 ( .A(n9393), .B(n9392), .Z(n9424) );
  NAND U9676 ( .A(n26), .B(n9394), .Z(n9396) );
  XOR U9677 ( .A(b[7]), .B(a[227]), .Z(n9435) );
  NAND U9678 ( .A(n10531), .B(n9435), .Z(n9395) );
  AND U9679 ( .A(n9396), .B(n9395), .Z(n9454) );
  NAND U9680 ( .A(n23), .B(n9397), .Z(n9399) );
  XOR U9681 ( .A(b[3]), .B(a[231]), .Z(n9438) );
  NAND U9682 ( .A(n24), .B(n9438), .Z(n9398) );
  NAND U9683 ( .A(n9399), .B(n9398), .Z(n9453) );
  XNOR U9684 ( .A(n9454), .B(n9453), .Z(n9456) );
  NAND U9685 ( .A(n25), .B(n9400), .Z(n9402) );
  XOR U9686 ( .A(b[5]), .B(a[229]), .Z(n9441) );
  NAND U9687 ( .A(n10456), .B(n9441), .Z(n9401) );
  AND U9688 ( .A(n9402), .B(n9401), .Z(n9448) );
  AND U9689 ( .A(b[7]), .B(a[225]), .Z(n9447) );
  XNOR U9690 ( .A(n9448), .B(n9447), .Z(n9449) );
  NAND U9691 ( .A(b[0]), .B(a[233]), .Z(n9403) );
  XNOR U9692 ( .A(b[1]), .B(n9403), .Z(n9405) );
  NANDN U9693 ( .A(b[0]), .B(a[232]), .Z(n9404) );
  NAND U9694 ( .A(n9405), .B(n9404), .Z(n9450) );
  XNOR U9695 ( .A(n9449), .B(n9450), .Z(n9455) );
  XOR U9696 ( .A(n9456), .B(n9455), .Z(n9430) );
  NANDN U9697 ( .A(n9407), .B(n9406), .Z(n9411) );
  NANDN U9698 ( .A(n9409), .B(n9408), .Z(n9410) );
  AND U9699 ( .A(n9411), .B(n9410), .Z(n9429) );
  XNOR U9700 ( .A(n9430), .B(n9429), .Z(n9431) );
  NANDN U9701 ( .A(n9413), .B(n9412), .Z(n9417) );
  NAND U9702 ( .A(n9415), .B(n9414), .Z(n9416) );
  NAND U9703 ( .A(n9417), .B(n9416), .Z(n9432) );
  XNOR U9704 ( .A(n9431), .B(n9432), .Z(n9423) );
  XNOR U9705 ( .A(n9424), .B(n9423), .Z(n9425) );
  XNOR U9706 ( .A(n9426), .B(n9425), .Z(n9459) );
  XNOR U9707 ( .A(sreg[481]), .B(n9459), .Z(n9461) );
  NANDN U9708 ( .A(sreg[480]), .B(n9418), .Z(n9422) );
  NAND U9709 ( .A(n9420), .B(n9419), .Z(n9421) );
  NAND U9710 ( .A(n9422), .B(n9421), .Z(n9460) );
  XNOR U9711 ( .A(n9461), .B(n9460), .Z(c[481]) );
  NANDN U9712 ( .A(n9424), .B(n9423), .Z(n9428) );
  NANDN U9713 ( .A(n9426), .B(n9425), .Z(n9427) );
  AND U9714 ( .A(n9428), .B(n9427), .Z(n9467) );
  NANDN U9715 ( .A(n9430), .B(n9429), .Z(n9434) );
  NANDN U9716 ( .A(n9432), .B(n9431), .Z(n9433) );
  AND U9717 ( .A(n9434), .B(n9433), .Z(n9465) );
  NAND U9718 ( .A(n26), .B(n9435), .Z(n9437) );
  XOR U9719 ( .A(b[7]), .B(a[228]), .Z(n9476) );
  NAND U9720 ( .A(n10531), .B(n9476), .Z(n9436) );
  AND U9721 ( .A(n9437), .B(n9436), .Z(n9495) );
  NAND U9722 ( .A(n23), .B(n9438), .Z(n9440) );
  XOR U9723 ( .A(b[3]), .B(a[232]), .Z(n9479) );
  NAND U9724 ( .A(n24), .B(n9479), .Z(n9439) );
  NAND U9725 ( .A(n9440), .B(n9439), .Z(n9494) );
  XNOR U9726 ( .A(n9495), .B(n9494), .Z(n9497) );
  NAND U9727 ( .A(n25), .B(n9441), .Z(n9443) );
  XOR U9728 ( .A(b[5]), .B(a[230]), .Z(n9485) );
  NAND U9729 ( .A(n10456), .B(n9485), .Z(n9442) );
  AND U9730 ( .A(n9443), .B(n9442), .Z(n9489) );
  AND U9731 ( .A(b[7]), .B(a[226]), .Z(n9488) );
  XNOR U9732 ( .A(n9489), .B(n9488), .Z(n9490) );
  NAND U9733 ( .A(b[0]), .B(a[234]), .Z(n9444) );
  XNOR U9734 ( .A(b[1]), .B(n9444), .Z(n9446) );
  NANDN U9735 ( .A(b[0]), .B(a[233]), .Z(n9445) );
  NAND U9736 ( .A(n9446), .B(n9445), .Z(n9491) );
  XNOR U9737 ( .A(n9490), .B(n9491), .Z(n9496) );
  XOR U9738 ( .A(n9497), .B(n9496), .Z(n9471) );
  NANDN U9739 ( .A(n9448), .B(n9447), .Z(n9452) );
  NANDN U9740 ( .A(n9450), .B(n9449), .Z(n9451) );
  AND U9741 ( .A(n9452), .B(n9451), .Z(n9470) );
  XNOR U9742 ( .A(n9471), .B(n9470), .Z(n9472) );
  NANDN U9743 ( .A(n9454), .B(n9453), .Z(n9458) );
  NAND U9744 ( .A(n9456), .B(n9455), .Z(n9457) );
  NAND U9745 ( .A(n9458), .B(n9457), .Z(n9473) );
  XNOR U9746 ( .A(n9472), .B(n9473), .Z(n9464) );
  XNOR U9747 ( .A(n9465), .B(n9464), .Z(n9466) );
  XNOR U9748 ( .A(n9467), .B(n9466), .Z(n9500) );
  XNOR U9749 ( .A(sreg[482]), .B(n9500), .Z(n9502) );
  NANDN U9750 ( .A(sreg[481]), .B(n9459), .Z(n9463) );
  NAND U9751 ( .A(n9461), .B(n9460), .Z(n9462) );
  NAND U9752 ( .A(n9463), .B(n9462), .Z(n9501) );
  XNOR U9753 ( .A(n9502), .B(n9501), .Z(c[482]) );
  NANDN U9754 ( .A(n9465), .B(n9464), .Z(n9469) );
  NANDN U9755 ( .A(n9467), .B(n9466), .Z(n9468) );
  AND U9756 ( .A(n9469), .B(n9468), .Z(n9508) );
  NANDN U9757 ( .A(n9471), .B(n9470), .Z(n9475) );
  NANDN U9758 ( .A(n9473), .B(n9472), .Z(n9474) );
  AND U9759 ( .A(n9475), .B(n9474), .Z(n9506) );
  NAND U9760 ( .A(n26), .B(n9476), .Z(n9478) );
  XOR U9761 ( .A(b[7]), .B(a[229]), .Z(n9517) );
  NAND U9762 ( .A(n10531), .B(n9517), .Z(n9477) );
  AND U9763 ( .A(n9478), .B(n9477), .Z(n9536) );
  NAND U9764 ( .A(n23), .B(n9479), .Z(n9481) );
  XOR U9765 ( .A(b[3]), .B(a[233]), .Z(n9520) );
  NAND U9766 ( .A(n24), .B(n9520), .Z(n9480) );
  NAND U9767 ( .A(n9481), .B(n9480), .Z(n9535) );
  XNOR U9768 ( .A(n9536), .B(n9535), .Z(n9538) );
  NAND U9769 ( .A(b[0]), .B(a[235]), .Z(n9482) );
  XNOR U9770 ( .A(b[1]), .B(n9482), .Z(n9484) );
  NANDN U9771 ( .A(b[0]), .B(a[234]), .Z(n9483) );
  NAND U9772 ( .A(n9484), .B(n9483), .Z(n9532) );
  NAND U9773 ( .A(n25), .B(n9485), .Z(n9487) );
  XOR U9774 ( .A(b[5]), .B(a[231]), .Z(n9526) );
  NAND U9775 ( .A(n10456), .B(n9526), .Z(n9486) );
  AND U9776 ( .A(n9487), .B(n9486), .Z(n9530) );
  AND U9777 ( .A(b[7]), .B(a[227]), .Z(n9529) );
  XNOR U9778 ( .A(n9530), .B(n9529), .Z(n9531) );
  XNOR U9779 ( .A(n9532), .B(n9531), .Z(n9537) );
  XOR U9780 ( .A(n9538), .B(n9537), .Z(n9512) );
  NANDN U9781 ( .A(n9489), .B(n9488), .Z(n9493) );
  NANDN U9782 ( .A(n9491), .B(n9490), .Z(n9492) );
  AND U9783 ( .A(n9493), .B(n9492), .Z(n9511) );
  XNOR U9784 ( .A(n9512), .B(n9511), .Z(n9513) );
  NANDN U9785 ( .A(n9495), .B(n9494), .Z(n9499) );
  NAND U9786 ( .A(n9497), .B(n9496), .Z(n9498) );
  NAND U9787 ( .A(n9499), .B(n9498), .Z(n9514) );
  XNOR U9788 ( .A(n9513), .B(n9514), .Z(n9505) );
  XNOR U9789 ( .A(n9506), .B(n9505), .Z(n9507) );
  XNOR U9790 ( .A(n9508), .B(n9507), .Z(n9541) );
  XNOR U9791 ( .A(sreg[483]), .B(n9541), .Z(n9543) );
  NANDN U9792 ( .A(sreg[482]), .B(n9500), .Z(n9504) );
  NAND U9793 ( .A(n9502), .B(n9501), .Z(n9503) );
  NAND U9794 ( .A(n9504), .B(n9503), .Z(n9542) );
  XNOR U9795 ( .A(n9543), .B(n9542), .Z(c[483]) );
  NANDN U9796 ( .A(n9506), .B(n9505), .Z(n9510) );
  NANDN U9797 ( .A(n9508), .B(n9507), .Z(n9509) );
  AND U9798 ( .A(n9510), .B(n9509), .Z(n9549) );
  NANDN U9799 ( .A(n9512), .B(n9511), .Z(n9516) );
  NANDN U9800 ( .A(n9514), .B(n9513), .Z(n9515) );
  AND U9801 ( .A(n9516), .B(n9515), .Z(n9547) );
  NAND U9802 ( .A(n26), .B(n9517), .Z(n9519) );
  XOR U9803 ( .A(b[7]), .B(a[230]), .Z(n9558) );
  NAND U9804 ( .A(n10531), .B(n9558), .Z(n9518) );
  AND U9805 ( .A(n9519), .B(n9518), .Z(n9577) );
  NAND U9806 ( .A(n23), .B(n9520), .Z(n9522) );
  XOR U9807 ( .A(b[3]), .B(a[234]), .Z(n9561) );
  NAND U9808 ( .A(n24), .B(n9561), .Z(n9521) );
  NAND U9809 ( .A(n9522), .B(n9521), .Z(n9576) );
  XNOR U9810 ( .A(n9577), .B(n9576), .Z(n9579) );
  NAND U9811 ( .A(b[0]), .B(a[236]), .Z(n9523) );
  XNOR U9812 ( .A(b[1]), .B(n9523), .Z(n9525) );
  NANDN U9813 ( .A(b[0]), .B(a[235]), .Z(n9524) );
  NAND U9814 ( .A(n9525), .B(n9524), .Z(n9573) );
  NAND U9815 ( .A(n25), .B(n9526), .Z(n9528) );
  XOR U9816 ( .A(b[5]), .B(a[232]), .Z(n9564) );
  NAND U9817 ( .A(n10456), .B(n9564), .Z(n9527) );
  AND U9818 ( .A(n9528), .B(n9527), .Z(n9571) );
  AND U9819 ( .A(b[7]), .B(a[228]), .Z(n9570) );
  XNOR U9820 ( .A(n9571), .B(n9570), .Z(n9572) );
  XNOR U9821 ( .A(n9573), .B(n9572), .Z(n9578) );
  XOR U9822 ( .A(n9579), .B(n9578), .Z(n9553) );
  NANDN U9823 ( .A(n9530), .B(n9529), .Z(n9534) );
  NANDN U9824 ( .A(n9532), .B(n9531), .Z(n9533) );
  AND U9825 ( .A(n9534), .B(n9533), .Z(n9552) );
  XNOR U9826 ( .A(n9553), .B(n9552), .Z(n9554) );
  NANDN U9827 ( .A(n9536), .B(n9535), .Z(n9540) );
  NAND U9828 ( .A(n9538), .B(n9537), .Z(n9539) );
  NAND U9829 ( .A(n9540), .B(n9539), .Z(n9555) );
  XNOR U9830 ( .A(n9554), .B(n9555), .Z(n9546) );
  XNOR U9831 ( .A(n9547), .B(n9546), .Z(n9548) );
  XNOR U9832 ( .A(n9549), .B(n9548), .Z(n9582) );
  XNOR U9833 ( .A(sreg[484]), .B(n9582), .Z(n9584) );
  NANDN U9834 ( .A(sreg[483]), .B(n9541), .Z(n9545) );
  NAND U9835 ( .A(n9543), .B(n9542), .Z(n9544) );
  NAND U9836 ( .A(n9545), .B(n9544), .Z(n9583) );
  XNOR U9837 ( .A(n9584), .B(n9583), .Z(c[484]) );
  NANDN U9838 ( .A(n9547), .B(n9546), .Z(n9551) );
  NANDN U9839 ( .A(n9549), .B(n9548), .Z(n9550) );
  AND U9840 ( .A(n9551), .B(n9550), .Z(n9590) );
  NANDN U9841 ( .A(n9553), .B(n9552), .Z(n9557) );
  NANDN U9842 ( .A(n9555), .B(n9554), .Z(n9556) );
  AND U9843 ( .A(n9557), .B(n9556), .Z(n9588) );
  NAND U9844 ( .A(n26), .B(n9558), .Z(n9560) );
  XOR U9845 ( .A(b[7]), .B(a[231]), .Z(n9599) );
  NAND U9846 ( .A(n10531), .B(n9599), .Z(n9559) );
  AND U9847 ( .A(n9560), .B(n9559), .Z(n9618) );
  NAND U9848 ( .A(n23), .B(n9561), .Z(n9563) );
  XOR U9849 ( .A(b[3]), .B(a[235]), .Z(n9602) );
  NAND U9850 ( .A(n24), .B(n9602), .Z(n9562) );
  NAND U9851 ( .A(n9563), .B(n9562), .Z(n9617) );
  XNOR U9852 ( .A(n9618), .B(n9617), .Z(n9620) );
  NAND U9853 ( .A(n25), .B(n9564), .Z(n9566) );
  XOR U9854 ( .A(b[5]), .B(a[233]), .Z(n9608) );
  NAND U9855 ( .A(n10456), .B(n9608), .Z(n9565) );
  AND U9856 ( .A(n9566), .B(n9565), .Z(n9612) );
  AND U9857 ( .A(b[7]), .B(a[229]), .Z(n9611) );
  XNOR U9858 ( .A(n9612), .B(n9611), .Z(n9613) );
  NAND U9859 ( .A(b[0]), .B(a[237]), .Z(n9567) );
  XNOR U9860 ( .A(b[1]), .B(n9567), .Z(n9569) );
  NANDN U9861 ( .A(b[0]), .B(a[236]), .Z(n9568) );
  NAND U9862 ( .A(n9569), .B(n9568), .Z(n9614) );
  XNOR U9863 ( .A(n9613), .B(n9614), .Z(n9619) );
  XOR U9864 ( .A(n9620), .B(n9619), .Z(n9594) );
  NANDN U9865 ( .A(n9571), .B(n9570), .Z(n9575) );
  NANDN U9866 ( .A(n9573), .B(n9572), .Z(n9574) );
  AND U9867 ( .A(n9575), .B(n9574), .Z(n9593) );
  XNOR U9868 ( .A(n9594), .B(n9593), .Z(n9595) );
  NANDN U9869 ( .A(n9577), .B(n9576), .Z(n9581) );
  NAND U9870 ( .A(n9579), .B(n9578), .Z(n9580) );
  NAND U9871 ( .A(n9581), .B(n9580), .Z(n9596) );
  XNOR U9872 ( .A(n9595), .B(n9596), .Z(n9587) );
  XNOR U9873 ( .A(n9588), .B(n9587), .Z(n9589) );
  XNOR U9874 ( .A(n9590), .B(n9589), .Z(n9623) );
  XNOR U9875 ( .A(sreg[485]), .B(n9623), .Z(n9625) );
  NANDN U9876 ( .A(sreg[484]), .B(n9582), .Z(n9586) );
  NAND U9877 ( .A(n9584), .B(n9583), .Z(n9585) );
  NAND U9878 ( .A(n9586), .B(n9585), .Z(n9624) );
  XNOR U9879 ( .A(n9625), .B(n9624), .Z(c[485]) );
  NANDN U9880 ( .A(n9588), .B(n9587), .Z(n9592) );
  NANDN U9881 ( .A(n9590), .B(n9589), .Z(n9591) );
  AND U9882 ( .A(n9592), .B(n9591), .Z(n9631) );
  NANDN U9883 ( .A(n9594), .B(n9593), .Z(n9598) );
  NANDN U9884 ( .A(n9596), .B(n9595), .Z(n9597) );
  AND U9885 ( .A(n9598), .B(n9597), .Z(n9629) );
  NAND U9886 ( .A(n26), .B(n9599), .Z(n9601) );
  XOR U9887 ( .A(b[7]), .B(a[232]), .Z(n9640) );
  NAND U9888 ( .A(n10531), .B(n9640), .Z(n9600) );
  AND U9889 ( .A(n9601), .B(n9600), .Z(n9659) );
  NAND U9890 ( .A(n23), .B(n9602), .Z(n9604) );
  XOR U9891 ( .A(b[3]), .B(a[236]), .Z(n9643) );
  NAND U9892 ( .A(n24), .B(n9643), .Z(n9603) );
  NAND U9893 ( .A(n9604), .B(n9603), .Z(n9658) );
  XNOR U9894 ( .A(n9659), .B(n9658), .Z(n9661) );
  NAND U9895 ( .A(b[0]), .B(a[238]), .Z(n9605) );
  XNOR U9896 ( .A(b[1]), .B(n9605), .Z(n9607) );
  NANDN U9897 ( .A(b[0]), .B(a[237]), .Z(n9606) );
  NAND U9898 ( .A(n9607), .B(n9606), .Z(n9655) );
  NAND U9899 ( .A(n25), .B(n9608), .Z(n9610) );
  XOR U9900 ( .A(b[5]), .B(a[234]), .Z(n9649) );
  NAND U9901 ( .A(n10456), .B(n9649), .Z(n9609) );
  AND U9902 ( .A(n9610), .B(n9609), .Z(n9653) );
  AND U9903 ( .A(b[7]), .B(a[230]), .Z(n9652) );
  XNOR U9904 ( .A(n9653), .B(n9652), .Z(n9654) );
  XNOR U9905 ( .A(n9655), .B(n9654), .Z(n9660) );
  XOR U9906 ( .A(n9661), .B(n9660), .Z(n9635) );
  NANDN U9907 ( .A(n9612), .B(n9611), .Z(n9616) );
  NANDN U9908 ( .A(n9614), .B(n9613), .Z(n9615) );
  AND U9909 ( .A(n9616), .B(n9615), .Z(n9634) );
  XNOR U9910 ( .A(n9635), .B(n9634), .Z(n9636) );
  NANDN U9911 ( .A(n9618), .B(n9617), .Z(n9622) );
  NAND U9912 ( .A(n9620), .B(n9619), .Z(n9621) );
  NAND U9913 ( .A(n9622), .B(n9621), .Z(n9637) );
  XNOR U9914 ( .A(n9636), .B(n9637), .Z(n9628) );
  XNOR U9915 ( .A(n9629), .B(n9628), .Z(n9630) );
  XNOR U9916 ( .A(n9631), .B(n9630), .Z(n9664) );
  XNOR U9917 ( .A(sreg[486]), .B(n9664), .Z(n9666) );
  NANDN U9918 ( .A(sreg[485]), .B(n9623), .Z(n9627) );
  NAND U9919 ( .A(n9625), .B(n9624), .Z(n9626) );
  NAND U9920 ( .A(n9627), .B(n9626), .Z(n9665) );
  XNOR U9921 ( .A(n9666), .B(n9665), .Z(c[486]) );
  NANDN U9922 ( .A(n9629), .B(n9628), .Z(n9633) );
  NANDN U9923 ( .A(n9631), .B(n9630), .Z(n9632) );
  AND U9924 ( .A(n9633), .B(n9632), .Z(n9672) );
  NANDN U9925 ( .A(n9635), .B(n9634), .Z(n9639) );
  NANDN U9926 ( .A(n9637), .B(n9636), .Z(n9638) );
  AND U9927 ( .A(n9639), .B(n9638), .Z(n9670) );
  NAND U9928 ( .A(n26), .B(n9640), .Z(n9642) );
  XOR U9929 ( .A(b[7]), .B(a[233]), .Z(n9681) );
  NAND U9930 ( .A(n10531), .B(n9681), .Z(n9641) );
  AND U9931 ( .A(n9642), .B(n9641), .Z(n9700) );
  NAND U9932 ( .A(n23), .B(n9643), .Z(n9645) );
  XOR U9933 ( .A(b[3]), .B(a[237]), .Z(n9684) );
  NAND U9934 ( .A(n24), .B(n9684), .Z(n9644) );
  NAND U9935 ( .A(n9645), .B(n9644), .Z(n9699) );
  XNOR U9936 ( .A(n9700), .B(n9699), .Z(n9702) );
  NAND U9937 ( .A(b[0]), .B(a[239]), .Z(n9646) );
  XNOR U9938 ( .A(b[1]), .B(n9646), .Z(n9648) );
  NANDN U9939 ( .A(b[0]), .B(a[238]), .Z(n9647) );
  NAND U9940 ( .A(n9648), .B(n9647), .Z(n9696) );
  NAND U9941 ( .A(n25), .B(n9649), .Z(n9651) );
  XOR U9942 ( .A(b[5]), .B(a[235]), .Z(n9690) );
  NAND U9943 ( .A(n10456), .B(n9690), .Z(n9650) );
  AND U9944 ( .A(n9651), .B(n9650), .Z(n9694) );
  AND U9945 ( .A(b[7]), .B(a[231]), .Z(n9693) );
  XNOR U9946 ( .A(n9694), .B(n9693), .Z(n9695) );
  XNOR U9947 ( .A(n9696), .B(n9695), .Z(n9701) );
  XOR U9948 ( .A(n9702), .B(n9701), .Z(n9676) );
  NANDN U9949 ( .A(n9653), .B(n9652), .Z(n9657) );
  NANDN U9950 ( .A(n9655), .B(n9654), .Z(n9656) );
  AND U9951 ( .A(n9657), .B(n9656), .Z(n9675) );
  XNOR U9952 ( .A(n9676), .B(n9675), .Z(n9677) );
  NANDN U9953 ( .A(n9659), .B(n9658), .Z(n9663) );
  NAND U9954 ( .A(n9661), .B(n9660), .Z(n9662) );
  NAND U9955 ( .A(n9663), .B(n9662), .Z(n9678) );
  XNOR U9956 ( .A(n9677), .B(n9678), .Z(n9669) );
  XNOR U9957 ( .A(n9670), .B(n9669), .Z(n9671) );
  XNOR U9958 ( .A(n9672), .B(n9671), .Z(n9705) );
  XNOR U9959 ( .A(sreg[487]), .B(n9705), .Z(n9707) );
  NANDN U9960 ( .A(sreg[486]), .B(n9664), .Z(n9668) );
  NAND U9961 ( .A(n9666), .B(n9665), .Z(n9667) );
  NAND U9962 ( .A(n9668), .B(n9667), .Z(n9706) );
  XNOR U9963 ( .A(n9707), .B(n9706), .Z(c[487]) );
  NANDN U9964 ( .A(n9670), .B(n9669), .Z(n9674) );
  NANDN U9965 ( .A(n9672), .B(n9671), .Z(n9673) );
  AND U9966 ( .A(n9674), .B(n9673), .Z(n9713) );
  NANDN U9967 ( .A(n9676), .B(n9675), .Z(n9680) );
  NANDN U9968 ( .A(n9678), .B(n9677), .Z(n9679) );
  AND U9969 ( .A(n9680), .B(n9679), .Z(n9711) );
  NAND U9970 ( .A(n26), .B(n9681), .Z(n9683) );
  XOR U9971 ( .A(b[7]), .B(a[234]), .Z(n9722) );
  NAND U9972 ( .A(n10531), .B(n9722), .Z(n9682) );
  AND U9973 ( .A(n9683), .B(n9682), .Z(n9741) );
  NAND U9974 ( .A(n23), .B(n9684), .Z(n9686) );
  XOR U9975 ( .A(b[3]), .B(a[238]), .Z(n9725) );
  NAND U9976 ( .A(n24), .B(n9725), .Z(n9685) );
  NAND U9977 ( .A(n9686), .B(n9685), .Z(n9740) );
  XNOR U9978 ( .A(n9741), .B(n9740), .Z(n9743) );
  NAND U9979 ( .A(b[0]), .B(a[240]), .Z(n9687) );
  XNOR U9980 ( .A(b[1]), .B(n9687), .Z(n9689) );
  NANDN U9981 ( .A(b[0]), .B(a[239]), .Z(n9688) );
  NAND U9982 ( .A(n9689), .B(n9688), .Z(n9737) );
  NAND U9983 ( .A(n25), .B(n9690), .Z(n9692) );
  XOR U9984 ( .A(b[5]), .B(a[236]), .Z(n9728) );
  NAND U9985 ( .A(n10456), .B(n9728), .Z(n9691) );
  AND U9986 ( .A(n9692), .B(n9691), .Z(n9735) );
  AND U9987 ( .A(b[7]), .B(a[232]), .Z(n9734) );
  XNOR U9988 ( .A(n9735), .B(n9734), .Z(n9736) );
  XNOR U9989 ( .A(n9737), .B(n9736), .Z(n9742) );
  XOR U9990 ( .A(n9743), .B(n9742), .Z(n9717) );
  NANDN U9991 ( .A(n9694), .B(n9693), .Z(n9698) );
  NANDN U9992 ( .A(n9696), .B(n9695), .Z(n9697) );
  AND U9993 ( .A(n9698), .B(n9697), .Z(n9716) );
  XNOR U9994 ( .A(n9717), .B(n9716), .Z(n9718) );
  NANDN U9995 ( .A(n9700), .B(n9699), .Z(n9704) );
  NAND U9996 ( .A(n9702), .B(n9701), .Z(n9703) );
  NAND U9997 ( .A(n9704), .B(n9703), .Z(n9719) );
  XNOR U9998 ( .A(n9718), .B(n9719), .Z(n9710) );
  XNOR U9999 ( .A(n9711), .B(n9710), .Z(n9712) );
  XNOR U10000 ( .A(n9713), .B(n9712), .Z(n9746) );
  XNOR U10001 ( .A(sreg[488]), .B(n9746), .Z(n9748) );
  NANDN U10002 ( .A(sreg[487]), .B(n9705), .Z(n9709) );
  NAND U10003 ( .A(n9707), .B(n9706), .Z(n9708) );
  NAND U10004 ( .A(n9709), .B(n9708), .Z(n9747) );
  XNOR U10005 ( .A(n9748), .B(n9747), .Z(c[488]) );
  NANDN U10006 ( .A(n9711), .B(n9710), .Z(n9715) );
  NANDN U10007 ( .A(n9713), .B(n9712), .Z(n9714) );
  AND U10008 ( .A(n9715), .B(n9714), .Z(n9758) );
  NANDN U10009 ( .A(n9717), .B(n9716), .Z(n9721) );
  NANDN U10010 ( .A(n9719), .B(n9718), .Z(n9720) );
  AND U10011 ( .A(n9721), .B(n9720), .Z(n9757) );
  NAND U10012 ( .A(n26), .B(n9722), .Z(n9724) );
  XOR U10013 ( .A(b[7]), .B(a[235]), .Z(n9768) );
  NAND U10014 ( .A(n10531), .B(n9768), .Z(n9723) );
  AND U10015 ( .A(n9724), .B(n9723), .Z(n9787) );
  NAND U10016 ( .A(n23), .B(n9725), .Z(n9727) );
  XOR U10017 ( .A(b[3]), .B(a[239]), .Z(n9771) );
  NAND U10018 ( .A(n24), .B(n9771), .Z(n9726) );
  NAND U10019 ( .A(n9727), .B(n9726), .Z(n9786) );
  XNOR U10020 ( .A(n9787), .B(n9786), .Z(n9789) );
  NAND U10021 ( .A(n25), .B(n9728), .Z(n9730) );
  XOR U10022 ( .A(b[5]), .B(a[237]), .Z(n9777) );
  NAND U10023 ( .A(n10456), .B(n9777), .Z(n9729) );
  AND U10024 ( .A(n9730), .B(n9729), .Z(n9781) );
  AND U10025 ( .A(b[7]), .B(a[233]), .Z(n9780) );
  XNOR U10026 ( .A(n9781), .B(n9780), .Z(n9782) );
  NAND U10027 ( .A(b[0]), .B(a[241]), .Z(n9731) );
  XNOR U10028 ( .A(b[1]), .B(n9731), .Z(n9733) );
  NANDN U10029 ( .A(b[0]), .B(a[240]), .Z(n9732) );
  NAND U10030 ( .A(n9733), .B(n9732), .Z(n9783) );
  XNOR U10031 ( .A(n9782), .B(n9783), .Z(n9788) );
  XOR U10032 ( .A(n9789), .B(n9788), .Z(n9763) );
  NANDN U10033 ( .A(n9735), .B(n9734), .Z(n9739) );
  NANDN U10034 ( .A(n9737), .B(n9736), .Z(n9738) );
  AND U10035 ( .A(n9739), .B(n9738), .Z(n9762) );
  XNOR U10036 ( .A(n9763), .B(n9762), .Z(n9764) );
  NANDN U10037 ( .A(n9741), .B(n9740), .Z(n9745) );
  NAND U10038 ( .A(n9743), .B(n9742), .Z(n9744) );
  NAND U10039 ( .A(n9745), .B(n9744), .Z(n9765) );
  XNOR U10040 ( .A(n9764), .B(n9765), .Z(n9756) );
  XOR U10041 ( .A(n9757), .B(n9756), .Z(n9759) );
  XOR U10042 ( .A(n9758), .B(n9759), .Z(n9751) );
  XNOR U10043 ( .A(n9751), .B(sreg[489]), .Z(n9753) );
  NANDN U10044 ( .A(sreg[488]), .B(n9746), .Z(n9750) );
  NAND U10045 ( .A(n9748), .B(n9747), .Z(n9749) );
  AND U10046 ( .A(n9750), .B(n9749), .Z(n9752) );
  XOR U10047 ( .A(n9753), .B(n9752), .Z(c[489]) );
  NANDN U10048 ( .A(n9751), .B(sreg[489]), .Z(n9755) );
  NAND U10049 ( .A(n9753), .B(n9752), .Z(n9754) );
  AND U10050 ( .A(n9755), .B(n9754), .Z(n9830) );
  NANDN U10051 ( .A(n9757), .B(n9756), .Z(n9761) );
  OR U10052 ( .A(n9759), .B(n9758), .Z(n9760) );
  AND U10053 ( .A(n9761), .B(n9760), .Z(n9795) );
  NANDN U10054 ( .A(n9763), .B(n9762), .Z(n9767) );
  NANDN U10055 ( .A(n9765), .B(n9764), .Z(n9766) );
  AND U10056 ( .A(n9767), .B(n9766), .Z(n9793) );
  NAND U10057 ( .A(n26), .B(n9768), .Z(n9770) );
  XOR U10058 ( .A(b[7]), .B(a[236]), .Z(n9804) );
  NAND U10059 ( .A(n10531), .B(n9804), .Z(n9769) );
  AND U10060 ( .A(n9770), .B(n9769), .Z(n9823) );
  NAND U10061 ( .A(n23), .B(n9771), .Z(n9773) );
  XOR U10062 ( .A(b[3]), .B(a[240]), .Z(n9807) );
  NAND U10063 ( .A(n24), .B(n9807), .Z(n9772) );
  NAND U10064 ( .A(n9773), .B(n9772), .Z(n9822) );
  XNOR U10065 ( .A(n9823), .B(n9822), .Z(n9825) );
  NAND U10066 ( .A(b[0]), .B(a[242]), .Z(n9774) );
  XNOR U10067 ( .A(b[1]), .B(n9774), .Z(n9776) );
  NANDN U10068 ( .A(b[0]), .B(a[241]), .Z(n9775) );
  NAND U10069 ( .A(n9776), .B(n9775), .Z(n9819) );
  NAND U10070 ( .A(n25), .B(n9777), .Z(n9779) );
  XOR U10071 ( .A(b[5]), .B(a[238]), .Z(n9810) );
  NAND U10072 ( .A(n10456), .B(n9810), .Z(n9778) );
  AND U10073 ( .A(n9779), .B(n9778), .Z(n9817) );
  AND U10074 ( .A(b[7]), .B(a[234]), .Z(n9816) );
  XNOR U10075 ( .A(n9817), .B(n9816), .Z(n9818) );
  XNOR U10076 ( .A(n9819), .B(n9818), .Z(n9824) );
  XOR U10077 ( .A(n9825), .B(n9824), .Z(n9799) );
  NANDN U10078 ( .A(n9781), .B(n9780), .Z(n9785) );
  NANDN U10079 ( .A(n9783), .B(n9782), .Z(n9784) );
  AND U10080 ( .A(n9785), .B(n9784), .Z(n9798) );
  XNOR U10081 ( .A(n9799), .B(n9798), .Z(n9800) );
  NANDN U10082 ( .A(n9787), .B(n9786), .Z(n9791) );
  NAND U10083 ( .A(n9789), .B(n9788), .Z(n9790) );
  NAND U10084 ( .A(n9791), .B(n9790), .Z(n9801) );
  XNOR U10085 ( .A(n9800), .B(n9801), .Z(n9792) );
  XNOR U10086 ( .A(n9793), .B(n9792), .Z(n9794) );
  XNOR U10087 ( .A(n9795), .B(n9794), .Z(n9828) );
  XNOR U10088 ( .A(sreg[490]), .B(n9828), .Z(n9829) );
  XNOR U10089 ( .A(n9830), .B(n9829), .Z(c[490]) );
  NANDN U10090 ( .A(n9793), .B(n9792), .Z(n9797) );
  NANDN U10091 ( .A(n9795), .B(n9794), .Z(n9796) );
  AND U10092 ( .A(n9797), .B(n9796), .Z(n9836) );
  NANDN U10093 ( .A(n9799), .B(n9798), .Z(n9803) );
  NANDN U10094 ( .A(n9801), .B(n9800), .Z(n9802) );
  AND U10095 ( .A(n9803), .B(n9802), .Z(n9834) );
  NAND U10096 ( .A(n26), .B(n9804), .Z(n9806) );
  XOR U10097 ( .A(b[7]), .B(a[237]), .Z(n9845) );
  NAND U10098 ( .A(n10531), .B(n9845), .Z(n9805) );
  AND U10099 ( .A(n9806), .B(n9805), .Z(n9864) );
  NAND U10100 ( .A(n23), .B(n9807), .Z(n9809) );
  XOR U10101 ( .A(b[3]), .B(a[241]), .Z(n9848) );
  NAND U10102 ( .A(n24), .B(n9848), .Z(n9808) );
  NAND U10103 ( .A(n9809), .B(n9808), .Z(n9863) );
  XNOR U10104 ( .A(n9864), .B(n9863), .Z(n9866) );
  NAND U10105 ( .A(n25), .B(n9810), .Z(n9812) );
  XOR U10106 ( .A(b[5]), .B(a[239]), .Z(n9854) );
  NAND U10107 ( .A(n10456), .B(n9854), .Z(n9811) );
  AND U10108 ( .A(n9812), .B(n9811), .Z(n9858) );
  AND U10109 ( .A(b[7]), .B(a[235]), .Z(n9857) );
  XNOR U10110 ( .A(n9858), .B(n9857), .Z(n9859) );
  NAND U10111 ( .A(b[0]), .B(a[243]), .Z(n9813) );
  XNOR U10112 ( .A(b[1]), .B(n9813), .Z(n9815) );
  NANDN U10113 ( .A(b[0]), .B(a[242]), .Z(n9814) );
  NAND U10114 ( .A(n9815), .B(n9814), .Z(n9860) );
  XNOR U10115 ( .A(n9859), .B(n9860), .Z(n9865) );
  XOR U10116 ( .A(n9866), .B(n9865), .Z(n9840) );
  NANDN U10117 ( .A(n9817), .B(n9816), .Z(n9821) );
  NANDN U10118 ( .A(n9819), .B(n9818), .Z(n9820) );
  AND U10119 ( .A(n9821), .B(n9820), .Z(n9839) );
  XNOR U10120 ( .A(n9840), .B(n9839), .Z(n9841) );
  NANDN U10121 ( .A(n9823), .B(n9822), .Z(n9827) );
  NAND U10122 ( .A(n9825), .B(n9824), .Z(n9826) );
  NAND U10123 ( .A(n9827), .B(n9826), .Z(n9842) );
  XNOR U10124 ( .A(n9841), .B(n9842), .Z(n9833) );
  XNOR U10125 ( .A(n9834), .B(n9833), .Z(n9835) );
  XNOR U10126 ( .A(n9836), .B(n9835), .Z(n9869) );
  XNOR U10127 ( .A(sreg[491]), .B(n9869), .Z(n9871) );
  NANDN U10128 ( .A(sreg[490]), .B(n9828), .Z(n9832) );
  NAND U10129 ( .A(n9830), .B(n9829), .Z(n9831) );
  NAND U10130 ( .A(n9832), .B(n9831), .Z(n9870) );
  XNOR U10131 ( .A(n9871), .B(n9870), .Z(c[491]) );
  NANDN U10132 ( .A(n9834), .B(n9833), .Z(n9838) );
  NANDN U10133 ( .A(n9836), .B(n9835), .Z(n9837) );
  AND U10134 ( .A(n9838), .B(n9837), .Z(n9877) );
  NANDN U10135 ( .A(n9840), .B(n9839), .Z(n9844) );
  NANDN U10136 ( .A(n9842), .B(n9841), .Z(n9843) );
  AND U10137 ( .A(n9844), .B(n9843), .Z(n9875) );
  NAND U10138 ( .A(n26), .B(n9845), .Z(n9847) );
  XOR U10139 ( .A(b[7]), .B(a[238]), .Z(n9886) );
  NAND U10140 ( .A(n10531), .B(n9886), .Z(n9846) );
  AND U10141 ( .A(n9847), .B(n9846), .Z(n9905) );
  NAND U10142 ( .A(n23), .B(n9848), .Z(n9850) );
  XOR U10143 ( .A(b[3]), .B(a[242]), .Z(n9889) );
  NAND U10144 ( .A(n24), .B(n9889), .Z(n9849) );
  NAND U10145 ( .A(n9850), .B(n9849), .Z(n9904) );
  XNOR U10146 ( .A(n9905), .B(n9904), .Z(n9907) );
  NAND U10147 ( .A(b[0]), .B(a[244]), .Z(n9851) );
  XNOR U10148 ( .A(b[1]), .B(n9851), .Z(n9853) );
  NANDN U10149 ( .A(b[0]), .B(a[243]), .Z(n9852) );
  NAND U10150 ( .A(n9853), .B(n9852), .Z(n9901) );
  NAND U10151 ( .A(n25), .B(n9854), .Z(n9856) );
  XOR U10152 ( .A(b[5]), .B(a[240]), .Z(n9895) );
  NAND U10153 ( .A(n10456), .B(n9895), .Z(n9855) );
  AND U10154 ( .A(n9856), .B(n9855), .Z(n9899) );
  AND U10155 ( .A(b[7]), .B(a[236]), .Z(n9898) );
  XNOR U10156 ( .A(n9899), .B(n9898), .Z(n9900) );
  XNOR U10157 ( .A(n9901), .B(n9900), .Z(n9906) );
  XOR U10158 ( .A(n9907), .B(n9906), .Z(n9881) );
  NANDN U10159 ( .A(n9858), .B(n9857), .Z(n9862) );
  NANDN U10160 ( .A(n9860), .B(n9859), .Z(n9861) );
  AND U10161 ( .A(n9862), .B(n9861), .Z(n9880) );
  XNOR U10162 ( .A(n9881), .B(n9880), .Z(n9882) );
  NANDN U10163 ( .A(n9864), .B(n9863), .Z(n9868) );
  NAND U10164 ( .A(n9866), .B(n9865), .Z(n9867) );
  NAND U10165 ( .A(n9868), .B(n9867), .Z(n9883) );
  XNOR U10166 ( .A(n9882), .B(n9883), .Z(n9874) );
  XNOR U10167 ( .A(n9875), .B(n9874), .Z(n9876) );
  XNOR U10168 ( .A(n9877), .B(n9876), .Z(n9910) );
  XNOR U10169 ( .A(sreg[492]), .B(n9910), .Z(n9912) );
  NANDN U10170 ( .A(sreg[491]), .B(n9869), .Z(n9873) );
  NAND U10171 ( .A(n9871), .B(n9870), .Z(n9872) );
  NAND U10172 ( .A(n9873), .B(n9872), .Z(n9911) );
  XNOR U10173 ( .A(n9912), .B(n9911), .Z(c[492]) );
  NANDN U10174 ( .A(n9875), .B(n9874), .Z(n9879) );
  NANDN U10175 ( .A(n9877), .B(n9876), .Z(n9878) );
  AND U10176 ( .A(n9879), .B(n9878), .Z(n9918) );
  NANDN U10177 ( .A(n9881), .B(n9880), .Z(n9885) );
  NANDN U10178 ( .A(n9883), .B(n9882), .Z(n9884) );
  AND U10179 ( .A(n9885), .B(n9884), .Z(n9916) );
  NAND U10180 ( .A(n26), .B(n9886), .Z(n9888) );
  XOR U10181 ( .A(b[7]), .B(a[239]), .Z(n9927) );
  NAND U10182 ( .A(n10531), .B(n9927), .Z(n9887) );
  AND U10183 ( .A(n9888), .B(n9887), .Z(n9946) );
  NAND U10184 ( .A(n23), .B(n9889), .Z(n9891) );
  XOR U10185 ( .A(b[3]), .B(a[243]), .Z(n9930) );
  NAND U10186 ( .A(n24), .B(n9930), .Z(n9890) );
  NAND U10187 ( .A(n9891), .B(n9890), .Z(n9945) );
  XNOR U10188 ( .A(n9946), .B(n9945), .Z(n9948) );
  NAND U10189 ( .A(b[0]), .B(a[245]), .Z(n9892) );
  XNOR U10190 ( .A(b[1]), .B(n9892), .Z(n9894) );
  NANDN U10191 ( .A(b[0]), .B(a[244]), .Z(n9893) );
  NAND U10192 ( .A(n9894), .B(n9893), .Z(n9942) );
  NAND U10193 ( .A(n25), .B(n9895), .Z(n9897) );
  XOR U10194 ( .A(b[5]), .B(a[241]), .Z(n9936) );
  NAND U10195 ( .A(n10456), .B(n9936), .Z(n9896) );
  AND U10196 ( .A(n9897), .B(n9896), .Z(n9940) );
  AND U10197 ( .A(b[7]), .B(a[237]), .Z(n9939) );
  XNOR U10198 ( .A(n9940), .B(n9939), .Z(n9941) );
  XNOR U10199 ( .A(n9942), .B(n9941), .Z(n9947) );
  XOR U10200 ( .A(n9948), .B(n9947), .Z(n9922) );
  NANDN U10201 ( .A(n9899), .B(n9898), .Z(n9903) );
  NANDN U10202 ( .A(n9901), .B(n9900), .Z(n9902) );
  AND U10203 ( .A(n9903), .B(n9902), .Z(n9921) );
  XNOR U10204 ( .A(n9922), .B(n9921), .Z(n9923) );
  NANDN U10205 ( .A(n9905), .B(n9904), .Z(n9909) );
  NAND U10206 ( .A(n9907), .B(n9906), .Z(n9908) );
  NAND U10207 ( .A(n9909), .B(n9908), .Z(n9924) );
  XNOR U10208 ( .A(n9923), .B(n9924), .Z(n9915) );
  XNOR U10209 ( .A(n9916), .B(n9915), .Z(n9917) );
  XNOR U10210 ( .A(n9918), .B(n9917), .Z(n9951) );
  XNOR U10211 ( .A(sreg[493]), .B(n9951), .Z(n9953) );
  NANDN U10212 ( .A(sreg[492]), .B(n9910), .Z(n9914) );
  NAND U10213 ( .A(n9912), .B(n9911), .Z(n9913) );
  NAND U10214 ( .A(n9914), .B(n9913), .Z(n9952) );
  XNOR U10215 ( .A(n9953), .B(n9952), .Z(c[493]) );
  NANDN U10216 ( .A(n9916), .B(n9915), .Z(n9920) );
  NANDN U10217 ( .A(n9918), .B(n9917), .Z(n9919) );
  AND U10218 ( .A(n9920), .B(n9919), .Z(n9959) );
  NANDN U10219 ( .A(n9922), .B(n9921), .Z(n9926) );
  NANDN U10220 ( .A(n9924), .B(n9923), .Z(n9925) );
  AND U10221 ( .A(n9926), .B(n9925), .Z(n9957) );
  NAND U10222 ( .A(n26), .B(n9927), .Z(n9929) );
  XOR U10223 ( .A(b[7]), .B(a[240]), .Z(n9968) );
  NAND U10224 ( .A(n10531), .B(n9968), .Z(n9928) );
  AND U10225 ( .A(n9929), .B(n9928), .Z(n9987) );
  NAND U10226 ( .A(n23), .B(n9930), .Z(n9932) );
  XOR U10227 ( .A(b[3]), .B(a[244]), .Z(n9971) );
  NAND U10228 ( .A(n24), .B(n9971), .Z(n9931) );
  NAND U10229 ( .A(n9932), .B(n9931), .Z(n9986) );
  XNOR U10230 ( .A(n9987), .B(n9986), .Z(n9989) );
  NAND U10231 ( .A(b[0]), .B(a[246]), .Z(n9933) );
  XNOR U10232 ( .A(b[1]), .B(n9933), .Z(n9935) );
  NANDN U10233 ( .A(b[0]), .B(a[245]), .Z(n9934) );
  NAND U10234 ( .A(n9935), .B(n9934), .Z(n9983) );
  NAND U10235 ( .A(n25), .B(n9936), .Z(n9938) );
  XOR U10236 ( .A(b[5]), .B(a[242]), .Z(n9977) );
  NAND U10237 ( .A(n10456), .B(n9977), .Z(n9937) );
  AND U10238 ( .A(n9938), .B(n9937), .Z(n9981) );
  AND U10239 ( .A(b[7]), .B(a[238]), .Z(n9980) );
  XNOR U10240 ( .A(n9981), .B(n9980), .Z(n9982) );
  XNOR U10241 ( .A(n9983), .B(n9982), .Z(n9988) );
  XOR U10242 ( .A(n9989), .B(n9988), .Z(n9963) );
  NANDN U10243 ( .A(n9940), .B(n9939), .Z(n9944) );
  NANDN U10244 ( .A(n9942), .B(n9941), .Z(n9943) );
  AND U10245 ( .A(n9944), .B(n9943), .Z(n9962) );
  XNOR U10246 ( .A(n9963), .B(n9962), .Z(n9964) );
  NANDN U10247 ( .A(n9946), .B(n9945), .Z(n9950) );
  NAND U10248 ( .A(n9948), .B(n9947), .Z(n9949) );
  NAND U10249 ( .A(n9950), .B(n9949), .Z(n9965) );
  XNOR U10250 ( .A(n9964), .B(n9965), .Z(n9956) );
  XNOR U10251 ( .A(n9957), .B(n9956), .Z(n9958) );
  XNOR U10252 ( .A(n9959), .B(n9958), .Z(n9992) );
  XNOR U10253 ( .A(sreg[494]), .B(n9992), .Z(n9994) );
  NANDN U10254 ( .A(sreg[493]), .B(n9951), .Z(n9955) );
  NAND U10255 ( .A(n9953), .B(n9952), .Z(n9954) );
  NAND U10256 ( .A(n9955), .B(n9954), .Z(n9993) );
  XNOR U10257 ( .A(n9994), .B(n9993), .Z(c[494]) );
  NANDN U10258 ( .A(n9957), .B(n9956), .Z(n9961) );
  NANDN U10259 ( .A(n9959), .B(n9958), .Z(n9960) );
  AND U10260 ( .A(n9961), .B(n9960), .Z(n10000) );
  NANDN U10261 ( .A(n9963), .B(n9962), .Z(n9967) );
  NANDN U10262 ( .A(n9965), .B(n9964), .Z(n9966) );
  AND U10263 ( .A(n9967), .B(n9966), .Z(n9998) );
  NAND U10264 ( .A(n26), .B(n9968), .Z(n9970) );
  XOR U10265 ( .A(b[7]), .B(a[241]), .Z(n10009) );
  NAND U10266 ( .A(n10531), .B(n10009), .Z(n9969) );
  AND U10267 ( .A(n9970), .B(n9969), .Z(n10028) );
  NAND U10268 ( .A(n23), .B(n9971), .Z(n9973) );
  XOR U10269 ( .A(b[3]), .B(a[245]), .Z(n10012) );
  NAND U10270 ( .A(n24), .B(n10012), .Z(n9972) );
  NAND U10271 ( .A(n9973), .B(n9972), .Z(n10027) );
  XNOR U10272 ( .A(n10028), .B(n10027), .Z(n10030) );
  NAND U10273 ( .A(b[0]), .B(a[247]), .Z(n9974) );
  XNOR U10274 ( .A(b[1]), .B(n9974), .Z(n9976) );
  NANDN U10275 ( .A(b[0]), .B(a[246]), .Z(n9975) );
  NAND U10276 ( .A(n9976), .B(n9975), .Z(n10024) );
  NAND U10277 ( .A(n25), .B(n9977), .Z(n9979) );
  XOR U10278 ( .A(b[5]), .B(a[243]), .Z(n10018) );
  NAND U10279 ( .A(n10456), .B(n10018), .Z(n9978) );
  AND U10280 ( .A(n9979), .B(n9978), .Z(n10022) );
  AND U10281 ( .A(b[7]), .B(a[239]), .Z(n10021) );
  XNOR U10282 ( .A(n10022), .B(n10021), .Z(n10023) );
  XNOR U10283 ( .A(n10024), .B(n10023), .Z(n10029) );
  XOR U10284 ( .A(n10030), .B(n10029), .Z(n10004) );
  NANDN U10285 ( .A(n9981), .B(n9980), .Z(n9985) );
  NANDN U10286 ( .A(n9983), .B(n9982), .Z(n9984) );
  AND U10287 ( .A(n9985), .B(n9984), .Z(n10003) );
  XNOR U10288 ( .A(n10004), .B(n10003), .Z(n10005) );
  NANDN U10289 ( .A(n9987), .B(n9986), .Z(n9991) );
  NAND U10290 ( .A(n9989), .B(n9988), .Z(n9990) );
  NAND U10291 ( .A(n9991), .B(n9990), .Z(n10006) );
  XNOR U10292 ( .A(n10005), .B(n10006), .Z(n9997) );
  XNOR U10293 ( .A(n9998), .B(n9997), .Z(n9999) );
  XNOR U10294 ( .A(n10000), .B(n9999), .Z(n10033) );
  XNOR U10295 ( .A(sreg[495]), .B(n10033), .Z(n10035) );
  NANDN U10296 ( .A(sreg[494]), .B(n9992), .Z(n9996) );
  NAND U10297 ( .A(n9994), .B(n9993), .Z(n9995) );
  NAND U10298 ( .A(n9996), .B(n9995), .Z(n10034) );
  XNOR U10299 ( .A(n10035), .B(n10034), .Z(c[495]) );
  NANDN U10300 ( .A(n9998), .B(n9997), .Z(n10002) );
  NANDN U10301 ( .A(n10000), .B(n9999), .Z(n10001) );
  AND U10302 ( .A(n10002), .B(n10001), .Z(n10041) );
  NANDN U10303 ( .A(n10004), .B(n10003), .Z(n10008) );
  NANDN U10304 ( .A(n10006), .B(n10005), .Z(n10007) );
  AND U10305 ( .A(n10008), .B(n10007), .Z(n10039) );
  NAND U10306 ( .A(n26), .B(n10009), .Z(n10011) );
  XOR U10307 ( .A(b[7]), .B(a[242]), .Z(n10050) );
  NAND U10308 ( .A(n10531), .B(n10050), .Z(n10010) );
  AND U10309 ( .A(n10011), .B(n10010), .Z(n10069) );
  NAND U10310 ( .A(n23), .B(n10012), .Z(n10014) );
  XOR U10311 ( .A(b[3]), .B(a[246]), .Z(n10053) );
  NAND U10312 ( .A(n24), .B(n10053), .Z(n10013) );
  NAND U10313 ( .A(n10014), .B(n10013), .Z(n10068) );
  XNOR U10314 ( .A(n10069), .B(n10068), .Z(n10071) );
  NAND U10315 ( .A(b[0]), .B(a[248]), .Z(n10015) );
  XNOR U10316 ( .A(b[1]), .B(n10015), .Z(n10017) );
  NANDN U10317 ( .A(b[0]), .B(a[247]), .Z(n10016) );
  NAND U10318 ( .A(n10017), .B(n10016), .Z(n10065) );
  NAND U10319 ( .A(n25), .B(n10018), .Z(n10020) );
  XOR U10320 ( .A(b[5]), .B(a[244]), .Z(n10059) );
  NAND U10321 ( .A(n10456), .B(n10059), .Z(n10019) );
  AND U10322 ( .A(n10020), .B(n10019), .Z(n10063) );
  AND U10323 ( .A(b[7]), .B(a[240]), .Z(n10062) );
  XNOR U10324 ( .A(n10063), .B(n10062), .Z(n10064) );
  XNOR U10325 ( .A(n10065), .B(n10064), .Z(n10070) );
  XOR U10326 ( .A(n10071), .B(n10070), .Z(n10045) );
  NANDN U10327 ( .A(n10022), .B(n10021), .Z(n10026) );
  NANDN U10328 ( .A(n10024), .B(n10023), .Z(n10025) );
  AND U10329 ( .A(n10026), .B(n10025), .Z(n10044) );
  XNOR U10330 ( .A(n10045), .B(n10044), .Z(n10046) );
  NANDN U10331 ( .A(n10028), .B(n10027), .Z(n10032) );
  NAND U10332 ( .A(n10030), .B(n10029), .Z(n10031) );
  NAND U10333 ( .A(n10032), .B(n10031), .Z(n10047) );
  XNOR U10334 ( .A(n10046), .B(n10047), .Z(n10038) );
  XNOR U10335 ( .A(n10039), .B(n10038), .Z(n10040) );
  XNOR U10336 ( .A(n10041), .B(n10040), .Z(n10074) );
  XNOR U10337 ( .A(sreg[496]), .B(n10074), .Z(n10076) );
  NANDN U10338 ( .A(sreg[495]), .B(n10033), .Z(n10037) );
  NAND U10339 ( .A(n10035), .B(n10034), .Z(n10036) );
  NAND U10340 ( .A(n10037), .B(n10036), .Z(n10075) );
  XNOR U10341 ( .A(n10076), .B(n10075), .Z(c[496]) );
  NANDN U10342 ( .A(n10039), .B(n10038), .Z(n10043) );
  NANDN U10343 ( .A(n10041), .B(n10040), .Z(n10042) );
  AND U10344 ( .A(n10043), .B(n10042), .Z(n10082) );
  NANDN U10345 ( .A(n10045), .B(n10044), .Z(n10049) );
  NANDN U10346 ( .A(n10047), .B(n10046), .Z(n10048) );
  AND U10347 ( .A(n10049), .B(n10048), .Z(n10080) );
  NAND U10348 ( .A(n26), .B(n10050), .Z(n10052) );
  XOR U10349 ( .A(b[7]), .B(a[243]), .Z(n10091) );
  NAND U10350 ( .A(n10531), .B(n10091), .Z(n10051) );
  AND U10351 ( .A(n10052), .B(n10051), .Z(n10110) );
  NAND U10352 ( .A(n23), .B(n10053), .Z(n10055) );
  XOR U10353 ( .A(b[3]), .B(a[247]), .Z(n10094) );
  NAND U10354 ( .A(n24), .B(n10094), .Z(n10054) );
  NAND U10355 ( .A(n10055), .B(n10054), .Z(n10109) );
  XNOR U10356 ( .A(n10110), .B(n10109), .Z(n10112) );
  NAND U10357 ( .A(b[0]), .B(a[249]), .Z(n10056) );
  XNOR U10358 ( .A(b[1]), .B(n10056), .Z(n10058) );
  NANDN U10359 ( .A(b[0]), .B(a[248]), .Z(n10057) );
  NAND U10360 ( .A(n10058), .B(n10057), .Z(n10106) );
  NAND U10361 ( .A(n25), .B(n10059), .Z(n10061) );
  XOR U10362 ( .A(b[5]), .B(a[245]), .Z(n10100) );
  NAND U10363 ( .A(n10456), .B(n10100), .Z(n10060) );
  AND U10364 ( .A(n10061), .B(n10060), .Z(n10104) );
  AND U10365 ( .A(b[7]), .B(a[241]), .Z(n10103) );
  XNOR U10366 ( .A(n10104), .B(n10103), .Z(n10105) );
  XNOR U10367 ( .A(n10106), .B(n10105), .Z(n10111) );
  XOR U10368 ( .A(n10112), .B(n10111), .Z(n10086) );
  NANDN U10369 ( .A(n10063), .B(n10062), .Z(n10067) );
  NANDN U10370 ( .A(n10065), .B(n10064), .Z(n10066) );
  AND U10371 ( .A(n10067), .B(n10066), .Z(n10085) );
  XNOR U10372 ( .A(n10086), .B(n10085), .Z(n10087) );
  NANDN U10373 ( .A(n10069), .B(n10068), .Z(n10073) );
  NAND U10374 ( .A(n10071), .B(n10070), .Z(n10072) );
  NAND U10375 ( .A(n10073), .B(n10072), .Z(n10088) );
  XNOR U10376 ( .A(n10087), .B(n10088), .Z(n10079) );
  XNOR U10377 ( .A(n10080), .B(n10079), .Z(n10081) );
  XNOR U10378 ( .A(n10082), .B(n10081), .Z(n10115) );
  XNOR U10379 ( .A(sreg[497]), .B(n10115), .Z(n10117) );
  NANDN U10380 ( .A(sreg[496]), .B(n10074), .Z(n10078) );
  NAND U10381 ( .A(n10076), .B(n10075), .Z(n10077) );
  NAND U10382 ( .A(n10078), .B(n10077), .Z(n10116) );
  XNOR U10383 ( .A(n10117), .B(n10116), .Z(c[497]) );
  NANDN U10384 ( .A(n10080), .B(n10079), .Z(n10084) );
  NANDN U10385 ( .A(n10082), .B(n10081), .Z(n10083) );
  AND U10386 ( .A(n10084), .B(n10083), .Z(n10123) );
  NANDN U10387 ( .A(n10086), .B(n10085), .Z(n10090) );
  NANDN U10388 ( .A(n10088), .B(n10087), .Z(n10089) );
  AND U10389 ( .A(n10090), .B(n10089), .Z(n10121) );
  NAND U10390 ( .A(n26), .B(n10091), .Z(n10093) );
  XOR U10391 ( .A(b[7]), .B(a[244]), .Z(n10132) );
  NAND U10392 ( .A(n10531), .B(n10132), .Z(n10092) );
  AND U10393 ( .A(n10093), .B(n10092), .Z(n10151) );
  NAND U10394 ( .A(n23), .B(n10094), .Z(n10096) );
  XOR U10395 ( .A(b[3]), .B(a[248]), .Z(n10135) );
  NAND U10396 ( .A(n24), .B(n10135), .Z(n10095) );
  NAND U10397 ( .A(n10096), .B(n10095), .Z(n10150) );
  XNOR U10398 ( .A(n10151), .B(n10150), .Z(n10153) );
  NAND U10399 ( .A(b[0]), .B(a[250]), .Z(n10097) );
  XNOR U10400 ( .A(b[1]), .B(n10097), .Z(n10099) );
  NANDN U10401 ( .A(b[0]), .B(a[249]), .Z(n10098) );
  NAND U10402 ( .A(n10099), .B(n10098), .Z(n10147) );
  NAND U10403 ( .A(n25), .B(n10100), .Z(n10102) );
  XOR U10404 ( .A(b[5]), .B(a[246]), .Z(n10138) );
  NAND U10405 ( .A(n10456), .B(n10138), .Z(n10101) );
  AND U10406 ( .A(n10102), .B(n10101), .Z(n10145) );
  AND U10407 ( .A(b[7]), .B(a[242]), .Z(n10144) );
  XNOR U10408 ( .A(n10145), .B(n10144), .Z(n10146) );
  XNOR U10409 ( .A(n10147), .B(n10146), .Z(n10152) );
  XOR U10410 ( .A(n10153), .B(n10152), .Z(n10127) );
  NANDN U10411 ( .A(n10104), .B(n10103), .Z(n10108) );
  NANDN U10412 ( .A(n10106), .B(n10105), .Z(n10107) );
  AND U10413 ( .A(n10108), .B(n10107), .Z(n10126) );
  XNOR U10414 ( .A(n10127), .B(n10126), .Z(n10128) );
  NANDN U10415 ( .A(n10110), .B(n10109), .Z(n10114) );
  NAND U10416 ( .A(n10112), .B(n10111), .Z(n10113) );
  NAND U10417 ( .A(n10114), .B(n10113), .Z(n10129) );
  XNOR U10418 ( .A(n10128), .B(n10129), .Z(n10120) );
  XNOR U10419 ( .A(n10121), .B(n10120), .Z(n10122) );
  XNOR U10420 ( .A(n10123), .B(n10122), .Z(n10156) );
  XNOR U10421 ( .A(sreg[498]), .B(n10156), .Z(n10158) );
  NANDN U10422 ( .A(sreg[497]), .B(n10115), .Z(n10119) );
  NAND U10423 ( .A(n10117), .B(n10116), .Z(n10118) );
  NAND U10424 ( .A(n10119), .B(n10118), .Z(n10157) );
  XNOR U10425 ( .A(n10158), .B(n10157), .Z(c[498]) );
  NANDN U10426 ( .A(n10121), .B(n10120), .Z(n10125) );
  NANDN U10427 ( .A(n10123), .B(n10122), .Z(n10124) );
  AND U10428 ( .A(n10125), .B(n10124), .Z(n10164) );
  NANDN U10429 ( .A(n10127), .B(n10126), .Z(n10131) );
  NANDN U10430 ( .A(n10129), .B(n10128), .Z(n10130) );
  AND U10431 ( .A(n10131), .B(n10130), .Z(n10162) );
  NAND U10432 ( .A(n26), .B(n10132), .Z(n10134) );
  XOR U10433 ( .A(b[7]), .B(a[245]), .Z(n10173) );
  NAND U10434 ( .A(n10531), .B(n10173), .Z(n10133) );
  AND U10435 ( .A(n10134), .B(n10133), .Z(n10192) );
  NAND U10436 ( .A(n23), .B(n10135), .Z(n10137) );
  XOR U10437 ( .A(b[3]), .B(a[249]), .Z(n10176) );
  NAND U10438 ( .A(n24), .B(n10176), .Z(n10136) );
  NAND U10439 ( .A(n10137), .B(n10136), .Z(n10191) );
  XNOR U10440 ( .A(n10192), .B(n10191), .Z(n10194) );
  NAND U10441 ( .A(n25), .B(n10138), .Z(n10140) );
  XOR U10442 ( .A(b[5]), .B(a[247]), .Z(n10182) );
  NAND U10443 ( .A(n10456), .B(n10182), .Z(n10139) );
  AND U10444 ( .A(n10140), .B(n10139), .Z(n10186) );
  AND U10445 ( .A(b[7]), .B(a[243]), .Z(n10185) );
  XNOR U10446 ( .A(n10186), .B(n10185), .Z(n10187) );
  NAND U10447 ( .A(b[0]), .B(a[251]), .Z(n10141) );
  XNOR U10448 ( .A(b[1]), .B(n10141), .Z(n10143) );
  NANDN U10449 ( .A(b[0]), .B(a[250]), .Z(n10142) );
  NAND U10450 ( .A(n10143), .B(n10142), .Z(n10188) );
  XNOR U10451 ( .A(n10187), .B(n10188), .Z(n10193) );
  XOR U10452 ( .A(n10194), .B(n10193), .Z(n10168) );
  NANDN U10453 ( .A(n10145), .B(n10144), .Z(n10149) );
  NANDN U10454 ( .A(n10147), .B(n10146), .Z(n10148) );
  AND U10455 ( .A(n10149), .B(n10148), .Z(n10167) );
  XNOR U10456 ( .A(n10168), .B(n10167), .Z(n10169) );
  NANDN U10457 ( .A(n10151), .B(n10150), .Z(n10155) );
  NAND U10458 ( .A(n10153), .B(n10152), .Z(n10154) );
  NAND U10459 ( .A(n10155), .B(n10154), .Z(n10170) );
  XNOR U10460 ( .A(n10169), .B(n10170), .Z(n10161) );
  XNOR U10461 ( .A(n10162), .B(n10161), .Z(n10163) );
  XNOR U10462 ( .A(n10164), .B(n10163), .Z(n10197) );
  XNOR U10463 ( .A(sreg[499]), .B(n10197), .Z(n10199) );
  NANDN U10464 ( .A(sreg[498]), .B(n10156), .Z(n10160) );
  NAND U10465 ( .A(n10158), .B(n10157), .Z(n10159) );
  NAND U10466 ( .A(n10160), .B(n10159), .Z(n10198) );
  XNOR U10467 ( .A(n10199), .B(n10198), .Z(c[499]) );
  NANDN U10468 ( .A(n10162), .B(n10161), .Z(n10166) );
  NANDN U10469 ( .A(n10164), .B(n10163), .Z(n10165) );
  AND U10470 ( .A(n10166), .B(n10165), .Z(n10205) );
  NANDN U10471 ( .A(n10168), .B(n10167), .Z(n10172) );
  NANDN U10472 ( .A(n10170), .B(n10169), .Z(n10171) );
  AND U10473 ( .A(n10172), .B(n10171), .Z(n10203) );
  NAND U10474 ( .A(n26), .B(n10173), .Z(n10175) );
  XOR U10475 ( .A(b[7]), .B(a[246]), .Z(n10214) );
  NAND U10476 ( .A(n10531), .B(n10214), .Z(n10174) );
  AND U10477 ( .A(n10175), .B(n10174), .Z(n10233) );
  NAND U10478 ( .A(n23), .B(n10176), .Z(n10178) );
  XOR U10479 ( .A(b[3]), .B(a[250]), .Z(n10217) );
  NAND U10480 ( .A(n24), .B(n10217), .Z(n10177) );
  NAND U10481 ( .A(n10178), .B(n10177), .Z(n10232) );
  XNOR U10482 ( .A(n10233), .B(n10232), .Z(n10235) );
  NAND U10483 ( .A(b[0]), .B(a[252]), .Z(n10179) );
  XNOR U10484 ( .A(b[1]), .B(n10179), .Z(n10181) );
  NANDN U10485 ( .A(b[0]), .B(a[251]), .Z(n10180) );
  NAND U10486 ( .A(n10181), .B(n10180), .Z(n10229) );
  NAND U10487 ( .A(n25), .B(n10182), .Z(n10184) );
  XOR U10488 ( .A(b[5]), .B(a[248]), .Z(n10223) );
  NAND U10489 ( .A(n10456), .B(n10223), .Z(n10183) );
  AND U10490 ( .A(n10184), .B(n10183), .Z(n10227) );
  AND U10491 ( .A(b[7]), .B(a[244]), .Z(n10226) );
  XNOR U10492 ( .A(n10227), .B(n10226), .Z(n10228) );
  XNOR U10493 ( .A(n10229), .B(n10228), .Z(n10234) );
  XOR U10494 ( .A(n10235), .B(n10234), .Z(n10209) );
  NANDN U10495 ( .A(n10186), .B(n10185), .Z(n10190) );
  NANDN U10496 ( .A(n10188), .B(n10187), .Z(n10189) );
  AND U10497 ( .A(n10190), .B(n10189), .Z(n10208) );
  XNOR U10498 ( .A(n10209), .B(n10208), .Z(n10210) );
  NANDN U10499 ( .A(n10192), .B(n10191), .Z(n10196) );
  NAND U10500 ( .A(n10194), .B(n10193), .Z(n10195) );
  NAND U10501 ( .A(n10196), .B(n10195), .Z(n10211) );
  XNOR U10502 ( .A(n10210), .B(n10211), .Z(n10202) );
  XNOR U10503 ( .A(n10203), .B(n10202), .Z(n10204) );
  XNOR U10504 ( .A(n10205), .B(n10204), .Z(n10238) );
  XNOR U10505 ( .A(sreg[500]), .B(n10238), .Z(n10240) );
  NANDN U10506 ( .A(sreg[499]), .B(n10197), .Z(n10201) );
  NAND U10507 ( .A(n10199), .B(n10198), .Z(n10200) );
  NAND U10508 ( .A(n10201), .B(n10200), .Z(n10239) );
  XNOR U10509 ( .A(n10240), .B(n10239), .Z(c[500]) );
  NANDN U10510 ( .A(n10203), .B(n10202), .Z(n10207) );
  NANDN U10511 ( .A(n10205), .B(n10204), .Z(n10206) );
  AND U10512 ( .A(n10207), .B(n10206), .Z(n10246) );
  NANDN U10513 ( .A(n10209), .B(n10208), .Z(n10213) );
  NANDN U10514 ( .A(n10211), .B(n10210), .Z(n10212) );
  AND U10515 ( .A(n10213), .B(n10212), .Z(n10244) );
  NAND U10516 ( .A(n26), .B(n10214), .Z(n10216) );
  XOR U10517 ( .A(b[7]), .B(a[247]), .Z(n10255) );
  NAND U10518 ( .A(n10531), .B(n10255), .Z(n10215) );
  AND U10519 ( .A(n10216), .B(n10215), .Z(n10274) );
  NAND U10520 ( .A(n23), .B(n10217), .Z(n10219) );
  XOR U10521 ( .A(b[3]), .B(a[251]), .Z(n10258) );
  NAND U10522 ( .A(n24), .B(n10258), .Z(n10218) );
  NAND U10523 ( .A(n10219), .B(n10218), .Z(n10273) );
  XNOR U10524 ( .A(n10274), .B(n10273), .Z(n10276) );
  NAND U10525 ( .A(b[0]), .B(a[253]), .Z(n10220) );
  XNOR U10526 ( .A(b[1]), .B(n10220), .Z(n10222) );
  NANDN U10527 ( .A(b[0]), .B(a[252]), .Z(n10221) );
  NAND U10528 ( .A(n10222), .B(n10221), .Z(n10270) );
  NAND U10529 ( .A(n25), .B(n10223), .Z(n10225) );
  XOR U10530 ( .A(b[5]), .B(a[249]), .Z(n10264) );
  NAND U10531 ( .A(n10456), .B(n10264), .Z(n10224) );
  AND U10532 ( .A(n10225), .B(n10224), .Z(n10268) );
  AND U10533 ( .A(b[7]), .B(a[245]), .Z(n10267) );
  XNOR U10534 ( .A(n10268), .B(n10267), .Z(n10269) );
  XNOR U10535 ( .A(n10270), .B(n10269), .Z(n10275) );
  XOR U10536 ( .A(n10276), .B(n10275), .Z(n10250) );
  NANDN U10537 ( .A(n10227), .B(n10226), .Z(n10231) );
  NANDN U10538 ( .A(n10229), .B(n10228), .Z(n10230) );
  AND U10539 ( .A(n10231), .B(n10230), .Z(n10249) );
  XNOR U10540 ( .A(n10250), .B(n10249), .Z(n10251) );
  NANDN U10541 ( .A(n10233), .B(n10232), .Z(n10237) );
  NAND U10542 ( .A(n10235), .B(n10234), .Z(n10236) );
  NAND U10543 ( .A(n10237), .B(n10236), .Z(n10252) );
  XNOR U10544 ( .A(n10251), .B(n10252), .Z(n10243) );
  XNOR U10545 ( .A(n10244), .B(n10243), .Z(n10245) );
  XNOR U10546 ( .A(n10246), .B(n10245), .Z(n10279) );
  XNOR U10547 ( .A(sreg[501]), .B(n10279), .Z(n10281) );
  NANDN U10548 ( .A(sreg[500]), .B(n10238), .Z(n10242) );
  NAND U10549 ( .A(n10240), .B(n10239), .Z(n10241) );
  NAND U10550 ( .A(n10242), .B(n10241), .Z(n10280) );
  XNOR U10551 ( .A(n10281), .B(n10280), .Z(c[501]) );
  NANDN U10552 ( .A(n10244), .B(n10243), .Z(n10248) );
  NANDN U10553 ( .A(n10246), .B(n10245), .Z(n10247) );
  AND U10554 ( .A(n10248), .B(n10247), .Z(n10287) );
  NANDN U10555 ( .A(n10250), .B(n10249), .Z(n10254) );
  NANDN U10556 ( .A(n10252), .B(n10251), .Z(n10253) );
  AND U10557 ( .A(n10254), .B(n10253), .Z(n10285) );
  NANDN U10558 ( .A(n21), .B(n10255), .Z(n10257) );
  XNOR U10559 ( .A(b[7]), .B(a[248]), .Z(n10308) );
  OR U10560 ( .A(n10308), .B(n10507), .Z(n10256) );
  NAND U10561 ( .A(n10257), .B(n10256), .Z(n10297) );
  NAND U10562 ( .A(n23), .B(n10258), .Z(n10260) );
  XNOR U10563 ( .A(a[252]), .B(b[3]), .Z(n10311) );
  OR U10564 ( .A(n10311), .B(n22), .Z(n10259) );
  NAND U10565 ( .A(n10260), .B(n10259), .Z(n10296) );
  XOR U10566 ( .A(n10297), .B(n10296), .Z(n10298) );
  NAND U10567 ( .A(b[0]), .B(a[254]), .Z(n10261) );
  XNOR U10568 ( .A(b[1]), .B(n10261), .Z(n10263) );
  NANDN U10569 ( .A(b[0]), .B(a[253]), .Z(n10262) );
  NAND U10570 ( .A(n10263), .B(n10262), .Z(n10305) );
  NANDN U10571 ( .A(n20), .B(n10264), .Z(n10266) );
  XNOR U10572 ( .A(b[5]), .B(a[250]), .Z(n10317) );
  OR U10573 ( .A(n10317), .B(n10424), .Z(n10265) );
  NAND U10574 ( .A(n10266), .B(n10265), .Z(n10302) );
  AND U10575 ( .A(b[7]), .B(a[246]), .Z(n10303) );
  XOR U10576 ( .A(n10302), .B(n10303), .Z(n10304) );
  NANDN U10577 ( .A(n10268), .B(n10267), .Z(n10272) );
  NANDN U10578 ( .A(n10270), .B(n10269), .Z(n10271) );
  AND U10579 ( .A(n10272), .B(n10271), .Z(n10290) );
  NANDN U10580 ( .A(n10274), .B(n10273), .Z(n10278) );
  NAND U10581 ( .A(n10276), .B(n10275), .Z(n10277) );
  AND U10582 ( .A(n10278), .B(n10277), .Z(n10292) );
  XOR U10583 ( .A(n10293), .B(n10292), .Z(n10284) );
  XNOR U10584 ( .A(n10285), .B(n10284), .Z(n10286) );
  XNOR U10585 ( .A(n10287), .B(n10286), .Z(n10320) );
  XNOR U10586 ( .A(sreg[502]), .B(n10320), .Z(n10322) );
  NANDN U10587 ( .A(sreg[501]), .B(n10279), .Z(n10283) );
  NAND U10588 ( .A(n10281), .B(n10280), .Z(n10282) );
  NAND U10589 ( .A(n10283), .B(n10282), .Z(n10321) );
  XNOR U10590 ( .A(n10322), .B(n10321), .Z(c[502]) );
  NANDN U10591 ( .A(n10285), .B(n10284), .Z(n10289) );
  NANDN U10592 ( .A(n10287), .B(n10286), .Z(n10288) );
  NAND U10593 ( .A(n10289), .B(n10288), .Z(n10332) );
  NAND U10594 ( .A(n10291), .B(n10290), .Z(n10295) );
  NAND U10595 ( .A(n10293), .B(n10292), .Z(n10294) );
  NAND U10596 ( .A(n10295), .B(n10294), .Z(n10331) );
  NAND U10597 ( .A(n10297), .B(n10296), .Z(n10301) );
  NAND U10598 ( .A(n10299), .B(n10298), .Z(n10300) );
  NAND U10599 ( .A(n10301), .B(n10300), .Z(n10359) );
  NAND U10600 ( .A(n10303), .B(n10302), .Z(n10307) );
  NANDN U10601 ( .A(n10305), .B(n10304), .Z(n10306) );
  NAND U10602 ( .A(n10307), .B(n10306), .Z(n10357) );
  OR U10603 ( .A(n10308), .B(n21), .Z(n10310) );
  XNOR U10604 ( .A(b[7]), .B(a[249]), .Z(n10348) );
  OR U10605 ( .A(n10348), .B(n10507), .Z(n10309) );
  NAND U10606 ( .A(n10310), .B(n10309), .Z(n10338) );
  OR U10607 ( .A(n10311), .B(n19), .Z(n10313) );
  XNOR U10608 ( .A(a[253]), .B(b[3]), .Z(n10351) );
  OR U10609 ( .A(n10351), .B(n22), .Z(n10312) );
  NAND U10610 ( .A(n10313), .B(n10312), .Z(n10336) );
  NAND U10611 ( .A(b[0]), .B(a[255]), .Z(n10314) );
  XNOR U10612 ( .A(b[1]), .B(n10314), .Z(n10316) );
  NANDN U10613 ( .A(b[0]), .B(a[254]), .Z(n10315) );
  NAND U10614 ( .A(n10316), .B(n10315), .Z(n10345) );
  OR U10615 ( .A(n10317), .B(n20), .Z(n10319) );
  XNOR U10616 ( .A(b[5]), .B(a[251]), .Z(n10354) );
  OR U10617 ( .A(n10354), .B(n10424), .Z(n10318) );
  NAND U10618 ( .A(n10319), .B(n10318), .Z(n10342) );
  AND U10619 ( .A(b[7]), .B(a[247]), .Z(n10343) );
  XOR U10620 ( .A(n10342), .B(n10343), .Z(n10344) );
  XOR U10621 ( .A(n10338), .B(n10339), .Z(n10358) );
  XOR U10622 ( .A(n10357), .B(n10358), .Z(n10360) );
  XOR U10623 ( .A(n10359), .B(n10360), .Z(n10330) );
  XOR U10624 ( .A(n10331), .B(n10330), .Z(n10333) );
  XOR U10625 ( .A(n10332), .B(n10333), .Z(n10325) );
  XNOR U10626 ( .A(sreg[503]), .B(n10325), .Z(n10327) );
  NANDN U10627 ( .A(sreg[502]), .B(n10320), .Z(n10324) );
  NAND U10628 ( .A(n10322), .B(n10321), .Z(n10323) );
  NAND U10629 ( .A(n10324), .B(n10323), .Z(n10326) );
  XNOR U10630 ( .A(n10327), .B(n10326), .Z(c[503]) );
  NANDN U10631 ( .A(sreg[503]), .B(n10325), .Z(n10329) );
  NAND U10632 ( .A(n10327), .B(n10326), .Z(n10328) );
  AND U10633 ( .A(n10329), .B(n10328), .Z(n10364) );
  NAND U10634 ( .A(n10331), .B(n10330), .Z(n10335) );
  NAND U10635 ( .A(n10333), .B(n10332), .Z(n10334) );
  NAND U10636 ( .A(n10335), .B(n10334), .Z(n10367) );
  NAND U10637 ( .A(n10337), .B(n10336), .Z(n10341) );
  NANDN U10638 ( .A(n10339), .B(n10338), .Z(n10340) );
  NAND U10639 ( .A(n10341), .B(n10340), .Z(n10394) );
  NAND U10640 ( .A(n10343), .B(n10342), .Z(n10347) );
  NANDN U10641 ( .A(n10345), .B(n10344), .Z(n10346) );
  NAND U10642 ( .A(n10347), .B(n10346), .Z(n10392) );
  OR U10643 ( .A(n10348), .B(n21), .Z(n10350) );
  XNOR U10644 ( .A(b[7]), .B(a[250]), .Z(n10377) );
  OR U10645 ( .A(n10377), .B(n10507), .Z(n10349) );
  NAND U10646 ( .A(n10350), .B(n10349), .Z(n10373) );
  OR U10647 ( .A(n10351), .B(n19), .Z(n10353) );
  XOR U10648 ( .A(b[3]), .B(a[254]), .Z(n10383) );
  NANDN U10649 ( .A(n22), .B(n10383), .Z(n10352) );
  NAND U10650 ( .A(n10353), .B(n10352), .Z(n10371) );
  OR U10651 ( .A(n10354), .B(n20), .Z(n10356) );
  XOR U10652 ( .A(b[5]), .B(a[252]), .Z(n10380) );
  NANDN U10653 ( .A(n10424), .B(n10380), .Z(n10355) );
  NAND U10654 ( .A(n10356), .B(n10355), .Z(n10388) );
  AND U10655 ( .A(b[7]), .B(a[248]), .Z(n10387) );
  XOR U10656 ( .A(n10386), .B(n10387), .Z(n10389) );
  XOR U10657 ( .A(n10388), .B(n10389), .Z(n10372) );
  XOR U10658 ( .A(n10371), .B(n10372), .Z(n10374) );
  XOR U10659 ( .A(n10373), .B(n10374), .Z(n10393) );
  XOR U10660 ( .A(n10392), .B(n10393), .Z(n10395) );
  XNOR U10661 ( .A(n10394), .B(n10395), .Z(n10366) );
  NANDN U10662 ( .A(n10358), .B(n10357), .Z(n10362) );
  NANDN U10663 ( .A(n10360), .B(n10359), .Z(n10361) );
  AND U10664 ( .A(n10362), .B(n10361), .Z(n10365) );
  XOR U10665 ( .A(n10367), .B(n10368), .Z(n10363) );
  XOR U10666 ( .A(n10364), .B(n10363), .Z(c[504]) );
  AND U10667 ( .A(n10364), .B(n10363), .Z(n10399) );
  NAND U10668 ( .A(n10366), .B(n10365), .Z(n10370) );
  NANDN U10669 ( .A(n10368), .B(n10367), .Z(n10369) );
  NAND U10670 ( .A(n10370), .B(n10369), .Z(n10402) );
  NAND U10671 ( .A(n10372), .B(n10371), .Z(n10376) );
  NAND U10672 ( .A(n10374), .B(n10373), .Z(n10375) );
  NAND U10673 ( .A(n10376), .B(n10375), .Z(n10408) );
  OR U10674 ( .A(n10377), .B(n21), .Z(n10379) );
  XNOR U10675 ( .A(b[7]), .B(a[251]), .Z(n10420) );
  OR U10676 ( .A(n10420), .B(n10507), .Z(n10378) );
  NAND U10677 ( .A(n10379), .B(n10378), .Z(n10428) );
  AND U10678 ( .A(b[7]), .B(a[249]), .Z(n10482) );
  NAND U10679 ( .A(n25), .B(n10380), .Z(n10382) );
  XNOR U10680 ( .A(b[5]), .B(a[253]), .Z(n10423) );
  OR U10681 ( .A(n10423), .B(n10424), .Z(n10381) );
  NAND U10682 ( .A(n10382), .B(n10381), .Z(n10427) );
  XNOR U10683 ( .A(n10482), .B(n10427), .Z(n10429) );
  XNOR U10684 ( .A(n10428), .B(n10429), .Z(n10414) );
  NAND U10685 ( .A(n23), .B(n10383), .Z(n10385) );
  XNOR U10686 ( .A(b[3]), .B(a[255]), .Z(n10417) );
  OR U10687 ( .A(n10417), .B(n22), .Z(n10384) );
  AND U10688 ( .A(n10385), .B(n10384), .Z(n10412) );
  XOR U10689 ( .A(b[1]), .B(n10412), .Z(n10413) );
  NAND U10690 ( .A(n10387), .B(n10386), .Z(n10391) );
  NAND U10691 ( .A(n10389), .B(n10388), .Z(n10390) );
  NAND U10692 ( .A(n10391), .B(n10390), .Z(n10406) );
  XNOR U10693 ( .A(n10408), .B(n10409), .Z(n10401) );
  NAND U10694 ( .A(n10393), .B(n10392), .Z(n10397) );
  NAND U10695 ( .A(n10395), .B(n10394), .Z(n10396) );
  AND U10696 ( .A(n10397), .B(n10396), .Z(n10400) );
  XOR U10697 ( .A(n10402), .B(n10403), .Z(n10398) );
  XOR U10698 ( .A(n10399), .B(n10398), .Z(c[505]) );
  AND U10699 ( .A(n10399), .B(n10398), .Z(n10433) );
  NAND U10700 ( .A(n10401), .B(n10400), .Z(n10405) );
  NANDN U10701 ( .A(n10403), .B(n10402), .Z(n10404) );
  NAND U10702 ( .A(n10405), .B(n10404), .Z(n10436) );
  NAND U10703 ( .A(n10407), .B(n10406), .Z(n10411) );
  NAND U10704 ( .A(n10409), .B(n10408), .Z(n10410) );
  AND U10705 ( .A(n10411), .B(n10410), .Z(n10435) );
  NAND U10706 ( .A(b[1]), .B(n10412), .Z(n10416) );
  NAND U10707 ( .A(n10414), .B(n10413), .Z(n10415) );
  NAND U10708 ( .A(n10416), .B(n10415), .Z(n10442) );
  NAND U10709 ( .A(n24), .B(b[3]), .Z(n10419) );
  OR U10710 ( .A(n10417), .B(n19), .Z(n10418) );
  AND U10711 ( .A(n10419), .B(n10418), .Z(n10459) );
  NAND U10712 ( .A(b[7]), .B(a[250]), .Z(n10460) );
  XOR U10713 ( .A(n10459), .B(n10460), .Z(n10461) );
  XNOR U10714 ( .A(n10482), .B(n10461), .Z(n10448) );
  OR U10715 ( .A(n10420), .B(n21), .Z(n10422) );
  XNOR U10716 ( .A(b[7]), .B(a[252]), .Z(n10452) );
  OR U10717 ( .A(n10452), .B(n10507), .Z(n10421) );
  NAND U10718 ( .A(n10422), .B(n10421), .Z(n10447) );
  OR U10719 ( .A(n10423), .B(n20), .Z(n10426) );
  XOR U10720 ( .A(b[5]), .B(a[254]), .Z(n10455) );
  NANDN U10721 ( .A(n10424), .B(n10455), .Z(n10425) );
  NAND U10722 ( .A(n10426), .B(n10425), .Z(n10446) );
  XOR U10723 ( .A(n10447), .B(n10446), .Z(n10449) );
  IV U10724 ( .A(n10482), .Z(n10462) );
  NAND U10725 ( .A(n10462), .B(n10427), .Z(n10431) );
  NAND U10726 ( .A(n10429), .B(n10428), .Z(n10430) );
  AND U10727 ( .A(n10431), .B(n10430), .Z(n10440) );
  XOR U10728 ( .A(n10442), .B(n10443), .Z(n10434) );
  XOR U10729 ( .A(n10435), .B(n10434), .Z(n10437) );
  XNOR U10730 ( .A(n10436), .B(n10437), .Z(n10432) );
  XOR U10731 ( .A(n10433), .B(n10432), .Z(c[506]) );
  AND U10732 ( .A(n10433), .B(n10432), .Z(n10466) );
  NAND U10733 ( .A(n10435), .B(n10434), .Z(n10439) );
  NAND U10734 ( .A(n10437), .B(n10436), .Z(n10438) );
  NAND U10735 ( .A(n10439), .B(n10438), .Z(n10469) );
  NAND U10736 ( .A(n10441), .B(n10440), .Z(n10445) );
  NAND U10737 ( .A(n10443), .B(n10442), .Z(n10444) );
  NAND U10738 ( .A(n10445), .B(n10444), .Z(n10467) );
  NAND U10739 ( .A(n10447), .B(n10446), .Z(n10451) );
  NAND U10740 ( .A(n10449), .B(n10448), .Z(n10450) );
  AND U10741 ( .A(n10451), .B(n10450), .Z(n10495) );
  OR U10742 ( .A(n10452), .B(n21), .Z(n10454) );
  XNOR U10743 ( .A(b[7]), .B(a[253]), .Z(n10485) );
  OR U10744 ( .A(n10485), .B(n10507), .Z(n10453) );
  NAND U10745 ( .A(n10454), .B(n10453), .Z(n10474) );
  NAND U10746 ( .A(n25), .B(n10455), .Z(n10458) );
  XOR U10747 ( .A(b[5]), .B(a[255]), .Z(n10488) );
  NAND U10748 ( .A(n10456), .B(n10488), .Z(n10457) );
  NAND U10749 ( .A(n10458), .B(n10457), .Z(n10473) );
  XOR U10750 ( .A(n10474), .B(n10473), .Z(n10475) );
  AND U10751 ( .A(b[7]), .B(a[251]), .Z(n10480) );
  XOR U10752 ( .A(n10479), .B(n10480), .Z(n10481) );
  XOR U10753 ( .A(n10482), .B(n10481), .Z(n10476) );
  OR U10754 ( .A(n10460), .B(n10459), .Z(n10464) );
  NAND U10755 ( .A(n10462), .B(n10461), .Z(n10463) );
  AND U10756 ( .A(n10464), .B(n10463), .Z(n10492) );
  XOR U10757 ( .A(n10495), .B(n10494), .Z(n10468) );
  XNOR U10758 ( .A(n10467), .B(n10468), .Z(n10470) );
  XOR U10759 ( .A(n10469), .B(n10470), .Z(n10465) );
  XOR U10760 ( .A(n10466), .B(n10465), .Z(c[507]) );
  AND U10761 ( .A(n10466), .B(n10465), .Z(n10499) );
  NAND U10762 ( .A(n10468), .B(n10467), .Z(n10472) );
  NANDN U10763 ( .A(n10470), .B(n10469), .Z(n10471) );
  NAND U10764 ( .A(n10472), .B(n10471), .Z(n10502) );
  NAND U10765 ( .A(n10474), .B(n10473), .Z(n10478) );
  NAND U10766 ( .A(n10476), .B(n10475), .Z(n10477) );
  NAND U10767 ( .A(n10478), .B(n10477), .Z(n10518) );
  NAND U10768 ( .A(n10480), .B(n10479), .Z(n10484) );
  NAND U10769 ( .A(n10482), .B(n10481), .Z(n10483) );
  NAND U10770 ( .A(n10484), .B(n10483), .Z(n10516) );
  OR U10771 ( .A(n10485), .B(n21), .Z(n10487) );
  XNOR U10772 ( .A(b[7]), .B(a[254]), .Z(n10506) );
  OR U10773 ( .A(n10506), .B(n10507), .Z(n10486) );
  NAND U10774 ( .A(n10487), .B(n10486), .Z(n10512) );
  AND U10775 ( .A(b[7]), .B(a[252]), .Z(n10527) );
  AND U10776 ( .A(n10488), .B(n25), .Z(n10491) );
  XOR U10777 ( .A(b[4]), .B(b[3]), .Z(n10489) );
  NAND U10778 ( .A(b[5]), .B(n10489), .Z(n10490) );
  NANDN U10779 ( .A(n10491), .B(n10490), .Z(n10510) );
  XNOR U10780 ( .A(n10527), .B(n10510), .Z(n10513) );
  XOR U10781 ( .A(n10512), .B(n10513), .Z(n10517) );
  XOR U10782 ( .A(n10516), .B(n10517), .Z(n10519) );
  XNOR U10783 ( .A(n10518), .B(n10519), .Z(n10501) );
  NAND U10784 ( .A(n10493), .B(n10492), .Z(n10497) );
  NAND U10785 ( .A(n10495), .B(n10494), .Z(n10496) );
  NAND U10786 ( .A(n10497), .B(n10496), .Z(n10500) );
  XOR U10787 ( .A(n10502), .B(n10503), .Z(n10498) );
  XOR U10788 ( .A(n10499), .B(n10498), .Z(c[508]) );
  AND U10789 ( .A(n10499), .B(n10498), .Z(n10523) );
  NAND U10790 ( .A(n10501), .B(n10500), .Z(n10505) );
  NANDN U10791 ( .A(n10503), .B(n10502), .Z(n10504) );
  NAND U10792 ( .A(n10505), .B(n10504), .Z(n10536) );
  IV U10793 ( .A(n10527), .Z(n10511) );
  AND U10794 ( .A(b[7]), .B(a[253]), .Z(n10525) );
  XOR U10795 ( .A(n10525), .B(n10524), .Z(n10526) );
  XNOR U10796 ( .A(n10511), .B(n10526), .Z(n10541) );
  OR U10797 ( .A(n10506), .B(n21), .Z(n10509) );
  XOR U10798 ( .A(b[7]), .B(a[255]), .Z(n10530) );
  NANDN U10799 ( .A(n10507), .B(n10530), .Z(n10508) );
  NAND U10800 ( .A(n10509), .B(n10508), .Z(n10540) );
  XOR U10801 ( .A(n10541), .B(n10540), .Z(n10543) );
  NAND U10802 ( .A(n10511), .B(n10510), .Z(n10515) );
  NAND U10803 ( .A(n10513), .B(n10512), .Z(n10514) );
  NAND U10804 ( .A(n10515), .B(n10514), .Z(n10542) );
  XNOR U10805 ( .A(n10543), .B(n10542), .Z(n10535) );
  NAND U10806 ( .A(n10517), .B(n10516), .Z(n10521) );
  NAND U10807 ( .A(n10519), .B(n10518), .Z(n10520) );
  AND U10808 ( .A(n10521), .B(n10520), .Z(n10534) );
  XOR U10809 ( .A(n10536), .B(n10537), .Z(n10522) );
  XOR U10810 ( .A(n10523), .B(n10522), .Z(c[509]) );
  AND U10811 ( .A(n10523), .B(n10522), .Z(n10548) );
  AND U10812 ( .A(n10525), .B(n10524), .Z(n10529) );
  NAND U10813 ( .A(n10527), .B(n10526), .Z(n10528) );
  NANDN U10814 ( .A(n10529), .B(n10528), .Z(n10563) );
  NAND U10815 ( .A(b[7]), .B(a[254]), .Z(n10562) );
  NAND U10816 ( .A(n26), .B(n10530), .Z(n10533) );
  NAND U10817 ( .A(n10531), .B(b[7]), .Z(n10532) );
  NAND U10818 ( .A(n10533), .B(n10532), .Z(n10561) );
  XOR U10819 ( .A(n10562), .B(n10561), .Z(n10564) );
  XOR U10820 ( .A(n10563), .B(n10564), .Z(n10547) );
  XNOR U10821 ( .A(n10548), .B(n10547), .Z(n10555) );
  NAND U10822 ( .A(n10535), .B(n10534), .Z(n10539) );
  NANDN U10823 ( .A(n10537), .B(n10536), .Z(n10538) );
  NAND U10824 ( .A(n10539), .B(n10538), .Z(n10552) );
  IV U10825 ( .A(n10552), .Z(n10549) );
  NAND U10826 ( .A(n10541), .B(n10540), .Z(n10545) );
  NAND U10827 ( .A(n10543), .B(n10542), .Z(n10544) );
  AND U10828 ( .A(n10545), .B(n10544), .Z(n10553) );
  XNOR U10829 ( .A(n10549), .B(n10553), .Z(n10546) );
  XNOR U10830 ( .A(n10555), .B(n10546), .Z(c[510]) );
  NAND U10831 ( .A(n10548), .B(n10547), .Z(n10551) );
  NANDN U10832 ( .A(n10553), .B(n10549), .Z(n10550) );
  AND U10833 ( .A(n10551), .B(n10550), .Z(n10557) );
  AND U10834 ( .A(n10553), .B(n10552), .Z(n10554) );
  OR U10835 ( .A(n10555), .B(n10554), .Z(n10556) );
  AND U10836 ( .A(n10557), .B(n10556), .Z(n10570) );
  XNOR U10837 ( .A(n10558), .B(a[254]), .Z(n10559) );
  XNOR U10838 ( .A(a[255]), .B(n10559), .Z(n10560) );
  ANDN U10839 ( .B(b[7]), .A(n10560), .Z(n10568) );
  AND U10840 ( .A(n10562), .B(n10561), .Z(n10566) );
  AND U10841 ( .A(n10564), .B(n10563), .Z(n10565) );
  OR U10842 ( .A(n10566), .B(n10565), .Z(n10567) );
  XNOR U10843 ( .A(n10568), .B(n10567), .Z(n10569) );
  XNOR U10844 ( .A(n10570), .B(n10569), .Z(c[511]) );
endmodule

