
module mult_N128_CC32 ( clk, rst, a, b, c );
  input [127:0] a;
  input [3:0] b;
  output [127:0] c;
  input clk, rst;
  wire   \mult_44/PROD1[3] , \mult_44/SUMB[1][1] , \mult_44/SUMB[1][2] ,
         \mult_44/SUMB[2][1] , \mult_44/SUMB[2][2] , \mult_44/SUMB[3][1] ,
         \mult_44/SUMB[3][2] , \mult_44/SUMB[4][1] , \mult_44/SUMB[4][2] ,
         \mult_44/SUMB[5][1] , \mult_44/SUMB[5][2] , \mult_44/SUMB[6][1] ,
         \mult_44/SUMB[6][2] , \mult_44/SUMB[7][1] , \mult_44/SUMB[7][2] ,
         \mult_44/SUMB[8][1] , \mult_44/SUMB[8][2] , \mult_44/SUMB[9][1] ,
         \mult_44/SUMB[9][2] , \mult_44/SUMB[10][1] , \mult_44/SUMB[10][2] ,
         \mult_44/SUMB[11][1] , \mult_44/SUMB[11][2] , \mult_44/SUMB[12][1] ,
         \mult_44/SUMB[12][2] , \mult_44/SUMB[13][1] , \mult_44/SUMB[13][2] ,
         \mult_44/SUMB[14][1] , \mult_44/SUMB[14][2] , \mult_44/SUMB[15][1] ,
         \mult_44/SUMB[15][2] , \mult_44/SUMB[16][1] , \mult_44/SUMB[16][2] ,
         \mult_44/SUMB[17][1] , \mult_44/SUMB[17][2] , \mult_44/SUMB[18][1] ,
         \mult_44/SUMB[18][2] , \mult_44/SUMB[19][1] , \mult_44/SUMB[19][2] ,
         \mult_44/SUMB[20][1] , \mult_44/SUMB[20][2] , \mult_44/SUMB[21][1] ,
         \mult_44/SUMB[21][2] , \mult_44/SUMB[22][1] , \mult_44/SUMB[22][2] ,
         \mult_44/SUMB[23][1] , \mult_44/SUMB[23][2] , \mult_44/SUMB[24][1] ,
         \mult_44/SUMB[24][2] , \mult_44/SUMB[25][1] , \mult_44/SUMB[25][2] ,
         \mult_44/SUMB[26][1] , \mult_44/SUMB[26][2] , \mult_44/SUMB[27][1] ,
         \mult_44/SUMB[27][2] , \mult_44/SUMB[28][1] , \mult_44/SUMB[28][2] ,
         \mult_44/SUMB[29][1] , \mult_44/SUMB[29][2] , \mult_44/SUMB[30][1] ,
         \mult_44/SUMB[30][2] , \mult_44/SUMB[31][1] , \mult_44/SUMB[31][2] ,
         \mult_44/SUMB[32][1] , \mult_44/SUMB[32][2] , \mult_44/SUMB[33][1] ,
         \mult_44/SUMB[33][2] , \mult_44/SUMB[34][1] , \mult_44/SUMB[34][2] ,
         \mult_44/SUMB[35][1] , \mult_44/SUMB[35][2] , \mult_44/SUMB[36][1] ,
         \mult_44/SUMB[36][2] , \mult_44/SUMB[37][1] , \mult_44/SUMB[37][2] ,
         \mult_44/SUMB[38][1] , \mult_44/SUMB[38][2] , \mult_44/SUMB[39][1] ,
         \mult_44/SUMB[39][2] , \mult_44/SUMB[40][1] , \mult_44/SUMB[40][2] ,
         \mult_44/SUMB[41][1] , \mult_44/SUMB[41][2] , \mult_44/SUMB[42][1] ,
         \mult_44/SUMB[42][2] , \mult_44/SUMB[43][1] , \mult_44/SUMB[43][2] ,
         \mult_44/SUMB[44][1] , \mult_44/SUMB[44][2] , \mult_44/SUMB[45][1] ,
         \mult_44/SUMB[45][2] , \mult_44/SUMB[46][1] , \mult_44/SUMB[46][2] ,
         \mult_44/SUMB[47][1] , \mult_44/SUMB[47][2] , \mult_44/SUMB[48][1] ,
         \mult_44/SUMB[48][2] , \mult_44/SUMB[49][1] , \mult_44/SUMB[49][2] ,
         \mult_44/SUMB[50][1] , \mult_44/SUMB[50][2] , \mult_44/SUMB[51][1] ,
         \mult_44/SUMB[51][2] , \mult_44/SUMB[52][1] , \mult_44/SUMB[52][2] ,
         \mult_44/SUMB[53][1] , \mult_44/SUMB[53][2] , \mult_44/SUMB[54][1] ,
         \mult_44/SUMB[54][2] , \mult_44/SUMB[55][1] , \mult_44/SUMB[55][2] ,
         \mult_44/SUMB[56][1] , \mult_44/SUMB[56][2] , \mult_44/SUMB[57][1] ,
         \mult_44/SUMB[57][2] , \mult_44/SUMB[58][1] , \mult_44/SUMB[58][2] ,
         \mult_44/SUMB[59][1] , \mult_44/SUMB[59][2] , \mult_44/SUMB[60][1] ,
         \mult_44/SUMB[60][2] , \mult_44/SUMB[61][1] , \mult_44/SUMB[61][2] ,
         \mult_44/SUMB[62][1] , \mult_44/SUMB[62][2] , \mult_44/SUMB[63][1] ,
         \mult_44/SUMB[63][2] , \mult_44/SUMB[64][1] , \mult_44/SUMB[64][2] ,
         \mult_44/SUMB[65][1] , \mult_44/SUMB[65][2] , \mult_44/SUMB[66][1] ,
         \mult_44/SUMB[66][2] , \mult_44/SUMB[67][1] , \mult_44/SUMB[67][2] ,
         \mult_44/SUMB[68][1] , \mult_44/SUMB[68][2] , \mult_44/SUMB[69][1] ,
         \mult_44/SUMB[69][2] , \mult_44/SUMB[70][1] , \mult_44/SUMB[70][2] ,
         \mult_44/SUMB[71][1] , \mult_44/SUMB[71][2] , \mult_44/SUMB[72][1] ,
         \mult_44/SUMB[72][2] , \mult_44/SUMB[73][1] , \mult_44/SUMB[73][2] ,
         \mult_44/SUMB[74][1] , \mult_44/SUMB[74][2] , \mult_44/SUMB[75][1] ,
         \mult_44/SUMB[75][2] , \mult_44/SUMB[76][1] , \mult_44/SUMB[76][2] ,
         \mult_44/SUMB[77][1] , \mult_44/SUMB[77][2] , \mult_44/SUMB[78][1] ,
         \mult_44/SUMB[78][2] , \mult_44/SUMB[79][1] , \mult_44/SUMB[79][2] ,
         \mult_44/SUMB[80][1] , \mult_44/SUMB[80][2] , \mult_44/SUMB[81][1] ,
         \mult_44/SUMB[81][2] , \mult_44/SUMB[82][1] , \mult_44/SUMB[82][2] ,
         \mult_44/SUMB[83][1] , \mult_44/SUMB[83][2] , \mult_44/SUMB[84][1] ,
         \mult_44/SUMB[84][2] , \mult_44/SUMB[85][1] , \mult_44/SUMB[85][2] ,
         \mult_44/SUMB[86][1] , \mult_44/SUMB[86][2] , \mult_44/SUMB[87][1] ,
         \mult_44/SUMB[87][2] , \mult_44/SUMB[88][1] , \mult_44/SUMB[88][2] ,
         \mult_44/SUMB[89][1] , \mult_44/SUMB[89][2] , \mult_44/SUMB[90][1] ,
         \mult_44/SUMB[90][2] , \mult_44/SUMB[91][1] , \mult_44/SUMB[91][2] ,
         \mult_44/SUMB[92][1] , \mult_44/SUMB[92][2] , \mult_44/SUMB[93][1] ,
         \mult_44/SUMB[93][2] , \mult_44/SUMB[94][1] , \mult_44/SUMB[94][2] ,
         \mult_44/SUMB[95][1] , \mult_44/SUMB[95][2] , \mult_44/SUMB[96][1] ,
         \mult_44/SUMB[96][2] , \mult_44/SUMB[97][1] , \mult_44/SUMB[97][2] ,
         \mult_44/SUMB[98][1] , \mult_44/SUMB[98][2] , \mult_44/SUMB[99][1] ,
         \mult_44/SUMB[99][2] , \mult_44/SUMB[100][1] , \mult_44/SUMB[100][2] ,
         \mult_44/SUMB[101][1] , \mult_44/SUMB[101][2] ,
         \mult_44/SUMB[102][1] , \mult_44/SUMB[102][2] ,
         \mult_44/SUMB[103][1] , \mult_44/SUMB[103][2] ,
         \mult_44/SUMB[104][1] , \mult_44/SUMB[104][2] ,
         \mult_44/SUMB[105][1] , \mult_44/SUMB[105][2] ,
         \mult_44/SUMB[106][1] , \mult_44/SUMB[106][2] ,
         \mult_44/SUMB[107][1] , \mult_44/SUMB[107][2] ,
         \mult_44/SUMB[108][1] , \mult_44/SUMB[108][2] ,
         \mult_44/SUMB[109][1] , \mult_44/SUMB[109][2] ,
         \mult_44/SUMB[110][1] , \mult_44/SUMB[110][2] ,
         \mult_44/SUMB[111][1] , \mult_44/SUMB[111][2] ,
         \mult_44/SUMB[112][1] , \mult_44/SUMB[112][2] ,
         \mult_44/SUMB[113][1] , \mult_44/SUMB[113][2] ,
         \mult_44/SUMB[114][1] , \mult_44/SUMB[114][2] ,
         \mult_44/SUMB[115][1] , \mult_44/SUMB[115][2] ,
         \mult_44/SUMB[116][1] , \mult_44/SUMB[116][2] ,
         \mult_44/SUMB[117][1] , \mult_44/SUMB[117][2] ,
         \mult_44/SUMB[118][1] , \mult_44/SUMB[118][2] ,
         \mult_44/SUMB[119][1] , \mult_44/SUMB[119][2] ,
         \mult_44/SUMB[120][1] , \mult_44/SUMB[120][2] ,
         \mult_44/SUMB[121][1] , \mult_44/SUMB[121][2] ,
         \mult_44/SUMB[122][1] , \mult_44/SUMB[122][2] ,
         \mult_44/SUMB[123][1] , \mult_44/SUMB[123][2] ,
         \mult_44/SUMB[124][1] , \mult_44/SUMB[124][2] ,
         \mult_44/SUMB[125][1] , \mult_44/SUMB[125][2] ,
         \mult_44/SUMB[126][1] , \mult_44/SUMB[127][0] ,
         \mult_44/CARRYB[1][0] , \mult_44/CARRYB[1][1] ,
         \mult_44/CARRYB[1][2] , \mult_44/CARRYB[2][0] ,
         \mult_44/CARRYB[2][1] , \mult_44/CARRYB[2][2] ,
         \mult_44/CARRYB[3][0] , \mult_44/CARRYB[3][1] ,
         \mult_44/CARRYB[3][2] , \mult_44/CARRYB[4][0] ,
         \mult_44/CARRYB[4][1] , \mult_44/CARRYB[4][2] ,
         \mult_44/CARRYB[5][0] , \mult_44/CARRYB[5][1] ,
         \mult_44/CARRYB[5][2] , \mult_44/CARRYB[6][0] ,
         \mult_44/CARRYB[6][1] , \mult_44/CARRYB[6][2] ,
         \mult_44/CARRYB[7][0] , \mult_44/CARRYB[7][1] ,
         \mult_44/CARRYB[7][2] , \mult_44/CARRYB[8][0] ,
         \mult_44/CARRYB[8][1] , \mult_44/CARRYB[8][2] ,
         \mult_44/CARRYB[9][0] , \mult_44/CARRYB[9][1] ,
         \mult_44/CARRYB[9][2] , \mult_44/CARRYB[10][0] ,
         \mult_44/CARRYB[10][1] , \mult_44/CARRYB[10][2] ,
         \mult_44/CARRYB[11][0] , \mult_44/CARRYB[11][1] ,
         \mult_44/CARRYB[11][2] , \mult_44/CARRYB[12][0] ,
         \mult_44/CARRYB[12][1] , \mult_44/CARRYB[12][2] ,
         \mult_44/CARRYB[13][0] , \mult_44/CARRYB[13][1] ,
         \mult_44/CARRYB[13][2] , \mult_44/CARRYB[14][0] ,
         \mult_44/CARRYB[14][1] , \mult_44/CARRYB[14][2] ,
         \mult_44/CARRYB[15][0] , \mult_44/CARRYB[15][1] ,
         \mult_44/CARRYB[15][2] , \mult_44/CARRYB[16][0] ,
         \mult_44/CARRYB[16][1] , \mult_44/CARRYB[16][2] ,
         \mult_44/CARRYB[17][0] , \mult_44/CARRYB[17][1] ,
         \mult_44/CARRYB[17][2] , \mult_44/CARRYB[18][0] ,
         \mult_44/CARRYB[18][1] , \mult_44/CARRYB[18][2] ,
         \mult_44/CARRYB[19][0] , \mult_44/CARRYB[19][1] ,
         \mult_44/CARRYB[19][2] , \mult_44/CARRYB[20][0] ,
         \mult_44/CARRYB[20][1] , \mult_44/CARRYB[20][2] ,
         \mult_44/CARRYB[21][0] , \mult_44/CARRYB[21][1] ,
         \mult_44/CARRYB[21][2] , \mult_44/CARRYB[22][0] ,
         \mult_44/CARRYB[22][1] , \mult_44/CARRYB[22][2] ,
         \mult_44/CARRYB[23][0] , \mult_44/CARRYB[23][1] ,
         \mult_44/CARRYB[23][2] , \mult_44/CARRYB[24][0] ,
         \mult_44/CARRYB[24][1] , \mult_44/CARRYB[24][2] ,
         \mult_44/CARRYB[25][0] , \mult_44/CARRYB[25][1] ,
         \mult_44/CARRYB[25][2] , \mult_44/CARRYB[26][0] ,
         \mult_44/CARRYB[26][1] , \mult_44/CARRYB[26][2] ,
         \mult_44/CARRYB[27][0] , \mult_44/CARRYB[27][1] ,
         \mult_44/CARRYB[27][2] , \mult_44/CARRYB[28][0] ,
         \mult_44/CARRYB[28][1] , \mult_44/CARRYB[28][2] ,
         \mult_44/CARRYB[29][0] , \mult_44/CARRYB[29][1] ,
         \mult_44/CARRYB[29][2] , \mult_44/CARRYB[30][0] ,
         \mult_44/CARRYB[30][1] , \mult_44/CARRYB[30][2] ,
         \mult_44/CARRYB[31][0] , \mult_44/CARRYB[31][1] ,
         \mult_44/CARRYB[31][2] , \mult_44/CARRYB[32][0] ,
         \mult_44/CARRYB[32][1] , \mult_44/CARRYB[32][2] ,
         \mult_44/CARRYB[33][0] , \mult_44/CARRYB[33][1] ,
         \mult_44/CARRYB[33][2] , \mult_44/CARRYB[34][0] ,
         \mult_44/CARRYB[34][1] , \mult_44/CARRYB[34][2] ,
         \mult_44/CARRYB[35][0] , \mult_44/CARRYB[35][1] ,
         \mult_44/CARRYB[35][2] , \mult_44/CARRYB[36][0] ,
         \mult_44/CARRYB[36][1] , \mult_44/CARRYB[36][2] ,
         \mult_44/CARRYB[37][0] , \mult_44/CARRYB[37][1] ,
         \mult_44/CARRYB[37][2] , \mult_44/CARRYB[38][0] ,
         \mult_44/CARRYB[38][1] , \mult_44/CARRYB[38][2] ,
         \mult_44/CARRYB[39][0] , \mult_44/CARRYB[39][1] ,
         \mult_44/CARRYB[39][2] , \mult_44/CARRYB[40][0] ,
         \mult_44/CARRYB[40][1] , \mult_44/CARRYB[40][2] ,
         \mult_44/CARRYB[41][0] , \mult_44/CARRYB[41][1] ,
         \mult_44/CARRYB[41][2] , \mult_44/CARRYB[42][0] ,
         \mult_44/CARRYB[42][1] , \mult_44/CARRYB[42][2] ,
         \mult_44/CARRYB[43][0] , \mult_44/CARRYB[43][1] ,
         \mult_44/CARRYB[43][2] , \mult_44/CARRYB[44][0] ,
         \mult_44/CARRYB[44][1] , \mult_44/CARRYB[44][2] ,
         \mult_44/CARRYB[45][0] , \mult_44/CARRYB[45][1] ,
         \mult_44/CARRYB[45][2] , \mult_44/CARRYB[46][0] ,
         \mult_44/CARRYB[46][1] , \mult_44/CARRYB[46][2] ,
         \mult_44/CARRYB[47][0] , \mult_44/CARRYB[47][1] ,
         \mult_44/CARRYB[47][2] , \mult_44/CARRYB[48][0] ,
         \mult_44/CARRYB[48][1] , \mult_44/CARRYB[48][2] ,
         \mult_44/CARRYB[49][0] , \mult_44/CARRYB[49][1] ,
         \mult_44/CARRYB[49][2] , \mult_44/CARRYB[50][0] ,
         \mult_44/CARRYB[50][1] , \mult_44/CARRYB[50][2] ,
         \mult_44/CARRYB[51][0] , \mult_44/CARRYB[51][1] ,
         \mult_44/CARRYB[51][2] , \mult_44/CARRYB[52][0] ,
         \mult_44/CARRYB[52][1] , \mult_44/CARRYB[52][2] ,
         \mult_44/CARRYB[53][0] , \mult_44/CARRYB[53][1] ,
         \mult_44/CARRYB[53][2] , \mult_44/CARRYB[54][0] ,
         \mult_44/CARRYB[54][1] , \mult_44/CARRYB[54][2] ,
         \mult_44/CARRYB[55][0] , \mult_44/CARRYB[55][1] ,
         \mult_44/CARRYB[55][2] , \mult_44/CARRYB[56][0] ,
         \mult_44/CARRYB[56][1] , \mult_44/CARRYB[56][2] ,
         \mult_44/CARRYB[57][0] , \mult_44/CARRYB[57][1] ,
         \mult_44/CARRYB[57][2] , \mult_44/CARRYB[58][0] ,
         \mult_44/CARRYB[58][1] , \mult_44/CARRYB[58][2] ,
         \mult_44/CARRYB[59][0] , \mult_44/CARRYB[59][1] ,
         \mult_44/CARRYB[59][2] , \mult_44/CARRYB[60][0] ,
         \mult_44/CARRYB[60][1] , \mult_44/CARRYB[60][2] ,
         \mult_44/CARRYB[61][0] , \mult_44/CARRYB[61][1] ,
         \mult_44/CARRYB[61][2] , \mult_44/CARRYB[62][0] ,
         \mult_44/CARRYB[62][1] , \mult_44/CARRYB[62][2] ,
         \mult_44/CARRYB[63][0] , \mult_44/CARRYB[63][1] ,
         \mult_44/CARRYB[63][2] , \mult_44/CARRYB[64][0] ,
         \mult_44/CARRYB[64][1] , \mult_44/CARRYB[64][2] ,
         \mult_44/CARRYB[65][0] , \mult_44/CARRYB[65][1] ,
         \mult_44/CARRYB[65][2] , \mult_44/CARRYB[66][0] ,
         \mult_44/CARRYB[66][1] , \mult_44/CARRYB[66][2] ,
         \mult_44/CARRYB[67][0] , \mult_44/CARRYB[67][1] ,
         \mult_44/CARRYB[67][2] , \mult_44/CARRYB[68][0] ,
         \mult_44/CARRYB[68][1] , \mult_44/CARRYB[68][2] ,
         \mult_44/CARRYB[69][0] , \mult_44/CARRYB[69][1] ,
         \mult_44/CARRYB[69][2] , \mult_44/CARRYB[70][0] ,
         \mult_44/CARRYB[70][1] , \mult_44/CARRYB[70][2] ,
         \mult_44/CARRYB[71][0] , \mult_44/CARRYB[71][1] ,
         \mult_44/CARRYB[71][2] , \mult_44/CARRYB[72][0] ,
         \mult_44/CARRYB[72][1] , \mult_44/CARRYB[72][2] ,
         \mult_44/CARRYB[73][0] , \mult_44/CARRYB[73][1] ,
         \mult_44/CARRYB[73][2] , \mult_44/CARRYB[74][0] ,
         \mult_44/CARRYB[74][1] , \mult_44/CARRYB[74][2] ,
         \mult_44/CARRYB[75][0] , \mult_44/CARRYB[75][1] ,
         \mult_44/CARRYB[75][2] , \mult_44/CARRYB[76][0] ,
         \mult_44/CARRYB[76][1] , \mult_44/CARRYB[76][2] ,
         \mult_44/CARRYB[77][0] , \mult_44/CARRYB[77][1] ,
         \mult_44/CARRYB[77][2] , \mult_44/CARRYB[78][0] ,
         \mult_44/CARRYB[78][1] , \mult_44/CARRYB[78][2] ,
         \mult_44/CARRYB[79][0] , \mult_44/CARRYB[79][1] ,
         \mult_44/CARRYB[79][2] , \mult_44/CARRYB[80][0] ,
         \mult_44/CARRYB[80][1] , \mult_44/CARRYB[80][2] ,
         \mult_44/CARRYB[81][0] , \mult_44/CARRYB[81][1] ,
         \mult_44/CARRYB[81][2] , \mult_44/CARRYB[82][0] ,
         \mult_44/CARRYB[82][1] , \mult_44/CARRYB[82][2] ,
         \mult_44/CARRYB[83][0] , \mult_44/CARRYB[83][1] ,
         \mult_44/CARRYB[83][2] , \mult_44/CARRYB[84][0] ,
         \mult_44/CARRYB[84][1] , \mult_44/CARRYB[84][2] ,
         \mult_44/CARRYB[85][0] , \mult_44/CARRYB[85][1] ,
         \mult_44/CARRYB[85][2] , \mult_44/CARRYB[86][0] ,
         \mult_44/CARRYB[86][1] , \mult_44/CARRYB[86][2] ,
         \mult_44/CARRYB[87][0] , \mult_44/CARRYB[87][1] ,
         \mult_44/CARRYB[87][2] , \mult_44/CARRYB[88][0] ,
         \mult_44/CARRYB[88][1] , \mult_44/CARRYB[88][2] ,
         \mult_44/CARRYB[89][0] , \mult_44/CARRYB[89][1] ,
         \mult_44/CARRYB[89][2] , \mult_44/CARRYB[90][0] ,
         \mult_44/CARRYB[90][1] , \mult_44/CARRYB[90][2] ,
         \mult_44/CARRYB[91][0] , \mult_44/CARRYB[91][1] ,
         \mult_44/CARRYB[91][2] , \mult_44/CARRYB[92][0] ,
         \mult_44/CARRYB[92][1] , \mult_44/CARRYB[92][2] ,
         \mult_44/CARRYB[93][0] , \mult_44/CARRYB[93][1] ,
         \mult_44/CARRYB[93][2] , \mult_44/CARRYB[94][0] ,
         \mult_44/CARRYB[94][1] , \mult_44/CARRYB[94][2] ,
         \mult_44/CARRYB[95][0] , \mult_44/CARRYB[95][1] ,
         \mult_44/CARRYB[95][2] , \mult_44/CARRYB[96][0] ,
         \mult_44/CARRYB[96][1] , \mult_44/CARRYB[96][2] ,
         \mult_44/CARRYB[97][0] , \mult_44/CARRYB[97][1] ,
         \mult_44/CARRYB[97][2] , \mult_44/CARRYB[98][0] ,
         \mult_44/CARRYB[98][1] , \mult_44/CARRYB[98][2] ,
         \mult_44/CARRYB[99][0] , \mult_44/CARRYB[99][1] ,
         \mult_44/CARRYB[99][2] , \mult_44/CARRYB[100][0] ,
         \mult_44/CARRYB[100][1] , \mult_44/CARRYB[100][2] ,
         \mult_44/CARRYB[101][0] , \mult_44/CARRYB[101][1] ,
         \mult_44/CARRYB[101][2] , \mult_44/CARRYB[102][0] ,
         \mult_44/CARRYB[102][1] , \mult_44/CARRYB[102][2] ,
         \mult_44/CARRYB[103][0] , \mult_44/CARRYB[103][1] ,
         \mult_44/CARRYB[103][2] , \mult_44/CARRYB[104][0] ,
         \mult_44/CARRYB[104][1] , \mult_44/CARRYB[104][2] ,
         \mult_44/CARRYB[105][0] , \mult_44/CARRYB[105][1] ,
         \mult_44/CARRYB[105][2] , \mult_44/CARRYB[106][0] ,
         \mult_44/CARRYB[106][1] , \mult_44/CARRYB[106][2] ,
         \mult_44/CARRYB[107][0] , \mult_44/CARRYB[107][1] ,
         \mult_44/CARRYB[107][2] , \mult_44/CARRYB[108][0] ,
         \mult_44/CARRYB[108][1] , \mult_44/CARRYB[108][2] ,
         \mult_44/CARRYB[109][0] , \mult_44/CARRYB[109][1] ,
         \mult_44/CARRYB[109][2] , \mult_44/CARRYB[110][0] ,
         \mult_44/CARRYB[110][1] , \mult_44/CARRYB[110][2] ,
         \mult_44/CARRYB[111][0] , \mult_44/CARRYB[111][1] ,
         \mult_44/CARRYB[111][2] , \mult_44/CARRYB[112][0] ,
         \mult_44/CARRYB[112][1] , \mult_44/CARRYB[112][2] ,
         \mult_44/CARRYB[113][0] , \mult_44/CARRYB[113][1] ,
         \mult_44/CARRYB[113][2] , \mult_44/CARRYB[114][0] ,
         \mult_44/CARRYB[114][1] , \mult_44/CARRYB[114][2] ,
         \mult_44/CARRYB[115][0] , \mult_44/CARRYB[115][1] ,
         \mult_44/CARRYB[115][2] , \mult_44/CARRYB[116][0] ,
         \mult_44/CARRYB[116][1] , \mult_44/CARRYB[116][2] ,
         \mult_44/CARRYB[117][0] , \mult_44/CARRYB[117][1] ,
         \mult_44/CARRYB[117][2] , \mult_44/CARRYB[118][0] ,
         \mult_44/CARRYB[118][1] , \mult_44/CARRYB[118][2] ,
         \mult_44/CARRYB[119][0] , \mult_44/CARRYB[119][1] ,
         \mult_44/CARRYB[119][2] , \mult_44/CARRYB[120][0] ,
         \mult_44/CARRYB[120][1] , \mult_44/CARRYB[120][2] ,
         \mult_44/CARRYB[121][0] , \mult_44/CARRYB[121][1] ,
         \mult_44/CARRYB[121][2] , \mult_44/CARRYB[122][0] ,
         \mult_44/CARRYB[122][1] , \mult_44/CARRYB[122][2] ,
         \mult_44/CARRYB[123][0] , \mult_44/CARRYB[123][1] ,
         \mult_44/CARRYB[123][2] , \mult_44/CARRYB[124][0] ,
         \mult_44/CARRYB[124][1] , \mult_44/CARRYB[124][2] ,
         \mult_44/CARRYB[125][0] , \mult_44/CARRYB[125][1] ,
         \mult_44/CARRYB[126][0] , \mult_44/ab[0][1] , \mult_44/ab[0][2] ,
         \mult_44/ab[0][3] , \mult_44/ab[1][0] , \mult_44/ab[1][1] ,
         \mult_44/ab[1][2] , \mult_44/ab[1][3] , \mult_44/ab[2][0] ,
         \mult_44/ab[2][1] , \mult_44/ab[2][2] , \mult_44/ab[2][3] ,
         \mult_44/ab[3][0] , \mult_44/ab[3][1] , \mult_44/ab[3][2] ,
         \mult_44/ab[3][3] , \mult_44/ab[4][0] , \mult_44/ab[4][1] ,
         \mult_44/ab[4][2] , \mult_44/ab[4][3] , \mult_44/ab[5][0] ,
         \mult_44/ab[5][1] , \mult_44/ab[5][2] , \mult_44/ab[5][3] ,
         \mult_44/ab[6][0] , \mult_44/ab[6][1] , \mult_44/ab[6][2] ,
         \mult_44/ab[6][3] , \mult_44/ab[7][0] , \mult_44/ab[7][1] ,
         \mult_44/ab[7][2] , \mult_44/ab[7][3] , \mult_44/ab[8][0] ,
         \mult_44/ab[8][1] , \mult_44/ab[8][2] , \mult_44/ab[8][3] ,
         \mult_44/ab[9][0] , \mult_44/ab[9][1] , \mult_44/ab[9][2] ,
         \mult_44/ab[9][3] , \mult_44/ab[10][0] , \mult_44/ab[10][1] ,
         \mult_44/ab[10][2] , \mult_44/ab[10][3] , \mult_44/ab[11][0] ,
         \mult_44/ab[11][1] , \mult_44/ab[11][2] , \mult_44/ab[11][3] ,
         \mult_44/ab[12][0] , \mult_44/ab[12][1] , \mult_44/ab[12][2] ,
         \mult_44/ab[12][3] , \mult_44/ab[13][0] , \mult_44/ab[13][1] ,
         \mult_44/ab[13][2] , \mult_44/ab[13][3] , \mult_44/ab[14][0] ,
         \mult_44/ab[14][1] , \mult_44/ab[14][2] , \mult_44/ab[14][3] ,
         \mult_44/ab[15][0] , \mult_44/ab[15][1] , \mult_44/ab[15][2] ,
         \mult_44/ab[15][3] , \mult_44/ab[16][0] , \mult_44/ab[16][1] ,
         \mult_44/ab[16][2] , \mult_44/ab[16][3] , \mult_44/ab[17][0] ,
         \mult_44/ab[17][1] , \mult_44/ab[17][2] , \mult_44/ab[17][3] ,
         \mult_44/ab[18][0] , \mult_44/ab[18][1] , \mult_44/ab[18][2] ,
         \mult_44/ab[18][3] , \mult_44/ab[19][0] , \mult_44/ab[19][1] ,
         \mult_44/ab[19][2] , \mult_44/ab[19][3] , \mult_44/ab[20][0] ,
         \mult_44/ab[20][1] , \mult_44/ab[20][2] , \mult_44/ab[20][3] ,
         \mult_44/ab[21][0] , \mult_44/ab[21][1] , \mult_44/ab[21][2] ,
         \mult_44/ab[21][3] , \mult_44/ab[22][0] , \mult_44/ab[22][1] ,
         \mult_44/ab[22][2] , \mult_44/ab[22][3] , \mult_44/ab[23][0] ,
         \mult_44/ab[23][1] , \mult_44/ab[23][2] , \mult_44/ab[23][3] ,
         \mult_44/ab[24][0] , \mult_44/ab[24][1] , \mult_44/ab[24][2] ,
         \mult_44/ab[24][3] , \mult_44/ab[25][0] , \mult_44/ab[25][1] ,
         \mult_44/ab[25][2] , \mult_44/ab[25][3] , \mult_44/ab[26][0] ,
         \mult_44/ab[26][1] , \mult_44/ab[26][2] , \mult_44/ab[26][3] ,
         \mult_44/ab[27][0] , \mult_44/ab[27][1] , \mult_44/ab[27][2] ,
         \mult_44/ab[27][3] , \mult_44/ab[28][0] , \mult_44/ab[28][1] ,
         \mult_44/ab[28][2] , \mult_44/ab[28][3] , \mult_44/ab[29][0] ,
         \mult_44/ab[29][1] , \mult_44/ab[29][2] , \mult_44/ab[29][3] ,
         \mult_44/ab[30][0] , \mult_44/ab[30][1] , \mult_44/ab[30][2] ,
         \mult_44/ab[30][3] , \mult_44/ab[31][0] , \mult_44/ab[31][1] ,
         \mult_44/ab[31][2] , \mult_44/ab[31][3] , \mult_44/ab[32][0] ,
         \mult_44/ab[32][1] , \mult_44/ab[32][2] , \mult_44/ab[32][3] ,
         \mult_44/ab[33][0] , \mult_44/ab[33][1] , \mult_44/ab[33][2] ,
         \mult_44/ab[33][3] , \mult_44/ab[34][0] , \mult_44/ab[34][1] ,
         \mult_44/ab[34][2] , \mult_44/ab[34][3] , \mult_44/ab[35][0] ,
         \mult_44/ab[35][1] , \mult_44/ab[35][2] , \mult_44/ab[35][3] ,
         \mult_44/ab[36][0] , \mult_44/ab[36][1] , \mult_44/ab[36][2] ,
         \mult_44/ab[36][3] , \mult_44/ab[37][0] , \mult_44/ab[37][1] ,
         \mult_44/ab[37][2] , \mult_44/ab[37][3] , \mult_44/ab[38][0] ,
         \mult_44/ab[38][1] , \mult_44/ab[38][2] , \mult_44/ab[38][3] ,
         \mult_44/ab[39][0] , \mult_44/ab[39][1] , \mult_44/ab[39][2] ,
         \mult_44/ab[39][3] , \mult_44/ab[40][0] , \mult_44/ab[40][1] ,
         \mult_44/ab[40][2] , \mult_44/ab[40][3] , \mult_44/ab[41][0] ,
         \mult_44/ab[41][1] , \mult_44/ab[41][2] , \mult_44/ab[41][3] ,
         \mult_44/ab[42][0] , \mult_44/ab[42][1] , \mult_44/ab[42][2] ,
         \mult_44/ab[42][3] , \mult_44/ab[43][0] , \mult_44/ab[43][1] ,
         \mult_44/ab[43][2] , \mult_44/ab[43][3] , \mult_44/ab[44][0] ,
         \mult_44/ab[44][1] , \mult_44/ab[44][2] , \mult_44/ab[44][3] ,
         \mult_44/ab[45][0] , \mult_44/ab[45][1] , \mult_44/ab[45][2] ,
         \mult_44/ab[45][3] , \mult_44/ab[46][0] , \mult_44/ab[46][1] ,
         \mult_44/ab[46][2] , \mult_44/ab[46][3] , \mult_44/ab[47][0] ,
         \mult_44/ab[47][1] , \mult_44/ab[47][2] , \mult_44/ab[47][3] ,
         \mult_44/ab[48][0] , \mult_44/ab[48][1] , \mult_44/ab[48][2] ,
         \mult_44/ab[48][3] , \mult_44/ab[49][0] , \mult_44/ab[49][1] ,
         \mult_44/ab[49][2] , \mult_44/ab[49][3] , \mult_44/ab[50][0] ,
         \mult_44/ab[50][1] , \mult_44/ab[50][2] , \mult_44/ab[50][3] ,
         \mult_44/ab[51][0] , \mult_44/ab[51][1] , \mult_44/ab[51][2] ,
         \mult_44/ab[51][3] , \mult_44/ab[52][0] , \mult_44/ab[52][1] ,
         \mult_44/ab[52][2] , \mult_44/ab[52][3] , \mult_44/ab[53][0] ,
         \mult_44/ab[53][1] , \mult_44/ab[53][2] , \mult_44/ab[53][3] ,
         \mult_44/ab[54][0] , \mult_44/ab[54][1] , \mult_44/ab[54][2] ,
         \mult_44/ab[54][3] , \mult_44/ab[55][0] , \mult_44/ab[55][1] ,
         \mult_44/ab[55][2] , \mult_44/ab[55][3] , \mult_44/ab[56][0] ,
         \mult_44/ab[56][1] , \mult_44/ab[56][2] , \mult_44/ab[56][3] ,
         \mult_44/ab[57][0] , \mult_44/ab[57][1] , \mult_44/ab[57][2] ,
         \mult_44/ab[57][3] , \mult_44/ab[58][0] , \mult_44/ab[58][1] ,
         \mult_44/ab[58][2] , \mult_44/ab[58][3] , \mult_44/ab[59][0] ,
         \mult_44/ab[59][1] , \mult_44/ab[59][2] , \mult_44/ab[59][3] ,
         \mult_44/ab[60][0] , \mult_44/ab[60][1] , \mult_44/ab[60][2] ,
         \mult_44/ab[60][3] , \mult_44/ab[61][0] , \mult_44/ab[61][1] ,
         \mult_44/ab[61][2] , \mult_44/ab[61][3] , \mult_44/ab[62][0] ,
         \mult_44/ab[62][1] , \mult_44/ab[62][2] , \mult_44/ab[62][3] ,
         \mult_44/ab[63][0] , \mult_44/ab[63][1] , \mult_44/ab[63][2] ,
         \mult_44/ab[63][3] , \mult_44/ab[64][0] , \mult_44/ab[64][1] ,
         \mult_44/ab[64][2] , \mult_44/ab[64][3] , \mult_44/ab[65][0] ,
         \mult_44/ab[65][1] , \mult_44/ab[65][2] , \mult_44/ab[65][3] ,
         \mult_44/ab[66][0] , \mult_44/ab[66][1] , \mult_44/ab[66][2] ,
         \mult_44/ab[66][3] , \mult_44/ab[67][0] , \mult_44/ab[67][1] ,
         \mult_44/ab[67][2] , \mult_44/ab[67][3] , \mult_44/ab[68][0] ,
         \mult_44/ab[68][1] , \mult_44/ab[68][2] , \mult_44/ab[68][3] ,
         \mult_44/ab[69][0] , \mult_44/ab[69][1] , \mult_44/ab[69][2] ,
         \mult_44/ab[69][3] , \mult_44/ab[70][0] , \mult_44/ab[70][1] ,
         \mult_44/ab[70][2] , \mult_44/ab[70][3] , \mult_44/ab[71][0] ,
         \mult_44/ab[71][1] , \mult_44/ab[71][2] , \mult_44/ab[71][3] ,
         \mult_44/ab[72][0] , \mult_44/ab[72][1] , \mult_44/ab[72][2] ,
         \mult_44/ab[72][3] , \mult_44/ab[73][0] , \mult_44/ab[73][1] ,
         \mult_44/ab[73][2] , \mult_44/ab[73][3] , \mult_44/ab[74][0] ,
         \mult_44/ab[74][1] , \mult_44/ab[74][2] , \mult_44/ab[74][3] ,
         \mult_44/ab[75][0] , \mult_44/ab[75][1] , \mult_44/ab[75][2] ,
         \mult_44/ab[75][3] , \mult_44/ab[76][0] , \mult_44/ab[76][1] ,
         \mult_44/ab[76][2] , \mult_44/ab[76][3] , \mult_44/ab[77][0] ,
         \mult_44/ab[77][1] , \mult_44/ab[77][2] , \mult_44/ab[77][3] ,
         \mult_44/ab[78][0] , \mult_44/ab[78][1] , \mult_44/ab[78][2] ,
         \mult_44/ab[78][3] , \mult_44/ab[79][0] , \mult_44/ab[79][1] ,
         \mult_44/ab[79][2] , \mult_44/ab[79][3] , \mult_44/ab[80][0] ,
         \mult_44/ab[80][1] , \mult_44/ab[80][2] , \mult_44/ab[80][3] ,
         \mult_44/ab[81][0] , \mult_44/ab[81][1] , \mult_44/ab[81][2] ,
         \mult_44/ab[81][3] , \mult_44/ab[82][0] , \mult_44/ab[82][1] ,
         \mult_44/ab[82][2] , \mult_44/ab[82][3] , \mult_44/ab[83][0] ,
         \mult_44/ab[83][1] , \mult_44/ab[83][2] , \mult_44/ab[83][3] ,
         \mult_44/ab[84][0] , \mult_44/ab[84][1] , \mult_44/ab[84][2] ,
         \mult_44/ab[84][3] , \mult_44/ab[85][0] , \mult_44/ab[85][1] ,
         \mult_44/ab[85][2] , \mult_44/ab[85][3] , \mult_44/ab[86][0] ,
         \mult_44/ab[86][1] , \mult_44/ab[86][2] , \mult_44/ab[86][3] ,
         \mult_44/ab[87][0] , \mult_44/ab[87][1] , \mult_44/ab[87][2] ,
         \mult_44/ab[87][3] , \mult_44/ab[88][0] , \mult_44/ab[88][1] ,
         \mult_44/ab[88][2] , \mult_44/ab[88][3] , \mult_44/ab[89][0] ,
         \mult_44/ab[89][1] , \mult_44/ab[89][2] , \mult_44/ab[89][3] ,
         \mult_44/ab[90][0] , \mult_44/ab[90][1] , \mult_44/ab[90][2] ,
         \mult_44/ab[90][3] , \mult_44/ab[91][0] , \mult_44/ab[91][1] ,
         \mult_44/ab[91][2] , \mult_44/ab[91][3] , \mult_44/ab[92][0] ,
         \mult_44/ab[92][1] , \mult_44/ab[92][2] , \mult_44/ab[92][3] ,
         \mult_44/ab[93][0] , \mult_44/ab[93][1] , \mult_44/ab[93][2] ,
         \mult_44/ab[93][3] , \mult_44/ab[94][0] , \mult_44/ab[94][1] ,
         \mult_44/ab[94][2] , \mult_44/ab[94][3] , \mult_44/ab[95][0] ,
         \mult_44/ab[95][1] , \mult_44/ab[95][2] , \mult_44/ab[95][3] ,
         \mult_44/ab[96][0] , \mult_44/ab[96][1] , \mult_44/ab[96][2] ,
         \mult_44/ab[96][3] , \mult_44/ab[97][0] , \mult_44/ab[97][1] ,
         \mult_44/ab[97][2] , \mult_44/ab[97][3] , \mult_44/ab[98][0] ,
         \mult_44/ab[98][1] , \mult_44/ab[98][2] , \mult_44/ab[98][3] ,
         \mult_44/ab[99][0] , \mult_44/ab[99][1] , \mult_44/ab[99][2] ,
         \mult_44/ab[99][3] , \mult_44/ab[100][0] , \mult_44/ab[100][1] ,
         \mult_44/ab[100][2] , \mult_44/ab[100][3] , \mult_44/ab[101][0] ,
         \mult_44/ab[101][1] , \mult_44/ab[101][2] , \mult_44/ab[101][3] ,
         \mult_44/ab[102][0] , \mult_44/ab[102][1] , \mult_44/ab[102][2] ,
         \mult_44/ab[102][3] , \mult_44/ab[103][0] , \mult_44/ab[103][1] ,
         \mult_44/ab[103][2] , \mult_44/ab[103][3] , \mult_44/ab[104][0] ,
         \mult_44/ab[104][1] , \mult_44/ab[104][2] , \mult_44/ab[104][3] ,
         \mult_44/ab[105][0] , \mult_44/ab[105][1] , \mult_44/ab[105][2] ,
         \mult_44/ab[105][3] , \mult_44/ab[106][0] , \mult_44/ab[106][1] ,
         \mult_44/ab[106][2] , \mult_44/ab[106][3] , \mult_44/ab[107][0] ,
         \mult_44/ab[107][1] , \mult_44/ab[107][2] , \mult_44/ab[107][3] ,
         \mult_44/ab[108][0] , \mult_44/ab[108][1] , \mult_44/ab[108][2] ,
         \mult_44/ab[108][3] , \mult_44/ab[109][0] , \mult_44/ab[109][1] ,
         \mult_44/ab[109][2] , \mult_44/ab[109][3] , \mult_44/ab[110][0] ,
         \mult_44/ab[110][1] , \mult_44/ab[110][2] , \mult_44/ab[110][3] ,
         \mult_44/ab[111][0] , \mult_44/ab[111][1] , \mult_44/ab[111][2] ,
         \mult_44/ab[111][3] , \mult_44/ab[112][0] , \mult_44/ab[112][1] ,
         \mult_44/ab[112][2] , \mult_44/ab[112][3] , \mult_44/ab[113][0] ,
         \mult_44/ab[113][1] , \mult_44/ab[113][2] , \mult_44/ab[113][3] ,
         \mult_44/ab[114][0] , \mult_44/ab[114][1] , \mult_44/ab[114][2] ,
         \mult_44/ab[114][3] , \mult_44/ab[115][0] , \mult_44/ab[115][1] ,
         \mult_44/ab[115][2] , \mult_44/ab[115][3] , \mult_44/ab[116][0] ,
         \mult_44/ab[116][1] , \mult_44/ab[116][2] , \mult_44/ab[116][3] ,
         \mult_44/ab[117][0] , \mult_44/ab[117][1] , \mult_44/ab[117][2] ,
         \mult_44/ab[117][3] , \mult_44/ab[118][0] , \mult_44/ab[118][1] ,
         \mult_44/ab[118][2] , \mult_44/ab[118][3] , \mult_44/ab[119][0] ,
         \mult_44/ab[119][1] , \mult_44/ab[119][2] , \mult_44/ab[119][3] ,
         \mult_44/ab[120][0] , \mult_44/ab[120][1] , \mult_44/ab[120][2] ,
         \mult_44/ab[120][3] , \mult_44/ab[121][0] , \mult_44/ab[121][1] ,
         \mult_44/ab[121][2] , \mult_44/ab[121][3] , \mult_44/ab[122][0] ,
         \mult_44/ab[122][1] , \mult_44/ab[122][2] , \mult_44/ab[122][3] ,
         \mult_44/ab[123][0] , \mult_44/ab[123][1] , \mult_44/ab[123][2] ,
         \mult_44/ab[123][3] , \mult_44/ab[124][0] , \mult_44/ab[124][1] ,
         \mult_44/ab[124][2] , \mult_44/ab[124][3] , \mult_44/ab[125][0] ,
         \mult_44/ab[125][1] , \mult_44/ab[125][2] , \mult_44/ab[126][0] ,
         \mult_44/ab[126][1] , \mult_44/ab[127][0] , n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625;
  wire   [127:4] swire;
  wire   [255:128] sreg;
  wire   [127:0] clocal;

  DFF \sreg_reg[128]  ( .D(swire[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[128]) );
  DFF \sreg_reg[129]  ( .D(swire[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[129]) );
  DFF \sreg_reg[130]  ( .D(swire[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[130]) );
  DFF \sreg_reg[131]  ( .D(swire[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[131]) );
  DFF \sreg_reg[132]  ( .D(swire[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[132]) );
  DFF \sreg_reg[133]  ( .D(swire[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[133]) );
  DFF \sreg_reg[134]  ( .D(swire[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[134]) );
  DFF \sreg_reg[135]  ( .D(swire[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[135]) );
  DFF \sreg_reg[136]  ( .D(swire[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[136]) );
  DFF \sreg_reg[137]  ( .D(swire[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[137]) );
  DFF \sreg_reg[138]  ( .D(swire[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[138]) );
  DFF \sreg_reg[139]  ( .D(swire[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[139]) );
  DFF \sreg_reg[140]  ( .D(swire[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[140]) );
  DFF \sreg_reg[141]  ( .D(swire[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[141]) );
  DFF \sreg_reg[142]  ( .D(swire[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[142]) );
  DFF \sreg_reg[143]  ( .D(swire[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[143]) );
  DFF \sreg_reg[144]  ( .D(swire[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[144]) );
  DFF \sreg_reg[145]  ( .D(swire[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[145]) );
  DFF \sreg_reg[146]  ( .D(swire[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[146]) );
  DFF \sreg_reg[147]  ( .D(swire[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[147]) );
  DFF \sreg_reg[148]  ( .D(swire[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[148]) );
  DFF \sreg_reg[149]  ( .D(swire[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[149]) );
  DFF \sreg_reg[150]  ( .D(swire[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[150]) );
  DFF \sreg_reg[151]  ( .D(swire[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[151]) );
  DFF \sreg_reg[152]  ( .D(swire[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[152]) );
  DFF \sreg_reg[153]  ( .D(swire[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[153]) );
  DFF \sreg_reg[154]  ( .D(swire[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[154]) );
  DFF \sreg_reg[155]  ( .D(swire[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[155]) );
  DFF \sreg_reg[156]  ( .D(swire[32]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[156]) );
  DFF \sreg_reg[157]  ( .D(swire[33]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[157]) );
  DFF \sreg_reg[158]  ( .D(swire[34]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[158]) );
  DFF \sreg_reg[159]  ( .D(swire[35]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[159]) );
  DFF \sreg_reg[160]  ( .D(swire[36]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[160]) );
  DFF \sreg_reg[161]  ( .D(swire[37]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[161]) );
  DFF \sreg_reg[162]  ( .D(swire[38]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[162]) );
  DFF \sreg_reg[163]  ( .D(swire[39]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[163]) );
  DFF \sreg_reg[164]  ( .D(swire[40]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[164]) );
  DFF \sreg_reg[165]  ( .D(swire[41]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[165]) );
  DFF \sreg_reg[166]  ( .D(swire[42]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[166]) );
  DFF \sreg_reg[167]  ( .D(swire[43]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[167]) );
  DFF \sreg_reg[168]  ( .D(swire[44]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[168]) );
  DFF \sreg_reg[169]  ( .D(swire[45]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[169]) );
  DFF \sreg_reg[170]  ( .D(swire[46]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[170]) );
  DFF \sreg_reg[171]  ( .D(swire[47]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[171]) );
  DFF \sreg_reg[172]  ( .D(swire[48]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[172]) );
  DFF \sreg_reg[173]  ( .D(swire[49]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[173]) );
  DFF \sreg_reg[174]  ( .D(swire[50]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[174]) );
  DFF \sreg_reg[175]  ( .D(swire[51]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[175]) );
  DFF \sreg_reg[176]  ( .D(swire[52]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[176]) );
  DFF \sreg_reg[177]  ( .D(swire[53]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[177]) );
  DFF \sreg_reg[178]  ( .D(swire[54]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[178]) );
  DFF \sreg_reg[179]  ( .D(swire[55]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[179]) );
  DFF \sreg_reg[180]  ( .D(swire[56]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[180]) );
  DFF \sreg_reg[181]  ( .D(swire[57]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[181]) );
  DFF \sreg_reg[182]  ( .D(swire[58]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[182]) );
  DFF \sreg_reg[183]  ( .D(swire[59]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[183]) );
  DFF \sreg_reg[184]  ( .D(swire[60]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[184]) );
  DFF \sreg_reg[185]  ( .D(swire[61]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[185]) );
  DFF \sreg_reg[186]  ( .D(swire[62]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[186]) );
  DFF \sreg_reg[187]  ( .D(swire[63]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[187]) );
  DFF \sreg_reg[188]  ( .D(swire[64]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[188]) );
  DFF \sreg_reg[189]  ( .D(swire[65]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[189]) );
  DFF \sreg_reg[190]  ( .D(swire[66]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[190]) );
  DFF \sreg_reg[191]  ( .D(swire[67]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[191]) );
  DFF \sreg_reg[192]  ( .D(swire[68]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[192]) );
  DFF \sreg_reg[193]  ( .D(swire[69]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[193]) );
  DFF \sreg_reg[194]  ( .D(swire[70]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[194]) );
  DFF \sreg_reg[195]  ( .D(swire[71]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[195]) );
  DFF \sreg_reg[196]  ( .D(swire[72]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[196]) );
  DFF \sreg_reg[197]  ( .D(swire[73]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[197]) );
  DFF \sreg_reg[198]  ( .D(swire[74]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[198]) );
  DFF \sreg_reg[199]  ( .D(swire[75]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[199]) );
  DFF \sreg_reg[200]  ( .D(swire[76]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[200]) );
  DFF \sreg_reg[201]  ( .D(swire[77]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[201]) );
  DFF \sreg_reg[202]  ( .D(swire[78]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[202]) );
  DFF \sreg_reg[203]  ( .D(swire[79]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[203]) );
  DFF \sreg_reg[204]  ( .D(swire[80]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[204]) );
  DFF \sreg_reg[205]  ( .D(swire[81]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[205]) );
  DFF \sreg_reg[206]  ( .D(swire[82]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[206]) );
  DFF \sreg_reg[207]  ( .D(swire[83]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[207]) );
  DFF \sreg_reg[208]  ( .D(swire[84]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[208]) );
  DFF \sreg_reg[209]  ( .D(swire[85]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[209]) );
  DFF \sreg_reg[210]  ( .D(swire[86]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[210]) );
  DFF \sreg_reg[211]  ( .D(swire[87]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[211]) );
  DFF \sreg_reg[212]  ( .D(swire[88]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[212]) );
  DFF \sreg_reg[213]  ( .D(swire[89]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[213]) );
  DFF \sreg_reg[214]  ( .D(swire[90]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[214]) );
  DFF \sreg_reg[215]  ( .D(swire[91]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[215]) );
  DFF \sreg_reg[216]  ( .D(swire[92]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[216]) );
  DFF \sreg_reg[217]  ( .D(swire[93]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[217]) );
  DFF \sreg_reg[218]  ( .D(swire[94]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[218]) );
  DFF \sreg_reg[219]  ( .D(swire[95]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[219]) );
  DFF \sreg_reg[220]  ( .D(swire[96]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[220]) );
  DFF \sreg_reg[221]  ( .D(swire[97]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[221]) );
  DFF \sreg_reg[222]  ( .D(swire[98]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[222]) );
  DFF \sreg_reg[223]  ( .D(swire[99]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[223]) );
  DFF \sreg_reg[224]  ( .D(swire[100]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[224]) );
  DFF \sreg_reg[225]  ( .D(swire[101]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[225]) );
  DFF \sreg_reg[226]  ( .D(swire[102]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[226]) );
  DFF \sreg_reg[227]  ( .D(swire[103]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[227]) );
  DFF \sreg_reg[228]  ( .D(swire[104]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[228]) );
  DFF \sreg_reg[229]  ( .D(swire[105]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[229]) );
  DFF \sreg_reg[230]  ( .D(swire[106]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[230]) );
  DFF \sreg_reg[231]  ( .D(swire[107]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[231]) );
  DFF \sreg_reg[232]  ( .D(swire[108]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[232]) );
  DFF \sreg_reg[233]  ( .D(swire[109]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[233]) );
  DFF \sreg_reg[234]  ( .D(swire[110]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[234]) );
  DFF \sreg_reg[235]  ( .D(swire[111]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[235]) );
  DFF \sreg_reg[236]  ( .D(swire[112]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[236]) );
  DFF \sreg_reg[237]  ( .D(swire[113]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[237]) );
  DFF \sreg_reg[238]  ( .D(swire[114]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[238]) );
  DFF \sreg_reg[239]  ( .D(swire[115]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[239]) );
  DFF \sreg_reg[240]  ( .D(swire[116]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[240]) );
  DFF \sreg_reg[241]  ( .D(swire[117]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[241]) );
  DFF \sreg_reg[242]  ( .D(swire[118]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[242]) );
  DFF \sreg_reg[243]  ( .D(swire[119]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[243]) );
  DFF \sreg_reg[244]  ( .D(swire[120]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[244]) );
  DFF \sreg_reg[245]  ( .D(swire[121]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[245]) );
  DFF \sreg_reg[246]  ( .D(swire[122]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[246]) );
  DFF \sreg_reg[247]  ( .D(swire[123]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[247]) );
  DFF \sreg_reg[248]  ( .D(swire[124]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[248]) );
  DFF \sreg_reg[249]  ( .D(swire[125]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[249]) );
  DFF \sreg_reg[250]  ( .D(swire[126]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[250]) );
  DFF \sreg_reg[251]  ( .D(swire[127]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[251]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[123])
         );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[122])
         );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[121])
         );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[120])
         );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[119])
         );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[118])
         );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[117])
         );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[116])
         );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[115])
         );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[114])
         );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[113])
         );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[112])
         );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[111])
         );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[110])
         );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[109])
         );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[108])
         );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[107])
         );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[106])
         );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[105])
         );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[104])
         );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[103])
         );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[102])
         );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[101])
         );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[100])
         );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[99])
         );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[98])
         );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[97])
         );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[96])
         );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[95]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[94]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[93]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[92]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[91]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[90]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[89]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[88]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[87]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[86]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[85]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[84]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[83]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[82]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[81]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[80]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[79]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[78]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[77]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[76]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[75]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[74]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[73]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[72]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[71]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[70]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[69]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[68]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[67]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[66]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[65]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[64]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[63]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[62]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[61]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[60]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[59]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[58]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[57]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[56]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[55]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[54]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[53]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[52]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[51]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[50]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[49]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[48]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[47]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[46]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[45]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[44]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[43]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[42]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[41]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[40]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[39]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[38]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[37]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[36]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[35]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[34]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[33]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[32]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[31]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[30]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[29]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[28]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[27]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[26]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[25]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[24]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[23]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[22]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[21]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[20]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[19]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[18]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[17]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[16]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[15]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[14]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[13]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[12]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[11]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[10]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[9]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[8]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[7]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[6]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[5]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[4]) );
  DFF \sreg_reg[7]  ( .D(c[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[3]) );
  DFF \sreg_reg[6]  ( .D(c[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[2]) );
  DFF \sreg_reg[5]  ( .D(c[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[1]) );
  DFF \sreg_reg[4]  ( .D(c[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[0]) );
  FADDER \mult_44/S3_2_2  ( .CIN(\mult_44/ab[2][2] ), .IN0(
        \mult_44/CARRYB[1][2] ), .IN1(\mult_44/ab[1][3] ), .COUT(
        \mult_44/CARRYB[2][2] ), .SUM(\mult_44/SUMB[2][2] ) );
  FADDER \mult_44/S2_2_1  ( .CIN(\mult_44/ab[2][1] ), .IN0(
        \mult_44/CARRYB[1][1] ), .IN1(\mult_44/SUMB[1][2] ), .COUT(
        \mult_44/CARRYB[2][1] ), .SUM(\mult_44/SUMB[2][1] ) );
  FADDER \mult_44/S1_2_0  ( .CIN(\mult_44/ab[2][0] ), .IN0(
        \mult_44/CARRYB[1][0] ), .IN1(\mult_44/SUMB[1][1] ), .COUT(
        \mult_44/CARRYB[2][0] ), .SUM(clocal[2]) );
  FADDER \mult_44/S3_3_2  ( .CIN(\mult_44/ab[3][2] ), .IN0(
        \mult_44/CARRYB[2][2] ), .IN1(\mult_44/ab[2][3] ), .COUT(
        \mult_44/CARRYB[3][2] ), .SUM(\mult_44/SUMB[3][2] ) );
  FADDER \mult_44/S2_3_1  ( .CIN(\mult_44/ab[3][1] ), .IN0(
        \mult_44/CARRYB[2][1] ), .IN1(\mult_44/SUMB[2][2] ), .COUT(
        \mult_44/CARRYB[3][1] ), .SUM(\mult_44/SUMB[3][1] ) );
  FADDER \mult_44/S1_3_0  ( .CIN(\mult_44/ab[3][0] ), .IN0(
        \mult_44/CARRYB[2][0] ), .IN1(\mult_44/SUMB[2][1] ), .COUT(
        \mult_44/CARRYB[3][0] ), .SUM(\mult_44/PROD1[3] ) );
  FADDER \mult_44/S3_4_2  ( .CIN(\mult_44/ab[4][2] ), .IN0(
        \mult_44/CARRYB[3][2] ), .IN1(\mult_44/ab[3][3] ), .COUT(
        \mult_44/CARRYB[4][2] ), .SUM(\mult_44/SUMB[4][2] ) );
  FADDER \mult_44/S2_4_1  ( .CIN(\mult_44/ab[4][1] ), .IN0(
        \mult_44/CARRYB[3][1] ), .IN1(\mult_44/SUMB[3][2] ), .COUT(
        \mult_44/CARRYB[4][1] ), .SUM(\mult_44/SUMB[4][1] ) );
  FADDER \mult_44/S1_4_0  ( .CIN(\mult_44/ab[4][0] ), .IN0(
        \mult_44/CARRYB[3][0] ), .IN1(\mult_44/SUMB[3][1] ), .COUT(
        \mult_44/CARRYB[4][0] ), .SUM(clocal[4]) );
  FADDER \mult_44/S3_5_2  ( .CIN(\mult_44/ab[5][2] ), .IN0(
        \mult_44/CARRYB[4][2] ), .IN1(\mult_44/ab[4][3] ), .COUT(
        \mult_44/CARRYB[5][2] ), .SUM(\mult_44/SUMB[5][2] ) );
  FADDER \mult_44/S2_5_1  ( .CIN(\mult_44/ab[5][1] ), .IN0(
        \mult_44/CARRYB[4][1] ), .IN1(\mult_44/SUMB[4][2] ), .COUT(
        \mult_44/CARRYB[5][1] ), .SUM(\mult_44/SUMB[5][1] ) );
  FADDER \mult_44/S1_5_0  ( .CIN(\mult_44/ab[5][0] ), .IN0(
        \mult_44/CARRYB[4][0] ), .IN1(\mult_44/SUMB[4][1] ), .COUT(
        \mult_44/CARRYB[5][0] ), .SUM(clocal[5]) );
  FADDER \mult_44/S3_6_2  ( .CIN(\mult_44/ab[6][2] ), .IN0(
        \mult_44/CARRYB[5][2] ), .IN1(\mult_44/ab[5][3] ), .COUT(
        \mult_44/CARRYB[6][2] ), .SUM(\mult_44/SUMB[6][2] ) );
  FADDER \mult_44/S2_6_1  ( .CIN(\mult_44/ab[6][1] ), .IN0(
        \mult_44/CARRYB[5][1] ), .IN1(\mult_44/SUMB[5][2] ), .COUT(
        \mult_44/CARRYB[6][1] ), .SUM(\mult_44/SUMB[6][1] ) );
  FADDER \mult_44/S1_6_0  ( .CIN(\mult_44/ab[6][0] ), .IN0(
        \mult_44/CARRYB[5][0] ), .IN1(\mult_44/SUMB[5][1] ), .COUT(
        \mult_44/CARRYB[6][0] ), .SUM(clocal[6]) );
  FADDER \mult_44/S3_7_2  ( .CIN(\mult_44/ab[7][2] ), .IN0(
        \mult_44/CARRYB[6][2] ), .IN1(\mult_44/ab[6][3] ), .COUT(
        \mult_44/CARRYB[7][2] ), .SUM(\mult_44/SUMB[7][2] ) );
  FADDER \mult_44/S2_7_1  ( .CIN(\mult_44/ab[7][1] ), .IN0(
        \mult_44/CARRYB[6][1] ), .IN1(\mult_44/SUMB[6][2] ), .COUT(
        \mult_44/CARRYB[7][1] ), .SUM(\mult_44/SUMB[7][1] ) );
  FADDER \mult_44/S1_7_0  ( .CIN(\mult_44/ab[7][0] ), .IN0(
        \mult_44/CARRYB[6][0] ), .IN1(\mult_44/SUMB[6][1] ), .COUT(
        \mult_44/CARRYB[7][0] ), .SUM(clocal[7]) );
  FADDER \mult_44/S3_8_2  ( .CIN(\mult_44/ab[8][2] ), .IN0(
        \mult_44/CARRYB[7][2] ), .IN1(\mult_44/ab[7][3] ), .COUT(
        \mult_44/CARRYB[8][2] ), .SUM(\mult_44/SUMB[8][2] ) );
  FADDER \mult_44/S2_8_1  ( .CIN(\mult_44/ab[8][1] ), .IN0(
        \mult_44/CARRYB[7][1] ), .IN1(\mult_44/SUMB[7][2] ), .COUT(
        \mult_44/CARRYB[8][1] ), .SUM(\mult_44/SUMB[8][1] ) );
  FADDER \mult_44/S1_8_0  ( .CIN(\mult_44/ab[8][0] ), .IN0(
        \mult_44/CARRYB[7][0] ), .IN1(\mult_44/SUMB[7][1] ), .COUT(
        \mult_44/CARRYB[8][0] ), .SUM(clocal[8]) );
  FADDER \mult_44/S3_9_2  ( .CIN(\mult_44/ab[9][2] ), .IN0(
        \mult_44/CARRYB[8][2] ), .IN1(\mult_44/ab[8][3] ), .COUT(
        \mult_44/CARRYB[9][2] ), .SUM(\mult_44/SUMB[9][2] ) );
  FADDER \mult_44/S2_9_1  ( .CIN(\mult_44/ab[9][1] ), .IN0(
        \mult_44/CARRYB[8][1] ), .IN1(\mult_44/SUMB[8][2] ), .COUT(
        \mult_44/CARRYB[9][1] ), .SUM(\mult_44/SUMB[9][1] ) );
  FADDER \mult_44/S1_9_0  ( .CIN(\mult_44/ab[9][0] ), .IN0(
        \mult_44/CARRYB[8][0] ), .IN1(\mult_44/SUMB[8][1] ), .COUT(
        \mult_44/CARRYB[9][0] ), .SUM(clocal[9]) );
  FADDER \mult_44/S3_10_2  ( .CIN(\mult_44/ab[10][2] ), .IN0(
        \mult_44/CARRYB[9][2] ), .IN1(\mult_44/ab[9][3] ), .COUT(
        \mult_44/CARRYB[10][2] ), .SUM(\mult_44/SUMB[10][2] ) );
  FADDER \mult_44/S2_10_1  ( .CIN(\mult_44/ab[10][1] ), .IN0(
        \mult_44/CARRYB[9][1] ), .IN1(\mult_44/SUMB[9][2] ), .COUT(
        \mult_44/CARRYB[10][1] ), .SUM(\mult_44/SUMB[10][1] ) );
  FADDER \mult_44/S1_10_0  ( .CIN(\mult_44/ab[10][0] ), .IN0(
        \mult_44/CARRYB[9][0] ), .IN1(\mult_44/SUMB[9][1] ), .COUT(
        \mult_44/CARRYB[10][0] ), .SUM(clocal[10]) );
  FADDER \mult_44/S3_11_2  ( .CIN(\mult_44/ab[11][2] ), .IN0(
        \mult_44/CARRYB[10][2] ), .IN1(\mult_44/ab[10][3] ), .COUT(
        \mult_44/CARRYB[11][2] ), .SUM(\mult_44/SUMB[11][2] ) );
  FADDER \mult_44/S2_11_1  ( .CIN(\mult_44/ab[11][1] ), .IN0(
        \mult_44/CARRYB[10][1] ), .IN1(\mult_44/SUMB[10][2] ), .COUT(
        \mult_44/CARRYB[11][1] ), .SUM(\mult_44/SUMB[11][1] ) );
  FADDER \mult_44/S1_11_0  ( .CIN(\mult_44/ab[11][0] ), .IN0(
        \mult_44/CARRYB[10][0] ), .IN1(\mult_44/SUMB[10][1] ), .COUT(
        \mult_44/CARRYB[11][0] ), .SUM(clocal[11]) );
  FADDER \mult_44/S3_12_2  ( .CIN(\mult_44/ab[12][2] ), .IN0(
        \mult_44/CARRYB[11][2] ), .IN1(\mult_44/ab[11][3] ), .COUT(
        \mult_44/CARRYB[12][2] ), .SUM(\mult_44/SUMB[12][2] ) );
  FADDER \mult_44/S2_12_1  ( .CIN(\mult_44/ab[12][1] ), .IN0(
        \mult_44/CARRYB[11][1] ), .IN1(\mult_44/SUMB[11][2] ), .COUT(
        \mult_44/CARRYB[12][1] ), .SUM(\mult_44/SUMB[12][1] ) );
  FADDER \mult_44/S1_12_0  ( .CIN(\mult_44/ab[12][0] ), .IN0(
        \mult_44/CARRYB[11][0] ), .IN1(\mult_44/SUMB[11][1] ), .COUT(
        \mult_44/CARRYB[12][0] ), .SUM(clocal[12]) );
  FADDER \mult_44/S3_13_2  ( .CIN(\mult_44/ab[13][2] ), .IN0(
        \mult_44/CARRYB[12][2] ), .IN1(\mult_44/ab[12][3] ), .COUT(
        \mult_44/CARRYB[13][2] ), .SUM(\mult_44/SUMB[13][2] ) );
  FADDER \mult_44/S2_13_1  ( .CIN(\mult_44/ab[13][1] ), .IN0(
        \mult_44/CARRYB[12][1] ), .IN1(\mult_44/SUMB[12][2] ), .COUT(
        \mult_44/CARRYB[13][1] ), .SUM(\mult_44/SUMB[13][1] ) );
  FADDER \mult_44/S1_13_0  ( .CIN(\mult_44/ab[13][0] ), .IN0(
        \mult_44/CARRYB[12][0] ), .IN1(\mult_44/SUMB[12][1] ), .COUT(
        \mult_44/CARRYB[13][0] ), .SUM(clocal[13]) );
  FADDER \mult_44/S3_14_2  ( .CIN(\mult_44/ab[14][2] ), .IN0(
        \mult_44/CARRYB[13][2] ), .IN1(\mult_44/ab[13][3] ), .COUT(
        \mult_44/CARRYB[14][2] ), .SUM(\mult_44/SUMB[14][2] ) );
  FADDER \mult_44/S2_14_1  ( .CIN(\mult_44/ab[14][1] ), .IN0(
        \mult_44/CARRYB[13][1] ), .IN1(\mult_44/SUMB[13][2] ), .COUT(
        \mult_44/CARRYB[14][1] ), .SUM(\mult_44/SUMB[14][1] ) );
  FADDER \mult_44/S1_14_0  ( .CIN(\mult_44/ab[14][0] ), .IN0(
        \mult_44/CARRYB[13][0] ), .IN1(\mult_44/SUMB[13][1] ), .COUT(
        \mult_44/CARRYB[14][0] ), .SUM(clocal[14]) );
  FADDER \mult_44/S3_15_2  ( .CIN(\mult_44/ab[15][2] ), .IN0(
        \mult_44/CARRYB[14][2] ), .IN1(\mult_44/ab[14][3] ), .COUT(
        \mult_44/CARRYB[15][2] ), .SUM(\mult_44/SUMB[15][2] ) );
  FADDER \mult_44/S2_15_1  ( .CIN(\mult_44/ab[15][1] ), .IN0(
        \mult_44/CARRYB[14][1] ), .IN1(\mult_44/SUMB[14][2] ), .COUT(
        \mult_44/CARRYB[15][1] ), .SUM(\mult_44/SUMB[15][1] ) );
  FADDER \mult_44/S1_15_0  ( .CIN(\mult_44/ab[15][0] ), .IN0(
        \mult_44/CARRYB[14][0] ), .IN1(\mult_44/SUMB[14][1] ), .COUT(
        \mult_44/CARRYB[15][0] ), .SUM(clocal[15]) );
  FADDER \mult_44/S3_16_2  ( .CIN(\mult_44/ab[16][2] ), .IN0(
        \mult_44/CARRYB[15][2] ), .IN1(\mult_44/ab[15][3] ), .COUT(
        \mult_44/CARRYB[16][2] ), .SUM(\mult_44/SUMB[16][2] ) );
  FADDER \mult_44/S2_16_1  ( .CIN(\mult_44/ab[16][1] ), .IN0(
        \mult_44/CARRYB[15][1] ), .IN1(\mult_44/SUMB[15][2] ), .COUT(
        \mult_44/CARRYB[16][1] ), .SUM(\mult_44/SUMB[16][1] ) );
  FADDER \mult_44/S1_16_0  ( .CIN(\mult_44/ab[16][0] ), .IN0(
        \mult_44/CARRYB[15][0] ), .IN1(\mult_44/SUMB[15][1] ), .COUT(
        \mult_44/CARRYB[16][0] ), .SUM(clocal[16]) );
  FADDER \mult_44/S3_17_2  ( .CIN(\mult_44/ab[17][2] ), .IN0(
        \mult_44/CARRYB[16][2] ), .IN1(\mult_44/ab[16][3] ), .COUT(
        \mult_44/CARRYB[17][2] ), .SUM(\mult_44/SUMB[17][2] ) );
  FADDER \mult_44/S2_17_1  ( .CIN(\mult_44/ab[17][1] ), .IN0(
        \mult_44/CARRYB[16][1] ), .IN1(\mult_44/SUMB[16][2] ), .COUT(
        \mult_44/CARRYB[17][1] ), .SUM(\mult_44/SUMB[17][1] ) );
  FADDER \mult_44/S1_17_0  ( .CIN(\mult_44/ab[17][0] ), .IN0(
        \mult_44/CARRYB[16][0] ), .IN1(\mult_44/SUMB[16][1] ), .COUT(
        \mult_44/CARRYB[17][0] ), .SUM(clocal[17]) );
  FADDER \mult_44/S3_18_2  ( .CIN(\mult_44/ab[18][2] ), .IN0(
        \mult_44/CARRYB[17][2] ), .IN1(\mult_44/ab[17][3] ), .COUT(
        \mult_44/CARRYB[18][2] ), .SUM(\mult_44/SUMB[18][2] ) );
  FADDER \mult_44/S2_18_1  ( .CIN(\mult_44/ab[18][1] ), .IN0(
        \mult_44/CARRYB[17][1] ), .IN1(\mult_44/SUMB[17][2] ), .COUT(
        \mult_44/CARRYB[18][1] ), .SUM(\mult_44/SUMB[18][1] ) );
  FADDER \mult_44/S1_18_0  ( .CIN(\mult_44/ab[18][0] ), .IN0(
        \mult_44/CARRYB[17][0] ), .IN1(\mult_44/SUMB[17][1] ), .COUT(
        \mult_44/CARRYB[18][0] ), .SUM(clocal[18]) );
  FADDER \mult_44/S3_19_2  ( .CIN(\mult_44/ab[19][2] ), .IN0(
        \mult_44/CARRYB[18][2] ), .IN1(\mult_44/ab[18][3] ), .COUT(
        \mult_44/CARRYB[19][2] ), .SUM(\mult_44/SUMB[19][2] ) );
  FADDER \mult_44/S2_19_1  ( .CIN(\mult_44/ab[19][1] ), .IN0(
        \mult_44/CARRYB[18][1] ), .IN1(\mult_44/SUMB[18][2] ), .COUT(
        \mult_44/CARRYB[19][1] ), .SUM(\mult_44/SUMB[19][1] ) );
  FADDER \mult_44/S1_19_0  ( .CIN(\mult_44/ab[19][0] ), .IN0(
        \mult_44/CARRYB[18][0] ), .IN1(\mult_44/SUMB[18][1] ), .COUT(
        \mult_44/CARRYB[19][0] ), .SUM(clocal[19]) );
  FADDER \mult_44/S3_20_2  ( .CIN(\mult_44/ab[20][2] ), .IN0(
        \mult_44/CARRYB[19][2] ), .IN1(\mult_44/ab[19][3] ), .COUT(
        \mult_44/CARRYB[20][2] ), .SUM(\mult_44/SUMB[20][2] ) );
  FADDER \mult_44/S2_20_1  ( .CIN(\mult_44/ab[20][1] ), .IN0(
        \mult_44/CARRYB[19][1] ), .IN1(\mult_44/SUMB[19][2] ), .COUT(
        \mult_44/CARRYB[20][1] ), .SUM(\mult_44/SUMB[20][1] ) );
  FADDER \mult_44/S1_20_0  ( .CIN(\mult_44/ab[20][0] ), .IN0(
        \mult_44/CARRYB[19][0] ), .IN1(\mult_44/SUMB[19][1] ), .COUT(
        \mult_44/CARRYB[20][0] ), .SUM(clocal[20]) );
  FADDER \mult_44/S3_21_2  ( .CIN(\mult_44/ab[21][2] ), .IN0(
        \mult_44/CARRYB[20][2] ), .IN1(\mult_44/ab[20][3] ), .COUT(
        \mult_44/CARRYB[21][2] ), .SUM(\mult_44/SUMB[21][2] ) );
  FADDER \mult_44/S2_21_1  ( .CIN(\mult_44/ab[21][1] ), .IN0(
        \mult_44/CARRYB[20][1] ), .IN1(\mult_44/SUMB[20][2] ), .COUT(
        \mult_44/CARRYB[21][1] ), .SUM(\mult_44/SUMB[21][1] ) );
  FADDER \mult_44/S1_21_0  ( .CIN(\mult_44/ab[21][0] ), .IN0(
        \mult_44/CARRYB[20][0] ), .IN1(\mult_44/SUMB[20][1] ), .COUT(
        \mult_44/CARRYB[21][0] ), .SUM(clocal[21]) );
  FADDER \mult_44/S3_22_2  ( .CIN(\mult_44/ab[22][2] ), .IN0(
        \mult_44/CARRYB[21][2] ), .IN1(\mult_44/ab[21][3] ), .COUT(
        \mult_44/CARRYB[22][2] ), .SUM(\mult_44/SUMB[22][2] ) );
  FADDER \mult_44/S2_22_1  ( .CIN(\mult_44/ab[22][1] ), .IN0(
        \mult_44/CARRYB[21][1] ), .IN1(\mult_44/SUMB[21][2] ), .COUT(
        \mult_44/CARRYB[22][1] ), .SUM(\mult_44/SUMB[22][1] ) );
  FADDER \mult_44/S1_22_0  ( .CIN(\mult_44/ab[22][0] ), .IN0(
        \mult_44/CARRYB[21][0] ), .IN1(\mult_44/SUMB[21][1] ), .COUT(
        \mult_44/CARRYB[22][0] ), .SUM(clocal[22]) );
  FADDER \mult_44/S3_23_2  ( .CIN(\mult_44/ab[23][2] ), .IN0(
        \mult_44/CARRYB[22][2] ), .IN1(\mult_44/ab[22][3] ), .COUT(
        \mult_44/CARRYB[23][2] ), .SUM(\mult_44/SUMB[23][2] ) );
  FADDER \mult_44/S2_23_1  ( .CIN(\mult_44/ab[23][1] ), .IN0(
        \mult_44/CARRYB[22][1] ), .IN1(\mult_44/SUMB[22][2] ), .COUT(
        \mult_44/CARRYB[23][1] ), .SUM(\mult_44/SUMB[23][1] ) );
  FADDER \mult_44/S1_23_0  ( .CIN(\mult_44/ab[23][0] ), .IN0(
        \mult_44/CARRYB[22][0] ), .IN1(\mult_44/SUMB[22][1] ), .COUT(
        \mult_44/CARRYB[23][0] ), .SUM(clocal[23]) );
  FADDER \mult_44/S3_24_2  ( .CIN(\mult_44/ab[24][2] ), .IN0(
        \mult_44/CARRYB[23][2] ), .IN1(\mult_44/ab[23][3] ), .COUT(
        \mult_44/CARRYB[24][2] ), .SUM(\mult_44/SUMB[24][2] ) );
  FADDER \mult_44/S2_24_1  ( .CIN(\mult_44/ab[24][1] ), .IN0(
        \mult_44/CARRYB[23][1] ), .IN1(\mult_44/SUMB[23][2] ), .COUT(
        \mult_44/CARRYB[24][1] ), .SUM(\mult_44/SUMB[24][1] ) );
  FADDER \mult_44/S1_24_0  ( .CIN(\mult_44/ab[24][0] ), .IN0(
        \mult_44/CARRYB[23][0] ), .IN1(\mult_44/SUMB[23][1] ), .COUT(
        \mult_44/CARRYB[24][0] ), .SUM(clocal[24]) );
  FADDER \mult_44/S3_25_2  ( .CIN(\mult_44/ab[25][2] ), .IN0(
        \mult_44/CARRYB[24][2] ), .IN1(\mult_44/ab[24][3] ), .COUT(
        \mult_44/CARRYB[25][2] ), .SUM(\mult_44/SUMB[25][2] ) );
  FADDER \mult_44/S2_25_1  ( .CIN(\mult_44/ab[25][1] ), .IN0(
        \mult_44/CARRYB[24][1] ), .IN1(\mult_44/SUMB[24][2] ), .COUT(
        \mult_44/CARRYB[25][1] ), .SUM(\mult_44/SUMB[25][1] ) );
  FADDER \mult_44/S1_25_0  ( .CIN(\mult_44/ab[25][0] ), .IN0(
        \mult_44/CARRYB[24][0] ), .IN1(\mult_44/SUMB[24][1] ), .COUT(
        \mult_44/CARRYB[25][0] ), .SUM(clocal[25]) );
  FADDER \mult_44/S3_26_2  ( .CIN(\mult_44/ab[26][2] ), .IN0(
        \mult_44/CARRYB[25][2] ), .IN1(\mult_44/ab[25][3] ), .COUT(
        \mult_44/CARRYB[26][2] ), .SUM(\mult_44/SUMB[26][2] ) );
  FADDER \mult_44/S2_26_1  ( .CIN(\mult_44/ab[26][1] ), .IN0(
        \mult_44/CARRYB[25][1] ), .IN1(\mult_44/SUMB[25][2] ), .COUT(
        \mult_44/CARRYB[26][1] ), .SUM(\mult_44/SUMB[26][1] ) );
  FADDER \mult_44/S1_26_0  ( .CIN(\mult_44/ab[26][0] ), .IN0(
        \mult_44/CARRYB[25][0] ), .IN1(\mult_44/SUMB[25][1] ), .COUT(
        \mult_44/CARRYB[26][0] ), .SUM(clocal[26]) );
  FADDER \mult_44/S3_27_2  ( .CIN(\mult_44/ab[27][2] ), .IN0(
        \mult_44/CARRYB[26][2] ), .IN1(\mult_44/ab[26][3] ), .COUT(
        \mult_44/CARRYB[27][2] ), .SUM(\mult_44/SUMB[27][2] ) );
  FADDER \mult_44/S2_27_1  ( .CIN(\mult_44/ab[27][1] ), .IN0(
        \mult_44/CARRYB[26][1] ), .IN1(\mult_44/SUMB[26][2] ), .COUT(
        \mult_44/CARRYB[27][1] ), .SUM(\mult_44/SUMB[27][1] ) );
  FADDER \mult_44/S1_27_0  ( .CIN(\mult_44/ab[27][0] ), .IN0(
        \mult_44/CARRYB[26][0] ), .IN1(\mult_44/SUMB[26][1] ), .COUT(
        \mult_44/CARRYB[27][0] ), .SUM(clocal[27]) );
  FADDER \mult_44/S3_28_2  ( .CIN(\mult_44/ab[28][2] ), .IN0(
        \mult_44/CARRYB[27][2] ), .IN1(\mult_44/ab[27][3] ), .COUT(
        \mult_44/CARRYB[28][2] ), .SUM(\mult_44/SUMB[28][2] ) );
  FADDER \mult_44/S2_28_1  ( .CIN(\mult_44/ab[28][1] ), .IN0(
        \mult_44/CARRYB[27][1] ), .IN1(\mult_44/SUMB[27][2] ), .COUT(
        \mult_44/CARRYB[28][1] ), .SUM(\mult_44/SUMB[28][1] ) );
  FADDER \mult_44/S1_28_0  ( .CIN(\mult_44/ab[28][0] ), .IN0(
        \mult_44/CARRYB[27][0] ), .IN1(\mult_44/SUMB[27][1] ), .COUT(
        \mult_44/CARRYB[28][0] ), .SUM(clocal[28]) );
  FADDER \mult_44/S3_29_2  ( .CIN(\mult_44/ab[29][2] ), .IN0(
        \mult_44/CARRYB[28][2] ), .IN1(\mult_44/ab[28][3] ), .COUT(
        \mult_44/CARRYB[29][2] ), .SUM(\mult_44/SUMB[29][2] ) );
  FADDER \mult_44/S2_29_1  ( .CIN(\mult_44/ab[29][1] ), .IN0(
        \mult_44/CARRYB[28][1] ), .IN1(\mult_44/SUMB[28][2] ), .COUT(
        \mult_44/CARRYB[29][1] ), .SUM(\mult_44/SUMB[29][1] ) );
  FADDER \mult_44/S1_29_0  ( .CIN(\mult_44/ab[29][0] ), .IN0(
        \mult_44/CARRYB[28][0] ), .IN1(\mult_44/SUMB[28][1] ), .COUT(
        \mult_44/CARRYB[29][0] ), .SUM(clocal[29]) );
  FADDER \mult_44/S3_30_2  ( .CIN(\mult_44/ab[30][2] ), .IN0(
        \mult_44/CARRYB[29][2] ), .IN1(\mult_44/ab[29][3] ), .COUT(
        \mult_44/CARRYB[30][2] ), .SUM(\mult_44/SUMB[30][2] ) );
  FADDER \mult_44/S2_30_1  ( .CIN(\mult_44/ab[30][1] ), .IN0(
        \mult_44/CARRYB[29][1] ), .IN1(\mult_44/SUMB[29][2] ), .COUT(
        \mult_44/CARRYB[30][1] ), .SUM(\mult_44/SUMB[30][1] ) );
  FADDER \mult_44/S1_30_0  ( .CIN(\mult_44/ab[30][0] ), .IN0(
        \mult_44/CARRYB[29][0] ), .IN1(\mult_44/SUMB[29][1] ), .COUT(
        \mult_44/CARRYB[30][0] ), .SUM(clocal[30]) );
  FADDER \mult_44/S3_31_2  ( .CIN(\mult_44/ab[31][2] ), .IN0(
        \mult_44/CARRYB[30][2] ), .IN1(\mult_44/ab[30][3] ), .COUT(
        \mult_44/CARRYB[31][2] ), .SUM(\mult_44/SUMB[31][2] ) );
  FADDER \mult_44/S2_31_1  ( .CIN(\mult_44/ab[31][1] ), .IN0(
        \mult_44/CARRYB[30][1] ), .IN1(\mult_44/SUMB[30][2] ), .COUT(
        \mult_44/CARRYB[31][1] ), .SUM(\mult_44/SUMB[31][1] ) );
  FADDER \mult_44/S1_31_0  ( .CIN(\mult_44/ab[31][0] ), .IN0(
        \mult_44/CARRYB[30][0] ), .IN1(\mult_44/SUMB[30][1] ), .COUT(
        \mult_44/CARRYB[31][0] ), .SUM(clocal[31]) );
  FADDER \mult_44/S3_32_2  ( .CIN(\mult_44/ab[32][2] ), .IN0(
        \mult_44/CARRYB[31][2] ), .IN1(\mult_44/ab[31][3] ), .COUT(
        \mult_44/CARRYB[32][2] ), .SUM(\mult_44/SUMB[32][2] ) );
  FADDER \mult_44/S2_32_1  ( .CIN(\mult_44/ab[32][1] ), .IN0(
        \mult_44/CARRYB[31][1] ), .IN1(\mult_44/SUMB[31][2] ), .COUT(
        \mult_44/CARRYB[32][1] ), .SUM(\mult_44/SUMB[32][1] ) );
  FADDER \mult_44/S1_32_0  ( .CIN(\mult_44/ab[32][0] ), .IN0(
        \mult_44/CARRYB[31][0] ), .IN1(\mult_44/SUMB[31][1] ), .COUT(
        \mult_44/CARRYB[32][0] ), .SUM(clocal[32]) );
  FADDER \mult_44/S3_33_2  ( .CIN(\mult_44/ab[33][2] ), .IN0(
        \mult_44/CARRYB[32][2] ), .IN1(\mult_44/ab[32][3] ), .COUT(
        \mult_44/CARRYB[33][2] ), .SUM(\mult_44/SUMB[33][2] ) );
  FADDER \mult_44/S2_33_1  ( .CIN(\mult_44/ab[33][1] ), .IN0(
        \mult_44/CARRYB[32][1] ), .IN1(\mult_44/SUMB[32][2] ), .COUT(
        \mult_44/CARRYB[33][1] ), .SUM(\mult_44/SUMB[33][1] ) );
  FADDER \mult_44/S1_33_0  ( .CIN(\mult_44/ab[33][0] ), .IN0(
        \mult_44/CARRYB[32][0] ), .IN1(\mult_44/SUMB[32][1] ), .COUT(
        \mult_44/CARRYB[33][0] ), .SUM(clocal[33]) );
  FADDER \mult_44/S3_34_2  ( .CIN(\mult_44/ab[34][2] ), .IN0(
        \mult_44/CARRYB[33][2] ), .IN1(\mult_44/ab[33][3] ), .COUT(
        \mult_44/CARRYB[34][2] ), .SUM(\mult_44/SUMB[34][2] ) );
  FADDER \mult_44/S2_34_1  ( .CIN(\mult_44/ab[34][1] ), .IN0(
        \mult_44/CARRYB[33][1] ), .IN1(\mult_44/SUMB[33][2] ), .COUT(
        \mult_44/CARRYB[34][1] ), .SUM(\mult_44/SUMB[34][1] ) );
  FADDER \mult_44/S1_34_0  ( .CIN(\mult_44/ab[34][0] ), .IN0(
        \mult_44/CARRYB[33][0] ), .IN1(\mult_44/SUMB[33][1] ), .COUT(
        \mult_44/CARRYB[34][0] ), .SUM(clocal[34]) );
  FADDER \mult_44/S3_35_2  ( .CIN(\mult_44/ab[35][2] ), .IN0(
        \mult_44/CARRYB[34][2] ), .IN1(\mult_44/ab[34][3] ), .COUT(
        \mult_44/CARRYB[35][2] ), .SUM(\mult_44/SUMB[35][2] ) );
  FADDER \mult_44/S2_35_1  ( .CIN(\mult_44/ab[35][1] ), .IN0(
        \mult_44/CARRYB[34][1] ), .IN1(\mult_44/SUMB[34][2] ), .COUT(
        \mult_44/CARRYB[35][1] ), .SUM(\mult_44/SUMB[35][1] ) );
  FADDER \mult_44/S1_35_0  ( .CIN(\mult_44/ab[35][0] ), .IN0(
        \mult_44/CARRYB[34][0] ), .IN1(\mult_44/SUMB[34][1] ), .COUT(
        \mult_44/CARRYB[35][0] ), .SUM(clocal[35]) );
  FADDER \mult_44/S3_36_2  ( .CIN(\mult_44/ab[36][2] ), .IN0(
        \mult_44/CARRYB[35][2] ), .IN1(\mult_44/ab[35][3] ), .COUT(
        \mult_44/CARRYB[36][2] ), .SUM(\mult_44/SUMB[36][2] ) );
  FADDER \mult_44/S2_36_1  ( .CIN(\mult_44/ab[36][1] ), .IN0(
        \mult_44/CARRYB[35][1] ), .IN1(\mult_44/SUMB[35][2] ), .COUT(
        \mult_44/CARRYB[36][1] ), .SUM(\mult_44/SUMB[36][1] ) );
  FADDER \mult_44/S1_36_0  ( .CIN(\mult_44/ab[36][0] ), .IN0(
        \mult_44/CARRYB[35][0] ), .IN1(\mult_44/SUMB[35][1] ), .COUT(
        \mult_44/CARRYB[36][0] ), .SUM(clocal[36]) );
  FADDER \mult_44/S3_37_2  ( .CIN(\mult_44/ab[37][2] ), .IN0(
        \mult_44/CARRYB[36][2] ), .IN1(\mult_44/ab[36][3] ), .COUT(
        \mult_44/CARRYB[37][2] ), .SUM(\mult_44/SUMB[37][2] ) );
  FADDER \mult_44/S2_37_1  ( .CIN(\mult_44/ab[37][1] ), .IN0(
        \mult_44/CARRYB[36][1] ), .IN1(\mult_44/SUMB[36][2] ), .COUT(
        \mult_44/CARRYB[37][1] ), .SUM(\mult_44/SUMB[37][1] ) );
  FADDER \mult_44/S1_37_0  ( .CIN(\mult_44/ab[37][0] ), .IN0(
        \mult_44/CARRYB[36][0] ), .IN1(\mult_44/SUMB[36][1] ), .COUT(
        \mult_44/CARRYB[37][0] ), .SUM(clocal[37]) );
  FADDER \mult_44/S3_38_2  ( .CIN(\mult_44/ab[38][2] ), .IN0(
        \mult_44/CARRYB[37][2] ), .IN1(\mult_44/ab[37][3] ), .COUT(
        \mult_44/CARRYB[38][2] ), .SUM(\mult_44/SUMB[38][2] ) );
  FADDER \mult_44/S2_38_1  ( .CIN(\mult_44/ab[38][1] ), .IN0(
        \mult_44/CARRYB[37][1] ), .IN1(\mult_44/SUMB[37][2] ), .COUT(
        \mult_44/CARRYB[38][1] ), .SUM(\mult_44/SUMB[38][1] ) );
  FADDER \mult_44/S1_38_0  ( .CIN(\mult_44/ab[38][0] ), .IN0(
        \mult_44/CARRYB[37][0] ), .IN1(\mult_44/SUMB[37][1] ), .COUT(
        \mult_44/CARRYB[38][0] ), .SUM(clocal[38]) );
  FADDER \mult_44/S3_39_2  ( .CIN(\mult_44/ab[39][2] ), .IN0(
        \mult_44/CARRYB[38][2] ), .IN1(\mult_44/ab[38][3] ), .COUT(
        \mult_44/CARRYB[39][2] ), .SUM(\mult_44/SUMB[39][2] ) );
  FADDER \mult_44/S2_39_1  ( .CIN(\mult_44/ab[39][1] ), .IN0(
        \mult_44/CARRYB[38][1] ), .IN1(\mult_44/SUMB[38][2] ), .COUT(
        \mult_44/CARRYB[39][1] ), .SUM(\mult_44/SUMB[39][1] ) );
  FADDER \mult_44/S1_39_0  ( .CIN(\mult_44/ab[39][0] ), .IN0(
        \mult_44/CARRYB[38][0] ), .IN1(\mult_44/SUMB[38][1] ), .COUT(
        \mult_44/CARRYB[39][0] ), .SUM(clocal[39]) );
  FADDER \mult_44/S3_40_2  ( .CIN(\mult_44/ab[40][2] ), .IN0(
        \mult_44/CARRYB[39][2] ), .IN1(\mult_44/ab[39][3] ), .COUT(
        \mult_44/CARRYB[40][2] ), .SUM(\mult_44/SUMB[40][2] ) );
  FADDER \mult_44/S2_40_1  ( .CIN(\mult_44/ab[40][1] ), .IN0(
        \mult_44/CARRYB[39][1] ), .IN1(\mult_44/SUMB[39][2] ), .COUT(
        \mult_44/CARRYB[40][1] ), .SUM(\mult_44/SUMB[40][1] ) );
  FADDER \mult_44/S1_40_0  ( .CIN(\mult_44/ab[40][0] ), .IN0(
        \mult_44/CARRYB[39][0] ), .IN1(\mult_44/SUMB[39][1] ), .COUT(
        \mult_44/CARRYB[40][0] ), .SUM(clocal[40]) );
  FADDER \mult_44/S3_41_2  ( .CIN(\mult_44/ab[41][2] ), .IN0(
        \mult_44/CARRYB[40][2] ), .IN1(\mult_44/ab[40][3] ), .COUT(
        \mult_44/CARRYB[41][2] ), .SUM(\mult_44/SUMB[41][2] ) );
  FADDER \mult_44/S2_41_1  ( .CIN(\mult_44/ab[41][1] ), .IN0(
        \mult_44/CARRYB[40][1] ), .IN1(\mult_44/SUMB[40][2] ), .COUT(
        \mult_44/CARRYB[41][1] ), .SUM(\mult_44/SUMB[41][1] ) );
  FADDER \mult_44/S1_41_0  ( .CIN(\mult_44/ab[41][0] ), .IN0(
        \mult_44/CARRYB[40][0] ), .IN1(\mult_44/SUMB[40][1] ), .COUT(
        \mult_44/CARRYB[41][0] ), .SUM(clocal[41]) );
  FADDER \mult_44/S3_42_2  ( .CIN(\mult_44/ab[42][2] ), .IN0(
        \mult_44/CARRYB[41][2] ), .IN1(\mult_44/ab[41][3] ), .COUT(
        \mult_44/CARRYB[42][2] ), .SUM(\mult_44/SUMB[42][2] ) );
  FADDER \mult_44/S2_42_1  ( .CIN(\mult_44/ab[42][1] ), .IN0(
        \mult_44/CARRYB[41][1] ), .IN1(\mult_44/SUMB[41][2] ), .COUT(
        \mult_44/CARRYB[42][1] ), .SUM(\mult_44/SUMB[42][1] ) );
  FADDER \mult_44/S1_42_0  ( .CIN(\mult_44/ab[42][0] ), .IN0(
        \mult_44/CARRYB[41][0] ), .IN1(\mult_44/SUMB[41][1] ), .COUT(
        \mult_44/CARRYB[42][0] ), .SUM(clocal[42]) );
  FADDER \mult_44/S3_43_2  ( .CIN(\mult_44/ab[43][2] ), .IN0(
        \mult_44/CARRYB[42][2] ), .IN1(\mult_44/ab[42][3] ), .COUT(
        \mult_44/CARRYB[43][2] ), .SUM(\mult_44/SUMB[43][2] ) );
  FADDER \mult_44/S2_43_1  ( .CIN(\mult_44/ab[43][1] ), .IN0(
        \mult_44/CARRYB[42][1] ), .IN1(\mult_44/SUMB[42][2] ), .COUT(
        \mult_44/CARRYB[43][1] ), .SUM(\mult_44/SUMB[43][1] ) );
  FADDER \mult_44/S1_43_0  ( .CIN(\mult_44/ab[43][0] ), .IN0(
        \mult_44/CARRYB[42][0] ), .IN1(\mult_44/SUMB[42][1] ), .COUT(
        \mult_44/CARRYB[43][0] ), .SUM(clocal[43]) );
  FADDER \mult_44/S3_44_2  ( .CIN(\mult_44/ab[44][2] ), .IN0(
        \mult_44/CARRYB[43][2] ), .IN1(\mult_44/ab[43][3] ), .COUT(
        \mult_44/CARRYB[44][2] ), .SUM(\mult_44/SUMB[44][2] ) );
  FADDER \mult_44/S2_44_1  ( .CIN(\mult_44/ab[44][1] ), .IN0(
        \mult_44/CARRYB[43][1] ), .IN1(\mult_44/SUMB[43][2] ), .COUT(
        \mult_44/CARRYB[44][1] ), .SUM(\mult_44/SUMB[44][1] ) );
  FADDER \mult_44/S1_44_0  ( .CIN(\mult_44/ab[44][0] ), .IN0(
        \mult_44/CARRYB[43][0] ), .IN1(\mult_44/SUMB[43][1] ), .COUT(
        \mult_44/CARRYB[44][0] ), .SUM(clocal[44]) );
  FADDER \mult_44/S3_45_2  ( .CIN(\mult_44/ab[45][2] ), .IN0(
        \mult_44/CARRYB[44][2] ), .IN1(\mult_44/ab[44][3] ), .COUT(
        \mult_44/CARRYB[45][2] ), .SUM(\mult_44/SUMB[45][2] ) );
  FADDER \mult_44/S2_45_1  ( .CIN(\mult_44/ab[45][1] ), .IN0(
        \mult_44/CARRYB[44][1] ), .IN1(\mult_44/SUMB[44][2] ), .COUT(
        \mult_44/CARRYB[45][1] ), .SUM(\mult_44/SUMB[45][1] ) );
  FADDER \mult_44/S1_45_0  ( .CIN(\mult_44/ab[45][0] ), .IN0(
        \mult_44/CARRYB[44][0] ), .IN1(\mult_44/SUMB[44][1] ), .COUT(
        \mult_44/CARRYB[45][0] ), .SUM(clocal[45]) );
  FADDER \mult_44/S3_46_2  ( .CIN(\mult_44/ab[46][2] ), .IN0(
        \mult_44/CARRYB[45][2] ), .IN1(\mult_44/ab[45][3] ), .COUT(
        \mult_44/CARRYB[46][2] ), .SUM(\mult_44/SUMB[46][2] ) );
  FADDER \mult_44/S2_46_1  ( .CIN(\mult_44/ab[46][1] ), .IN0(
        \mult_44/CARRYB[45][1] ), .IN1(\mult_44/SUMB[45][2] ), .COUT(
        \mult_44/CARRYB[46][1] ), .SUM(\mult_44/SUMB[46][1] ) );
  FADDER \mult_44/S1_46_0  ( .CIN(\mult_44/ab[46][0] ), .IN0(
        \mult_44/CARRYB[45][0] ), .IN1(\mult_44/SUMB[45][1] ), .COUT(
        \mult_44/CARRYB[46][0] ), .SUM(clocal[46]) );
  FADDER \mult_44/S3_47_2  ( .CIN(\mult_44/ab[47][2] ), .IN0(
        \mult_44/CARRYB[46][2] ), .IN1(\mult_44/ab[46][3] ), .COUT(
        \mult_44/CARRYB[47][2] ), .SUM(\mult_44/SUMB[47][2] ) );
  FADDER \mult_44/S2_47_1  ( .CIN(\mult_44/ab[47][1] ), .IN0(
        \mult_44/CARRYB[46][1] ), .IN1(\mult_44/SUMB[46][2] ), .COUT(
        \mult_44/CARRYB[47][1] ), .SUM(\mult_44/SUMB[47][1] ) );
  FADDER \mult_44/S1_47_0  ( .CIN(\mult_44/ab[47][0] ), .IN0(
        \mult_44/CARRYB[46][0] ), .IN1(\mult_44/SUMB[46][1] ), .COUT(
        \mult_44/CARRYB[47][0] ), .SUM(clocal[47]) );
  FADDER \mult_44/S3_48_2  ( .CIN(\mult_44/ab[48][2] ), .IN0(
        \mult_44/CARRYB[47][2] ), .IN1(\mult_44/ab[47][3] ), .COUT(
        \mult_44/CARRYB[48][2] ), .SUM(\mult_44/SUMB[48][2] ) );
  FADDER \mult_44/S2_48_1  ( .CIN(\mult_44/ab[48][1] ), .IN0(
        \mult_44/CARRYB[47][1] ), .IN1(\mult_44/SUMB[47][2] ), .COUT(
        \mult_44/CARRYB[48][1] ), .SUM(\mult_44/SUMB[48][1] ) );
  FADDER \mult_44/S1_48_0  ( .CIN(\mult_44/ab[48][0] ), .IN0(
        \mult_44/CARRYB[47][0] ), .IN1(\mult_44/SUMB[47][1] ), .COUT(
        \mult_44/CARRYB[48][0] ), .SUM(clocal[48]) );
  FADDER \mult_44/S3_49_2  ( .CIN(\mult_44/ab[49][2] ), .IN0(
        \mult_44/CARRYB[48][2] ), .IN1(\mult_44/ab[48][3] ), .COUT(
        \mult_44/CARRYB[49][2] ), .SUM(\mult_44/SUMB[49][2] ) );
  FADDER \mult_44/S2_49_1  ( .CIN(\mult_44/ab[49][1] ), .IN0(
        \mult_44/CARRYB[48][1] ), .IN1(\mult_44/SUMB[48][2] ), .COUT(
        \mult_44/CARRYB[49][1] ), .SUM(\mult_44/SUMB[49][1] ) );
  FADDER \mult_44/S1_49_0  ( .CIN(\mult_44/ab[49][0] ), .IN0(
        \mult_44/CARRYB[48][0] ), .IN1(\mult_44/SUMB[48][1] ), .COUT(
        \mult_44/CARRYB[49][0] ), .SUM(clocal[49]) );
  FADDER \mult_44/S3_50_2  ( .CIN(\mult_44/ab[50][2] ), .IN0(
        \mult_44/CARRYB[49][2] ), .IN1(\mult_44/ab[49][3] ), .COUT(
        \mult_44/CARRYB[50][2] ), .SUM(\mult_44/SUMB[50][2] ) );
  FADDER \mult_44/S2_50_1  ( .CIN(\mult_44/ab[50][1] ), .IN0(
        \mult_44/CARRYB[49][1] ), .IN1(\mult_44/SUMB[49][2] ), .COUT(
        \mult_44/CARRYB[50][1] ), .SUM(\mult_44/SUMB[50][1] ) );
  FADDER \mult_44/S1_50_0  ( .CIN(\mult_44/ab[50][0] ), .IN0(
        \mult_44/CARRYB[49][0] ), .IN1(\mult_44/SUMB[49][1] ), .COUT(
        \mult_44/CARRYB[50][0] ), .SUM(clocal[50]) );
  FADDER \mult_44/S3_51_2  ( .CIN(\mult_44/ab[51][2] ), .IN0(
        \mult_44/CARRYB[50][2] ), .IN1(\mult_44/ab[50][3] ), .COUT(
        \mult_44/CARRYB[51][2] ), .SUM(\mult_44/SUMB[51][2] ) );
  FADDER \mult_44/S2_51_1  ( .CIN(\mult_44/ab[51][1] ), .IN0(
        \mult_44/CARRYB[50][1] ), .IN1(\mult_44/SUMB[50][2] ), .COUT(
        \mult_44/CARRYB[51][1] ), .SUM(\mult_44/SUMB[51][1] ) );
  FADDER \mult_44/S1_51_0  ( .CIN(\mult_44/ab[51][0] ), .IN0(
        \mult_44/CARRYB[50][0] ), .IN1(\mult_44/SUMB[50][1] ), .COUT(
        \mult_44/CARRYB[51][0] ), .SUM(clocal[51]) );
  FADDER \mult_44/S3_52_2  ( .CIN(\mult_44/ab[52][2] ), .IN0(
        \mult_44/CARRYB[51][2] ), .IN1(\mult_44/ab[51][3] ), .COUT(
        \mult_44/CARRYB[52][2] ), .SUM(\mult_44/SUMB[52][2] ) );
  FADDER \mult_44/S2_52_1  ( .CIN(\mult_44/ab[52][1] ), .IN0(
        \mult_44/CARRYB[51][1] ), .IN1(\mult_44/SUMB[51][2] ), .COUT(
        \mult_44/CARRYB[52][1] ), .SUM(\mult_44/SUMB[52][1] ) );
  FADDER \mult_44/S1_52_0  ( .CIN(\mult_44/ab[52][0] ), .IN0(
        \mult_44/CARRYB[51][0] ), .IN1(\mult_44/SUMB[51][1] ), .COUT(
        \mult_44/CARRYB[52][0] ), .SUM(clocal[52]) );
  FADDER \mult_44/S3_53_2  ( .CIN(\mult_44/ab[53][2] ), .IN0(
        \mult_44/CARRYB[52][2] ), .IN1(\mult_44/ab[52][3] ), .COUT(
        \mult_44/CARRYB[53][2] ), .SUM(\mult_44/SUMB[53][2] ) );
  FADDER \mult_44/S2_53_1  ( .CIN(\mult_44/ab[53][1] ), .IN0(
        \mult_44/CARRYB[52][1] ), .IN1(\mult_44/SUMB[52][2] ), .COUT(
        \mult_44/CARRYB[53][1] ), .SUM(\mult_44/SUMB[53][1] ) );
  FADDER \mult_44/S1_53_0  ( .CIN(\mult_44/ab[53][0] ), .IN0(
        \mult_44/CARRYB[52][0] ), .IN1(\mult_44/SUMB[52][1] ), .COUT(
        \mult_44/CARRYB[53][0] ), .SUM(clocal[53]) );
  FADDER \mult_44/S3_54_2  ( .CIN(\mult_44/ab[54][2] ), .IN0(
        \mult_44/CARRYB[53][2] ), .IN1(\mult_44/ab[53][3] ), .COUT(
        \mult_44/CARRYB[54][2] ), .SUM(\mult_44/SUMB[54][2] ) );
  FADDER \mult_44/S2_54_1  ( .CIN(\mult_44/ab[54][1] ), .IN0(
        \mult_44/CARRYB[53][1] ), .IN1(\mult_44/SUMB[53][2] ), .COUT(
        \mult_44/CARRYB[54][1] ), .SUM(\mult_44/SUMB[54][1] ) );
  FADDER \mult_44/S1_54_0  ( .CIN(\mult_44/ab[54][0] ), .IN0(
        \mult_44/CARRYB[53][0] ), .IN1(\mult_44/SUMB[53][1] ), .COUT(
        \mult_44/CARRYB[54][0] ), .SUM(clocal[54]) );
  FADDER \mult_44/S3_55_2  ( .CIN(\mult_44/ab[55][2] ), .IN0(
        \mult_44/CARRYB[54][2] ), .IN1(\mult_44/ab[54][3] ), .COUT(
        \mult_44/CARRYB[55][2] ), .SUM(\mult_44/SUMB[55][2] ) );
  FADDER \mult_44/S2_55_1  ( .CIN(\mult_44/ab[55][1] ), .IN0(
        \mult_44/CARRYB[54][1] ), .IN1(\mult_44/SUMB[54][2] ), .COUT(
        \mult_44/CARRYB[55][1] ), .SUM(\mult_44/SUMB[55][1] ) );
  FADDER \mult_44/S1_55_0  ( .CIN(\mult_44/ab[55][0] ), .IN0(
        \mult_44/CARRYB[54][0] ), .IN1(\mult_44/SUMB[54][1] ), .COUT(
        \mult_44/CARRYB[55][0] ), .SUM(clocal[55]) );
  FADDER \mult_44/S3_56_2  ( .CIN(\mult_44/ab[56][2] ), .IN0(
        \mult_44/CARRYB[55][2] ), .IN1(\mult_44/ab[55][3] ), .COUT(
        \mult_44/CARRYB[56][2] ), .SUM(\mult_44/SUMB[56][2] ) );
  FADDER \mult_44/S2_56_1  ( .CIN(\mult_44/ab[56][1] ), .IN0(
        \mult_44/CARRYB[55][1] ), .IN1(\mult_44/SUMB[55][2] ), .COUT(
        \mult_44/CARRYB[56][1] ), .SUM(\mult_44/SUMB[56][1] ) );
  FADDER \mult_44/S1_56_0  ( .CIN(\mult_44/ab[56][0] ), .IN0(
        \mult_44/CARRYB[55][0] ), .IN1(\mult_44/SUMB[55][1] ), .COUT(
        \mult_44/CARRYB[56][0] ), .SUM(clocal[56]) );
  FADDER \mult_44/S3_57_2  ( .CIN(\mult_44/ab[57][2] ), .IN0(
        \mult_44/CARRYB[56][2] ), .IN1(\mult_44/ab[56][3] ), .COUT(
        \mult_44/CARRYB[57][2] ), .SUM(\mult_44/SUMB[57][2] ) );
  FADDER \mult_44/S2_57_1  ( .CIN(\mult_44/ab[57][1] ), .IN0(
        \mult_44/CARRYB[56][1] ), .IN1(\mult_44/SUMB[56][2] ), .COUT(
        \mult_44/CARRYB[57][1] ), .SUM(\mult_44/SUMB[57][1] ) );
  FADDER \mult_44/S1_57_0  ( .CIN(\mult_44/ab[57][0] ), .IN0(
        \mult_44/CARRYB[56][0] ), .IN1(\mult_44/SUMB[56][1] ), .COUT(
        \mult_44/CARRYB[57][0] ), .SUM(clocal[57]) );
  FADDER \mult_44/S3_58_2  ( .CIN(\mult_44/ab[58][2] ), .IN0(
        \mult_44/CARRYB[57][2] ), .IN1(\mult_44/ab[57][3] ), .COUT(
        \mult_44/CARRYB[58][2] ), .SUM(\mult_44/SUMB[58][2] ) );
  FADDER \mult_44/S2_58_1  ( .CIN(\mult_44/ab[58][1] ), .IN0(
        \mult_44/CARRYB[57][1] ), .IN1(\mult_44/SUMB[57][2] ), .COUT(
        \mult_44/CARRYB[58][1] ), .SUM(\mult_44/SUMB[58][1] ) );
  FADDER \mult_44/S1_58_0  ( .CIN(\mult_44/ab[58][0] ), .IN0(
        \mult_44/CARRYB[57][0] ), .IN1(\mult_44/SUMB[57][1] ), .COUT(
        \mult_44/CARRYB[58][0] ), .SUM(clocal[58]) );
  FADDER \mult_44/S3_59_2  ( .CIN(\mult_44/ab[59][2] ), .IN0(
        \mult_44/CARRYB[58][2] ), .IN1(\mult_44/ab[58][3] ), .COUT(
        \mult_44/CARRYB[59][2] ), .SUM(\mult_44/SUMB[59][2] ) );
  FADDER \mult_44/S2_59_1  ( .CIN(\mult_44/ab[59][1] ), .IN0(
        \mult_44/CARRYB[58][1] ), .IN1(\mult_44/SUMB[58][2] ), .COUT(
        \mult_44/CARRYB[59][1] ), .SUM(\mult_44/SUMB[59][1] ) );
  FADDER \mult_44/S1_59_0  ( .CIN(\mult_44/ab[59][0] ), .IN0(
        \mult_44/CARRYB[58][0] ), .IN1(\mult_44/SUMB[58][1] ), .COUT(
        \mult_44/CARRYB[59][0] ), .SUM(clocal[59]) );
  FADDER \mult_44/S3_60_2  ( .CIN(\mult_44/ab[60][2] ), .IN0(
        \mult_44/CARRYB[59][2] ), .IN1(\mult_44/ab[59][3] ), .COUT(
        \mult_44/CARRYB[60][2] ), .SUM(\mult_44/SUMB[60][2] ) );
  FADDER \mult_44/S2_60_1  ( .CIN(\mult_44/ab[60][1] ), .IN0(
        \mult_44/CARRYB[59][1] ), .IN1(\mult_44/SUMB[59][2] ), .COUT(
        \mult_44/CARRYB[60][1] ), .SUM(\mult_44/SUMB[60][1] ) );
  FADDER \mult_44/S1_60_0  ( .CIN(\mult_44/ab[60][0] ), .IN0(
        \mult_44/CARRYB[59][0] ), .IN1(\mult_44/SUMB[59][1] ), .COUT(
        \mult_44/CARRYB[60][0] ), .SUM(clocal[60]) );
  FADDER \mult_44/S3_61_2  ( .CIN(\mult_44/ab[61][2] ), .IN0(
        \mult_44/CARRYB[60][2] ), .IN1(\mult_44/ab[60][3] ), .COUT(
        \mult_44/CARRYB[61][2] ), .SUM(\mult_44/SUMB[61][2] ) );
  FADDER \mult_44/S2_61_1  ( .CIN(\mult_44/ab[61][1] ), .IN0(
        \mult_44/CARRYB[60][1] ), .IN1(\mult_44/SUMB[60][2] ), .COUT(
        \mult_44/CARRYB[61][1] ), .SUM(\mult_44/SUMB[61][1] ) );
  FADDER \mult_44/S1_61_0  ( .CIN(\mult_44/ab[61][0] ), .IN0(
        \mult_44/CARRYB[60][0] ), .IN1(\mult_44/SUMB[60][1] ), .COUT(
        \mult_44/CARRYB[61][0] ), .SUM(clocal[61]) );
  FADDER \mult_44/S3_62_2  ( .CIN(\mult_44/ab[62][2] ), .IN0(
        \mult_44/CARRYB[61][2] ), .IN1(\mult_44/ab[61][3] ), .COUT(
        \mult_44/CARRYB[62][2] ), .SUM(\mult_44/SUMB[62][2] ) );
  FADDER \mult_44/S2_62_1  ( .CIN(\mult_44/ab[62][1] ), .IN0(
        \mult_44/CARRYB[61][1] ), .IN1(\mult_44/SUMB[61][2] ), .COUT(
        \mult_44/CARRYB[62][1] ), .SUM(\mult_44/SUMB[62][1] ) );
  FADDER \mult_44/S1_62_0  ( .CIN(\mult_44/ab[62][0] ), .IN0(
        \mult_44/CARRYB[61][0] ), .IN1(\mult_44/SUMB[61][1] ), .COUT(
        \mult_44/CARRYB[62][0] ), .SUM(clocal[62]) );
  FADDER \mult_44/S3_63_2  ( .CIN(\mult_44/ab[63][2] ), .IN0(
        \mult_44/CARRYB[62][2] ), .IN1(\mult_44/ab[62][3] ), .COUT(
        \mult_44/CARRYB[63][2] ), .SUM(\mult_44/SUMB[63][2] ) );
  FADDER \mult_44/S2_63_1  ( .CIN(\mult_44/ab[63][1] ), .IN0(
        \mult_44/CARRYB[62][1] ), .IN1(\mult_44/SUMB[62][2] ), .COUT(
        \mult_44/CARRYB[63][1] ), .SUM(\mult_44/SUMB[63][1] ) );
  FADDER \mult_44/S1_63_0  ( .CIN(\mult_44/ab[63][0] ), .IN0(
        \mult_44/CARRYB[62][0] ), .IN1(\mult_44/SUMB[62][1] ), .COUT(
        \mult_44/CARRYB[63][0] ), .SUM(clocal[63]) );
  FADDER \mult_44/S3_64_2  ( .CIN(\mult_44/ab[64][2] ), .IN0(
        \mult_44/CARRYB[63][2] ), .IN1(\mult_44/ab[63][3] ), .COUT(
        \mult_44/CARRYB[64][2] ), .SUM(\mult_44/SUMB[64][2] ) );
  FADDER \mult_44/S2_64_1  ( .CIN(\mult_44/ab[64][1] ), .IN0(
        \mult_44/CARRYB[63][1] ), .IN1(\mult_44/SUMB[63][2] ), .COUT(
        \mult_44/CARRYB[64][1] ), .SUM(\mult_44/SUMB[64][1] ) );
  FADDER \mult_44/S1_64_0  ( .CIN(\mult_44/ab[64][0] ), .IN0(
        \mult_44/CARRYB[63][0] ), .IN1(\mult_44/SUMB[63][1] ), .COUT(
        \mult_44/CARRYB[64][0] ), .SUM(clocal[64]) );
  FADDER \mult_44/S3_65_2  ( .CIN(\mult_44/ab[65][2] ), .IN0(
        \mult_44/CARRYB[64][2] ), .IN1(\mult_44/ab[64][3] ), .COUT(
        \mult_44/CARRYB[65][2] ), .SUM(\mult_44/SUMB[65][2] ) );
  FADDER \mult_44/S2_65_1  ( .CIN(\mult_44/ab[65][1] ), .IN0(
        \mult_44/CARRYB[64][1] ), .IN1(\mult_44/SUMB[64][2] ), .COUT(
        \mult_44/CARRYB[65][1] ), .SUM(\mult_44/SUMB[65][1] ) );
  FADDER \mult_44/S1_65_0  ( .CIN(\mult_44/ab[65][0] ), .IN0(
        \mult_44/CARRYB[64][0] ), .IN1(\mult_44/SUMB[64][1] ), .COUT(
        \mult_44/CARRYB[65][0] ), .SUM(clocal[65]) );
  FADDER \mult_44/S3_66_2  ( .CIN(\mult_44/ab[66][2] ), .IN0(
        \mult_44/CARRYB[65][2] ), .IN1(\mult_44/ab[65][3] ), .COUT(
        \mult_44/CARRYB[66][2] ), .SUM(\mult_44/SUMB[66][2] ) );
  FADDER \mult_44/S2_66_1  ( .CIN(\mult_44/ab[66][1] ), .IN0(
        \mult_44/CARRYB[65][1] ), .IN1(\mult_44/SUMB[65][2] ), .COUT(
        \mult_44/CARRYB[66][1] ), .SUM(\mult_44/SUMB[66][1] ) );
  FADDER \mult_44/S1_66_0  ( .CIN(\mult_44/ab[66][0] ), .IN0(
        \mult_44/CARRYB[65][0] ), .IN1(\mult_44/SUMB[65][1] ), .COUT(
        \mult_44/CARRYB[66][0] ), .SUM(clocal[66]) );
  FADDER \mult_44/S3_67_2  ( .CIN(\mult_44/ab[67][2] ), .IN0(
        \mult_44/CARRYB[66][2] ), .IN1(\mult_44/ab[66][3] ), .COUT(
        \mult_44/CARRYB[67][2] ), .SUM(\mult_44/SUMB[67][2] ) );
  FADDER \mult_44/S2_67_1  ( .CIN(\mult_44/ab[67][1] ), .IN0(
        \mult_44/CARRYB[66][1] ), .IN1(\mult_44/SUMB[66][2] ), .COUT(
        \mult_44/CARRYB[67][1] ), .SUM(\mult_44/SUMB[67][1] ) );
  FADDER \mult_44/S1_67_0  ( .CIN(\mult_44/ab[67][0] ), .IN0(
        \mult_44/CARRYB[66][0] ), .IN1(\mult_44/SUMB[66][1] ), .COUT(
        \mult_44/CARRYB[67][0] ), .SUM(clocal[67]) );
  FADDER \mult_44/S3_68_2  ( .CIN(\mult_44/ab[68][2] ), .IN0(
        \mult_44/CARRYB[67][2] ), .IN1(\mult_44/ab[67][3] ), .COUT(
        \mult_44/CARRYB[68][2] ), .SUM(\mult_44/SUMB[68][2] ) );
  FADDER \mult_44/S2_68_1  ( .CIN(\mult_44/ab[68][1] ), .IN0(
        \mult_44/CARRYB[67][1] ), .IN1(\mult_44/SUMB[67][2] ), .COUT(
        \mult_44/CARRYB[68][1] ), .SUM(\mult_44/SUMB[68][1] ) );
  FADDER \mult_44/S1_68_0  ( .CIN(\mult_44/ab[68][0] ), .IN0(
        \mult_44/CARRYB[67][0] ), .IN1(\mult_44/SUMB[67][1] ), .COUT(
        \mult_44/CARRYB[68][0] ), .SUM(clocal[68]) );
  FADDER \mult_44/S3_69_2  ( .CIN(\mult_44/ab[69][2] ), .IN0(
        \mult_44/CARRYB[68][2] ), .IN1(\mult_44/ab[68][3] ), .COUT(
        \mult_44/CARRYB[69][2] ), .SUM(\mult_44/SUMB[69][2] ) );
  FADDER \mult_44/S2_69_1  ( .CIN(\mult_44/ab[69][1] ), .IN0(
        \mult_44/CARRYB[68][1] ), .IN1(\mult_44/SUMB[68][2] ), .COUT(
        \mult_44/CARRYB[69][1] ), .SUM(\mult_44/SUMB[69][1] ) );
  FADDER \mult_44/S1_69_0  ( .CIN(\mult_44/ab[69][0] ), .IN0(
        \mult_44/CARRYB[68][0] ), .IN1(\mult_44/SUMB[68][1] ), .COUT(
        \mult_44/CARRYB[69][0] ), .SUM(clocal[69]) );
  FADDER \mult_44/S3_70_2  ( .CIN(\mult_44/ab[70][2] ), .IN0(
        \mult_44/CARRYB[69][2] ), .IN1(\mult_44/ab[69][3] ), .COUT(
        \mult_44/CARRYB[70][2] ), .SUM(\mult_44/SUMB[70][2] ) );
  FADDER \mult_44/S2_70_1  ( .CIN(\mult_44/ab[70][1] ), .IN0(
        \mult_44/CARRYB[69][1] ), .IN1(\mult_44/SUMB[69][2] ), .COUT(
        \mult_44/CARRYB[70][1] ), .SUM(\mult_44/SUMB[70][1] ) );
  FADDER \mult_44/S1_70_0  ( .CIN(\mult_44/ab[70][0] ), .IN0(
        \mult_44/CARRYB[69][0] ), .IN1(\mult_44/SUMB[69][1] ), .COUT(
        \mult_44/CARRYB[70][0] ), .SUM(clocal[70]) );
  FADDER \mult_44/S3_71_2  ( .CIN(\mult_44/ab[71][2] ), .IN0(
        \mult_44/CARRYB[70][2] ), .IN1(\mult_44/ab[70][3] ), .COUT(
        \mult_44/CARRYB[71][2] ), .SUM(\mult_44/SUMB[71][2] ) );
  FADDER \mult_44/S2_71_1  ( .CIN(\mult_44/ab[71][1] ), .IN0(
        \mult_44/CARRYB[70][1] ), .IN1(\mult_44/SUMB[70][2] ), .COUT(
        \mult_44/CARRYB[71][1] ), .SUM(\mult_44/SUMB[71][1] ) );
  FADDER \mult_44/S1_71_0  ( .CIN(\mult_44/ab[71][0] ), .IN0(
        \mult_44/CARRYB[70][0] ), .IN1(\mult_44/SUMB[70][1] ), .COUT(
        \mult_44/CARRYB[71][0] ), .SUM(clocal[71]) );
  FADDER \mult_44/S3_72_2  ( .CIN(\mult_44/ab[72][2] ), .IN0(
        \mult_44/CARRYB[71][2] ), .IN1(\mult_44/ab[71][3] ), .COUT(
        \mult_44/CARRYB[72][2] ), .SUM(\mult_44/SUMB[72][2] ) );
  FADDER \mult_44/S2_72_1  ( .CIN(\mult_44/ab[72][1] ), .IN0(
        \mult_44/CARRYB[71][1] ), .IN1(\mult_44/SUMB[71][2] ), .COUT(
        \mult_44/CARRYB[72][1] ), .SUM(\mult_44/SUMB[72][1] ) );
  FADDER \mult_44/S1_72_0  ( .CIN(\mult_44/ab[72][0] ), .IN0(
        \mult_44/CARRYB[71][0] ), .IN1(\mult_44/SUMB[71][1] ), .COUT(
        \mult_44/CARRYB[72][0] ), .SUM(clocal[72]) );
  FADDER \mult_44/S3_73_2  ( .CIN(\mult_44/ab[73][2] ), .IN0(
        \mult_44/CARRYB[72][2] ), .IN1(\mult_44/ab[72][3] ), .COUT(
        \mult_44/CARRYB[73][2] ), .SUM(\mult_44/SUMB[73][2] ) );
  FADDER \mult_44/S2_73_1  ( .CIN(\mult_44/ab[73][1] ), .IN0(
        \mult_44/CARRYB[72][1] ), .IN1(\mult_44/SUMB[72][2] ), .COUT(
        \mult_44/CARRYB[73][1] ), .SUM(\mult_44/SUMB[73][1] ) );
  FADDER \mult_44/S1_73_0  ( .CIN(\mult_44/ab[73][0] ), .IN0(
        \mult_44/CARRYB[72][0] ), .IN1(\mult_44/SUMB[72][1] ), .COUT(
        \mult_44/CARRYB[73][0] ), .SUM(clocal[73]) );
  FADDER \mult_44/S3_74_2  ( .CIN(\mult_44/ab[74][2] ), .IN0(
        \mult_44/CARRYB[73][2] ), .IN1(\mult_44/ab[73][3] ), .COUT(
        \mult_44/CARRYB[74][2] ), .SUM(\mult_44/SUMB[74][2] ) );
  FADDER \mult_44/S2_74_1  ( .CIN(\mult_44/ab[74][1] ), .IN0(
        \mult_44/CARRYB[73][1] ), .IN1(\mult_44/SUMB[73][2] ), .COUT(
        \mult_44/CARRYB[74][1] ), .SUM(\mult_44/SUMB[74][1] ) );
  FADDER \mult_44/S1_74_0  ( .CIN(\mult_44/ab[74][0] ), .IN0(
        \mult_44/CARRYB[73][0] ), .IN1(\mult_44/SUMB[73][1] ), .COUT(
        \mult_44/CARRYB[74][0] ), .SUM(clocal[74]) );
  FADDER \mult_44/S3_75_2  ( .CIN(\mult_44/ab[75][2] ), .IN0(
        \mult_44/CARRYB[74][2] ), .IN1(\mult_44/ab[74][3] ), .COUT(
        \mult_44/CARRYB[75][2] ), .SUM(\mult_44/SUMB[75][2] ) );
  FADDER \mult_44/S2_75_1  ( .CIN(\mult_44/ab[75][1] ), .IN0(
        \mult_44/CARRYB[74][1] ), .IN1(\mult_44/SUMB[74][2] ), .COUT(
        \mult_44/CARRYB[75][1] ), .SUM(\mult_44/SUMB[75][1] ) );
  FADDER \mult_44/S1_75_0  ( .CIN(\mult_44/ab[75][0] ), .IN0(
        \mult_44/CARRYB[74][0] ), .IN1(\mult_44/SUMB[74][1] ), .COUT(
        \mult_44/CARRYB[75][0] ), .SUM(clocal[75]) );
  FADDER \mult_44/S3_76_2  ( .CIN(\mult_44/ab[76][2] ), .IN0(
        \mult_44/CARRYB[75][2] ), .IN1(\mult_44/ab[75][3] ), .COUT(
        \mult_44/CARRYB[76][2] ), .SUM(\mult_44/SUMB[76][2] ) );
  FADDER \mult_44/S2_76_1  ( .CIN(\mult_44/ab[76][1] ), .IN0(
        \mult_44/CARRYB[75][1] ), .IN1(\mult_44/SUMB[75][2] ), .COUT(
        \mult_44/CARRYB[76][1] ), .SUM(\mult_44/SUMB[76][1] ) );
  FADDER \mult_44/S1_76_0  ( .CIN(\mult_44/ab[76][0] ), .IN0(
        \mult_44/CARRYB[75][0] ), .IN1(\mult_44/SUMB[75][1] ), .COUT(
        \mult_44/CARRYB[76][0] ), .SUM(clocal[76]) );
  FADDER \mult_44/S3_77_2  ( .CIN(\mult_44/ab[77][2] ), .IN0(
        \mult_44/CARRYB[76][2] ), .IN1(\mult_44/ab[76][3] ), .COUT(
        \mult_44/CARRYB[77][2] ), .SUM(\mult_44/SUMB[77][2] ) );
  FADDER \mult_44/S2_77_1  ( .CIN(\mult_44/ab[77][1] ), .IN0(
        \mult_44/CARRYB[76][1] ), .IN1(\mult_44/SUMB[76][2] ), .COUT(
        \mult_44/CARRYB[77][1] ), .SUM(\mult_44/SUMB[77][1] ) );
  FADDER \mult_44/S1_77_0  ( .CIN(\mult_44/ab[77][0] ), .IN0(
        \mult_44/CARRYB[76][0] ), .IN1(\mult_44/SUMB[76][1] ), .COUT(
        \mult_44/CARRYB[77][0] ), .SUM(clocal[77]) );
  FADDER \mult_44/S3_78_2  ( .CIN(\mult_44/ab[78][2] ), .IN0(
        \mult_44/CARRYB[77][2] ), .IN1(\mult_44/ab[77][3] ), .COUT(
        \mult_44/CARRYB[78][2] ), .SUM(\mult_44/SUMB[78][2] ) );
  FADDER \mult_44/S2_78_1  ( .CIN(\mult_44/ab[78][1] ), .IN0(
        \mult_44/CARRYB[77][1] ), .IN1(\mult_44/SUMB[77][2] ), .COUT(
        \mult_44/CARRYB[78][1] ), .SUM(\mult_44/SUMB[78][1] ) );
  FADDER \mult_44/S1_78_0  ( .CIN(\mult_44/ab[78][0] ), .IN0(
        \mult_44/CARRYB[77][0] ), .IN1(\mult_44/SUMB[77][1] ), .COUT(
        \mult_44/CARRYB[78][0] ), .SUM(clocal[78]) );
  FADDER \mult_44/S3_79_2  ( .CIN(\mult_44/ab[79][2] ), .IN0(
        \mult_44/CARRYB[78][2] ), .IN1(\mult_44/ab[78][3] ), .COUT(
        \mult_44/CARRYB[79][2] ), .SUM(\mult_44/SUMB[79][2] ) );
  FADDER \mult_44/S2_79_1  ( .CIN(\mult_44/ab[79][1] ), .IN0(
        \mult_44/CARRYB[78][1] ), .IN1(\mult_44/SUMB[78][2] ), .COUT(
        \mult_44/CARRYB[79][1] ), .SUM(\mult_44/SUMB[79][1] ) );
  FADDER \mult_44/S1_79_0  ( .CIN(\mult_44/ab[79][0] ), .IN0(
        \mult_44/CARRYB[78][0] ), .IN1(\mult_44/SUMB[78][1] ), .COUT(
        \mult_44/CARRYB[79][0] ), .SUM(clocal[79]) );
  FADDER \mult_44/S3_80_2  ( .CIN(\mult_44/ab[80][2] ), .IN0(
        \mult_44/CARRYB[79][2] ), .IN1(\mult_44/ab[79][3] ), .COUT(
        \mult_44/CARRYB[80][2] ), .SUM(\mult_44/SUMB[80][2] ) );
  FADDER \mult_44/S2_80_1  ( .CIN(\mult_44/ab[80][1] ), .IN0(
        \mult_44/CARRYB[79][1] ), .IN1(\mult_44/SUMB[79][2] ), .COUT(
        \mult_44/CARRYB[80][1] ), .SUM(\mult_44/SUMB[80][1] ) );
  FADDER \mult_44/S1_80_0  ( .CIN(\mult_44/ab[80][0] ), .IN0(
        \mult_44/CARRYB[79][0] ), .IN1(\mult_44/SUMB[79][1] ), .COUT(
        \mult_44/CARRYB[80][0] ), .SUM(clocal[80]) );
  FADDER \mult_44/S3_81_2  ( .CIN(\mult_44/ab[81][2] ), .IN0(
        \mult_44/CARRYB[80][2] ), .IN1(\mult_44/ab[80][3] ), .COUT(
        \mult_44/CARRYB[81][2] ), .SUM(\mult_44/SUMB[81][2] ) );
  FADDER \mult_44/S2_81_1  ( .CIN(\mult_44/ab[81][1] ), .IN0(
        \mult_44/CARRYB[80][1] ), .IN1(\mult_44/SUMB[80][2] ), .COUT(
        \mult_44/CARRYB[81][1] ), .SUM(\mult_44/SUMB[81][1] ) );
  FADDER \mult_44/S1_81_0  ( .CIN(\mult_44/ab[81][0] ), .IN0(
        \mult_44/CARRYB[80][0] ), .IN1(\mult_44/SUMB[80][1] ), .COUT(
        \mult_44/CARRYB[81][0] ), .SUM(clocal[81]) );
  FADDER \mult_44/S3_82_2  ( .CIN(\mult_44/ab[82][2] ), .IN0(
        \mult_44/CARRYB[81][2] ), .IN1(\mult_44/ab[81][3] ), .COUT(
        \mult_44/CARRYB[82][2] ), .SUM(\mult_44/SUMB[82][2] ) );
  FADDER \mult_44/S2_82_1  ( .CIN(\mult_44/ab[82][1] ), .IN0(
        \mult_44/CARRYB[81][1] ), .IN1(\mult_44/SUMB[81][2] ), .COUT(
        \mult_44/CARRYB[82][1] ), .SUM(\mult_44/SUMB[82][1] ) );
  FADDER \mult_44/S1_82_0  ( .CIN(\mult_44/ab[82][0] ), .IN0(
        \mult_44/CARRYB[81][0] ), .IN1(\mult_44/SUMB[81][1] ), .COUT(
        \mult_44/CARRYB[82][0] ), .SUM(clocal[82]) );
  FADDER \mult_44/S3_83_2  ( .CIN(\mult_44/ab[83][2] ), .IN0(
        \mult_44/CARRYB[82][2] ), .IN1(\mult_44/ab[82][3] ), .COUT(
        \mult_44/CARRYB[83][2] ), .SUM(\mult_44/SUMB[83][2] ) );
  FADDER \mult_44/S2_83_1  ( .CIN(\mult_44/ab[83][1] ), .IN0(
        \mult_44/CARRYB[82][1] ), .IN1(\mult_44/SUMB[82][2] ), .COUT(
        \mult_44/CARRYB[83][1] ), .SUM(\mult_44/SUMB[83][1] ) );
  FADDER \mult_44/S1_83_0  ( .CIN(\mult_44/ab[83][0] ), .IN0(
        \mult_44/CARRYB[82][0] ), .IN1(\mult_44/SUMB[82][1] ), .COUT(
        \mult_44/CARRYB[83][0] ), .SUM(clocal[83]) );
  FADDER \mult_44/S3_84_2  ( .CIN(\mult_44/ab[84][2] ), .IN0(
        \mult_44/CARRYB[83][2] ), .IN1(\mult_44/ab[83][3] ), .COUT(
        \mult_44/CARRYB[84][2] ), .SUM(\mult_44/SUMB[84][2] ) );
  FADDER \mult_44/S2_84_1  ( .CIN(\mult_44/ab[84][1] ), .IN0(
        \mult_44/CARRYB[83][1] ), .IN1(\mult_44/SUMB[83][2] ), .COUT(
        \mult_44/CARRYB[84][1] ), .SUM(\mult_44/SUMB[84][1] ) );
  FADDER \mult_44/S1_84_0  ( .CIN(\mult_44/ab[84][0] ), .IN0(
        \mult_44/CARRYB[83][0] ), .IN1(\mult_44/SUMB[83][1] ), .COUT(
        \mult_44/CARRYB[84][0] ), .SUM(clocal[84]) );
  FADDER \mult_44/S3_85_2  ( .CIN(\mult_44/ab[85][2] ), .IN0(
        \mult_44/CARRYB[84][2] ), .IN1(\mult_44/ab[84][3] ), .COUT(
        \mult_44/CARRYB[85][2] ), .SUM(\mult_44/SUMB[85][2] ) );
  FADDER \mult_44/S2_85_1  ( .CIN(\mult_44/ab[85][1] ), .IN0(
        \mult_44/CARRYB[84][1] ), .IN1(\mult_44/SUMB[84][2] ), .COUT(
        \mult_44/CARRYB[85][1] ), .SUM(\mult_44/SUMB[85][1] ) );
  FADDER \mult_44/S1_85_0  ( .CIN(\mult_44/ab[85][0] ), .IN0(
        \mult_44/CARRYB[84][0] ), .IN1(\mult_44/SUMB[84][1] ), .COUT(
        \mult_44/CARRYB[85][0] ), .SUM(clocal[85]) );
  FADDER \mult_44/S3_86_2  ( .CIN(\mult_44/ab[86][2] ), .IN0(
        \mult_44/CARRYB[85][2] ), .IN1(\mult_44/ab[85][3] ), .COUT(
        \mult_44/CARRYB[86][2] ), .SUM(\mult_44/SUMB[86][2] ) );
  FADDER \mult_44/S2_86_1  ( .CIN(\mult_44/ab[86][1] ), .IN0(
        \mult_44/CARRYB[85][1] ), .IN1(\mult_44/SUMB[85][2] ), .COUT(
        \mult_44/CARRYB[86][1] ), .SUM(\mult_44/SUMB[86][1] ) );
  FADDER \mult_44/S1_86_0  ( .CIN(\mult_44/ab[86][0] ), .IN0(
        \mult_44/CARRYB[85][0] ), .IN1(\mult_44/SUMB[85][1] ), .COUT(
        \mult_44/CARRYB[86][0] ), .SUM(clocal[86]) );
  FADDER \mult_44/S3_87_2  ( .CIN(\mult_44/ab[87][2] ), .IN0(
        \mult_44/CARRYB[86][2] ), .IN1(\mult_44/ab[86][3] ), .COUT(
        \mult_44/CARRYB[87][2] ), .SUM(\mult_44/SUMB[87][2] ) );
  FADDER \mult_44/S2_87_1  ( .CIN(\mult_44/ab[87][1] ), .IN0(
        \mult_44/CARRYB[86][1] ), .IN1(\mult_44/SUMB[86][2] ), .COUT(
        \mult_44/CARRYB[87][1] ), .SUM(\mult_44/SUMB[87][1] ) );
  FADDER \mult_44/S1_87_0  ( .CIN(\mult_44/ab[87][0] ), .IN0(
        \mult_44/CARRYB[86][0] ), .IN1(\mult_44/SUMB[86][1] ), .COUT(
        \mult_44/CARRYB[87][0] ), .SUM(clocal[87]) );
  FADDER \mult_44/S3_88_2  ( .CIN(\mult_44/ab[88][2] ), .IN0(
        \mult_44/CARRYB[87][2] ), .IN1(\mult_44/ab[87][3] ), .COUT(
        \mult_44/CARRYB[88][2] ), .SUM(\mult_44/SUMB[88][2] ) );
  FADDER \mult_44/S2_88_1  ( .CIN(\mult_44/ab[88][1] ), .IN0(
        \mult_44/CARRYB[87][1] ), .IN1(\mult_44/SUMB[87][2] ), .COUT(
        \mult_44/CARRYB[88][1] ), .SUM(\mult_44/SUMB[88][1] ) );
  FADDER \mult_44/S1_88_0  ( .CIN(\mult_44/ab[88][0] ), .IN0(
        \mult_44/CARRYB[87][0] ), .IN1(\mult_44/SUMB[87][1] ), .COUT(
        \mult_44/CARRYB[88][0] ), .SUM(clocal[88]) );
  FADDER \mult_44/S3_89_2  ( .CIN(\mult_44/ab[89][2] ), .IN0(
        \mult_44/CARRYB[88][2] ), .IN1(\mult_44/ab[88][3] ), .COUT(
        \mult_44/CARRYB[89][2] ), .SUM(\mult_44/SUMB[89][2] ) );
  FADDER \mult_44/S2_89_1  ( .CIN(\mult_44/ab[89][1] ), .IN0(
        \mult_44/CARRYB[88][1] ), .IN1(\mult_44/SUMB[88][2] ), .COUT(
        \mult_44/CARRYB[89][1] ), .SUM(\mult_44/SUMB[89][1] ) );
  FADDER \mult_44/S1_89_0  ( .CIN(\mult_44/ab[89][0] ), .IN0(
        \mult_44/CARRYB[88][0] ), .IN1(\mult_44/SUMB[88][1] ), .COUT(
        \mult_44/CARRYB[89][0] ), .SUM(clocal[89]) );
  FADDER \mult_44/S3_90_2  ( .CIN(\mult_44/ab[90][2] ), .IN0(
        \mult_44/CARRYB[89][2] ), .IN1(\mult_44/ab[89][3] ), .COUT(
        \mult_44/CARRYB[90][2] ), .SUM(\mult_44/SUMB[90][2] ) );
  FADDER \mult_44/S2_90_1  ( .CIN(\mult_44/ab[90][1] ), .IN0(
        \mult_44/CARRYB[89][1] ), .IN1(\mult_44/SUMB[89][2] ), .COUT(
        \mult_44/CARRYB[90][1] ), .SUM(\mult_44/SUMB[90][1] ) );
  FADDER \mult_44/S1_90_0  ( .CIN(\mult_44/ab[90][0] ), .IN0(
        \mult_44/CARRYB[89][0] ), .IN1(\mult_44/SUMB[89][1] ), .COUT(
        \mult_44/CARRYB[90][0] ), .SUM(clocal[90]) );
  FADDER \mult_44/S3_91_2  ( .CIN(\mult_44/ab[91][2] ), .IN0(
        \mult_44/CARRYB[90][2] ), .IN1(\mult_44/ab[90][3] ), .COUT(
        \mult_44/CARRYB[91][2] ), .SUM(\mult_44/SUMB[91][2] ) );
  FADDER \mult_44/S2_91_1  ( .CIN(\mult_44/ab[91][1] ), .IN0(
        \mult_44/CARRYB[90][1] ), .IN1(\mult_44/SUMB[90][2] ), .COUT(
        \mult_44/CARRYB[91][1] ), .SUM(\mult_44/SUMB[91][1] ) );
  FADDER \mult_44/S1_91_0  ( .CIN(\mult_44/ab[91][0] ), .IN0(
        \mult_44/CARRYB[90][0] ), .IN1(\mult_44/SUMB[90][1] ), .COUT(
        \mult_44/CARRYB[91][0] ), .SUM(clocal[91]) );
  FADDER \mult_44/S3_92_2  ( .CIN(\mult_44/ab[92][2] ), .IN0(
        \mult_44/CARRYB[91][2] ), .IN1(\mult_44/ab[91][3] ), .COUT(
        \mult_44/CARRYB[92][2] ), .SUM(\mult_44/SUMB[92][2] ) );
  FADDER \mult_44/S2_92_1  ( .CIN(\mult_44/ab[92][1] ), .IN0(
        \mult_44/CARRYB[91][1] ), .IN1(\mult_44/SUMB[91][2] ), .COUT(
        \mult_44/CARRYB[92][1] ), .SUM(\mult_44/SUMB[92][1] ) );
  FADDER \mult_44/S1_92_0  ( .CIN(\mult_44/ab[92][0] ), .IN0(
        \mult_44/CARRYB[91][0] ), .IN1(\mult_44/SUMB[91][1] ), .COUT(
        \mult_44/CARRYB[92][0] ), .SUM(clocal[92]) );
  FADDER \mult_44/S3_93_2  ( .CIN(\mult_44/ab[93][2] ), .IN0(
        \mult_44/CARRYB[92][2] ), .IN1(\mult_44/ab[92][3] ), .COUT(
        \mult_44/CARRYB[93][2] ), .SUM(\mult_44/SUMB[93][2] ) );
  FADDER \mult_44/S2_93_1  ( .CIN(\mult_44/ab[93][1] ), .IN0(
        \mult_44/CARRYB[92][1] ), .IN1(\mult_44/SUMB[92][2] ), .COUT(
        \mult_44/CARRYB[93][1] ), .SUM(\mult_44/SUMB[93][1] ) );
  FADDER \mult_44/S1_93_0  ( .CIN(\mult_44/ab[93][0] ), .IN0(
        \mult_44/CARRYB[92][0] ), .IN1(\mult_44/SUMB[92][1] ), .COUT(
        \mult_44/CARRYB[93][0] ), .SUM(clocal[93]) );
  FADDER \mult_44/S3_94_2  ( .CIN(\mult_44/ab[94][2] ), .IN0(
        \mult_44/CARRYB[93][2] ), .IN1(\mult_44/ab[93][3] ), .COUT(
        \mult_44/CARRYB[94][2] ), .SUM(\mult_44/SUMB[94][2] ) );
  FADDER \mult_44/S2_94_1  ( .CIN(\mult_44/ab[94][1] ), .IN0(
        \mult_44/CARRYB[93][1] ), .IN1(\mult_44/SUMB[93][2] ), .COUT(
        \mult_44/CARRYB[94][1] ), .SUM(\mult_44/SUMB[94][1] ) );
  FADDER \mult_44/S1_94_0  ( .CIN(\mult_44/ab[94][0] ), .IN0(
        \mult_44/CARRYB[93][0] ), .IN1(\mult_44/SUMB[93][1] ), .COUT(
        \mult_44/CARRYB[94][0] ), .SUM(clocal[94]) );
  FADDER \mult_44/S3_95_2  ( .CIN(\mult_44/ab[95][2] ), .IN0(
        \mult_44/CARRYB[94][2] ), .IN1(\mult_44/ab[94][3] ), .COUT(
        \mult_44/CARRYB[95][2] ), .SUM(\mult_44/SUMB[95][2] ) );
  FADDER \mult_44/S2_95_1  ( .CIN(\mult_44/ab[95][1] ), .IN0(
        \mult_44/CARRYB[94][1] ), .IN1(\mult_44/SUMB[94][2] ), .COUT(
        \mult_44/CARRYB[95][1] ), .SUM(\mult_44/SUMB[95][1] ) );
  FADDER \mult_44/S1_95_0  ( .CIN(\mult_44/ab[95][0] ), .IN0(
        \mult_44/CARRYB[94][0] ), .IN1(\mult_44/SUMB[94][1] ), .COUT(
        \mult_44/CARRYB[95][0] ), .SUM(clocal[95]) );
  FADDER \mult_44/S3_96_2  ( .CIN(\mult_44/ab[96][2] ), .IN0(
        \mult_44/CARRYB[95][2] ), .IN1(\mult_44/ab[95][3] ), .COUT(
        \mult_44/CARRYB[96][2] ), .SUM(\mult_44/SUMB[96][2] ) );
  FADDER \mult_44/S2_96_1  ( .CIN(\mult_44/ab[96][1] ), .IN0(
        \mult_44/CARRYB[95][1] ), .IN1(\mult_44/SUMB[95][2] ), .COUT(
        \mult_44/CARRYB[96][1] ), .SUM(\mult_44/SUMB[96][1] ) );
  FADDER \mult_44/S1_96_0  ( .CIN(\mult_44/ab[96][0] ), .IN0(
        \mult_44/CARRYB[95][0] ), .IN1(\mult_44/SUMB[95][1] ), .COUT(
        \mult_44/CARRYB[96][0] ), .SUM(clocal[96]) );
  FADDER \mult_44/S3_97_2  ( .CIN(\mult_44/ab[97][2] ), .IN0(
        \mult_44/CARRYB[96][2] ), .IN1(\mult_44/ab[96][3] ), .COUT(
        \mult_44/CARRYB[97][2] ), .SUM(\mult_44/SUMB[97][2] ) );
  FADDER \mult_44/S2_97_1  ( .CIN(\mult_44/ab[97][1] ), .IN0(
        \mult_44/CARRYB[96][1] ), .IN1(\mult_44/SUMB[96][2] ), .COUT(
        \mult_44/CARRYB[97][1] ), .SUM(\mult_44/SUMB[97][1] ) );
  FADDER \mult_44/S1_97_0  ( .CIN(\mult_44/ab[97][0] ), .IN0(
        \mult_44/CARRYB[96][0] ), .IN1(\mult_44/SUMB[96][1] ), .COUT(
        \mult_44/CARRYB[97][0] ), .SUM(clocal[97]) );
  FADDER \mult_44/S3_98_2  ( .CIN(\mult_44/ab[98][2] ), .IN0(
        \mult_44/CARRYB[97][2] ), .IN1(\mult_44/ab[97][3] ), .COUT(
        \mult_44/CARRYB[98][2] ), .SUM(\mult_44/SUMB[98][2] ) );
  FADDER \mult_44/S2_98_1  ( .CIN(\mult_44/ab[98][1] ), .IN0(
        \mult_44/CARRYB[97][1] ), .IN1(\mult_44/SUMB[97][2] ), .COUT(
        \mult_44/CARRYB[98][1] ), .SUM(\mult_44/SUMB[98][1] ) );
  FADDER \mult_44/S1_98_0  ( .CIN(\mult_44/ab[98][0] ), .IN0(
        \mult_44/CARRYB[97][0] ), .IN1(\mult_44/SUMB[97][1] ), .COUT(
        \mult_44/CARRYB[98][0] ), .SUM(clocal[98]) );
  FADDER \mult_44/S3_99_2  ( .CIN(\mult_44/ab[99][2] ), .IN0(
        \mult_44/CARRYB[98][2] ), .IN1(\mult_44/ab[98][3] ), .COUT(
        \mult_44/CARRYB[99][2] ), .SUM(\mult_44/SUMB[99][2] ) );
  FADDER \mult_44/S2_99_1  ( .CIN(\mult_44/ab[99][1] ), .IN0(
        \mult_44/CARRYB[98][1] ), .IN1(\mult_44/SUMB[98][2] ), .COUT(
        \mult_44/CARRYB[99][1] ), .SUM(\mult_44/SUMB[99][1] ) );
  FADDER \mult_44/S1_99_0  ( .CIN(\mult_44/ab[99][0] ), .IN0(
        \mult_44/CARRYB[98][0] ), .IN1(\mult_44/SUMB[98][1] ), .COUT(
        \mult_44/CARRYB[99][0] ), .SUM(clocal[99]) );
  FADDER \mult_44/S3_100_2  ( .CIN(\mult_44/ab[100][2] ), .IN0(
        \mult_44/CARRYB[99][2] ), .IN1(\mult_44/ab[99][3] ), .COUT(
        \mult_44/CARRYB[100][2] ), .SUM(\mult_44/SUMB[100][2] ) );
  FADDER \mult_44/S2_100_1  ( .CIN(\mult_44/ab[100][1] ), .IN0(
        \mult_44/CARRYB[99][1] ), .IN1(\mult_44/SUMB[99][2] ), .COUT(
        \mult_44/CARRYB[100][1] ), .SUM(\mult_44/SUMB[100][1] ) );
  FADDER \mult_44/S1_100_0  ( .CIN(\mult_44/ab[100][0] ), .IN0(
        \mult_44/CARRYB[99][0] ), .IN1(\mult_44/SUMB[99][1] ), .COUT(
        \mult_44/CARRYB[100][0] ), .SUM(clocal[100]) );
  FADDER \mult_44/S3_101_2  ( .CIN(\mult_44/ab[101][2] ), .IN0(
        \mult_44/CARRYB[100][2] ), .IN1(\mult_44/ab[100][3] ), .COUT(
        \mult_44/CARRYB[101][2] ), .SUM(\mult_44/SUMB[101][2] ) );
  FADDER \mult_44/S2_101_1  ( .CIN(\mult_44/ab[101][1] ), .IN0(
        \mult_44/CARRYB[100][1] ), .IN1(\mult_44/SUMB[100][2] ), .COUT(
        \mult_44/CARRYB[101][1] ), .SUM(\mult_44/SUMB[101][1] ) );
  FADDER \mult_44/S1_101_0  ( .CIN(\mult_44/ab[101][0] ), .IN0(
        \mult_44/CARRYB[100][0] ), .IN1(\mult_44/SUMB[100][1] ), .COUT(
        \mult_44/CARRYB[101][0] ), .SUM(clocal[101]) );
  FADDER \mult_44/S3_102_2  ( .CIN(\mult_44/ab[102][2] ), .IN0(
        \mult_44/CARRYB[101][2] ), .IN1(\mult_44/ab[101][3] ), .COUT(
        \mult_44/CARRYB[102][2] ), .SUM(\mult_44/SUMB[102][2] ) );
  FADDER \mult_44/S2_102_1  ( .CIN(\mult_44/ab[102][1] ), .IN0(
        \mult_44/CARRYB[101][1] ), .IN1(\mult_44/SUMB[101][2] ), .COUT(
        \mult_44/CARRYB[102][1] ), .SUM(\mult_44/SUMB[102][1] ) );
  FADDER \mult_44/S1_102_0  ( .CIN(\mult_44/ab[102][0] ), .IN0(
        \mult_44/CARRYB[101][0] ), .IN1(\mult_44/SUMB[101][1] ), .COUT(
        \mult_44/CARRYB[102][0] ), .SUM(clocal[102]) );
  FADDER \mult_44/S3_103_2  ( .CIN(\mult_44/ab[103][2] ), .IN0(
        \mult_44/CARRYB[102][2] ), .IN1(\mult_44/ab[102][3] ), .COUT(
        \mult_44/CARRYB[103][2] ), .SUM(\mult_44/SUMB[103][2] ) );
  FADDER \mult_44/S2_103_1  ( .CIN(\mult_44/ab[103][1] ), .IN0(
        \mult_44/CARRYB[102][1] ), .IN1(\mult_44/SUMB[102][2] ), .COUT(
        \mult_44/CARRYB[103][1] ), .SUM(\mult_44/SUMB[103][1] ) );
  FADDER \mult_44/S1_103_0  ( .CIN(\mult_44/ab[103][0] ), .IN0(
        \mult_44/CARRYB[102][0] ), .IN1(\mult_44/SUMB[102][1] ), .COUT(
        \mult_44/CARRYB[103][0] ), .SUM(clocal[103]) );
  FADDER \mult_44/S3_104_2  ( .CIN(\mult_44/ab[104][2] ), .IN0(
        \mult_44/CARRYB[103][2] ), .IN1(\mult_44/ab[103][3] ), .COUT(
        \mult_44/CARRYB[104][2] ), .SUM(\mult_44/SUMB[104][2] ) );
  FADDER \mult_44/S2_104_1  ( .CIN(\mult_44/ab[104][1] ), .IN0(
        \mult_44/CARRYB[103][1] ), .IN1(\mult_44/SUMB[103][2] ), .COUT(
        \mult_44/CARRYB[104][1] ), .SUM(\mult_44/SUMB[104][1] ) );
  FADDER \mult_44/S1_104_0  ( .CIN(\mult_44/ab[104][0] ), .IN0(
        \mult_44/CARRYB[103][0] ), .IN1(\mult_44/SUMB[103][1] ), .COUT(
        \mult_44/CARRYB[104][0] ), .SUM(clocal[104]) );
  FADDER \mult_44/S3_105_2  ( .CIN(\mult_44/ab[105][2] ), .IN0(
        \mult_44/CARRYB[104][2] ), .IN1(\mult_44/ab[104][3] ), .COUT(
        \mult_44/CARRYB[105][2] ), .SUM(\mult_44/SUMB[105][2] ) );
  FADDER \mult_44/S2_105_1  ( .CIN(\mult_44/ab[105][1] ), .IN0(
        \mult_44/CARRYB[104][1] ), .IN1(\mult_44/SUMB[104][2] ), .COUT(
        \mult_44/CARRYB[105][1] ), .SUM(\mult_44/SUMB[105][1] ) );
  FADDER \mult_44/S1_105_0  ( .CIN(\mult_44/ab[105][0] ), .IN0(
        \mult_44/CARRYB[104][0] ), .IN1(\mult_44/SUMB[104][1] ), .COUT(
        \mult_44/CARRYB[105][0] ), .SUM(clocal[105]) );
  FADDER \mult_44/S3_106_2  ( .CIN(\mult_44/ab[106][2] ), .IN0(
        \mult_44/CARRYB[105][2] ), .IN1(\mult_44/ab[105][3] ), .COUT(
        \mult_44/CARRYB[106][2] ), .SUM(\mult_44/SUMB[106][2] ) );
  FADDER \mult_44/S2_106_1  ( .CIN(\mult_44/ab[106][1] ), .IN0(
        \mult_44/CARRYB[105][1] ), .IN1(\mult_44/SUMB[105][2] ), .COUT(
        \mult_44/CARRYB[106][1] ), .SUM(\mult_44/SUMB[106][1] ) );
  FADDER \mult_44/S1_106_0  ( .CIN(\mult_44/ab[106][0] ), .IN0(
        \mult_44/CARRYB[105][0] ), .IN1(\mult_44/SUMB[105][1] ), .COUT(
        \mult_44/CARRYB[106][0] ), .SUM(clocal[106]) );
  FADDER \mult_44/S3_107_2  ( .CIN(\mult_44/ab[107][2] ), .IN0(
        \mult_44/CARRYB[106][2] ), .IN1(\mult_44/ab[106][3] ), .COUT(
        \mult_44/CARRYB[107][2] ), .SUM(\mult_44/SUMB[107][2] ) );
  FADDER \mult_44/S2_107_1  ( .CIN(\mult_44/ab[107][1] ), .IN0(
        \mult_44/CARRYB[106][1] ), .IN1(\mult_44/SUMB[106][2] ), .COUT(
        \mult_44/CARRYB[107][1] ), .SUM(\mult_44/SUMB[107][1] ) );
  FADDER \mult_44/S1_107_0  ( .CIN(\mult_44/ab[107][0] ), .IN0(
        \mult_44/CARRYB[106][0] ), .IN1(\mult_44/SUMB[106][1] ), .COUT(
        \mult_44/CARRYB[107][0] ), .SUM(clocal[107]) );
  FADDER \mult_44/S3_108_2  ( .CIN(\mult_44/ab[108][2] ), .IN0(
        \mult_44/CARRYB[107][2] ), .IN1(\mult_44/ab[107][3] ), .COUT(
        \mult_44/CARRYB[108][2] ), .SUM(\mult_44/SUMB[108][2] ) );
  FADDER \mult_44/S2_108_1  ( .CIN(\mult_44/ab[108][1] ), .IN0(
        \mult_44/CARRYB[107][1] ), .IN1(\mult_44/SUMB[107][2] ), .COUT(
        \mult_44/CARRYB[108][1] ), .SUM(\mult_44/SUMB[108][1] ) );
  FADDER \mult_44/S1_108_0  ( .CIN(\mult_44/ab[108][0] ), .IN0(
        \mult_44/CARRYB[107][0] ), .IN1(\mult_44/SUMB[107][1] ), .COUT(
        \mult_44/CARRYB[108][0] ), .SUM(clocal[108]) );
  FADDER \mult_44/S3_109_2  ( .CIN(\mult_44/ab[109][2] ), .IN0(
        \mult_44/CARRYB[108][2] ), .IN1(\mult_44/ab[108][3] ), .COUT(
        \mult_44/CARRYB[109][2] ), .SUM(\mult_44/SUMB[109][2] ) );
  FADDER \mult_44/S2_109_1  ( .CIN(\mult_44/ab[109][1] ), .IN0(
        \mult_44/CARRYB[108][1] ), .IN1(\mult_44/SUMB[108][2] ), .COUT(
        \mult_44/CARRYB[109][1] ), .SUM(\mult_44/SUMB[109][1] ) );
  FADDER \mult_44/S1_109_0  ( .CIN(\mult_44/ab[109][0] ), .IN0(
        \mult_44/CARRYB[108][0] ), .IN1(\mult_44/SUMB[108][1] ), .COUT(
        \mult_44/CARRYB[109][0] ), .SUM(clocal[109]) );
  FADDER \mult_44/S3_110_2  ( .CIN(\mult_44/ab[110][2] ), .IN0(
        \mult_44/CARRYB[109][2] ), .IN1(\mult_44/ab[109][3] ), .COUT(
        \mult_44/CARRYB[110][2] ), .SUM(\mult_44/SUMB[110][2] ) );
  FADDER \mult_44/S2_110_1  ( .CIN(\mult_44/ab[110][1] ), .IN0(
        \mult_44/CARRYB[109][1] ), .IN1(\mult_44/SUMB[109][2] ), .COUT(
        \mult_44/CARRYB[110][1] ), .SUM(\mult_44/SUMB[110][1] ) );
  FADDER \mult_44/S1_110_0  ( .CIN(\mult_44/ab[110][0] ), .IN0(
        \mult_44/CARRYB[109][0] ), .IN1(\mult_44/SUMB[109][1] ), .COUT(
        \mult_44/CARRYB[110][0] ), .SUM(clocal[110]) );
  FADDER \mult_44/S3_111_2  ( .CIN(\mult_44/ab[111][2] ), .IN0(
        \mult_44/CARRYB[110][2] ), .IN1(\mult_44/ab[110][3] ), .COUT(
        \mult_44/CARRYB[111][2] ), .SUM(\mult_44/SUMB[111][2] ) );
  FADDER \mult_44/S2_111_1  ( .CIN(\mult_44/ab[111][1] ), .IN0(
        \mult_44/CARRYB[110][1] ), .IN1(\mult_44/SUMB[110][2] ), .COUT(
        \mult_44/CARRYB[111][1] ), .SUM(\mult_44/SUMB[111][1] ) );
  FADDER \mult_44/S1_111_0  ( .CIN(\mult_44/ab[111][0] ), .IN0(
        \mult_44/CARRYB[110][0] ), .IN1(\mult_44/SUMB[110][1] ), .COUT(
        \mult_44/CARRYB[111][0] ), .SUM(clocal[111]) );
  FADDER \mult_44/S3_112_2  ( .CIN(\mult_44/ab[112][2] ), .IN0(
        \mult_44/CARRYB[111][2] ), .IN1(\mult_44/ab[111][3] ), .COUT(
        \mult_44/CARRYB[112][2] ), .SUM(\mult_44/SUMB[112][2] ) );
  FADDER \mult_44/S2_112_1  ( .CIN(\mult_44/ab[112][1] ), .IN0(
        \mult_44/CARRYB[111][1] ), .IN1(\mult_44/SUMB[111][2] ), .COUT(
        \mult_44/CARRYB[112][1] ), .SUM(\mult_44/SUMB[112][1] ) );
  FADDER \mult_44/S1_112_0  ( .CIN(\mult_44/ab[112][0] ), .IN0(
        \mult_44/CARRYB[111][0] ), .IN1(\mult_44/SUMB[111][1] ), .COUT(
        \mult_44/CARRYB[112][0] ), .SUM(clocal[112]) );
  FADDER \mult_44/S3_113_2  ( .CIN(\mult_44/ab[113][2] ), .IN0(
        \mult_44/CARRYB[112][2] ), .IN1(\mult_44/ab[112][3] ), .COUT(
        \mult_44/CARRYB[113][2] ), .SUM(\mult_44/SUMB[113][2] ) );
  FADDER \mult_44/S2_113_1  ( .CIN(\mult_44/ab[113][1] ), .IN0(
        \mult_44/CARRYB[112][1] ), .IN1(\mult_44/SUMB[112][2] ), .COUT(
        \mult_44/CARRYB[113][1] ), .SUM(\mult_44/SUMB[113][1] ) );
  FADDER \mult_44/S1_113_0  ( .CIN(\mult_44/ab[113][0] ), .IN0(
        \mult_44/CARRYB[112][0] ), .IN1(\mult_44/SUMB[112][1] ), .COUT(
        \mult_44/CARRYB[113][0] ), .SUM(clocal[113]) );
  FADDER \mult_44/S3_114_2  ( .CIN(\mult_44/ab[114][2] ), .IN0(
        \mult_44/CARRYB[113][2] ), .IN1(\mult_44/ab[113][3] ), .COUT(
        \mult_44/CARRYB[114][2] ), .SUM(\mult_44/SUMB[114][2] ) );
  FADDER \mult_44/S2_114_1  ( .CIN(\mult_44/ab[114][1] ), .IN0(
        \mult_44/CARRYB[113][1] ), .IN1(\mult_44/SUMB[113][2] ), .COUT(
        \mult_44/CARRYB[114][1] ), .SUM(\mult_44/SUMB[114][1] ) );
  FADDER \mult_44/S1_114_0  ( .CIN(\mult_44/ab[114][0] ), .IN0(
        \mult_44/CARRYB[113][0] ), .IN1(\mult_44/SUMB[113][1] ), .COUT(
        \mult_44/CARRYB[114][0] ), .SUM(clocal[114]) );
  FADDER \mult_44/S3_115_2  ( .CIN(\mult_44/ab[115][2] ), .IN0(
        \mult_44/CARRYB[114][2] ), .IN1(\mult_44/ab[114][3] ), .COUT(
        \mult_44/CARRYB[115][2] ), .SUM(\mult_44/SUMB[115][2] ) );
  FADDER \mult_44/S2_115_1  ( .CIN(\mult_44/ab[115][1] ), .IN0(
        \mult_44/CARRYB[114][1] ), .IN1(\mult_44/SUMB[114][2] ), .COUT(
        \mult_44/CARRYB[115][1] ), .SUM(\mult_44/SUMB[115][1] ) );
  FADDER \mult_44/S1_115_0  ( .CIN(\mult_44/ab[115][0] ), .IN0(
        \mult_44/CARRYB[114][0] ), .IN1(\mult_44/SUMB[114][1] ), .COUT(
        \mult_44/CARRYB[115][0] ), .SUM(clocal[115]) );
  FADDER \mult_44/S3_116_2  ( .CIN(\mult_44/ab[116][2] ), .IN0(
        \mult_44/CARRYB[115][2] ), .IN1(\mult_44/ab[115][3] ), .COUT(
        \mult_44/CARRYB[116][2] ), .SUM(\mult_44/SUMB[116][2] ) );
  FADDER \mult_44/S2_116_1  ( .CIN(\mult_44/ab[116][1] ), .IN0(
        \mult_44/CARRYB[115][1] ), .IN1(\mult_44/SUMB[115][2] ), .COUT(
        \mult_44/CARRYB[116][1] ), .SUM(\mult_44/SUMB[116][1] ) );
  FADDER \mult_44/S1_116_0  ( .CIN(\mult_44/ab[116][0] ), .IN0(
        \mult_44/CARRYB[115][0] ), .IN1(\mult_44/SUMB[115][1] ), .COUT(
        \mult_44/CARRYB[116][0] ), .SUM(clocal[116]) );
  FADDER \mult_44/S3_117_2  ( .CIN(\mult_44/ab[117][2] ), .IN0(
        \mult_44/CARRYB[116][2] ), .IN1(\mult_44/ab[116][3] ), .COUT(
        \mult_44/CARRYB[117][2] ), .SUM(\mult_44/SUMB[117][2] ) );
  FADDER \mult_44/S2_117_1  ( .CIN(\mult_44/ab[117][1] ), .IN0(
        \mult_44/CARRYB[116][1] ), .IN1(\mult_44/SUMB[116][2] ), .COUT(
        \mult_44/CARRYB[117][1] ), .SUM(\mult_44/SUMB[117][1] ) );
  FADDER \mult_44/S1_117_0  ( .CIN(\mult_44/ab[117][0] ), .IN0(
        \mult_44/CARRYB[116][0] ), .IN1(\mult_44/SUMB[116][1] ), .COUT(
        \mult_44/CARRYB[117][0] ), .SUM(clocal[117]) );
  FADDER \mult_44/S3_118_2  ( .CIN(\mult_44/ab[118][2] ), .IN0(
        \mult_44/CARRYB[117][2] ), .IN1(\mult_44/ab[117][3] ), .COUT(
        \mult_44/CARRYB[118][2] ), .SUM(\mult_44/SUMB[118][2] ) );
  FADDER \mult_44/S2_118_1  ( .CIN(\mult_44/ab[118][1] ), .IN0(
        \mult_44/CARRYB[117][1] ), .IN1(\mult_44/SUMB[117][2] ), .COUT(
        \mult_44/CARRYB[118][1] ), .SUM(\mult_44/SUMB[118][1] ) );
  FADDER \mult_44/S1_118_0  ( .CIN(\mult_44/ab[118][0] ), .IN0(
        \mult_44/CARRYB[117][0] ), .IN1(\mult_44/SUMB[117][1] ), .COUT(
        \mult_44/CARRYB[118][0] ), .SUM(clocal[118]) );
  FADDER \mult_44/S3_119_2  ( .CIN(\mult_44/ab[119][2] ), .IN0(
        \mult_44/CARRYB[118][2] ), .IN1(\mult_44/ab[118][3] ), .COUT(
        \mult_44/CARRYB[119][2] ), .SUM(\mult_44/SUMB[119][2] ) );
  FADDER \mult_44/S2_119_1  ( .CIN(\mult_44/ab[119][1] ), .IN0(
        \mult_44/CARRYB[118][1] ), .IN1(\mult_44/SUMB[118][2] ), .COUT(
        \mult_44/CARRYB[119][1] ), .SUM(\mult_44/SUMB[119][1] ) );
  FADDER \mult_44/S1_119_0  ( .CIN(\mult_44/ab[119][0] ), .IN0(
        \mult_44/CARRYB[118][0] ), .IN1(\mult_44/SUMB[118][1] ), .COUT(
        \mult_44/CARRYB[119][0] ), .SUM(clocal[119]) );
  FADDER \mult_44/S3_120_2  ( .CIN(\mult_44/ab[120][2] ), .IN0(
        \mult_44/CARRYB[119][2] ), .IN1(\mult_44/ab[119][3] ), .COUT(
        \mult_44/CARRYB[120][2] ), .SUM(\mult_44/SUMB[120][2] ) );
  FADDER \mult_44/S2_120_1  ( .CIN(\mult_44/ab[120][1] ), .IN0(
        \mult_44/CARRYB[119][1] ), .IN1(\mult_44/SUMB[119][2] ), .COUT(
        \mult_44/CARRYB[120][1] ), .SUM(\mult_44/SUMB[120][1] ) );
  FADDER \mult_44/S1_120_0  ( .CIN(\mult_44/ab[120][0] ), .IN0(
        \mult_44/CARRYB[119][0] ), .IN1(\mult_44/SUMB[119][1] ), .COUT(
        \mult_44/CARRYB[120][0] ), .SUM(clocal[120]) );
  FADDER \mult_44/S3_121_2  ( .CIN(\mult_44/ab[121][2] ), .IN0(
        \mult_44/CARRYB[120][2] ), .IN1(\mult_44/ab[120][3] ), .COUT(
        \mult_44/CARRYB[121][2] ), .SUM(\mult_44/SUMB[121][2] ) );
  FADDER \mult_44/S2_121_1  ( .CIN(\mult_44/ab[121][1] ), .IN0(
        \mult_44/CARRYB[120][1] ), .IN1(\mult_44/SUMB[120][2] ), .COUT(
        \mult_44/CARRYB[121][1] ), .SUM(\mult_44/SUMB[121][1] ) );
  FADDER \mult_44/S1_121_0  ( .CIN(\mult_44/ab[121][0] ), .IN0(
        \mult_44/CARRYB[120][0] ), .IN1(\mult_44/SUMB[120][1] ), .COUT(
        \mult_44/CARRYB[121][0] ), .SUM(clocal[121]) );
  FADDER \mult_44/S3_122_2  ( .CIN(\mult_44/ab[122][2] ), .IN0(
        \mult_44/CARRYB[121][2] ), .IN1(\mult_44/ab[121][3] ), .COUT(
        \mult_44/CARRYB[122][2] ), .SUM(\mult_44/SUMB[122][2] ) );
  FADDER \mult_44/S2_122_1  ( .CIN(\mult_44/ab[122][1] ), .IN0(
        \mult_44/CARRYB[121][1] ), .IN1(\mult_44/SUMB[121][2] ), .COUT(
        \mult_44/CARRYB[122][1] ), .SUM(\mult_44/SUMB[122][1] ) );
  FADDER \mult_44/S1_122_0  ( .CIN(\mult_44/ab[122][0] ), .IN0(
        \mult_44/CARRYB[121][0] ), .IN1(\mult_44/SUMB[121][1] ), .COUT(
        \mult_44/CARRYB[122][0] ), .SUM(clocal[122]) );
  FADDER \mult_44/S3_123_2  ( .CIN(\mult_44/ab[123][2] ), .IN0(
        \mult_44/CARRYB[122][2] ), .IN1(\mult_44/ab[122][3] ), .COUT(
        \mult_44/CARRYB[123][2] ), .SUM(\mult_44/SUMB[123][2] ) );
  FADDER \mult_44/S2_123_1  ( .CIN(\mult_44/ab[123][1] ), .IN0(
        \mult_44/CARRYB[122][1] ), .IN1(\mult_44/SUMB[122][2] ), .COUT(
        \mult_44/CARRYB[123][1] ), .SUM(\mult_44/SUMB[123][1] ) );
  FADDER \mult_44/S1_123_0  ( .CIN(\mult_44/ab[123][0] ), .IN0(
        \mult_44/CARRYB[122][0] ), .IN1(\mult_44/SUMB[122][1] ), .COUT(
        \mult_44/CARRYB[123][0] ), .SUM(clocal[123]) );
  FADDER \mult_44/S3_124_2  ( .CIN(\mult_44/ab[124][2] ), .IN0(
        \mult_44/CARRYB[123][2] ), .IN1(\mult_44/ab[123][3] ), .COUT(
        \mult_44/CARRYB[124][2] ), .SUM(\mult_44/SUMB[124][2] ) );
  FADDER \mult_44/S2_124_1  ( .CIN(\mult_44/ab[124][1] ), .IN0(
        \mult_44/CARRYB[123][1] ), .IN1(\mult_44/SUMB[123][2] ), .COUT(
        \mult_44/CARRYB[124][1] ), .SUM(\mult_44/SUMB[124][1] ) );
  FADDER \mult_44/S1_124_0  ( .CIN(\mult_44/ab[124][0] ), .IN0(
        \mult_44/CARRYB[123][0] ), .IN1(\mult_44/SUMB[123][1] ), .COUT(
        \mult_44/CARRYB[124][0] ), .SUM(clocal[124]) );
  FADDER \mult_44/S3_125_2  ( .CIN(\mult_44/ab[125][2] ), .IN0(
        \mult_44/CARRYB[124][2] ), .IN1(\mult_44/ab[124][3] ), .SUM(
        \mult_44/SUMB[125][2] ) );
  FADDER \mult_44/S2_125_1  ( .CIN(\mult_44/ab[125][1] ), .IN0(
        \mult_44/CARRYB[124][1] ), .IN1(\mult_44/SUMB[124][2] ), .COUT(
        \mult_44/CARRYB[125][1] ), .SUM(\mult_44/SUMB[125][1] ) );
  FADDER \mult_44/S1_125_0  ( .CIN(\mult_44/ab[125][0] ), .IN0(
        \mult_44/CARRYB[124][0] ), .IN1(\mult_44/SUMB[124][1] ), .COUT(
        \mult_44/CARRYB[125][0] ), .SUM(clocal[125]) );
  FADDER \mult_44/S2_126_1  ( .CIN(\mult_44/ab[126][1] ), .IN0(
        \mult_44/CARRYB[125][1] ), .IN1(\mult_44/SUMB[125][2] ), .SUM(
        \mult_44/SUMB[126][1] ) );
  FADDER \mult_44/S1_126_0  ( .CIN(\mult_44/ab[126][0] ), .IN0(
        \mult_44/CARRYB[125][0] ), .IN1(\mult_44/SUMB[125][1] ), .COUT(
        \mult_44/CARRYB[126][0] ), .SUM(clocal[126]) );
  FADDER \mult_44/S4_0  ( .CIN(\mult_44/ab[127][0] ), .IN0(
        \mult_44/CARRYB[126][0] ), .IN1(\mult_44/SUMB[126][1] ), .SUM(
        \mult_44/SUMB[127][0] ) );
  MUX U256 ( .IN0(clocal[120]), .IN1(n359), .SEL(n360), .F(n355) );
  MUX U257 ( .IN0(clocal[116]), .IN1(n372), .SEL(n373), .F(n368) );
  MUX U258 ( .IN0(clocal[112]), .IN1(n384), .SEL(n385), .F(n380) );
  MUX U259 ( .IN0(clocal[108]), .IN1(n397), .SEL(n398), .F(n392) );
  MUX U260 ( .IN0(clocal[104]), .IN1(n409), .SEL(n410), .F(n405) );
  MUX U261 ( .IN0(clocal[100]), .IN1(n421), .SEL(n422), .F(n417) );
  MUX U262 ( .IN0(clocal[96]), .IN1(n430), .SEL(n254), .F(n427) );
  MUX U263 ( .IN0(clocal[92]), .IN1(n438), .SEL(n258), .F(n435) );
  MUX U264 ( .IN0(clocal[88]), .IN1(n446), .SEL(n263), .F(n443) );
  MUX U265 ( .IN0(clocal[84]), .IN1(n454), .SEL(n267), .F(n451) );
  MUX U266 ( .IN0(clocal[80]), .IN1(n462), .SEL(n271), .F(n459) );
  MUX U267 ( .IN0(clocal[76]), .IN1(n470), .SEL(n276), .F(n467) );
  MUX U268 ( .IN0(clocal[72]), .IN1(n478), .SEL(n280), .F(n475) );
  MUX U269 ( .IN0(clocal[68]), .IN1(n486), .SEL(n285), .F(n483) );
  MUX U270 ( .IN0(clocal[64]), .IN1(n494), .SEL(n289), .F(n491) );
  MUX U271 ( .IN0(clocal[60]), .IN1(n502), .SEL(n293), .F(n499) );
  MUX U272 ( .IN0(clocal[56]), .IN1(n510), .SEL(n298), .F(n507) );
  MUX U273 ( .IN0(clocal[52]), .IN1(n518), .SEL(n302), .F(n515) );
  MUX U274 ( .IN0(clocal[48]), .IN1(n526), .SEL(n307), .F(n523) );
  MUX U275 ( .IN0(clocal[44]), .IN1(n534), .SEL(n311), .F(n531) );
  MUX U276 ( .IN0(clocal[40]), .IN1(n542), .SEL(n315), .F(n539) );
  MUX U277 ( .IN0(clocal[36]), .IN1(n550), .SEL(n319), .F(n547) );
  MUX U278 ( .IN0(clocal[32]), .IN1(n558), .SEL(n323), .F(n555) );
  MUX U279 ( .IN0(clocal[28]), .IN1(n566), .SEL(n327), .F(n563) );
  MUX U280 ( .IN0(clocal[24]), .IN1(n574), .SEL(n331), .F(n571) );
  MUX U281 ( .IN0(clocal[20]), .IN1(n582), .SEL(n335), .F(n579) );
  MUX U282 ( .IN0(clocal[16]), .IN1(n590), .SEL(n339), .F(n587) );
  MUX U283 ( .IN0(clocal[12]), .IN1(n598), .SEL(n343), .F(n595) );
  MUX U284 ( .IN0(clocal[8]), .IN1(n606), .SEL(n261), .F(n603) );
  MUX U285 ( .IN0(clocal[4]), .IN1(n614), .SEL(n305), .F(n611) );
  MUX U286 ( .IN0(clocal[119]), .IN1(n361), .SEL(n362), .F(n359) );
  MUX U287 ( .IN0(clocal[115]), .IN1(n374), .SEL(n375), .F(n372) );
  MUX U288 ( .IN0(clocal[111]), .IN1(n386), .SEL(n387), .F(n384) );
  MUX U289 ( .IN0(clocal[107]), .IN1(n399), .SEL(n400), .F(n397) );
  MUX U290 ( .IN0(clocal[103]), .IN1(n411), .SEL(n412), .F(n409) );
  MUX U291 ( .IN0(clocal[99]), .IN1(n423), .SEL(n251), .F(n421) );
  MUX U292 ( .IN0(clocal[95]), .IN1(n431), .SEL(n255), .F(n430) );
  MUX U293 ( .IN0(clocal[91]), .IN1(n439), .SEL(n259), .F(n438) );
  MUX U294 ( .IN0(clocal[87]), .IN1(n447), .SEL(n264), .F(n446) );
  MUX U295 ( .IN0(clocal[83]), .IN1(n455), .SEL(n268), .F(n454) );
  MUX U296 ( .IN0(clocal[79]), .IN1(n463), .SEL(n273), .F(n462) );
  MUX U297 ( .IN0(clocal[75]), .IN1(n471), .SEL(n277), .F(n470) );
  MUX U298 ( .IN0(clocal[71]), .IN1(n479), .SEL(n281), .F(n478) );
  MUX U299 ( .IN0(clocal[67]), .IN1(n487), .SEL(n286), .F(n486) );
  MUX U300 ( .IN0(clocal[63]), .IN1(n495), .SEL(n290), .F(n494) );
  MUX U301 ( .IN0(clocal[59]), .IN1(n503), .SEL(n295), .F(n502) );
  MUX U302 ( .IN0(clocal[55]), .IN1(n511), .SEL(n299), .F(n510) );
  MUX U303 ( .IN0(clocal[51]), .IN1(n519), .SEL(n303), .F(n518) );
  MUX U304 ( .IN0(clocal[47]), .IN1(n527), .SEL(n308), .F(n526) );
  MUX U305 ( .IN0(clocal[43]), .IN1(n535), .SEL(n312), .F(n534) );
  MUX U306 ( .IN0(clocal[39]), .IN1(n543), .SEL(n316), .F(n542) );
  MUX U307 ( .IN0(clocal[35]), .IN1(n551), .SEL(n320), .F(n550) );
  MUX U308 ( .IN0(clocal[31]), .IN1(n559), .SEL(n324), .F(n558) );
  MUX U309 ( .IN0(clocal[27]), .IN1(n567), .SEL(n328), .F(n566) );
  MUX U310 ( .IN0(clocal[23]), .IN1(n575), .SEL(n332), .F(n574) );
  MUX U311 ( .IN0(clocal[19]), .IN1(n583), .SEL(n336), .F(n582) );
  MUX U312 ( .IN0(clocal[15]), .IN1(n591), .SEL(n340), .F(n590) );
  MUX U313 ( .IN0(clocal[11]), .IN1(n599), .SEL(n363), .F(n598) );
  MUX U314 ( .IN0(clocal[7]), .IN1(n607), .SEL(n272), .F(n606) );
  MUX U315 ( .IN0(\mult_44/PROD1[3] ), .IN1(n615), .SEL(n616), .F(n614) );
  MUX U316 ( .IN0(clocal[123]), .IN1(n349), .SEL(n350), .F(n348) );
  XNOR U317 ( .A(n615), .B(sreg[131]), .Z(n616) );
  XNOR U318 ( .A(n349), .B(sreg[251]), .Z(n350) );
  XNOR U319 ( .A(n359), .B(sreg[248]), .Z(n360) );
  XNOR U320 ( .A(n368), .B(sreg[245]), .Z(n371) );
  XNOR U321 ( .A(n376), .B(sreg[242]), .Z(n379) );
  XNOR U322 ( .A(n386), .B(sreg[239]), .Z(n387) );
  XNOR U323 ( .A(n397), .B(sreg[236]), .Z(n398) );
  XNOR U324 ( .A(n405), .B(sreg[233]), .Z(n408) );
  XNOR U325 ( .A(n413), .B(sreg[230]), .Z(n416) );
  XNOR U326 ( .A(n423), .B(sreg[227]), .Z(n251) );
  XNOR U327 ( .A(n430), .B(sreg[224]), .Z(n254) );
  XNOR U328 ( .A(n435), .B(sreg[221]), .Z(n257) );
  XNOR U329 ( .A(n440), .B(sreg[218]), .Z(n260) );
  XNOR U330 ( .A(n447), .B(sreg[215]), .Z(n264) );
  XNOR U331 ( .A(n454), .B(sreg[212]), .Z(n267) );
  XNOR U332 ( .A(n459), .B(sreg[209]), .Z(n270) );
  XNOR U333 ( .A(n464), .B(sreg[206]), .Z(n274) );
  XNOR U334 ( .A(n471), .B(sreg[203]), .Z(n277) );
  XNOR U335 ( .A(n478), .B(sreg[200]), .Z(n280) );
  XNOR U336 ( .A(n483), .B(sreg[197]), .Z(n284) );
  XNOR U337 ( .A(n488), .B(sreg[194]), .Z(n287) );
  XNOR U338 ( .A(n495), .B(sreg[191]), .Z(n290) );
  XNOR U339 ( .A(n502), .B(sreg[188]), .Z(n293) );
  XNOR U340 ( .A(n507), .B(sreg[185]), .Z(n297) );
  XNOR U341 ( .A(n512), .B(sreg[182]), .Z(n300) );
  XNOR U342 ( .A(n519), .B(sreg[179]), .Z(n303) );
  XNOR U343 ( .A(n526), .B(sreg[176]), .Z(n307) );
  XNOR U344 ( .A(n531), .B(sreg[173]), .Z(n310) );
  XNOR U345 ( .A(n536), .B(sreg[170]), .Z(n313) );
  XNOR U346 ( .A(n543), .B(sreg[167]), .Z(n316) );
  XNOR U347 ( .A(n550), .B(sreg[164]), .Z(n319) );
  XNOR U348 ( .A(n555), .B(sreg[161]), .Z(n322) );
  XNOR U349 ( .A(n560), .B(sreg[158]), .Z(n325) );
  XNOR U350 ( .A(n567), .B(sreg[155]), .Z(n328) );
  XNOR U351 ( .A(n574), .B(sreg[152]), .Z(n331) );
  XNOR U352 ( .A(n579), .B(sreg[149]), .Z(n334) );
  XNOR U353 ( .A(n584), .B(sreg[146]), .Z(n337) );
  XNOR U354 ( .A(n591), .B(sreg[143]), .Z(n340) );
  XNOR U355 ( .A(n598), .B(sreg[140]), .Z(n343) );
  XNOR U356 ( .A(n603), .B(sreg[137]), .Z(n250) );
  XNOR U357 ( .A(n608), .B(sreg[134]), .Z(n283) );
  XNOR U358 ( .A(n617), .B(sreg[130]), .Z(n620) );
  XNOR U359 ( .A(n351), .B(sreg[250]), .Z(n354) );
  XNOR U360 ( .A(n361), .B(sreg[247]), .Z(n362) );
  XNOR U361 ( .A(n372), .B(sreg[244]), .Z(n373) );
  XNOR U362 ( .A(n380), .B(sreg[241]), .Z(n383) );
  XNOR U363 ( .A(n388), .B(sreg[238]), .Z(n391) );
  XNOR U364 ( .A(n399), .B(sreg[235]), .Z(n400) );
  XNOR U365 ( .A(n409), .B(sreg[232]), .Z(n410) );
  XNOR U366 ( .A(n417), .B(sreg[229]), .Z(n420) );
  XNOR U367 ( .A(n424), .B(sreg[226]), .Z(n252) );
  XNOR U368 ( .A(n431), .B(sreg[223]), .Z(n255) );
  XNOR U369 ( .A(n438), .B(sreg[220]), .Z(n258) );
  XNOR U370 ( .A(n443), .B(sreg[217]), .Z(n262) );
  XNOR U371 ( .A(n448), .B(sreg[214]), .Z(n265) );
  XNOR U372 ( .A(n455), .B(sreg[211]), .Z(n268) );
  XNOR U373 ( .A(n462), .B(sreg[208]), .Z(n271) );
  XNOR U374 ( .A(n467), .B(sreg[205]), .Z(n275) );
  XNOR U375 ( .A(n472), .B(sreg[202]), .Z(n278) );
  XNOR U376 ( .A(n479), .B(sreg[199]), .Z(n281) );
  XNOR U377 ( .A(n486), .B(sreg[196]), .Z(n285) );
  XNOR U378 ( .A(n491), .B(sreg[193]), .Z(n288) );
  XNOR U379 ( .A(n496), .B(sreg[190]), .Z(n291) );
  XNOR U380 ( .A(n503), .B(sreg[187]), .Z(n295) );
  XNOR U381 ( .A(n510), .B(sreg[184]), .Z(n298) );
  XNOR U382 ( .A(n515), .B(sreg[181]), .Z(n301) );
  XNOR U383 ( .A(n520), .B(sreg[178]), .Z(n304) );
  XNOR U384 ( .A(n527), .B(sreg[175]), .Z(n308) );
  XNOR U385 ( .A(n534), .B(sreg[172]), .Z(n311) );
  XNOR U386 ( .A(n539), .B(sreg[169]), .Z(n314) );
  XNOR U387 ( .A(n544), .B(sreg[166]), .Z(n317) );
  XNOR U388 ( .A(n551), .B(sreg[163]), .Z(n320) );
  XNOR U389 ( .A(n558), .B(sreg[160]), .Z(n323) );
  XNOR U390 ( .A(n563), .B(sreg[157]), .Z(n326) );
  XNOR U391 ( .A(n568), .B(sreg[154]), .Z(n329) );
  XNOR U392 ( .A(n575), .B(sreg[151]), .Z(n332) );
  XNOR U393 ( .A(n582), .B(sreg[148]), .Z(n335) );
  XNOR U394 ( .A(n587), .B(sreg[145]), .Z(n338) );
  XNOR U395 ( .A(n592), .B(sreg[142]), .Z(n341) );
  XNOR U396 ( .A(n599), .B(sreg[139]), .Z(n363) );
  XNOR U397 ( .A(n606), .B(sreg[136]), .Z(n261) );
  XNOR U398 ( .A(n611), .B(sreg[133]), .Z(n294) );
  XNOR U399 ( .A(n355), .B(sreg[249]), .Z(n358) );
  XNOR U400 ( .A(n364), .B(sreg[246]), .Z(n367) );
  XNOR U401 ( .A(n374), .B(sreg[243]), .Z(n375) );
  XNOR U402 ( .A(n384), .B(sreg[240]), .Z(n385) );
  XNOR U403 ( .A(n392), .B(sreg[237]), .Z(n395) );
  XNOR U404 ( .A(n401), .B(sreg[234]), .Z(n404) );
  XNOR U405 ( .A(n411), .B(sreg[231]), .Z(n412) );
  XNOR U406 ( .A(n421), .B(sreg[228]), .Z(n422) );
  XNOR U407 ( .A(n427), .B(sreg[225]), .Z(n253) );
  XNOR U408 ( .A(n432), .B(sreg[222]), .Z(n256) );
  XNOR U409 ( .A(n439), .B(sreg[219]), .Z(n259) );
  XNOR U410 ( .A(n446), .B(sreg[216]), .Z(n263) );
  XNOR U411 ( .A(n451), .B(sreg[213]), .Z(n266) );
  XNOR U412 ( .A(n456), .B(sreg[210]), .Z(n269) );
  XNOR U413 ( .A(n463), .B(sreg[207]), .Z(n273) );
  XNOR U414 ( .A(n470), .B(sreg[204]), .Z(n276) );
  XNOR U415 ( .A(n475), .B(sreg[201]), .Z(n279) );
  XNOR U416 ( .A(n480), .B(sreg[198]), .Z(n282) );
  XNOR U417 ( .A(n487), .B(sreg[195]), .Z(n286) );
  XNOR U418 ( .A(n494), .B(sreg[192]), .Z(n289) );
  XNOR U419 ( .A(n499), .B(sreg[189]), .Z(n292) );
  XNOR U420 ( .A(n504), .B(sreg[186]), .Z(n296) );
  XNOR U421 ( .A(n511), .B(sreg[183]), .Z(n299) );
  XNOR U422 ( .A(n518), .B(sreg[180]), .Z(n302) );
  XNOR U423 ( .A(n523), .B(sreg[177]), .Z(n306) );
  XNOR U424 ( .A(n528), .B(sreg[174]), .Z(n309) );
  XNOR U425 ( .A(n535), .B(sreg[171]), .Z(n312) );
  XNOR U426 ( .A(n542), .B(sreg[168]), .Z(n315) );
  XNOR U427 ( .A(n547), .B(sreg[165]), .Z(n318) );
  XNOR U428 ( .A(n552), .B(sreg[162]), .Z(n321) );
  XNOR U429 ( .A(n559), .B(sreg[159]), .Z(n324) );
  XNOR U430 ( .A(n566), .B(sreg[156]), .Z(n327) );
  XNOR U431 ( .A(n571), .B(sreg[153]), .Z(n330) );
  XNOR U432 ( .A(n576), .B(sreg[150]), .Z(n333) );
  XNOR U433 ( .A(n583), .B(sreg[147]), .Z(n336) );
  XNOR U434 ( .A(n590), .B(sreg[144]), .Z(n339) );
  XNOR U435 ( .A(n595), .B(sreg[141]), .Z(n342) );
  XNOR U436 ( .A(n600), .B(sreg[138]), .Z(n396) );
  XNOR U437 ( .A(n607), .B(sreg[135]), .Z(n272) );
  XNOR U438 ( .A(n614), .B(sreg[132]), .Z(n305) );
  AND U439 ( .A(\mult_44/ab[0][1] ), .B(\mult_44/ab[1][0] ), .Z(
        \mult_44/CARRYB[1][0] ) );
  XOR U440 ( .A(\mult_44/ab[0][1] ), .B(\mult_44/ab[1][0] ), .Z(clocal[1]) );
  AND U441 ( .A(\mult_44/ab[1][1] ), .B(\mult_44/ab[0][2] ), .Z(
        \mult_44/CARRYB[1][1] ) );
  XOR U442 ( .A(\mult_44/ab[0][2] ), .B(\mult_44/ab[1][1] ), .Z(
        \mult_44/SUMB[1][1] ) );
  AND U443 ( .A(\mult_44/ab[1][2] ), .B(\mult_44/ab[0][3] ), .Z(
        \mult_44/CARRYB[1][2] ) );
  XOR U444 ( .A(\mult_44/ab[0][3] ), .B(\mult_44/ab[1][2] ), .Z(
        \mult_44/SUMB[1][2] ) );
  XNOR U445 ( .A(clocal[9]), .B(n250), .Z(swire[9]) );
  XNOR U446 ( .A(clocal[99]), .B(n251), .Z(swire[99]) );
  XNOR U447 ( .A(clocal[98]), .B(n252), .Z(swire[98]) );
  XNOR U448 ( .A(clocal[97]), .B(n253), .Z(swire[97]) );
  XNOR U449 ( .A(clocal[96]), .B(n254), .Z(swire[96]) );
  XNOR U450 ( .A(clocal[95]), .B(n255), .Z(swire[95]) );
  XNOR U451 ( .A(clocal[94]), .B(n256), .Z(swire[94]) );
  XNOR U452 ( .A(clocal[93]), .B(n257), .Z(swire[93]) );
  XNOR U453 ( .A(clocal[92]), .B(n258), .Z(swire[92]) );
  XNOR U454 ( .A(clocal[91]), .B(n259), .Z(swire[91]) );
  XNOR U455 ( .A(clocal[90]), .B(n260), .Z(swire[90]) );
  XNOR U456 ( .A(clocal[8]), .B(n261), .Z(swire[8]) );
  XNOR U457 ( .A(clocal[89]), .B(n262), .Z(swire[89]) );
  XNOR U458 ( .A(clocal[88]), .B(n263), .Z(swire[88]) );
  XNOR U459 ( .A(clocal[87]), .B(n264), .Z(swire[87]) );
  XNOR U460 ( .A(clocal[86]), .B(n265), .Z(swire[86]) );
  XNOR U461 ( .A(clocal[85]), .B(n266), .Z(swire[85]) );
  XNOR U462 ( .A(clocal[84]), .B(n267), .Z(swire[84]) );
  XNOR U463 ( .A(clocal[83]), .B(n268), .Z(swire[83]) );
  XNOR U464 ( .A(clocal[82]), .B(n269), .Z(swire[82]) );
  XNOR U465 ( .A(clocal[81]), .B(n270), .Z(swire[81]) );
  XNOR U466 ( .A(clocal[80]), .B(n271), .Z(swire[80]) );
  XNOR U467 ( .A(clocal[7]), .B(n272), .Z(swire[7]) );
  XNOR U468 ( .A(clocal[79]), .B(n273), .Z(swire[79]) );
  XNOR U469 ( .A(clocal[78]), .B(n274), .Z(swire[78]) );
  XNOR U470 ( .A(clocal[77]), .B(n275), .Z(swire[77]) );
  XNOR U471 ( .A(clocal[76]), .B(n276), .Z(swire[76]) );
  XNOR U472 ( .A(clocal[75]), .B(n277), .Z(swire[75]) );
  XNOR U473 ( .A(clocal[74]), .B(n278), .Z(swire[74]) );
  XNOR U474 ( .A(clocal[73]), .B(n279), .Z(swire[73]) );
  XNOR U475 ( .A(clocal[72]), .B(n280), .Z(swire[72]) );
  XNOR U476 ( .A(clocal[71]), .B(n281), .Z(swire[71]) );
  XNOR U477 ( .A(clocal[70]), .B(n282), .Z(swire[70]) );
  XNOR U478 ( .A(clocal[6]), .B(n283), .Z(swire[6]) );
  XNOR U479 ( .A(clocal[69]), .B(n284), .Z(swire[69]) );
  XNOR U480 ( .A(clocal[68]), .B(n285), .Z(swire[68]) );
  XNOR U481 ( .A(clocal[67]), .B(n286), .Z(swire[67]) );
  XNOR U482 ( .A(clocal[66]), .B(n287), .Z(swire[66]) );
  XNOR U483 ( .A(clocal[65]), .B(n288), .Z(swire[65]) );
  XNOR U484 ( .A(clocal[64]), .B(n289), .Z(swire[64]) );
  XNOR U485 ( .A(clocal[63]), .B(n290), .Z(swire[63]) );
  XNOR U486 ( .A(clocal[62]), .B(n291), .Z(swire[62]) );
  XNOR U487 ( .A(clocal[61]), .B(n292), .Z(swire[61]) );
  XNOR U488 ( .A(clocal[60]), .B(n293), .Z(swire[60]) );
  XNOR U489 ( .A(clocal[5]), .B(n294), .Z(swire[5]) );
  XNOR U490 ( .A(clocal[59]), .B(n295), .Z(swire[59]) );
  XNOR U491 ( .A(clocal[58]), .B(n296), .Z(swire[58]) );
  XNOR U492 ( .A(clocal[57]), .B(n297), .Z(swire[57]) );
  XNOR U493 ( .A(clocal[56]), .B(n298), .Z(swire[56]) );
  XNOR U494 ( .A(clocal[55]), .B(n299), .Z(swire[55]) );
  XNOR U495 ( .A(clocal[54]), .B(n300), .Z(swire[54]) );
  XNOR U496 ( .A(clocal[53]), .B(n301), .Z(swire[53]) );
  XNOR U497 ( .A(clocal[52]), .B(n302), .Z(swire[52]) );
  XNOR U498 ( .A(clocal[51]), .B(n303), .Z(swire[51]) );
  XNOR U499 ( .A(clocal[50]), .B(n304), .Z(swire[50]) );
  XNOR U500 ( .A(clocal[4]), .B(n305), .Z(swire[4]) );
  XNOR U501 ( .A(clocal[49]), .B(n306), .Z(swire[49]) );
  XNOR U502 ( .A(clocal[48]), .B(n307), .Z(swire[48]) );
  XNOR U503 ( .A(clocal[47]), .B(n308), .Z(swire[47]) );
  XNOR U504 ( .A(clocal[46]), .B(n309), .Z(swire[46]) );
  XNOR U505 ( .A(clocal[45]), .B(n310), .Z(swire[45]) );
  XNOR U506 ( .A(clocal[44]), .B(n311), .Z(swire[44]) );
  XNOR U507 ( .A(clocal[43]), .B(n312), .Z(swire[43]) );
  XNOR U508 ( .A(clocal[42]), .B(n313), .Z(swire[42]) );
  XNOR U509 ( .A(clocal[41]), .B(n314), .Z(swire[41]) );
  XNOR U510 ( .A(clocal[40]), .B(n315), .Z(swire[40]) );
  XNOR U511 ( .A(clocal[39]), .B(n316), .Z(swire[39]) );
  XNOR U512 ( .A(clocal[38]), .B(n317), .Z(swire[38]) );
  XNOR U513 ( .A(clocal[37]), .B(n318), .Z(swire[37]) );
  XNOR U514 ( .A(clocal[36]), .B(n319), .Z(swire[36]) );
  XNOR U515 ( .A(clocal[35]), .B(n320), .Z(swire[35]) );
  XNOR U516 ( .A(clocal[34]), .B(n321), .Z(swire[34]) );
  XNOR U517 ( .A(clocal[33]), .B(n322), .Z(swire[33]) );
  XNOR U518 ( .A(clocal[32]), .B(n323), .Z(swire[32]) );
  XNOR U519 ( .A(clocal[31]), .B(n324), .Z(swire[31]) );
  XNOR U520 ( .A(clocal[30]), .B(n325), .Z(swire[30]) );
  XNOR U521 ( .A(clocal[29]), .B(n326), .Z(swire[29]) );
  XNOR U522 ( .A(clocal[28]), .B(n327), .Z(swire[28]) );
  XNOR U523 ( .A(clocal[27]), .B(n328), .Z(swire[27]) );
  XNOR U524 ( .A(clocal[26]), .B(n329), .Z(swire[26]) );
  XNOR U525 ( .A(clocal[25]), .B(n330), .Z(swire[25]) );
  XNOR U526 ( .A(clocal[24]), .B(n331), .Z(swire[24]) );
  XNOR U527 ( .A(clocal[23]), .B(n332), .Z(swire[23]) );
  XNOR U528 ( .A(clocal[22]), .B(n333), .Z(swire[22]) );
  XNOR U529 ( .A(clocal[21]), .B(n334), .Z(swire[21]) );
  XNOR U530 ( .A(clocal[20]), .B(n335), .Z(swire[20]) );
  XNOR U531 ( .A(clocal[19]), .B(n336), .Z(swire[19]) );
  XNOR U532 ( .A(clocal[18]), .B(n337), .Z(swire[18]) );
  XNOR U533 ( .A(clocal[17]), .B(n338), .Z(swire[17]) );
  XNOR U534 ( .A(clocal[16]), .B(n339), .Z(swire[16]) );
  XNOR U535 ( .A(clocal[15]), .B(n340), .Z(swire[15]) );
  XNOR U536 ( .A(clocal[14]), .B(n341), .Z(swire[14]) );
  XNOR U537 ( .A(clocal[13]), .B(n342), .Z(swire[13]) );
  XNOR U538 ( .A(clocal[12]), .B(n343), .Z(swire[12]) );
  XOR U539 ( .A(n344), .B(n345), .Z(swire[127]) );
  XOR U540 ( .A(\mult_44/SUMB[127][0] ), .B(n346), .Z(n345) );
  ANDN U541 ( .B(n344), .A(clocal[126]), .Z(n346) );
  XOR U542 ( .A(clocal[126]), .B(n344), .Z(swire[126]) );
  ANDN U543 ( .B(clocal[125]), .A(n347), .Z(n344) );
  XNOR U544 ( .A(clocal[125]), .B(n347), .Z(swire[125]) );
  NAND U545 ( .A(n348), .B(clocal[124]), .Z(n347) );
  XOR U546 ( .A(clocal[124]), .B(n348), .Z(swire[124]) );
  XNOR U547 ( .A(clocal[123]), .B(n350), .Z(swire[123]) );
  XOR U548 ( .A(n351), .B(n352), .Z(n349) );
  ANDN U549 ( .B(n353), .A(n354), .Z(n352) );
  XOR U550 ( .A(clocal[122]), .B(n351), .Z(n353) );
  XNOR U551 ( .A(clocal[122]), .B(n354), .Z(swire[122]) );
  XOR U552 ( .A(n355), .B(n356), .Z(n351) );
  ANDN U553 ( .B(n357), .A(n358), .Z(n356) );
  XOR U554 ( .A(clocal[121]), .B(n355), .Z(n357) );
  XNOR U555 ( .A(clocal[121]), .B(n358), .Z(swire[121]) );
  XNOR U556 ( .A(clocal[120]), .B(n360), .Z(swire[120]) );
  XNOR U557 ( .A(clocal[11]), .B(n363), .Z(swire[11]) );
  XNOR U558 ( .A(clocal[119]), .B(n362), .Z(swire[119]) );
  XOR U559 ( .A(n364), .B(n365), .Z(n361) );
  ANDN U560 ( .B(n366), .A(n367), .Z(n365) );
  XOR U561 ( .A(clocal[118]), .B(n364), .Z(n366) );
  XNOR U562 ( .A(clocal[118]), .B(n367), .Z(swire[118]) );
  XOR U563 ( .A(n368), .B(n369), .Z(n364) );
  ANDN U564 ( .B(n370), .A(n371), .Z(n369) );
  XOR U565 ( .A(clocal[117]), .B(n368), .Z(n370) );
  XNOR U566 ( .A(clocal[117]), .B(n371), .Z(swire[117]) );
  XNOR U567 ( .A(clocal[116]), .B(n373), .Z(swire[116]) );
  XNOR U568 ( .A(clocal[115]), .B(n375), .Z(swire[115]) );
  XOR U569 ( .A(n376), .B(n377), .Z(n374) );
  ANDN U570 ( .B(n378), .A(n379), .Z(n377) );
  XOR U571 ( .A(clocal[114]), .B(n376), .Z(n378) );
  XNOR U572 ( .A(clocal[114]), .B(n379), .Z(swire[114]) );
  XOR U573 ( .A(n380), .B(n381), .Z(n376) );
  ANDN U574 ( .B(n382), .A(n383), .Z(n381) );
  XOR U575 ( .A(clocal[113]), .B(n380), .Z(n382) );
  XNOR U576 ( .A(clocal[113]), .B(n383), .Z(swire[113]) );
  XNOR U577 ( .A(clocal[112]), .B(n385), .Z(swire[112]) );
  XNOR U578 ( .A(clocal[111]), .B(n387), .Z(swire[111]) );
  XOR U579 ( .A(n388), .B(n389), .Z(n386) );
  ANDN U580 ( .B(n390), .A(n391), .Z(n389) );
  XOR U581 ( .A(clocal[110]), .B(n388), .Z(n390) );
  XNOR U582 ( .A(clocal[110]), .B(n391), .Z(swire[110]) );
  XOR U583 ( .A(n392), .B(n393), .Z(n388) );
  ANDN U584 ( .B(n394), .A(n395), .Z(n393) );
  XOR U585 ( .A(clocal[109]), .B(n392), .Z(n394) );
  XNOR U586 ( .A(clocal[10]), .B(n396), .Z(swire[10]) );
  XNOR U587 ( .A(clocal[109]), .B(n395), .Z(swire[109]) );
  XNOR U588 ( .A(clocal[108]), .B(n398), .Z(swire[108]) );
  XNOR U589 ( .A(clocal[107]), .B(n400), .Z(swire[107]) );
  XOR U590 ( .A(n401), .B(n402), .Z(n399) );
  ANDN U591 ( .B(n403), .A(n404), .Z(n402) );
  XOR U592 ( .A(clocal[106]), .B(n401), .Z(n403) );
  XNOR U593 ( .A(clocal[106]), .B(n404), .Z(swire[106]) );
  XOR U594 ( .A(n405), .B(n406), .Z(n401) );
  ANDN U595 ( .B(n407), .A(n408), .Z(n406) );
  XOR U596 ( .A(clocal[105]), .B(n405), .Z(n407) );
  XNOR U597 ( .A(clocal[105]), .B(n408), .Z(swire[105]) );
  XNOR U598 ( .A(clocal[104]), .B(n410), .Z(swire[104]) );
  XNOR U599 ( .A(clocal[103]), .B(n412), .Z(swire[103]) );
  XOR U600 ( .A(n413), .B(n414), .Z(n411) );
  ANDN U601 ( .B(n415), .A(n416), .Z(n414) );
  XOR U602 ( .A(clocal[102]), .B(n413), .Z(n415) );
  XNOR U603 ( .A(clocal[102]), .B(n416), .Z(swire[102]) );
  XOR U604 ( .A(n417), .B(n418), .Z(n413) );
  ANDN U605 ( .B(n419), .A(n420), .Z(n418) );
  XOR U606 ( .A(clocal[101]), .B(n417), .Z(n419) );
  XNOR U607 ( .A(clocal[101]), .B(n420), .Z(swire[101]) );
  XNOR U608 ( .A(clocal[100]), .B(n422), .Z(swire[100]) );
  XOR U609 ( .A(n424), .B(n425), .Z(n423) );
  ANDN U610 ( .B(n426), .A(n252), .Z(n425) );
  XOR U611 ( .A(clocal[98]), .B(n424), .Z(n426) );
  XOR U612 ( .A(n427), .B(n428), .Z(n424) );
  ANDN U613 ( .B(n429), .A(n253), .Z(n428) );
  XOR U614 ( .A(clocal[97]), .B(n427), .Z(n429) );
  XOR U615 ( .A(n432), .B(n433), .Z(n431) );
  ANDN U616 ( .B(n434), .A(n256), .Z(n433) );
  XOR U617 ( .A(clocal[94]), .B(n432), .Z(n434) );
  XOR U618 ( .A(n435), .B(n436), .Z(n432) );
  ANDN U619 ( .B(n437), .A(n257), .Z(n436) );
  XOR U620 ( .A(clocal[93]), .B(n435), .Z(n437) );
  XOR U621 ( .A(n440), .B(n441), .Z(n439) );
  ANDN U622 ( .B(n442), .A(n260), .Z(n441) );
  XOR U623 ( .A(clocal[90]), .B(n440), .Z(n442) );
  XOR U624 ( .A(n443), .B(n444), .Z(n440) );
  ANDN U625 ( .B(n445), .A(n262), .Z(n444) );
  XOR U626 ( .A(clocal[89]), .B(n443), .Z(n445) );
  XOR U627 ( .A(n448), .B(n449), .Z(n447) );
  ANDN U628 ( .B(n450), .A(n265), .Z(n449) );
  XOR U629 ( .A(clocal[86]), .B(n448), .Z(n450) );
  XOR U630 ( .A(n451), .B(n452), .Z(n448) );
  ANDN U631 ( .B(n453), .A(n266), .Z(n452) );
  XOR U632 ( .A(clocal[85]), .B(n451), .Z(n453) );
  XOR U633 ( .A(n456), .B(n457), .Z(n455) );
  ANDN U634 ( .B(n458), .A(n269), .Z(n457) );
  XOR U635 ( .A(clocal[82]), .B(n456), .Z(n458) );
  XOR U636 ( .A(n459), .B(n460), .Z(n456) );
  ANDN U637 ( .B(n461), .A(n270), .Z(n460) );
  XOR U638 ( .A(clocal[81]), .B(n459), .Z(n461) );
  XOR U639 ( .A(n464), .B(n465), .Z(n463) );
  ANDN U640 ( .B(n466), .A(n274), .Z(n465) );
  XOR U641 ( .A(clocal[78]), .B(n464), .Z(n466) );
  XOR U642 ( .A(n467), .B(n468), .Z(n464) );
  ANDN U643 ( .B(n469), .A(n275), .Z(n468) );
  XOR U644 ( .A(clocal[77]), .B(n467), .Z(n469) );
  XOR U645 ( .A(n472), .B(n473), .Z(n471) );
  ANDN U646 ( .B(n474), .A(n278), .Z(n473) );
  XOR U647 ( .A(clocal[74]), .B(n472), .Z(n474) );
  XOR U648 ( .A(n475), .B(n476), .Z(n472) );
  ANDN U649 ( .B(n477), .A(n279), .Z(n476) );
  XOR U650 ( .A(clocal[73]), .B(n475), .Z(n477) );
  XOR U651 ( .A(n480), .B(n481), .Z(n479) );
  ANDN U652 ( .B(n482), .A(n282), .Z(n481) );
  XOR U653 ( .A(clocal[70]), .B(n480), .Z(n482) );
  XOR U654 ( .A(n483), .B(n484), .Z(n480) );
  ANDN U655 ( .B(n485), .A(n284), .Z(n484) );
  XOR U656 ( .A(clocal[69]), .B(n483), .Z(n485) );
  XOR U657 ( .A(n488), .B(n489), .Z(n487) );
  ANDN U658 ( .B(n490), .A(n287), .Z(n489) );
  XOR U659 ( .A(clocal[66]), .B(n488), .Z(n490) );
  XOR U660 ( .A(n491), .B(n492), .Z(n488) );
  ANDN U661 ( .B(n493), .A(n288), .Z(n492) );
  XOR U662 ( .A(clocal[65]), .B(n491), .Z(n493) );
  XOR U663 ( .A(n496), .B(n497), .Z(n495) );
  ANDN U664 ( .B(n498), .A(n291), .Z(n497) );
  XOR U665 ( .A(clocal[62]), .B(n496), .Z(n498) );
  XOR U666 ( .A(n499), .B(n500), .Z(n496) );
  ANDN U667 ( .B(n501), .A(n292), .Z(n500) );
  XOR U668 ( .A(clocal[61]), .B(n499), .Z(n501) );
  XOR U669 ( .A(n504), .B(n505), .Z(n503) );
  ANDN U670 ( .B(n506), .A(n296), .Z(n505) );
  XOR U671 ( .A(clocal[58]), .B(n504), .Z(n506) );
  XOR U672 ( .A(n507), .B(n508), .Z(n504) );
  ANDN U673 ( .B(n509), .A(n297), .Z(n508) );
  XOR U674 ( .A(clocal[57]), .B(n507), .Z(n509) );
  XOR U675 ( .A(n512), .B(n513), .Z(n511) );
  ANDN U676 ( .B(n514), .A(n300), .Z(n513) );
  XOR U677 ( .A(clocal[54]), .B(n512), .Z(n514) );
  XOR U678 ( .A(n515), .B(n516), .Z(n512) );
  ANDN U679 ( .B(n517), .A(n301), .Z(n516) );
  XOR U680 ( .A(clocal[53]), .B(n515), .Z(n517) );
  XOR U681 ( .A(n520), .B(n521), .Z(n519) );
  ANDN U682 ( .B(n522), .A(n304), .Z(n521) );
  XOR U683 ( .A(clocal[50]), .B(n520), .Z(n522) );
  XOR U684 ( .A(n523), .B(n524), .Z(n520) );
  ANDN U685 ( .B(n525), .A(n306), .Z(n524) );
  XOR U686 ( .A(clocal[49]), .B(n523), .Z(n525) );
  XOR U687 ( .A(n528), .B(n529), .Z(n527) );
  ANDN U688 ( .B(n530), .A(n309), .Z(n529) );
  XOR U689 ( .A(clocal[46]), .B(n528), .Z(n530) );
  XOR U690 ( .A(n531), .B(n532), .Z(n528) );
  ANDN U691 ( .B(n533), .A(n310), .Z(n532) );
  XOR U692 ( .A(clocal[45]), .B(n531), .Z(n533) );
  XOR U693 ( .A(n536), .B(n537), .Z(n535) );
  ANDN U694 ( .B(n538), .A(n313), .Z(n537) );
  XOR U695 ( .A(clocal[42]), .B(n536), .Z(n538) );
  XOR U696 ( .A(n539), .B(n540), .Z(n536) );
  ANDN U697 ( .B(n541), .A(n314), .Z(n540) );
  XOR U698 ( .A(clocal[41]), .B(n539), .Z(n541) );
  XOR U699 ( .A(n544), .B(n545), .Z(n543) );
  ANDN U700 ( .B(n546), .A(n317), .Z(n545) );
  XOR U701 ( .A(clocal[38]), .B(n544), .Z(n546) );
  XOR U702 ( .A(n547), .B(n548), .Z(n544) );
  ANDN U703 ( .B(n549), .A(n318), .Z(n548) );
  XOR U704 ( .A(clocal[37]), .B(n547), .Z(n549) );
  XOR U705 ( .A(n552), .B(n553), .Z(n551) );
  ANDN U706 ( .B(n554), .A(n321), .Z(n553) );
  XOR U707 ( .A(clocal[34]), .B(n552), .Z(n554) );
  XOR U708 ( .A(n555), .B(n556), .Z(n552) );
  ANDN U709 ( .B(n557), .A(n322), .Z(n556) );
  XOR U710 ( .A(clocal[33]), .B(n555), .Z(n557) );
  XOR U711 ( .A(n560), .B(n561), .Z(n559) );
  ANDN U712 ( .B(n562), .A(n325), .Z(n561) );
  XOR U713 ( .A(clocal[30]), .B(n560), .Z(n562) );
  XOR U714 ( .A(n563), .B(n564), .Z(n560) );
  ANDN U715 ( .B(n565), .A(n326), .Z(n564) );
  XOR U716 ( .A(clocal[29]), .B(n563), .Z(n565) );
  XOR U717 ( .A(n568), .B(n569), .Z(n567) );
  ANDN U718 ( .B(n570), .A(n329), .Z(n569) );
  XOR U719 ( .A(clocal[26]), .B(n568), .Z(n570) );
  XOR U720 ( .A(n571), .B(n572), .Z(n568) );
  ANDN U721 ( .B(n573), .A(n330), .Z(n572) );
  XOR U722 ( .A(clocal[25]), .B(n571), .Z(n573) );
  XOR U723 ( .A(n576), .B(n577), .Z(n575) );
  ANDN U724 ( .B(n578), .A(n333), .Z(n577) );
  XOR U725 ( .A(clocal[22]), .B(n576), .Z(n578) );
  XOR U726 ( .A(n579), .B(n580), .Z(n576) );
  ANDN U727 ( .B(n581), .A(n334), .Z(n580) );
  XOR U728 ( .A(clocal[21]), .B(n579), .Z(n581) );
  XOR U729 ( .A(n584), .B(n585), .Z(n583) );
  ANDN U730 ( .B(n586), .A(n337), .Z(n585) );
  XOR U731 ( .A(clocal[18]), .B(n584), .Z(n586) );
  XOR U732 ( .A(n587), .B(n588), .Z(n584) );
  ANDN U733 ( .B(n589), .A(n338), .Z(n588) );
  XOR U734 ( .A(clocal[17]), .B(n587), .Z(n589) );
  XOR U735 ( .A(n592), .B(n593), .Z(n591) );
  ANDN U736 ( .B(n594), .A(n341), .Z(n593) );
  XOR U737 ( .A(clocal[14]), .B(n592), .Z(n594) );
  XOR U738 ( .A(n595), .B(n596), .Z(n592) );
  ANDN U739 ( .B(n597), .A(n342), .Z(n596) );
  XOR U740 ( .A(clocal[13]), .B(n595), .Z(n597) );
  XOR U741 ( .A(n600), .B(n601), .Z(n599) );
  ANDN U742 ( .B(n602), .A(n396), .Z(n601) );
  XOR U743 ( .A(clocal[10]), .B(n600), .Z(n602) );
  XOR U744 ( .A(n603), .B(n604), .Z(n600) );
  ANDN U745 ( .B(n605), .A(n250), .Z(n604) );
  XOR U746 ( .A(clocal[9]), .B(n603), .Z(n605) );
  XOR U747 ( .A(n608), .B(n609), .Z(n607) );
  ANDN U748 ( .B(n610), .A(n283), .Z(n609) );
  XOR U749 ( .A(clocal[6]), .B(n608), .Z(n610) );
  XOR U750 ( .A(n611), .B(n612), .Z(n608) );
  ANDN U751 ( .B(n613), .A(n294), .Z(n612) );
  XOR U752 ( .A(clocal[5]), .B(n611), .Z(n613) );
  AND U753 ( .A(a[9]), .B(b[3]), .Z(\mult_44/ab[9][3] ) );
  AND U754 ( .A(a[9]), .B(b[2]), .Z(\mult_44/ab[9][2] ) );
  AND U755 ( .A(a[9]), .B(b[1]), .Z(\mult_44/ab[9][1] ) );
  AND U756 ( .A(b[0]), .B(a[9]), .Z(\mult_44/ab[9][0] ) );
  AND U757 ( .A(b[3]), .B(a[99]), .Z(\mult_44/ab[99][3] ) );
  AND U758 ( .A(b[2]), .B(a[99]), .Z(\mult_44/ab[99][2] ) );
  AND U759 ( .A(b[1]), .B(a[99]), .Z(\mult_44/ab[99][1] ) );
  AND U760 ( .A(a[99]), .B(b[0]), .Z(\mult_44/ab[99][0] ) );
  AND U761 ( .A(b[3]), .B(a[98]), .Z(\mult_44/ab[98][3] ) );
  AND U762 ( .A(b[2]), .B(a[98]), .Z(\mult_44/ab[98][2] ) );
  AND U763 ( .A(b[1]), .B(a[98]), .Z(\mult_44/ab[98][1] ) );
  AND U764 ( .A(a[98]), .B(b[0]), .Z(\mult_44/ab[98][0] ) );
  AND U765 ( .A(b[3]), .B(a[97]), .Z(\mult_44/ab[97][3] ) );
  AND U766 ( .A(b[2]), .B(a[97]), .Z(\mult_44/ab[97][2] ) );
  AND U767 ( .A(b[1]), .B(a[97]), .Z(\mult_44/ab[97][1] ) );
  AND U768 ( .A(a[97]), .B(b[0]), .Z(\mult_44/ab[97][0] ) );
  AND U769 ( .A(b[3]), .B(a[96]), .Z(\mult_44/ab[96][3] ) );
  AND U770 ( .A(b[2]), .B(a[96]), .Z(\mult_44/ab[96][2] ) );
  AND U771 ( .A(b[1]), .B(a[96]), .Z(\mult_44/ab[96][1] ) );
  AND U772 ( .A(a[96]), .B(b[0]), .Z(\mult_44/ab[96][0] ) );
  AND U773 ( .A(b[3]), .B(a[95]), .Z(\mult_44/ab[95][3] ) );
  AND U774 ( .A(b[2]), .B(a[95]), .Z(\mult_44/ab[95][2] ) );
  AND U775 ( .A(b[1]), .B(a[95]), .Z(\mult_44/ab[95][1] ) );
  AND U776 ( .A(a[95]), .B(b[0]), .Z(\mult_44/ab[95][0] ) );
  AND U777 ( .A(b[3]), .B(a[94]), .Z(\mult_44/ab[94][3] ) );
  AND U778 ( .A(b[2]), .B(a[94]), .Z(\mult_44/ab[94][2] ) );
  AND U779 ( .A(b[1]), .B(a[94]), .Z(\mult_44/ab[94][1] ) );
  AND U780 ( .A(a[94]), .B(b[0]), .Z(\mult_44/ab[94][0] ) );
  AND U781 ( .A(b[3]), .B(a[93]), .Z(\mult_44/ab[93][3] ) );
  AND U782 ( .A(b[2]), .B(a[93]), .Z(\mult_44/ab[93][2] ) );
  AND U783 ( .A(b[1]), .B(a[93]), .Z(\mult_44/ab[93][1] ) );
  AND U784 ( .A(a[93]), .B(b[0]), .Z(\mult_44/ab[93][0] ) );
  AND U785 ( .A(b[3]), .B(a[92]), .Z(\mult_44/ab[92][3] ) );
  AND U786 ( .A(b[2]), .B(a[92]), .Z(\mult_44/ab[92][2] ) );
  AND U787 ( .A(b[1]), .B(a[92]), .Z(\mult_44/ab[92][1] ) );
  AND U788 ( .A(a[92]), .B(b[0]), .Z(\mult_44/ab[92][0] ) );
  AND U789 ( .A(b[3]), .B(a[91]), .Z(\mult_44/ab[91][3] ) );
  AND U790 ( .A(b[2]), .B(a[91]), .Z(\mult_44/ab[91][2] ) );
  AND U791 ( .A(b[1]), .B(a[91]), .Z(\mult_44/ab[91][1] ) );
  AND U792 ( .A(a[91]), .B(b[0]), .Z(\mult_44/ab[91][0] ) );
  AND U793 ( .A(b[3]), .B(a[90]), .Z(\mult_44/ab[90][3] ) );
  AND U794 ( .A(b[2]), .B(a[90]), .Z(\mult_44/ab[90][2] ) );
  AND U795 ( .A(b[1]), .B(a[90]), .Z(\mult_44/ab[90][1] ) );
  AND U796 ( .A(a[90]), .B(b[0]), .Z(\mult_44/ab[90][0] ) );
  AND U797 ( .A(b[3]), .B(a[8]), .Z(\mult_44/ab[8][3] ) );
  AND U798 ( .A(b[2]), .B(a[8]), .Z(\mult_44/ab[8][2] ) );
  AND U799 ( .A(b[1]), .B(a[8]), .Z(\mult_44/ab[8][1] ) );
  AND U800 ( .A(a[8]), .B(b[0]), .Z(\mult_44/ab[8][0] ) );
  AND U801 ( .A(b[3]), .B(a[89]), .Z(\mult_44/ab[89][3] ) );
  AND U802 ( .A(b[2]), .B(a[89]), .Z(\mult_44/ab[89][2] ) );
  AND U803 ( .A(b[1]), .B(a[89]), .Z(\mult_44/ab[89][1] ) );
  AND U804 ( .A(a[89]), .B(b[0]), .Z(\mult_44/ab[89][0] ) );
  AND U805 ( .A(b[3]), .B(a[88]), .Z(\mult_44/ab[88][3] ) );
  AND U806 ( .A(b[2]), .B(a[88]), .Z(\mult_44/ab[88][2] ) );
  AND U807 ( .A(b[1]), .B(a[88]), .Z(\mult_44/ab[88][1] ) );
  AND U808 ( .A(a[88]), .B(b[0]), .Z(\mult_44/ab[88][0] ) );
  AND U809 ( .A(b[3]), .B(a[87]), .Z(\mult_44/ab[87][3] ) );
  AND U810 ( .A(b[2]), .B(a[87]), .Z(\mult_44/ab[87][2] ) );
  AND U811 ( .A(b[1]), .B(a[87]), .Z(\mult_44/ab[87][1] ) );
  AND U812 ( .A(a[87]), .B(b[0]), .Z(\mult_44/ab[87][0] ) );
  AND U813 ( .A(b[3]), .B(a[86]), .Z(\mult_44/ab[86][3] ) );
  AND U814 ( .A(b[2]), .B(a[86]), .Z(\mult_44/ab[86][2] ) );
  AND U815 ( .A(b[1]), .B(a[86]), .Z(\mult_44/ab[86][1] ) );
  AND U816 ( .A(a[86]), .B(b[0]), .Z(\mult_44/ab[86][0] ) );
  AND U817 ( .A(b[3]), .B(a[85]), .Z(\mult_44/ab[85][3] ) );
  AND U818 ( .A(b[2]), .B(a[85]), .Z(\mult_44/ab[85][2] ) );
  AND U819 ( .A(b[1]), .B(a[85]), .Z(\mult_44/ab[85][1] ) );
  AND U820 ( .A(a[85]), .B(b[0]), .Z(\mult_44/ab[85][0] ) );
  AND U821 ( .A(b[3]), .B(a[84]), .Z(\mult_44/ab[84][3] ) );
  AND U822 ( .A(b[2]), .B(a[84]), .Z(\mult_44/ab[84][2] ) );
  AND U823 ( .A(b[1]), .B(a[84]), .Z(\mult_44/ab[84][1] ) );
  AND U824 ( .A(a[84]), .B(b[0]), .Z(\mult_44/ab[84][0] ) );
  AND U825 ( .A(b[3]), .B(a[83]), .Z(\mult_44/ab[83][3] ) );
  AND U826 ( .A(b[2]), .B(a[83]), .Z(\mult_44/ab[83][2] ) );
  AND U827 ( .A(b[1]), .B(a[83]), .Z(\mult_44/ab[83][1] ) );
  AND U828 ( .A(a[83]), .B(b[0]), .Z(\mult_44/ab[83][0] ) );
  AND U829 ( .A(b[3]), .B(a[82]), .Z(\mult_44/ab[82][3] ) );
  AND U830 ( .A(b[2]), .B(a[82]), .Z(\mult_44/ab[82][2] ) );
  AND U831 ( .A(b[1]), .B(a[82]), .Z(\mult_44/ab[82][1] ) );
  AND U832 ( .A(a[82]), .B(b[0]), .Z(\mult_44/ab[82][0] ) );
  AND U833 ( .A(b[3]), .B(a[81]), .Z(\mult_44/ab[81][3] ) );
  AND U834 ( .A(b[2]), .B(a[81]), .Z(\mult_44/ab[81][2] ) );
  AND U835 ( .A(b[1]), .B(a[81]), .Z(\mult_44/ab[81][1] ) );
  AND U836 ( .A(a[81]), .B(b[0]), .Z(\mult_44/ab[81][0] ) );
  AND U837 ( .A(b[3]), .B(a[80]), .Z(\mult_44/ab[80][3] ) );
  AND U838 ( .A(b[2]), .B(a[80]), .Z(\mult_44/ab[80][2] ) );
  AND U839 ( .A(b[1]), .B(a[80]), .Z(\mult_44/ab[80][1] ) );
  AND U840 ( .A(a[80]), .B(b[0]), .Z(\mult_44/ab[80][0] ) );
  AND U841 ( .A(b[3]), .B(a[7]), .Z(\mult_44/ab[7][3] ) );
  AND U842 ( .A(b[2]), .B(a[7]), .Z(\mult_44/ab[7][2] ) );
  AND U843 ( .A(b[1]), .B(a[7]), .Z(\mult_44/ab[7][1] ) );
  AND U844 ( .A(a[7]), .B(b[0]), .Z(\mult_44/ab[7][0] ) );
  AND U845 ( .A(b[3]), .B(a[79]), .Z(\mult_44/ab[79][3] ) );
  AND U846 ( .A(b[2]), .B(a[79]), .Z(\mult_44/ab[79][2] ) );
  AND U847 ( .A(b[1]), .B(a[79]), .Z(\mult_44/ab[79][1] ) );
  AND U848 ( .A(a[79]), .B(b[0]), .Z(\mult_44/ab[79][0] ) );
  AND U849 ( .A(b[3]), .B(a[78]), .Z(\mult_44/ab[78][3] ) );
  AND U850 ( .A(b[2]), .B(a[78]), .Z(\mult_44/ab[78][2] ) );
  AND U851 ( .A(b[1]), .B(a[78]), .Z(\mult_44/ab[78][1] ) );
  AND U852 ( .A(a[78]), .B(b[0]), .Z(\mult_44/ab[78][0] ) );
  AND U853 ( .A(b[3]), .B(a[77]), .Z(\mult_44/ab[77][3] ) );
  AND U854 ( .A(b[2]), .B(a[77]), .Z(\mult_44/ab[77][2] ) );
  AND U855 ( .A(b[1]), .B(a[77]), .Z(\mult_44/ab[77][1] ) );
  AND U856 ( .A(a[77]), .B(b[0]), .Z(\mult_44/ab[77][0] ) );
  AND U857 ( .A(b[3]), .B(a[76]), .Z(\mult_44/ab[76][3] ) );
  AND U858 ( .A(b[2]), .B(a[76]), .Z(\mult_44/ab[76][2] ) );
  AND U859 ( .A(b[1]), .B(a[76]), .Z(\mult_44/ab[76][1] ) );
  AND U860 ( .A(a[76]), .B(b[0]), .Z(\mult_44/ab[76][0] ) );
  AND U861 ( .A(b[3]), .B(a[75]), .Z(\mult_44/ab[75][3] ) );
  AND U862 ( .A(b[2]), .B(a[75]), .Z(\mult_44/ab[75][2] ) );
  AND U863 ( .A(b[1]), .B(a[75]), .Z(\mult_44/ab[75][1] ) );
  AND U864 ( .A(a[75]), .B(b[0]), .Z(\mult_44/ab[75][0] ) );
  AND U865 ( .A(b[3]), .B(a[74]), .Z(\mult_44/ab[74][3] ) );
  AND U866 ( .A(b[2]), .B(a[74]), .Z(\mult_44/ab[74][2] ) );
  AND U867 ( .A(b[1]), .B(a[74]), .Z(\mult_44/ab[74][1] ) );
  AND U868 ( .A(a[74]), .B(b[0]), .Z(\mult_44/ab[74][0] ) );
  AND U869 ( .A(b[3]), .B(a[73]), .Z(\mult_44/ab[73][3] ) );
  AND U870 ( .A(b[2]), .B(a[73]), .Z(\mult_44/ab[73][2] ) );
  AND U871 ( .A(b[1]), .B(a[73]), .Z(\mult_44/ab[73][1] ) );
  AND U872 ( .A(a[73]), .B(b[0]), .Z(\mult_44/ab[73][0] ) );
  AND U873 ( .A(b[3]), .B(a[72]), .Z(\mult_44/ab[72][3] ) );
  AND U874 ( .A(b[2]), .B(a[72]), .Z(\mult_44/ab[72][2] ) );
  AND U875 ( .A(b[1]), .B(a[72]), .Z(\mult_44/ab[72][1] ) );
  AND U876 ( .A(a[72]), .B(b[0]), .Z(\mult_44/ab[72][0] ) );
  AND U877 ( .A(b[3]), .B(a[71]), .Z(\mult_44/ab[71][3] ) );
  AND U878 ( .A(b[2]), .B(a[71]), .Z(\mult_44/ab[71][2] ) );
  AND U879 ( .A(b[1]), .B(a[71]), .Z(\mult_44/ab[71][1] ) );
  AND U880 ( .A(a[71]), .B(b[0]), .Z(\mult_44/ab[71][0] ) );
  AND U881 ( .A(b[3]), .B(a[70]), .Z(\mult_44/ab[70][3] ) );
  AND U882 ( .A(b[2]), .B(a[70]), .Z(\mult_44/ab[70][2] ) );
  AND U883 ( .A(b[1]), .B(a[70]), .Z(\mult_44/ab[70][1] ) );
  AND U884 ( .A(a[70]), .B(b[0]), .Z(\mult_44/ab[70][0] ) );
  AND U885 ( .A(b[3]), .B(a[6]), .Z(\mult_44/ab[6][3] ) );
  AND U886 ( .A(b[2]), .B(a[6]), .Z(\mult_44/ab[6][2] ) );
  AND U887 ( .A(b[1]), .B(a[6]), .Z(\mult_44/ab[6][1] ) );
  AND U888 ( .A(a[6]), .B(b[0]), .Z(\mult_44/ab[6][0] ) );
  AND U889 ( .A(b[3]), .B(a[69]), .Z(\mult_44/ab[69][3] ) );
  AND U890 ( .A(b[2]), .B(a[69]), .Z(\mult_44/ab[69][2] ) );
  AND U891 ( .A(b[1]), .B(a[69]), .Z(\mult_44/ab[69][1] ) );
  AND U892 ( .A(a[69]), .B(b[0]), .Z(\mult_44/ab[69][0] ) );
  AND U893 ( .A(b[3]), .B(a[68]), .Z(\mult_44/ab[68][3] ) );
  AND U894 ( .A(b[2]), .B(a[68]), .Z(\mult_44/ab[68][2] ) );
  AND U895 ( .A(b[1]), .B(a[68]), .Z(\mult_44/ab[68][1] ) );
  AND U896 ( .A(a[68]), .B(b[0]), .Z(\mult_44/ab[68][0] ) );
  AND U897 ( .A(b[3]), .B(a[67]), .Z(\mult_44/ab[67][3] ) );
  AND U898 ( .A(b[2]), .B(a[67]), .Z(\mult_44/ab[67][2] ) );
  AND U899 ( .A(b[1]), .B(a[67]), .Z(\mult_44/ab[67][1] ) );
  AND U900 ( .A(a[67]), .B(b[0]), .Z(\mult_44/ab[67][0] ) );
  AND U901 ( .A(b[3]), .B(a[66]), .Z(\mult_44/ab[66][3] ) );
  AND U902 ( .A(b[2]), .B(a[66]), .Z(\mult_44/ab[66][2] ) );
  AND U903 ( .A(b[1]), .B(a[66]), .Z(\mult_44/ab[66][1] ) );
  AND U904 ( .A(a[66]), .B(b[0]), .Z(\mult_44/ab[66][0] ) );
  AND U905 ( .A(b[3]), .B(a[65]), .Z(\mult_44/ab[65][3] ) );
  AND U906 ( .A(b[2]), .B(a[65]), .Z(\mult_44/ab[65][2] ) );
  AND U907 ( .A(b[1]), .B(a[65]), .Z(\mult_44/ab[65][1] ) );
  AND U908 ( .A(a[65]), .B(b[0]), .Z(\mult_44/ab[65][0] ) );
  AND U909 ( .A(b[3]), .B(a[64]), .Z(\mult_44/ab[64][3] ) );
  AND U910 ( .A(b[2]), .B(a[64]), .Z(\mult_44/ab[64][2] ) );
  AND U911 ( .A(b[1]), .B(a[64]), .Z(\mult_44/ab[64][1] ) );
  AND U912 ( .A(a[64]), .B(b[0]), .Z(\mult_44/ab[64][0] ) );
  AND U913 ( .A(b[3]), .B(a[63]), .Z(\mult_44/ab[63][3] ) );
  AND U914 ( .A(b[2]), .B(a[63]), .Z(\mult_44/ab[63][2] ) );
  AND U915 ( .A(b[1]), .B(a[63]), .Z(\mult_44/ab[63][1] ) );
  AND U916 ( .A(a[63]), .B(b[0]), .Z(\mult_44/ab[63][0] ) );
  AND U917 ( .A(b[3]), .B(a[62]), .Z(\mult_44/ab[62][3] ) );
  AND U918 ( .A(b[2]), .B(a[62]), .Z(\mult_44/ab[62][2] ) );
  AND U919 ( .A(b[1]), .B(a[62]), .Z(\mult_44/ab[62][1] ) );
  AND U920 ( .A(a[62]), .B(b[0]), .Z(\mult_44/ab[62][0] ) );
  AND U921 ( .A(b[3]), .B(a[61]), .Z(\mult_44/ab[61][3] ) );
  AND U922 ( .A(b[2]), .B(a[61]), .Z(\mult_44/ab[61][2] ) );
  AND U923 ( .A(b[1]), .B(a[61]), .Z(\mult_44/ab[61][1] ) );
  AND U924 ( .A(a[61]), .B(b[0]), .Z(\mult_44/ab[61][0] ) );
  AND U925 ( .A(b[3]), .B(a[60]), .Z(\mult_44/ab[60][3] ) );
  AND U926 ( .A(b[2]), .B(a[60]), .Z(\mult_44/ab[60][2] ) );
  AND U927 ( .A(b[1]), .B(a[60]), .Z(\mult_44/ab[60][1] ) );
  AND U928 ( .A(a[60]), .B(b[0]), .Z(\mult_44/ab[60][0] ) );
  AND U929 ( .A(b[3]), .B(a[5]), .Z(\mult_44/ab[5][3] ) );
  AND U930 ( .A(b[2]), .B(a[5]), .Z(\mult_44/ab[5][2] ) );
  AND U931 ( .A(b[1]), .B(a[5]), .Z(\mult_44/ab[5][1] ) );
  AND U932 ( .A(a[5]), .B(b[0]), .Z(\mult_44/ab[5][0] ) );
  AND U933 ( .A(b[3]), .B(a[59]), .Z(\mult_44/ab[59][3] ) );
  AND U934 ( .A(b[2]), .B(a[59]), .Z(\mult_44/ab[59][2] ) );
  AND U935 ( .A(b[1]), .B(a[59]), .Z(\mult_44/ab[59][1] ) );
  AND U936 ( .A(a[59]), .B(b[0]), .Z(\mult_44/ab[59][0] ) );
  AND U937 ( .A(b[3]), .B(a[58]), .Z(\mult_44/ab[58][3] ) );
  AND U938 ( .A(b[2]), .B(a[58]), .Z(\mult_44/ab[58][2] ) );
  AND U939 ( .A(b[1]), .B(a[58]), .Z(\mult_44/ab[58][1] ) );
  AND U940 ( .A(a[58]), .B(b[0]), .Z(\mult_44/ab[58][0] ) );
  AND U941 ( .A(b[3]), .B(a[57]), .Z(\mult_44/ab[57][3] ) );
  AND U942 ( .A(b[2]), .B(a[57]), .Z(\mult_44/ab[57][2] ) );
  AND U943 ( .A(b[1]), .B(a[57]), .Z(\mult_44/ab[57][1] ) );
  AND U944 ( .A(a[57]), .B(b[0]), .Z(\mult_44/ab[57][0] ) );
  AND U945 ( .A(b[3]), .B(a[56]), .Z(\mult_44/ab[56][3] ) );
  AND U946 ( .A(b[2]), .B(a[56]), .Z(\mult_44/ab[56][2] ) );
  AND U947 ( .A(b[1]), .B(a[56]), .Z(\mult_44/ab[56][1] ) );
  AND U948 ( .A(a[56]), .B(b[0]), .Z(\mult_44/ab[56][0] ) );
  AND U949 ( .A(b[3]), .B(a[55]), .Z(\mult_44/ab[55][3] ) );
  AND U950 ( .A(b[2]), .B(a[55]), .Z(\mult_44/ab[55][2] ) );
  AND U951 ( .A(b[1]), .B(a[55]), .Z(\mult_44/ab[55][1] ) );
  AND U952 ( .A(a[55]), .B(b[0]), .Z(\mult_44/ab[55][0] ) );
  AND U953 ( .A(b[3]), .B(a[54]), .Z(\mult_44/ab[54][3] ) );
  AND U954 ( .A(b[2]), .B(a[54]), .Z(\mult_44/ab[54][2] ) );
  AND U955 ( .A(b[1]), .B(a[54]), .Z(\mult_44/ab[54][1] ) );
  AND U956 ( .A(a[54]), .B(b[0]), .Z(\mult_44/ab[54][0] ) );
  AND U957 ( .A(b[3]), .B(a[53]), .Z(\mult_44/ab[53][3] ) );
  AND U958 ( .A(b[2]), .B(a[53]), .Z(\mult_44/ab[53][2] ) );
  AND U959 ( .A(b[1]), .B(a[53]), .Z(\mult_44/ab[53][1] ) );
  AND U960 ( .A(a[53]), .B(b[0]), .Z(\mult_44/ab[53][0] ) );
  AND U961 ( .A(b[3]), .B(a[52]), .Z(\mult_44/ab[52][3] ) );
  AND U962 ( .A(b[2]), .B(a[52]), .Z(\mult_44/ab[52][2] ) );
  AND U963 ( .A(b[1]), .B(a[52]), .Z(\mult_44/ab[52][1] ) );
  AND U964 ( .A(a[52]), .B(b[0]), .Z(\mult_44/ab[52][0] ) );
  AND U965 ( .A(b[3]), .B(a[51]), .Z(\mult_44/ab[51][3] ) );
  AND U966 ( .A(b[2]), .B(a[51]), .Z(\mult_44/ab[51][2] ) );
  AND U967 ( .A(b[1]), .B(a[51]), .Z(\mult_44/ab[51][1] ) );
  AND U968 ( .A(a[51]), .B(b[0]), .Z(\mult_44/ab[51][0] ) );
  AND U969 ( .A(b[3]), .B(a[50]), .Z(\mult_44/ab[50][3] ) );
  AND U970 ( .A(b[2]), .B(a[50]), .Z(\mult_44/ab[50][2] ) );
  AND U971 ( .A(b[1]), .B(a[50]), .Z(\mult_44/ab[50][1] ) );
  AND U972 ( .A(a[50]), .B(b[0]), .Z(\mult_44/ab[50][0] ) );
  AND U973 ( .A(b[3]), .B(a[4]), .Z(\mult_44/ab[4][3] ) );
  AND U974 ( .A(b[2]), .B(a[4]), .Z(\mult_44/ab[4][2] ) );
  AND U975 ( .A(b[1]), .B(a[4]), .Z(\mult_44/ab[4][1] ) );
  AND U976 ( .A(a[4]), .B(b[0]), .Z(\mult_44/ab[4][0] ) );
  AND U977 ( .A(b[3]), .B(a[49]), .Z(\mult_44/ab[49][3] ) );
  AND U978 ( .A(b[2]), .B(a[49]), .Z(\mult_44/ab[49][2] ) );
  AND U979 ( .A(b[1]), .B(a[49]), .Z(\mult_44/ab[49][1] ) );
  AND U980 ( .A(a[49]), .B(b[0]), .Z(\mult_44/ab[49][0] ) );
  AND U981 ( .A(b[3]), .B(a[48]), .Z(\mult_44/ab[48][3] ) );
  AND U982 ( .A(b[2]), .B(a[48]), .Z(\mult_44/ab[48][2] ) );
  AND U983 ( .A(b[1]), .B(a[48]), .Z(\mult_44/ab[48][1] ) );
  AND U984 ( .A(a[48]), .B(b[0]), .Z(\mult_44/ab[48][0] ) );
  AND U985 ( .A(b[3]), .B(a[47]), .Z(\mult_44/ab[47][3] ) );
  AND U986 ( .A(b[2]), .B(a[47]), .Z(\mult_44/ab[47][2] ) );
  AND U987 ( .A(b[1]), .B(a[47]), .Z(\mult_44/ab[47][1] ) );
  AND U988 ( .A(a[47]), .B(b[0]), .Z(\mult_44/ab[47][0] ) );
  AND U989 ( .A(b[3]), .B(a[46]), .Z(\mult_44/ab[46][3] ) );
  AND U990 ( .A(b[2]), .B(a[46]), .Z(\mult_44/ab[46][2] ) );
  AND U991 ( .A(b[1]), .B(a[46]), .Z(\mult_44/ab[46][1] ) );
  AND U992 ( .A(a[46]), .B(b[0]), .Z(\mult_44/ab[46][0] ) );
  AND U993 ( .A(b[3]), .B(a[45]), .Z(\mult_44/ab[45][3] ) );
  AND U994 ( .A(b[2]), .B(a[45]), .Z(\mult_44/ab[45][2] ) );
  AND U995 ( .A(b[1]), .B(a[45]), .Z(\mult_44/ab[45][1] ) );
  AND U996 ( .A(a[45]), .B(b[0]), .Z(\mult_44/ab[45][0] ) );
  AND U997 ( .A(b[3]), .B(a[44]), .Z(\mult_44/ab[44][3] ) );
  AND U998 ( .A(b[2]), .B(a[44]), .Z(\mult_44/ab[44][2] ) );
  AND U999 ( .A(b[1]), .B(a[44]), .Z(\mult_44/ab[44][1] ) );
  AND U1000 ( .A(a[44]), .B(b[0]), .Z(\mult_44/ab[44][0] ) );
  AND U1001 ( .A(b[3]), .B(a[43]), .Z(\mult_44/ab[43][3] ) );
  AND U1002 ( .A(b[2]), .B(a[43]), .Z(\mult_44/ab[43][2] ) );
  AND U1003 ( .A(b[1]), .B(a[43]), .Z(\mult_44/ab[43][1] ) );
  AND U1004 ( .A(a[43]), .B(b[0]), .Z(\mult_44/ab[43][0] ) );
  AND U1005 ( .A(b[3]), .B(a[42]), .Z(\mult_44/ab[42][3] ) );
  AND U1006 ( .A(b[2]), .B(a[42]), .Z(\mult_44/ab[42][2] ) );
  AND U1007 ( .A(b[1]), .B(a[42]), .Z(\mult_44/ab[42][1] ) );
  AND U1008 ( .A(a[42]), .B(b[0]), .Z(\mult_44/ab[42][0] ) );
  AND U1009 ( .A(b[3]), .B(a[41]), .Z(\mult_44/ab[41][3] ) );
  AND U1010 ( .A(b[2]), .B(a[41]), .Z(\mult_44/ab[41][2] ) );
  AND U1011 ( .A(b[1]), .B(a[41]), .Z(\mult_44/ab[41][1] ) );
  AND U1012 ( .A(a[41]), .B(b[0]), .Z(\mult_44/ab[41][0] ) );
  AND U1013 ( .A(b[3]), .B(a[40]), .Z(\mult_44/ab[40][3] ) );
  AND U1014 ( .A(b[2]), .B(a[40]), .Z(\mult_44/ab[40][2] ) );
  AND U1015 ( .A(b[1]), .B(a[40]), .Z(\mult_44/ab[40][1] ) );
  AND U1016 ( .A(a[40]), .B(b[0]), .Z(\mult_44/ab[40][0] ) );
  AND U1017 ( .A(b[3]), .B(a[3]), .Z(\mult_44/ab[3][3] ) );
  AND U1018 ( .A(b[2]), .B(a[3]), .Z(\mult_44/ab[3][2] ) );
  AND U1019 ( .A(b[1]), .B(a[3]), .Z(\mult_44/ab[3][1] ) );
  AND U1020 ( .A(a[3]), .B(b[0]), .Z(\mult_44/ab[3][0] ) );
  AND U1021 ( .A(b[3]), .B(a[39]), .Z(\mult_44/ab[39][3] ) );
  AND U1022 ( .A(b[2]), .B(a[39]), .Z(\mult_44/ab[39][2] ) );
  AND U1023 ( .A(b[1]), .B(a[39]), .Z(\mult_44/ab[39][1] ) );
  AND U1024 ( .A(a[39]), .B(b[0]), .Z(\mult_44/ab[39][0] ) );
  AND U1025 ( .A(b[3]), .B(a[38]), .Z(\mult_44/ab[38][3] ) );
  AND U1026 ( .A(b[2]), .B(a[38]), .Z(\mult_44/ab[38][2] ) );
  AND U1027 ( .A(b[1]), .B(a[38]), .Z(\mult_44/ab[38][1] ) );
  AND U1028 ( .A(a[38]), .B(b[0]), .Z(\mult_44/ab[38][0] ) );
  AND U1029 ( .A(b[3]), .B(a[37]), .Z(\mult_44/ab[37][3] ) );
  AND U1030 ( .A(b[2]), .B(a[37]), .Z(\mult_44/ab[37][2] ) );
  AND U1031 ( .A(b[1]), .B(a[37]), .Z(\mult_44/ab[37][1] ) );
  AND U1032 ( .A(a[37]), .B(b[0]), .Z(\mult_44/ab[37][0] ) );
  AND U1033 ( .A(b[3]), .B(a[36]), .Z(\mult_44/ab[36][3] ) );
  AND U1034 ( .A(b[2]), .B(a[36]), .Z(\mult_44/ab[36][2] ) );
  AND U1035 ( .A(b[1]), .B(a[36]), .Z(\mult_44/ab[36][1] ) );
  AND U1036 ( .A(a[36]), .B(b[0]), .Z(\mult_44/ab[36][0] ) );
  AND U1037 ( .A(b[3]), .B(a[35]), .Z(\mult_44/ab[35][3] ) );
  AND U1038 ( .A(b[2]), .B(a[35]), .Z(\mult_44/ab[35][2] ) );
  AND U1039 ( .A(b[1]), .B(a[35]), .Z(\mult_44/ab[35][1] ) );
  AND U1040 ( .A(a[35]), .B(b[0]), .Z(\mult_44/ab[35][0] ) );
  AND U1041 ( .A(b[3]), .B(a[34]), .Z(\mult_44/ab[34][3] ) );
  AND U1042 ( .A(b[2]), .B(a[34]), .Z(\mult_44/ab[34][2] ) );
  AND U1043 ( .A(b[1]), .B(a[34]), .Z(\mult_44/ab[34][1] ) );
  AND U1044 ( .A(a[34]), .B(b[0]), .Z(\mult_44/ab[34][0] ) );
  AND U1045 ( .A(b[3]), .B(a[33]), .Z(\mult_44/ab[33][3] ) );
  AND U1046 ( .A(b[2]), .B(a[33]), .Z(\mult_44/ab[33][2] ) );
  AND U1047 ( .A(b[1]), .B(a[33]), .Z(\mult_44/ab[33][1] ) );
  AND U1048 ( .A(a[33]), .B(b[0]), .Z(\mult_44/ab[33][0] ) );
  AND U1049 ( .A(b[3]), .B(a[32]), .Z(\mult_44/ab[32][3] ) );
  AND U1050 ( .A(b[2]), .B(a[32]), .Z(\mult_44/ab[32][2] ) );
  AND U1051 ( .A(b[1]), .B(a[32]), .Z(\mult_44/ab[32][1] ) );
  AND U1052 ( .A(a[32]), .B(b[0]), .Z(\mult_44/ab[32][0] ) );
  AND U1053 ( .A(b[3]), .B(a[31]), .Z(\mult_44/ab[31][3] ) );
  AND U1054 ( .A(b[2]), .B(a[31]), .Z(\mult_44/ab[31][2] ) );
  AND U1055 ( .A(b[1]), .B(a[31]), .Z(\mult_44/ab[31][1] ) );
  AND U1056 ( .A(a[31]), .B(b[0]), .Z(\mult_44/ab[31][0] ) );
  AND U1057 ( .A(b[3]), .B(a[30]), .Z(\mult_44/ab[30][3] ) );
  AND U1058 ( .A(b[2]), .B(a[30]), .Z(\mult_44/ab[30][2] ) );
  AND U1059 ( .A(b[1]), .B(a[30]), .Z(\mult_44/ab[30][1] ) );
  AND U1060 ( .A(a[30]), .B(b[0]), .Z(\mult_44/ab[30][0] ) );
  AND U1061 ( .A(b[3]), .B(a[2]), .Z(\mult_44/ab[2][3] ) );
  AND U1062 ( .A(b[2]), .B(a[2]), .Z(\mult_44/ab[2][2] ) );
  AND U1063 ( .A(b[1]), .B(a[2]), .Z(\mult_44/ab[2][1] ) );
  AND U1064 ( .A(a[2]), .B(b[0]), .Z(\mult_44/ab[2][0] ) );
  AND U1065 ( .A(b[3]), .B(a[29]), .Z(\mult_44/ab[29][3] ) );
  AND U1066 ( .A(b[2]), .B(a[29]), .Z(\mult_44/ab[29][2] ) );
  AND U1067 ( .A(b[1]), .B(a[29]), .Z(\mult_44/ab[29][1] ) );
  AND U1068 ( .A(a[29]), .B(b[0]), .Z(\mult_44/ab[29][0] ) );
  AND U1069 ( .A(b[3]), .B(a[28]), .Z(\mult_44/ab[28][3] ) );
  AND U1070 ( .A(b[2]), .B(a[28]), .Z(\mult_44/ab[28][2] ) );
  AND U1071 ( .A(b[1]), .B(a[28]), .Z(\mult_44/ab[28][1] ) );
  AND U1072 ( .A(a[28]), .B(b[0]), .Z(\mult_44/ab[28][0] ) );
  AND U1073 ( .A(b[3]), .B(a[27]), .Z(\mult_44/ab[27][3] ) );
  AND U1074 ( .A(b[2]), .B(a[27]), .Z(\mult_44/ab[27][2] ) );
  AND U1075 ( .A(b[1]), .B(a[27]), .Z(\mult_44/ab[27][1] ) );
  AND U1076 ( .A(a[27]), .B(b[0]), .Z(\mult_44/ab[27][0] ) );
  AND U1077 ( .A(b[3]), .B(a[26]), .Z(\mult_44/ab[26][3] ) );
  AND U1078 ( .A(b[2]), .B(a[26]), .Z(\mult_44/ab[26][2] ) );
  AND U1079 ( .A(b[1]), .B(a[26]), .Z(\mult_44/ab[26][1] ) );
  AND U1080 ( .A(a[26]), .B(b[0]), .Z(\mult_44/ab[26][0] ) );
  AND U1081 ( .A(b[3]), .B(a[25]), .Z(\mult_44/ab[25][3] ) );
  AND U1082 ( .A(b[2]), .B(a[25]), .Z(\mult_44/ab[25][2] ) );
  AND U1083 ( .A(b[1]), .B(a[25]), .Z(\mult_44/ab[25][1] ) );
  AND U1084 ( .A(a[25]), .B(b[0]), .Z(\mult_44/ab[25][0] ) );
  AND U1085 ( .A(b[3]), .B(a[24]), .Z(\mult_44/ab[24][3] ) );
  AND U1086 ( .A(b[2]), .B(a[24]), .Z(\mult_44/ab[24][2] ) );
  AND U1087 ( .A(b[1]), .B(a[24]), .Z(\mult_44/ab[24][1] ) );
  AND U1088 ( .A(a[24]), .B(b[0]), .Z(\mult_44/ab[24][0] ) );
  AND U1089 ( .A(b[3]), .B(a[23]), .Z(\mult_44/ab[23][3] ) );
  AND U1090 ( .A(b[2]), .B(a[23]), .Z(\mult_44/ab[23][2] ) );
  AND U1091 ( .A(b[1]), .B(a[23]), .Z(\mult_44/ab[23][1] ) );
  AND U1092 ( .A(a[23]), .B(b[0]), .Z(\mult_44/ab[23][0] ) );
  AND U1093 ( .A(b[3]), .B(a[22]), .Z(\mult_44/ab[22][3] ) );
  AND U1094 ( .A(b[2]), .B(a[22]), .Z(\mult_44/ab[22][2] ) );
  AND U1095 ( .A(b[1]), .B(a[22]), .Z(\mult_44/ab[22][1] ) );
  AND U1096 ( .A(a[22]), .B(b[0]), .Z(\mult_44/ab[22][0] ) );
  AND U1097 ( .A(b[3]), .B(a[21]), .Z(\mult_44/ab[21][3] ) );
  AND U1098 ( .A(b[2]), .B(a[21]), .Z(\mult_44/ab[21][2] ) );
  AND U1099 ( .A(b[1]), .B(a[21]), .Z(\mult_44/ab[21][1] ) );
  AND U1100 ( .A(a[21]), .B(b[0]), .Z(\mult_44/ab[21][0] ) );
  AND U1101 ( .A(b[3]), .B(a[20]), .Z(\mult_44/ab[20][3] ) );
  AND U1102 ( .A(b[2]), .B(a[20]), .Z(\mult_44/ab[20][2] ) );
  AND U1103 ( .A(b[1]), .B(a[20]), .Z(\mult_44/ab[20][1] ) );
  AND U1104 ( .A(a[20]), .B(b[0]), .Z(\mult_44/ab[20][0] ) );
  AND U1105 ( .A(b[3]), .B(a[1]), .Z(\mult_44/ab[1][3] ) );
  AND U1106 ( .A(b[2]), .B(a[1]), .Z(\mult_44/ab[1][2] ) );
  AND U1107 ( .A(b[1]), .B(a[1]), .Z(\mult_44/ab[1][1] ) );
  AND U1108 ( .A(a[1]), .B(b[0]), .Z(\mult_44/ab[1][0] ) );
  AND U1109 ( .A(b[3]), .B(a[19]), .Z(\mult_44/ab[19][3] ) );
  AND U1110 ( .A(b[2]), .B(a[19]), .Z(\mult_44/ab[19][2] ) );
  AND U1111 ( .A(b[1]), .B(a[19]), .Z(\mult_44/ab[19][1] ) );
  AND U1112 ( .A(a[19]), .B(b[0]), .Z(\mult_44/ab[19][0] ) );
  AND U1113 ( .A(b[3]), .B(a[18]), .Z(\mult_44/ab[18][3] ) );
  AND U1114 ( .A(b[2]), .B(a[18]), .Z(\mult_44/ab[18][2] ) );
  AND U1115 ( .A(b[1]), .B(a[18]), .Z(\mult_44/ab[18][1] ) );
  AND U1116 ( .A(a[18]), .B(b[0]), .Z(\mult_44/ab[18][0] ) );
  AND U1117 ( .A(b[3]), .B(a[17]), .Z(\mult_44/ab[17][3] ) );
  AND U1118 ( .A(b[2]), .B(a[17]), .Z(\mult_44/ab[17][2] ) );
  AND U1119 ( .A(b[1]), .B(a[17]), .Z(\mult_44/ab[17][1] ) );
  AND U1120 ( .A(a[17]), .B(b[0]), .Z(\mult_44/ab[17][0] ) );
  AND U1121 ( .A(b[3]), .B(a[16]), .Z(\mult_44/ab[16][3] ) );
  AND U1122 ( .A(b[2]), .B(a[16]), .Z(\mult_44/ab[16][2] ) );
  AND U1123 ( .A(b[1]), .B(a[16]), .Z(\mult_44/ab[16][1] ) );
  AND U1124 ( .A(a[16]), .B(b[0]), .Z(\mult_44/ab[16][0] ) );
  AND U1125 ( .A(b[3]), .B(a[15]), .Z(\mult_44/ab[15][3] ) );
  AND U1126 ( .A(b[2]), .B(a[15]), .Z(\mult_44/ab[15][2] ) );
  AND U1127 ( .A(b[1]), .B(a[15]), .Z(\mult_44/ab[15][1] ) );
  AND U1128 ( .A(a[15]), .B(b[0]), .Z(\mult_44/ab[15][0] ) );
  AND U1129 ( .A(b[3]), .B(a[14]), .Z(\mult_44/ab[14][3] ) );
  AND U1130 ( .A(b[2]), .B(a[14]), .Z(\mult_44/ab[14][2] ) );
  AND U1131 ( .A(b[1]), .B(a[14]), .Z(\mult_44/ab[14][1] ) );
  AND U1132 ( .A(a[14]), .B(b[0]), .Z(\mult_44/ab[14][0] ) );
  AND U1133 ( .A(b[3]), .B(a[13]), .Z(\mult_44/ab[13][3] ) );
  AND U1134 ( .A(b[2]), .B(a[13]), .Z(\mult_44/ab[13][2] ) );
  AND U1135 ( .A(b[1]), .B(a[13]), .Z(\mult_44/ab[13][1] ) );
  AND U1136 ( .A(a[13]), .B(b[0]), .Z(\mult_44/ab[13][0] ) );
  AND U1137 ( .A(b[3]), .B(a[12]), .Z(\mult_44/ab[12][3] ) );
  AND U1138 ( .A(b[2]), .B(a[12]), .Z(\mult_44/ab[12][2] ) );
  AND U1139 ( .A(b[1]), .B(a[12]), .Z(\mult_44/ab[12][1] ) );
  AND U1140 ( .A(a[12]), .B(b[0]), .Z(\mult_44/ab[12][0] ) );
  AND U1141 ( .A(a[127]), .B(b[0]), .Z(\mult_44/ab[127][0] ) );
  AND U1142 ( .A(b[1]), .B(a[126]), .Z(\mult_44/ab[126][1] ) );
  AND U1143 ( .A(a[126]), .B(b[0]), .Z(\mult_44/ab[126][0] ) );
  AND U1144 ( .A(b[2]), .B(a[125]), .Z(\mult_44/ab[125][2] ) );
  AND U1145 ( .A(b[1]), .B(a[125]), .Z(\mult_44/ab[125][1] ) );
  AND U1146 ( .A(a[125]), .B(b[0]), .Z(\mult_44/ab[125][0] ) );
  AND U1147 ( .A(b[3]), .B(a[124]), .Z(\mult_44/ab[124][3] ) );
  AND U1148 ( .A(b[2]), .B(a[124]), .Z(\mult_44/ab[124][2] ) );
  AND U1149 ( .A(b[1]), .B(a[124]), .Z(\mult_44/ab[124][1] ) );
  AND U1150 ( .A(a[124]), .B(b[0]), .Z(\mult_44/ab[124][0] ) );
  AND U1151 ( .A(b[3]), .B(a[123]), .Z(\mult_44/ab[123][3] ) );
  AND U1152 ( .A(b[2]), .B(a[123]), .Z(\mult_44/ab[123][2] ) );
  AND U1153 ( .A(b[1]), .B(a[123]), .Z(\mult_44/ab[123][1] ) );
  AND U1154 ( .A(a[123]), .B(b[0]), .Z(\mult_44/ab[123][0] ) );
  AND U1155 ( .A(b[3]), .B(a[122]), .Z(\mult_44/ab[122][3] ) );
  AND U1156 ( .A(b[2]), .B(a[122]), .Z(\mult_44/ab[122][2] ) );
  AND U1157 ( .A(b[1]), .B(a[122]), .Z(\mult_44/ab[122][1] ) );
  AND U1158 ( .A(a[122]), .B(b[0]), .Z(\mult_44/ab[122][0] ) );
  AND U1159 ( .A(b[3]), .B(a[121]), .Z(\mult_44/ab[121][3] ) );
  AND U1160 ( .A(b[2]), .B(a[121]), .Z(\mult_44/ab[121][2] ) );
  AND U1161 ( .A(b[1]), .B(a[121]), .Z(\mult_44/ab[121][1] ) );
  AND U1162 ( .A(a[121]), .B(b[0]), .Z(\mult_44/ab[121][0] ) );
  AND U1163 ( .A(b[3]), .B(a[120]), .Z(\mult_44/ab[120][3] ) );
  AND U1164 ( .A(b[2]), .B(a[120]), .Z(\mult_44/ab[120][2] ) );
  AND U1165 ( .A(b[1]), .B(a[120]), .Z(\mult_44/ab[120][1] ) );
  AND U1166 ( .A(a[120]), .B(b[0]), .Z(\mult_44/ab[120][0] ) );
  AND U1167 ( .A(b[3]), .B(a[11]), .Z(\mult_44/ab[11][3] ) );
  AND U1168 ( .A(b[2]), .B(a[11]), .Z(\mult_44/ab[11][2] ) );
  AND U1169 ( .A(b[1]), .B(a[11]), .Z(\mult_44/ab[11][1] ) );
  AND U1170 ( .A(a[11]), .B(b[0]), .Z(\mult_44/ab[11][0] ) );
  AND U1171 ( .A(b[3]), .B(a[119]), .Z(\mult_44/ab[119][3] ) );
  AND U1172 ( .A(b[2]), .B(a[119]), .Z(\mult_44/ab[119][2] ) );
  AND U1173 ( .A(b[1]), .B(a[119]), .Z(\mult_44/ab[119][1] ) );
  AND U1174 ( .A(a[119]), .B(b[0]), .Z(\mult_44/ab[119][0] ) );
  AND U1175 ( .A(b[3]), .B(a[118]), .Z(\mult_44/ab[118][3] ) );
  AND U1176 ( .A(b[2]), .B(a[118]), .Z(\mult_44/ab[118][2] ) );
  AND U1177 ( .A(b[1]), .B(a[118]), .Z(\mult_44/ab[118][1] ) );
  AND U1178 ( .A(a[118]), .B(b[0]), .Z(\mult_44/ab[118][0] ) );
  AND U1179 ( .A(b[3]), .B(a[117]), .Z(\mult_44/ab[117][3] ) );
  AND U1180 ( .A(b[2]), .B(a[117]), .Z(\mult_44/ab[117][2] ) );
  AND U1181 ( .A(b[1]), .B(a[117]), .Z(\mult_44/ab[117][1] ) );
  AND U1182 ( .A(a[117]), .B(b[0]), .Z(\mult_44/ab[117][0] ) );
  AND U1183 ( .A(b[3]), .B(a[116]), .Z(\mult_44/ab[116][3] ) );
  AND U1184 ( .A(b[2]), .B(a[116]), .Z(\mult_44/ab[116][2] ) );
  AND U1185 ( .A(b[1]), .B(a[116]), .Z(\mult_44/ab[116][1] ) );
  AND U1186 ( .A(a[116]), .B(b[0]), .Z(\mult_44/ab[116][0] ) );
  AND U1187 ( .A(b[3]), .B(a[115]), .Z(\mult_44/ab[115][3] ) );
  AND U1188 ( .A(b[2]), .B(a[115]), .Z(\mult_44/ab[115][2] ) );
  AND U1189 ( .A(b[1]), .B(a[115]), .Z(\mult_44/ab[115][1] ) );
  AND U1190 ( .A(a[115]), .B(b[0]), .Z(\mult_44/ab[115][0] ) );
  AND U1191 ( .A(b[3]), .B(a[114]), .Z(\mult_44/ab[114][3] ) );
  AND U1192 ( .A(b[2]), .B(a[114]), .Z(\mult_44/ab[114][2] ) );
  AND U1193 ( .A(b[1]), .B(a[114]), .Z(\mult_44/ab[114][1] ) );
  AND U1194 ( .A(a[114]), .B(b[0]), .Z(\mult_44/ab[114][0] ) );
  AND U1195 ( .A(b[3]), .B(a[113]), .Z(\mult_44/ab[113][3] ) );
  AND U1196 ( .A(b[2]), .B(a[113]), .Z(\mult_44/ab[113][2] ) );
  AND U1197 ( .A(b[1]), .B(a[113]), .Z(\mult_44/ab[113][1] ) );
  AND U1198 ( .A(a[113]), .B(b[0]), .Z(\mult_44/ab[113][0] ) );
  AND U1199 ( .A(b[3]), .B(a[112]), .Z(\mult_44/ab[112][3] ) );
  AND U1200 ( .A(b[2]), .B(a[112]), .Z(\mult_44/ab[112][2] ) );
  AND U1201 ( .A(b[1]), .B(a[112]), .Z(\mult_44/ab[112][1] ) );
  AND U1202 ( .A(a[112]), .B(b[0]), .Z(\mult_44/ab[112][0] ) );
  AND U1203 ( .A(b[3]), .B(a[111]), .Z(\mult_44/ab[111][3] ) );
  AND U1204 ( .A(b[2]), .B(a[111]), .Z(\mult_44/ab[111][2] ) );
  AND U1205 ( .A(b[1]), .B(a[111]), .Z(\mult_44/ab[111][1] ) );
  AND U1206 ( .A(a[111]), .B(b[0]), .Z(\mult_44/ab[111][0] ) );
  AND U1207 ( .A(b[3]), .B(a[110]), .Z(\mult_44/ab[110][3] ) );
  AND U1208 ( .A(b[2]), .B(a[110]), .Z(\mult_44/ab[110][2] ) );
  AND U1209 ( .A(b[1]), .B(a[110]), .Z(\mult_44/ab[110][1] ) );
  AND U1210 ( .A(a[110]), .B(b[0]), .Z(\mult_44/ab[110][0] ) );
  AND U1211 ( .A(b[3]), .B(a[10]), .Z(\mult_44/ab[10][3] ) );
  AND U1212 ( .A(b[2]), .B(a[10]), .Z(\mult_44/ab[10][2] ) );
  AND U1213 ( .A(b[1]), .B(a[10]), .Z(\mult_44/ab[10][1] ) );
  AND U1214 ( .A(a[10]), .B(b[0]), .Z(\mult_44/ab[10][0] ) );
  AND U1215 ( .A(b[3]), .B(a[109]), .Z(\mult_44/ab[109][3] ) );
  AND U1216 ( .A(b[2]), .B(a[109]), .Z(\mult_44/ab[109][2] ) );
  AND U1217 ( .A(b[1]), .B(a[109]), .Z(\mult_44/ab[109][1] ) );
  AND U1218 ( .A(a[109]), .B(b[0]), .Z(\mult_44/ab[109][0] ) );
  AND U1219 ( .A(b[3]), .B(a[108]), .Z(\mult_44/ab[108][3] ) );
  AND U1220 ( .A(b[2]), .B(a[108]), .Z(\mult_44/ab[108][2] ) );
  AND U1221 ( .A(b[1]), .B(a[108]), .Z(\mult_44/ab[108][1] ) );
  AND U1222 ( .A(a[108]), .B(b[0]), .Z(\mult_44/ab[108][0] ) );
  AND U1223 ( .A(b[3]), .B(a[107]), .Z(\mult_44/ab[107][3] ) );
  AND U1224 ( .A(b[2]), .B(a[107]), .Z(\mult_44/ab[107][2] ) );
  AND U1225 ( .A(b[1]), .B(a[107]), .Z(\mult_44/ab[107][1] ) );
  AND U1226 ( .A(a[107]), .B(b[0]), .Z(\mult_44/ab[107][0] ) );
  AND U1227 ( .A(b[3]), .B(a[106]), .Z(\mult_44/ab[106][3] ) );
  AND U1228 ( .A(b[2]), .B(a[106]), .Z(\mult_44/ab[106][2] ) );
  AND U1229 ( .A(b[1]), .B(a[106]), .Z(\mult_44/ab[106][1] ) );
  AND U1230 ( .A(a[106]), .B(b[0]), .Z(\mult_44/ab[106][0] ) );
  AND U1231 ( .A(b[3]), .B(a[105]), .Z(\mult_44/ab[105][3] ) );
  AND U1232 ( .A(b[2]), .B(a[105]), .Z(\mult_44/ab[105][2] ) );
  AND U1233 ( .A(b[1]), .B(a[105]), .Z(\mult_44/ab[105][1] ) );
  AND U1234 ( .A(a[105]), .B(b[0]), .Z(\mult_44/ab[105][0] ) );
  AND U1235 ( .A(b[3]), .B(a[104]), .Z(\mult_44/ab[104][3] ) );
  AND U1236 ( .A(b[2]), .B(a[104]), .Z(\mult_44/ab[104][2] ) );
  AND U1237 ( .A(b[1]), .B(a[104]), .Z(\mult_44/ab[104][1] ) );
  AND U1238 ( .A(a[104]), .B(b[0]), .Z(\mult_44/ab[104][0] ) );
  AND U1239 ( .A(b[3]), .B(a[103]), .Z(\mult_44/ab[103][3] ) );
  AND U1240 ( .A(b[2]), .B(a[103]), .Z(\mult_44/ab[103][2] ) );
  AND U1241 ( .A(b[1]), .B(a[103]), .Z(\mult_44/ab[103][1] ) );
  AND U1242 ( .A(a[103]), .B(b[0]), .Z(\mult_44/ab[103][0] ) );
  AND U1243 ( .A(b[3]), .B(a[102]), .Z(\mult_44/ab[102][3] ) );
  AND U1244 ( .A(b[2]), .B(a[102]), .Z(\mult_44/ab[102][2] ) );
  AND U1245 ( .A(b[1]), .B(a[102]), .Z(\mult_44/ab[102][1] ) );
  AND U1246 ( .A(a[102]), .B(b[0]), .Z(\mult_44/ab[102][0] ) );
  AND U1247 ( .A(b[3]), .B(a[101]), .Z(\mult_44/ab[101][3] ) );
  AND U1248 ( .A(b[2]), .B(a[101]), .Z(\mult_44/ab[101][2] ) );
  AND U1249 ( .A(b[1]), .B(a[101]), .Z(\mult_44/ab[101][1] ) );
  AND U1250 ( .A(a[101]), .B(b[0]), .Z(\mult_44/ab[101][0] ) );
  AND U1251 ( .A(b[3]), .B(a[100]), .Z(\mult_44/ab[100][3] ) );
  AND U1252 ( .A(b[2]), .B(a[100]), .Z(\mult_44/ab[100][2] ) );
  AND U1253 ( .A(b[1]), .B(a[100]), .Z(\mult_44/ab[100][1] ) );
  AND U1254 ( .A(a[100]), .B(b[0]), .Z(\mult_44/ab[100][0] ) );
  AND U1255 ( .A(a[0]), .B(b[3]), .Z(\mult_44/ab[0][3] ) );
  AND U1256 ( .A(a[0]), .B(b[2]), .Z(\mult_44/ab[0][2] ) );
  AND U1257 ( .A(a[0]), .B(b[1]), .Z(\mult_44/ab[0][1] ) );
  XNOR U1258 ( .A(\mult_44/PROD1[3] ), .B(n616), .Z(c[127]) );
  XOR U1259 ( .A(n617), .B(n618), .Z(n615) );
  ANDN U1260 ( .B(n619), .A(n620), .Z(n618) );
  XOR U1261 ( .A(clocal[2]), .B(n617), .Z(n619) );
  XNOR U1262 ( .A(clocal[2]), .B(n620), .Z(c[126]) );
  XNOR U1263 ( .A(n621), .B(n622), .Z(n617) );
  NANDN U1264 ( .A(n623), .B(n624), .Z(n621) );
  XOR U1265 ( .A(clocal[1]), .B(n622), .Z(n624) );
  XNOR U1266 ( .A(clocal[1]), .B(n623), .Z(c[125]) );
  XNOR U1267 ( .A(n622), .B(sreg[129]), .Z(n623) );
  ANDN U1268 ( .B(sreg[128]), .A(n625), .Z(n622) );
  XNOR U1269 ( .A(sreg[128]), .B(n625), .Z(c[124]) );
  NAND U1270 ( .A(b[0]), .B(a[0]), .Z(n625) );
endmodule

