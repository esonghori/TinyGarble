
module sum_N128_CC1 ( clk, rst, a, b, c );
  input [127:0] a;
  input [127:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634;

  XOR U2 ( .A(a[24]), .B(b[24]), .Z(n2) );
  NANDN U3 ( .A(n467), .B(n2), .Z(n3) );
  NAND U4 ( .A(a[24]), .B(b[24]), .Z(n4) );
  AND U5 ( .A(n3), .B(n4), .Z(n379) );
  XOR U6 ( .A(a[3]), .B(b[3]), .Z(n5) );
  NANDN U7 ( .A(n501), .B(n5), .Z(n6) );
  NAND U8 ( .A(a[3]), .B(b[3]), .Z(n7) );
  AND U9 ( .A(n6), .B(n7), .Z(n523) );
  XOR U10 ( .A(a[6]), .B(b[6]), .Z(n8) );
  NANDN U11 ( .A(n567), .B(n8), .Z(n9) );
  NAND U12 ( .A(a[6]), .B(b[6]), .Z(n10) );
  AND U13 ( .A(n9), .B(n10), .Z(n589) );
  XOR U14 ( .A(b[9]), .B(a[9]), .Z(n11) );
  NANDN U15 ( .A(n633), .B(n11), .Z(n12) );
  NAND U16 ( .A(b[9]), .B(a[9]), .Z(n13) );
  AND U17 ( .A(n12), .B(n13), .Z(n402) );
  XOR U18 ( .A(a[12]), .B(b[12]), .Z(n14) );
  NANDN U19 ( .A(n441), .B(n14), .Z(n15) );
  NAND U20 ( .A(a[12]), .B(b[12]), .Z(n16) );
  AND U21 ( .A(n15), .B(n16), .Z(n443) );
  XOR U22 ( .A(a[15]), .B(b[15]), .Z(n17) );
  NANDN U23 ( .A(n447), .B(n17), .Z(n18) );
  NAND U24 ( .A(a[15]), .B(b[15]), .Z(n19) );
  AND U25 ( .A(n18), .B(n19), .Z(n449) );
  XOR U26 ( .A(a[18]), .B(b[18]), .Z(n20) );
  NANDN U27 ( .A(n453), .B(n20), .Z(n21) );
  NAND U28 ( .A(a[18]), .B(b[18]), .Z(n22) );
  AND U29 ( .A(n21), .B(n22), .Z(n455) );
  XOR U30 ( .A(a[21]), .B(b[21]), .Z(n23) );
  NANDN U31 ( .A(n461), .B(n23), .Z(n24) );
  NAND U32 ( .A(a[21]), .B(b[21]), .Z(n25) );
  AND U33 ( .A(n24), .B(n25), .Z(n463) );
  XOR U34 ( .A(a[28]), .B(b[28]), .Z(n26) );
  NANDN U35 ( .A(n475), .B(n26), .Z(n27) );
  NAND U36 ( .A(a[28]), .B(b[28]), .Z(n28) );
  AND U37 ( .A(n27), .B(n28), .Z(n477) );
  XOR U38 ( .A(a[31]), .B(b[31]), .Z(n29) );
  NANDN U39 ( .A(n483), .B(n29), .Z(n30) );
  NAND U40 ( .A(a[31]), .B(b[31]), .Z(n31) );
  AND U41 ( .A(n30), .B(n31), .Z(n485) );
  XOR U42 ( .A(a[34]), .B(b[34]), .Z(n32) );
  NANDN U43 ( .A(n489), .B(n32), .Z(n33) );
  NAND U44 ( .A(a[34]), .B(b[34]), .Z(n34) );
  AND U45 ( .A(n33), .B(n34), .Z(n491) );
  XOR U46 ( .A(a[37]), .B(b[37]), .Z(n35) );
  NANDN U47 ( .A(n495), .B(n35), .Z(n36) );
  NAND U48 ( .A(a[37]), .B(b[37]), .Z(n37) );
  AND U49 ( .A(n36), .B(n37), .Z(n497) );
  XOR U50 ( .A(a[40]), .B(b[40]), .Z(n38) );
  NANDN U51 ( .A(n503), .B(n38), .Z(n39) );
  NAND U52 ( .A(a[40]), .B(b[40]), .Z(n40) );
  AND U53 ( .A(n39), .B(n40), .Z(n505) );
  XOR U54 ( .A(a[43]), .B(b[43]), .Z(n41) );
  NANDN U55 ( .A(n509), .B(n41), .Z(n42) );
  NAND U56 ( .A(a[43]), .B(b[43]), .Z(n43) );
  AND U57 ( .A(n42), .B(n43), .Z(n511) );
  XOR U58 ( .A(a[46]), .B(b[46]), .Z(n44) );
  NANDN U59 ( .A(n515), .B(n44), .Z(n45) );
  NAND U60 ( .A(a[46]), .B(b[46]), .Z(n46) );
  AND U61 ( .A(n45), .B(n46), .Z(n517) );
  XOR U62 ( .A(a[49]), .B(b[49]), .Z(n47) );
  NANDN U63 ( .A(n521), .B(n47), .Z(n48) );
  NAND U64 ( .A(a[49]), .B(b[49]), .Z(n49) );
  AND U65 ( .A(n48), .B(n49), .Z(n525) );
  XOR U66 ( .A(a[52]), .B(b[52]), .Z(n50) );
  NANDN U67 ( .A(n529), .B(n50), .Z(n51) );
  NAND U68 ( .A(a[52]), .B(b[52]), .Z(n52) );
  AND U69 ( .A(n51), .B(n52), .Z(n531) );
  XOR U70 ( .A(a[55]), .B(b[55]), .Z(n53) );
  NANDN U71 ( .A(n535), .B(n53), .Z(n54) );
  NAND U72 ( .A(a[55]), .B(b[55]), .Z(n55) );
  AND U73 ( .A(n54), .B(n55), .Z(n537) );
  XOR U74 ( .A(a[58]), .B(b[58]), .Z(n56) );
  NANDN U75 ( .A(n541), .B(n56), .Z(n57) );
  NAND U76 ( .A(a[58]), .B(b[58]), .Z(n58) );
  AND U77 ( .A(n57), .B(n58), .Z(n543) );
  XOR U78 ( .A(a[61]), .B(b[61]), .Z(n59) );
  NANDN U79 ( .A(n549), .B(n59), .Z(n60) );
  NAND U80 ( .A(a[61]), .B(b[61]), .Z(n61) );
  AND U81 ( .A(n60), .B(n61), .Z(n551) );
  XOR U82 ( .A(a[64]), .B(b[64]), .Z(n62) );
  NANDN U83 ( .A(n555), .B(n62), .Z(n63) );
  NAND U84 ( .A(a[64]), .B(b[64]), .Z(n64) );
  AND U85 ( .A(n63), .B(n64), .Z(n557) );
  XOR U86 ( .A(a[67]), .B(b[67]), .Z(n65) );
  NANDN U87 ( .A(n561), .B(n65), .Z(n66) );
  NAND U88 ( .A(a[67]), .B(b[67]), .Z(n67) );
  AND U89 ( .A(n66), .B(n67), .Z(n563) );
  XOR U90 ( .A(a[70]), .B(b[70]), .Z(n68) );
  NANDN U91 ( .A(n569), .B(n68), .Z(n69) );
  NAND U92 ( .A(a[70]), .B(b[70]), .Z(n70) );
  AND U93 ( .A(n69), .B(n70), .Z(n571) );
  XOR U94 ( .A(a[73]), .B(b[73]), .Z(n71) );
  NANDN U95 ( .A(n575), .B(n71), .Z(n72) );
  NAND U96 ( .A(a[73]), .B(b[73]), .Z(n73) );
  AND U97 ( .A(n72), .B(n73), .Z(n577) );
  XOR U98 ( .A(a[76]), .B(b[76]), .Z(n74) );
  NANDN U99 ( .A(n581), .B(n74), .Z(n75) );
  NAND U100 ( .A(a[76]), .B(b[76]), .Z(n76) );
  AND U101 ( .A(n75), .B(n76), .Z(n583) );
  XOR U102 ( .A(a[79]), .B(b[79]), .Z(n77) );
  NANDN U103 ( .A(n587), .B(n77), .Z(n78) );
  NAND U104 ( .A(a[79]), .B(b[79]), .Z(n79) );
  AND U105 ( .A(n78), .B(n79), .Z(n591) );
  XOR U106 ( .A(a[82]), .B(b[82]), .Z(n80) );
  NANDN U107 ( .A(n595), .B(n80), .Z(n81) );
  NAND U108 ( .A(a[82]), .B(b[82]), .Z(n82) );
  AND U109 ( .A(n81), .B(n82), .Z(n597) );
  XOR U110 ( .A(a[85]), .B(b[85]), .Z(n83) );
  NANDN U111 ( .A(n601), .B(n83), .Z(n84) );
  NAND U112 ( .A(a[85]), .B(b[85]), .Z(n85) );
  AND U113 ( .A(n84), .B(n85), .Z(n603) );
  XOR U114 ( .A(a[88]), .B(b[88]), .Z(n86) );
  NANDN U115 ( .A(n607), .B(n86), .Z(n87) );
  NAND U116 ( .A(a[88]), .B(b[88]), .Z(n88) );
  AND U117 ( .A(n87), .B(n88), .Z(n609) );
  XOR U118 ( .A(a[91]), .B(b[91]), .Z(n89) );
  NANDN U119 ( .A(n615), .B(n89), .Z(n90) );
  NAND U120 ( .A(a[91]), .B(b[91]), .Z(n91) );
  AND U121 ( .A(n90), .B(n91), .Z(n617) );
  XOR U122 ( .A(a[94]), .B(b[94]), .Z(n92) );
  NANDN U123 ( .A(n621), .B(n92), .Z(n93) );
  NAND U124 ( .A(a[94]), .B(b[94]), .Z(n94) );
  AND U125 ( .A(n93), .B(n94), .Z(n623) );
  XOR U126 ( .A(a[97]), .B(b[97]), .Z(n95) );
  NANDN U127 ( .A(n627), .B(n95), .Z(n96) );
  NAND U128 ( .A(a[97]), .B(b[97]), .Z(n97) );
  AND U129 ( .A(n96), .B(n97), .Z(n629) );
  XOR U130 ( .A(b[100]), .B(a[100]), .Z(n98) );
  NANDN U131 ( .A(n384), .B(n98), .Z(n99) );
  NAND U132 ( .A(b[100]), .B(a[100]), .Z(n100) );
  AND U133 ( .A(n99), .B(n100), .Z(n386) );
  XOR U134 ( .A(b[103]), .B(a[103]), .Z(n101) );
  NANDN U135 ( .A(n390), .B(n101), .Z(n102) );
  NAND U136 ( .A(b[103]), .B(a[103]), .Z(n103) );
  AND U137 ( .A(n102), .B(n103), .Z(n392) );
  XOR U138 ( .A(b[106]), .B(a[106]), .Z(n104) );
  NANDN U139 ( .A(n396), .B(n104), .Z(n105) );
  NAND U140 ( .A(b[106]), .B(a[106]), .Z(n106) );
  AND U141 ( .A(n105), .B(n106), .Z(n398) );
  XOR U142 ( .A(b[109]), .B(a[109]), .Z(n107) );
  NANDN U143 ( .A(n404), .B(n107), .Z(n108) );
  NAND U144 ( .A(b[109]), .B(a[109]), .Z(n109) );
  AND U145 ( .A(n108), .B(n109), .Z(n406) );
  XOR U146 ( .A(b[112]), .B(a[112]), .Z(n110) );
  NANDN U147 ( .A(n410), .B(n110), .Z(n111) );
  NAND U148 ( .A(b[112]), .B(a[112]), .Z(n112) );
  AND U149 ( .A(n111), .B(n112), .Z(n412) );
  XOR U150 ( .A(b[115]), .B(a[115]), .Z(n113) );
  NANDN U151 ( .A(n416), .B(n113), .Z(n114) );
  NAND U152 ( .A(b[115]), .B(a[115]), .Z(n115) );
  AND U153 ( .A(n114), .B(n115), .Z(n418) );
  XOR U154 ( .A(b[118]), .B(a[118]), .Z(n116) );
  NANDN U155 ( .A(n422), .B(n116), .Z(n117) );
  NAND U156 ( .A(b[118]), .B(a[118]), .Z(n118) );
  AND U157 ( .A(n117), .B(n118), .Z(n426) );
  XOR U158 ( .A(b[121]), .B(a[121]), .Z(n119) );
  NANDN U159 ( .A(n430), .B(n119), .Z(n120) );
  NAND U160 ( .A(b[121]), .B(a[121]), .Z(n121) );
  AND U161 ( .A(n120), .B(n121), .Z(n432) );
  XOR U162 ( .A(b[124]), .B(a[124]), .Z(n122) );
  NANDN U163 ( .A(n436), .B(n122), .Z(n123) );
  NAND U164 ( .A(b[124]), .B(a[124]), .Z(n124) );
  AND U165 ( .A(n123), .B(n124), .Z(n438) );
  XOR U166 ( .A(b[1]), .B(a[1]), .Z(n125) );
  NANDN U167 ( .A(n458), .B(n125), .Z(n126) );
  NAND U168 ( .A(b[1]), .B(a[1]), .Z(n127) );
  AND U169 ( .A(n126), .B(n127), .Z(n479) );
  XOR U170 ( .A(a[4]), .B(b[4]), .Z(n128) );
  NANDN U171 ( .A(n523), .B(n128), .Z(n129) );
  NAND U172 ( .A(a[4]), .B(b[4]), .Z(n130) );
  AND U173 ( .A(n129), .B(n130), .Z(n545) );
  XOR U174 ( .A(a[7]), .B(b[7]), .Z(n131) );
  NANDN U175 ( .A(n589), .B(n131), .Z(n132) );
  NAND U176 ( .A(a[7]), .B(b[7]), .Z(n133) );
  AND U177 ( .A(n132), .B(n133), .Z(n611) );
  XOR U178 ( .A(a[10]), .B(b[10]), .Z(n134) );
  NANDN U179 ( .A(n402), .B(n134), .Z(n135) );
  NAND U180 ( .A(a[10]), .B(b[10]), .Z(n136) );
  AND U181 ( .A(n135), .B(n136), .Z(n424) );
  XOR U182 ( .A(a[13]), .B(b[13]), .Z(n137) );
  NANDN U183 ( .A(n443), .B(n137), .Z(n138) );
  NAND U184 ( .A(a[13]), .B(b[13]), .Z(n139) );
  AND U185 ( .A(n138), .B(n139), .Z(n445) );
  XOR U186 ( .A(a[16]), .B(b[16]), .Z(n140) );
  NANDN U187 ( .A(n449), .B(n140), .Z(n141) );
  NAND U188 ( .A(a[16]), .B(b[16]), .Z(n142) );
  AND U189 ( .A(n141), .B(n142), .Z(n451) );
  XOR U190 ( .A(a[19]), .B(b[19]), .Z(n143) );
  NANDN U191 ( .A(n455), .B(n143), .Z(n144) );
  NAND U192 ( .A(a[19]), .B(b[19]), .Z(n145) );
  AND U193 ( .A(n144), .B(n145), .Z(n459) );
  XOR U194 ( .A(a[22]), .B(b[22]), .Z(n146) );
  NANDN U195 ( .A(n463), .B(n146), .Z(n147) );
  NAND U196 ( .A(a[22]), .B(b[22]), .Z(n148) );
  AND U197 ( .A(n147), .B(n148), .Z(n465) );
  XOR U198 ( .A(a[26]), .B(b[26]), .Z(n149) );
  NANDN U199 ( .A(n471), .B(n149), .Z(n150) );
  NAND U200 ( .A(a[26]), .B(b[26]), .Z(n151) );
  AND U201 ( .A(n150), .B(n151), .Z(n473) );
  XOR U202 ( .A(a[29]), .B(b[29]), .Z(n152) );
  NANDN U203 ( .A(n477), .B(n152), .Z(n153) );
  NAND U204 ( .A(a[29]), .B(b[29]), .Z(n154) );
  AND U205 ( .A(n153), .B(n154), .Z(n481) );
  XOR U206 ( .A(a[32]), .B(b[32]), .Z(n155) );
  NANDN U207 ( .A(n485), .B(n155), .Z(n156) );
  NAND U208 ( .A(a[32]), .B(b[32]), .Z(n157) );
  AND U209 ( .A(n156), .B(n157), .Z(n487) );
  XOR U210 ( .A(a[35]), .B(b[35]), .Z(n158) );
  NANDN U211 ( .A(n491), .B(n158), .Z(n159) );
  NAND U212 ( .A(a[35]), .B(b[35]), .Z(n160) );
  AND U213 ( .A(n159), .B(n160), .Z(n493) );
  XOR U214 ( .A(a[38]), .B(b[38]), .Z(n161) );
  NANDN U215 ( .A(n497), .B(n161), .Z(n162) );
  NAND U216 ( .A(a[38]), .B(b[38]), .Z(n163) );
  AND U217 ( .A(n162), .B(n163), .Z(n499) );
  XOR U218 ( .A(a[41]), .B(b[41]), .Z(n164) );
  NANDN U219 ( .A(n505), .B(n164), .Z(n165) );
  NAND U220 ( .A(a[41]), .B(b[41]), .Z(n166) );
  AND U221 ( .A(n165), .B(n166), .Z(n507) );
  XOR U222 ( .A(a[44]), .B(b[44]), .Z(n167) );
  NANDN U223 ( .A(n511), .B(n167), .Z(n168) );
  NAND U224 ( .A(a[44]), .B(b[44]), .Z(n169) );
  AND U225 ( .A(n168), .B(n169), .Z(n513) );
  XOR U226 ( .A(a[47]), .B(b[47]), .Z(n170) );
  NANDN U227 ( .A(n517), .B(n170), .Z(n171) );
  NAND U228 ( .A(a[47]), .B(b[47]), .Z(n172) );
  AND U229 ( .A(n171), .B(n172), .Z(n519) );
  XOR U230 ( .A(a[50]), .B(b[50]), .Z(n173) );
  NANDN U231 ( .A(n525), .B(n173), .Z(n174) );
  NAND U232 ( .A(a[50]), .B(b[50]), .Z(n175) );
  AND U233 ( .A(n174), .B(n175), .Z(n527) );
  XOR U234 ( .A(a[53]), .B(b[53]), .Z(n176) );
  NANDN U235 ( .A(n531), .B(n176), .Z(n177) );
  NAND U236 ( .A(a[53]), .B(b[53]), .Z(n178) );
  AND U237 ( .A(n177), .B(n178), .Z(n533) );
  XOR U238 ( .A(a[56]), .B(b[56]), .Z(n179) );
  NANDN U239 ( .A(n537), .B(n179), .Z(n180) );
  NAND U240 ( .A(a[56]), .B(b[56]), .Z(n181) );
  AND U241 ( .A(n180), .B(n181), .Z(n539) );
  XOR U242 ( .A(a[59]), .B(b[59]), .Z(n182) );
  NANDN U243 ( .A(n543), .B(n182), .Z(n183) );
  NAND U244 ( .A(a[59]), .B(b[59]), .Z(n184) );
  AND U245 ( .A(n183), .B(n184), .Z(n547) );
  XOR U246 ( .A(a[62]), .B(b[62]), .Z(n185) );
  NANDN U247 ( .A(n551), .B(n185), .Z(n186) );
  NAND U248 ( .A(a[62]), .B(b[62]), .Z(n187) );
  AND U249 ( .A(n186), .B(n187), .Z(n553) );
  XOR U250 ( .A(a[65]), .B(b[65]), .Z(n188) );
  NANDN U251 ( .A(n557), .B(n188), .Z(n189) );
  NAND U252 ( .A(a[65]), .B(b[65]), .Z(n190) );
  AND U253 ( .A(n189), .B(n190), .Z(n559) );
  XOR U254 ( .A(a[68]), .B(b[68]), .Z(n191) );
  NANDN U255 ( .A(n563), .B(n191), .Z(n192) );
  NAND U256 ( .A(a[68]), .B(b[68]), .Z(n193) );
  AND U257 ( .A(n192), .B(n193), .Z(n565) );
  XOR U258 ( .A(a[71]), .B(b[71]), .Z(n194) );
  NANDN U259 ( .A(n571), .B(n194), .Z(n195) );
  NAND U260 ( .A(a[71]), .B(b[71]), .Z(n196) );
  AND U261 ( .A(n195), .B(n196), .Z(n573) );
  XOR U262 ( .A(a[74]), .B(b[74]), .Z(n197) );
  NANDN U263 ( .A(n577), .B(n197), .Z(n198) );
  NAND U264 ( .A(a[74]), .B(b[74]), .Z(n199) );
  AND U265 ( .A(n198), .B(n199), .Z(n579) );
  XOR U266 ( .A(a[77]), .B(b[77]), .Z(n200) );
  NANDN U267 ( .A(n583), .B(n200), .Z(n201) );
  NAND U268 ( .A(a[77]), .B(b[77]), .Z(n202) );
  AND U269 ( .A(n201), .B(n202), .Z(n585) );
  XOR U270 ( .A(a[80]), .B(b[80]), .Z(n203) );
  NANDN U271 ( .A(n591), .B(n203), .Z(n204) );
  NAND U272 ( .A(a[80]), .B(b[80]), .Z(n205) );
  AND U273 ( .A(n204), .B(n205), .Z(n593) );
  XOR U274 ( .A(a[83]), .B(b[83]), .Z(n206) );
  NANDN U275 ( .A(n597), .B(n206), .Z(n207) );
  NAND U276 ( .A(a[83]), .B(b[83]), .Z(n208) );
  AND U277 ( .A(n207), .B(n208), .Z(n599) );
  XOR U278 ( .A(a[86]), .B(b[86]), .Z(n209) );
  NANDN U279 ( .A(n603), .B(n209), .Z(n210) );
  NAND U280 ( .A(a[86]), .B(b[86]), .Z(n211) );
  AND U281 ( .A(n210), .B(n211), .Z(n605) );
  XOR U282 ( .A(a[89]), .B(b[89]), .Z(n212) );
  NANDN U283 ( .A(n609), .B(n212), .Z(n213) );
  NAND U284 ( .A(a[89]), .B(b[89]), .Z(n214) );
  AND U285 ( .A(n213), .B(n214), .Z(n613) );
  XOR U286 ( .A(a[92]), .B(b[92]), .Z(n215) );
  NANDN U287 ( .A(n617), .B(n215), .Z(n216) );
  NAND U288 ( .A(a[92]), .B(b[92]), .Z(n217) );
  AND U289 ( .A(n216), .B(n217), .Z(n619) );
  XOR U290 ( .A(a[95]), .B(b[95]), .Z(n218) );
  NANDN U291 ( .A(n623), .B(n218), .Z(n219) );
  NAND U292 ( .A(a[95]), .B(b[95]), .Z(n220) );
  AND U293 ( .A(n219), .B(n220), .Z(n625) );
  XOR U294 ( .A(a[98]), .B(b[98]), .Z(n221) );
  NANDN U295 ( .A(n629), .B(n221), .Z(n222) );
  NAND U296 ( .A(a[98]), .B(b[98]), .Z(n223) );
  AND U297 ( .A(n222), .B(n223), .Z(n631) );
  XOR U298 ( .A(b[101]), .B(a[101]), .Z(n224) );
  NANDN U299 ( .A(n386), .B(n224), .Z(n225) );
  NAND U300 ( .A(b[101]), .B(a[101]), .Z(n226) );
  AND U301 ( .A(n225), .B(n226), .Z(n388) );
  XOR U302 ( .A(b[104]), .B(a[104]), .Z(n227) );
  NANDN U303 ( .A(n392), .B(n227), .Z(n228) );
  NAND U304 ( .A(b[104]), .B(a[104]), .Z(n229) );
  AND U305 ( .A(n228), .B(n229), .Z(n394) );
  XOR U306 ( .A(b[107]), .B(a[107]), .Z(n230) );
  NANDN U307 ( .A(n398), .B(n230), .Z(n231) );
  NAND U308 ( .A(b[107]), .B(a[107]), .Z(n232) );
  AND U309 ( .A(n231), .B(n232), .Z(n400) );
  XOR U310 ( .A(b[110]), .B(a[110]), .Z(n233) );
  NANDN U311 ( .A(n406), .B(n233), .Z(n234) );
  NAND U312 ( .A(b[110]), .B(a[110]), .Z(n235) );
  AND U313 ( .A(n234), .B(n235), .Z(n408) );
  XOR U314 ( .A(b[113]), .B(a[113]), .Z(n236) );
  NANDN U315 ( .A(n412), .B(n236), .Z(n237) );
  NAND U316 ( .A(b[113]), .B(a[113]), .Z(n238) );
  AND U317 ( .A(n237), .B(n238), .Z(n414) );
  XOR U318 ( .A(b[116]), .B(a[116]), .Z(n239) );
  NANDN U319 ( .A(n418), .B(n239), .Z(n240) );
  NAND U320 ( .A(b[116]), .B(a[116]), .Z(n241) );
  AND U321 ( .A(n240), .B(n241), .Z(n420) );
  XOR U322 ( .A(b[119]), .B(a[119]), .Z(n242) );
  NANDN U323 ( .A(n426), .B(n242), .Z(n243) );
  NAND U324 ( .A(b[119]), .B(a[119]), .Z(n244) );
  AND U325 ( .A(n243), .B(n244), .Z(n428) );
  XOR U326 ( .A(b[122]), .B(a[122]), .Z(n245) );
  NANDN U327 ( .A(n432), .B(n245), .Z(n246) );
  NAND U328 ( .A(b[122]), .B(a[122]), .Z(n247) );
  AND U329 ( .A(n246), .B(n247), .Z(n434) );
  XOR U330 ( .A(b[125]), .B(a[125]), .Z(n248) );
  NANDN U331 ( .A(n438), .B(n248), .Z(n249) );
  NAND U332 ( .A(b[125]), .B(a[125]), .Z(n250) );
  AND U333 ( .A(n249), .B(n250), .Z(n440) );
  XOR U334 ( .A(a[2]), .B(b[2]), .Z(n251) );
  NANDN U335 ( .A(n479), .B(n251), .Z(n252) );
  NAND U336 ( .A(a[2]), .B(b[2]), .Z(n253) );
  AND U337 ( .A(n252), .B(n253), .Z(n501) );
  XOR U338 ( .A(a[5]), .B(b[5]), .Z(n254) );
  NANDN U339 ( .A(n545), .B(n254), .Z(n255) );
  NAND U340 ( .A(a[5]), .B(b[5]), .Z(n256) );
  AND U341 ( .A(n255), .B(n256), .Z(n567) );
  XOR U342 ( .A(a[8]), .B(b[8]), .Z(n257) );
  NANDN U343 ( .A(n611), .B(n257), .Z(n258) );
  NAND U344 ( .A(a[8]), .B(b[8]), .Z(n259) );
  AND U345 ( .A(n258), .B(n259), .Z(n633) );
  XOR U346 ( .A(a[11]), .B(b[11]), .Z(n260) );
  NANDN U347 ( .A(n424), .B(n260), .Z(n261) );
  NAND U348 ( .A(a[11]), .B(b[11]), .Z(n262) );
  AND U349 ( .A(n261), .B(n262), .Z(n441) );
  XOR U350 ( .A(a[14]), .B(b[14]), .Z(n263) );
  NANDN U351 ( .A(n445), .B(n263), .Z(n264) );
  NAND U352 ( .A(a[14]), .B(b[14]), .Z(n265) );
  AND U353 ( .A(n264), .B(n265), .Z(n447) );
  XOR U354 ( .A(a[17]), .B(b[17]), .Z(n266) );
  NANDN U355 ( .A(n451), .B(n266), .Z(n267) );
  NAND U356 ( .A(a[17]), .B(b[17]), .Z(n268) );
  AND U357 ( .A(n267), .B(n268), .Z(n453) );
  XOR U358 ( .A(a[20]), .B(b[20]), .Z(n269) );
  NANDN U359 ( .A(n459), .B(n269), .Z(n270) );
  NAND U360 ( .A(a[20]), .B(b[20]), .Z(n271) );
  AND U361 ( .A(n270), .B(n271), .Z(n461) );
  XOR U362 ( .A(a[23]), .B(b[23]), .Z(n272) );
  NANDN U363 ( .A(n465), .B(n272), .Z(n273) );
  NAND U364 ( .A(a[23]), .B(b[23]), .Z(n274) );
  AND U365 ( .A(n273), .B(n274), .Z(n467) );
  XOR U366 ( .A(a[27]), .B(b[27]), .Z(n275) );
  NANDN U367 ( .A(n473), .B(n275), .Z(n276) );
  NAND U368 ( .A(a[27]), .B(b[27]), .Z(n277) );
  AND U369 ( .A(n276), .B(n277), .Z(n475) );
  XOR U370 ( .A(a[30]), .B(b[30]), .Z(n278) );
  NANDN U371 ( .A(n481), .B(n278), .Z(n279) );
  NAND U372 ( .A(a[30]), .B(b[30]), .Z(n280) );
  AND U373 ( .A(n279), .B(n280), .Z(n483) );
  XOR U374 ( .A(a[33]), .B(b[33]), .Z(n281) );
  NANDN U375 ( .A(n487), .B(n281), .Z(n282) );
  NAND U376 ( .A(a[33]), .B(b[33]), .Z(n283) );
  AND U377 ( .A(n282), .B(n283), .Z(n489) );
  XOR U378 ( .A(a[36]), .B(b[36]), .Z(n284) );
  NANDN U379 ( .A(n493), .B(n284), .Z(n285) );
  NAND U380 ( .A(a[36]), .B(b[36]), .Z(n286) );
  AND U381 ( .A(n285), .B(n286), .Z(n495) );
  XOR U382 ( .A(a[39]), .B(b[39]), .Z(n287) );
  NANDN U383 ( .A(n499), .B(n287), .Z(n288) );
  NAND U384 ( .A(a[39]), .B(b[39]), .Z(n289) );
  AND U385 ( .A(n288), .B(n289), .Z(n503) );
  XOR U386 ( .A(a[42]), .B(b[42]), .Z(n290) );
  NANDN U387 ( .A(n507), .B(n290), .Z(n291) );
  NAND U388 ( .A(a[42]), .B(b[42]), .Z(n292) );
  AND U389 ( .A(n291), .B(n292), .Z(n509) );
  XOR U390 ( .A(a[45]), .B(b[45]), .Z(n293) );
  NANDN U391 ( .A(n513), .B(n293), .Z(n294) );
  NAND U392 ( .A(a[45]), .B(b[45]), .Z(n295) );
  AND U393 ( .A(n294), .B(n295), .Z(n515) );
  XOR U394 ( .A(a[48]), .B(b[48]), .Z(n296) );
  NANDN U395 ( .A(n519), .B(n296), .Z(n297) );
  NAND U396 ( .A(a[48]), .B(b[48]), .Z(n298) );
  AND U397 ( .A(n297), .B(n298), .Z(n521) );
  XOR U398 ( .A(a[51]), .B(b[51]), .Z(n299) );
  NANDN U399 ( .A(n527), .B(n299), .Z(n300) );
  NAND U400 ( .A(a[51]), .B(b[51]), .Z(n301) );
  AND U401 ( .A(n300), .B(n301), .Z(n529) );
  XOR U402 ( .A(a[54]), .B(b[54]), .Z(n302) );
  NANDN U403 ( .A(n533), .B(n302), .Z(n303) );
  NAND U404 ( .A(a[54]), .B(b[54]), .Z(n304) );
  AND U405 ( .A(n303), .B(n304), .Z(n535) );
  XOR U406 ( .A(a[57]), .B(b[57]), .Z(n305) );
  NANDN U407 ( .A(n539), .B(n305), .Z(n306) );
  NAND U408 ( .A(a[57]), .B(b[57]), .Z(n307) );
  AND U409 ( .A(n306), .B(n307), .Z(n541) );
  XOR U410 ( .A(a[60]), .B(b[60]), .Z(n308) );
  NANDN U411 ( .A(n547), .B(n308), .Z(n309) );
  NAND U412 ( .A(a[60]), .B(b[60]), .Z(n310) );
  AND U413 ( .A(n309), .B(n310), .Z(n549) );
  XOR U414 ( .A(a[63]), .B(b[63]), .Z(n311) );
  NANDN U415 ( .A(n553), .B(n311), .Z(n312) );
  NAND U416 ( .A(a[63]), .B(b[63]), .Z(n313) );
  AND U417 ( .A(n312), .B(n313), .Z(n555) );
  XOR U418 ( .A(a[66]), .B(b[66]), .Z(n314) );
  NANDN U419 ( .A(n559), .B(n314), .Z(n315) );
  NAND U420 ( .A(a[66]), .B(b[66]), .Z(n316) );
  AND U421 ( .A(n315), .B(n316), .Z(n561) );
  XOR U422 ( .A(a[69]), .B(b[69]), .Z(n317) );
  NANDN U423 ( .A(n565), .B(n317), .Z(n318) );
  NAND U424 ( .A(a[69]), .B(b[69]), .Z(n319) );
  AND U425 ( .A(n318), .B(n319), .Z(n569) );
  XOR U426 ( .A(a[72]), .B(b[72]), .Z(n320) );
  NANDN U427 ( .A(n573), .B(n320), .Z(n321) );
  NAND U428 ( .A(a[72]), .B(b[72]), .Z(n322) );
  AND U429 ( .A(n321), .B(n322), .Z(n575) );
  XOR U430 ( .A(a[75]), .B(b[75]), .Z(n323) );
  NANDN U431 ( .A(n579), .B(n323), .Z(n324) );
  NAND U432 ( .A(a[75]), .B(b[75]), .Z(n325) );
  AND U433 ( .A(n324), .B(n325), .Z(n581) );
  XOR U434 ( .A(a[78]), .B(b[78]), .Z(n326) );
  NANDN U435 ( .A(n585), .B(n326), .Z(n327) );
  NAND U436 ( .A(a[78]), .B(b[78]), .Z(n328) );
  AND U437 ( .A(n327), .B(n328), .Z(n587) );
  XOR U438 ( .A(a[81]), .B(b[81]), .Z(n329) );
  NANDN U439 ( .A(n593), .B(n329), .Z(n330) );
  NAND U440 ( .A(a[81]), .B(b[81]), .Z(n331) );
  AND U441 ( .A(n330), .B(n331), .Z(n595) );
  XOR U442 ( .A(a[84]), .B(b[84]), .Z(n332) );
  NANDN U443 ( .A(n599), .B(n332), .Z(n333) );
  NAND U444 ( .A(a[84]), .B(b[84]), .Z(n334) );
  AND U445 ( .A(n333), .B(n334), .Z(n601) );
  XOR U446 ( .A(a[87]), .B(b[87]), .Z(n335) );
  NANDN U447 ( .A(n605), .B(n335), .Z(n336) );
  NAND U448 ( .A(a[87]), .B(b[87]), .Z(n337) );
  AND U449 ( .A(n336), .B(n337), .Z(n607) );
  XOR U450 ( .A(a[90]), .B(b[90]), .Z(n338) );
  NANDN U451 ( .A(n613), .B(n338), .Z(n339) );
  NAND U452 ( .A(a[90]), .B(b[90]), .Z(n340) );
  AND U453 ( .A(n339), .B(n340), .Z(n615) );
  XOR U454 ( .A(a[93]), .B(b[93]), .Z(n341) );
  NANDN U455 ( .A(n619), .B(n341), .Z(n342) );
  NAND U456 ( .A(a[93]), .B(b[93]), .Z(n343) );
  AND U457 ( .A(n342), .B(n343), .Z(n621) );
  XOR U458 ( .A(a[96]), .B(b[96]), .Z(n344) );
  NANDN U459 ( .A(n625), .B(n344), .Z(n345) );
  NAND U460 ( .A(a[96]), .B(b[96]), .Z(n346) );
  AND U461 ( .A(n345), .B(n346), .Z(n627) );
  XOR U462 ( .A(b[99]), .B(a[99]), .Z(n347) );
  NANDN U463 ( .A(n631), .B(n347), .Z(n348) );
  NAND U464 ( .A(b[99]), .B(a[99]), .Z(n349) );
  AND U465 ( .A(n348), .B(n349), .Z(n384) );
  XOR U466 ( .A(b[102]), .B(a[102]), .Z(n350) );
  NANDN U467 ( .A(n388), .B(n350), .Z(n351) );
  NAND U468 ( .A(b[102]), .B(a[102]), .Z(n352) );
  AND U469 ( .A(n351), .B(n352), .Z(n390) );
  XOR U470 ( .A(b[105]), .B(a[105]), .Z(n353) );
  NANDN U471 ( .A(n394), .B(n353), .Z(n354) );
  NAND U472 ( .A(b[105]), .B(a[105]), .Z(n355) );
  AND U473 ( .A(n354), .B(n355), .Z(n396) );
  XOR U474 ( .A(b[108]), .B(a[108]), .Z(n356) );
  NANDN U475 ( .A(n400), .B(n356), .Z(n357) );
  NAND U476 ( .A(b[108]), .B(a[108]), .Z(n358) );
  AND U477 ( .A(n357), .B(n358), .Z(n404) );
  XOR U478 ( .A(b[111]), .B(a[111]), .Z(n359) );
  NANDN U479 ( .A(n408), .B(n359), .Z(n360) );
  NAND U480 ( .A(b[111]), .B(a[111]), .Z(n361) );
  AND U481 ( .A(n360), .B(n361), .Z(n410) );
  XOR U482 ( .A(b[114]), .B(a[114]), .Z(n362) );
  NANDN U483 ( .A(n414), .B(n362), .Z(n363) );
  NAND U484 ( .A(b[114]), .B(a[114]), .Z(n364) );
  AND U485 ( .A(n363), .B(n364), .Z(n416) );
  XOR U486 ( .A(b[117]), .B(a[117]), .Z(n365) );
  NANDN U487 ( .A(n420), .B(n365), .Z(n366) );
  NAND U488 ( .A(b[117]), .B(a[117]), .Z(n367) );
  AND U489 ( .A(n366), .B(n367), .Z(n422) );
  XOR U490 ( .A(b[120]), .B(a[120]), .Z(n368) );
  NANDN U491 ( .A(n428), .B(n368), .Z(n369) );
  NAND U492 ( .A(b[120]), .B(a[120]), .Z(n370) );
  AND U493 ( .A(n369), .B(n370), .Z(n430) );
  XOR U494 ( .A(b[123]), .B(a[123]), .Z(n371) );
  NANDN U495 ( .A(n434), .B(n371), .Z(n372) );
  NAND U496 ( .A(b[123]), .B(a[123]), .Z(n373) );
  AND U497 ( .A(n372), .B(n373), .Z(n436) );
  NANDN U498 ( .A(n440), .B(b[126]), .Z(n374) );
  XNOR U499 ( .A(n440), .B(b[126]), .Z(n375) );
  NAND U500 ( .A(a[126]), .B(n375), .Z(n376) );
  NAND U501 ( .A(n374), .B(n376), .Z(n377) );
  XNOR U502 ( .A(a[127]), .B(n377), .Z(n378) );
  XNOR U503 ( .A(b[127]), .B(n378), .Z(c[127]) );
  XOR U504 ( .A(a[0]), .B(b[0]), .Z(c[0]) );
  NAND U505 ( .A(a[0]), .B(b[0]), .Z(n458) );
  IV U506 ( .A(n379), .Z(n470) );
  NAND U507 ( .A(n470), .B(b[25]), .Z(n382) );
  ANDN U508 ( .B(n379), .A(b[25]), .Z(n380) );
  NANDN U509 ( .A(n380), .B(a[25]), .Z(n381) );
  AND U510 ( .A(n382), .B(n381), .Z(n471) );
  XOR U511 ( .A(a[100]), .B(n384), .Z(n383) );
  XNOR U512 ( .A(b[100]), .B(n383), .Z(c[100]) );
  XOR U513 ( .A(a[101]), .B(n386), .Z(n385) );
  XNOR U514 ( .A(b[101]), .B(n385), .Z(c[101]) );
  XOR U515 ( .A(a[102]), .B(n388), .Z(n387) );
  XNOR U516 ( .A(b[102]), .B(n387), .Z(c[102]) );
  XOR U517 ( .A(a[103]), .B(n390), .Z(n389) );
  XNOR U518 ( .A(b[103]), .B(n389), .Z(c[103]) );
  XOR U519 ( .A(a[104]), .B(n392), .Z(n391) );
  XNOR U520 ( .A(b[104]), .B(n391), .Z(c[104]) );
  XOR U521 ( .A(a[105]), .B(n394), .Z(n393) );
  XNOR U522 ( .A(b[105]), .B(n393), .Z(c[105]) );
  XOR U523 ( .A(a[106]), .B(n396), .Z(n395) );
  XNOR U524 ( .A(b[106]), .B(n395), .Z(c[106]) );
  XOR U525 ( .A(a[107]), .B(n398), .Z(n397) );
  XNOR U526 ( .A(b[107]), .B(n397), .Z(c[107]) );
  XOR U527 ( .A(a[108]), .B(n400), .Z(n399) );
  XNOR U528 ( .A(b[108]), .B(n399), .Z(c[108]) );
  XOR U529 ( .A(a[109]), .B(n404), .Z(n401) );
  XNOR U530 ( .A(b[109]), .B(n401), .Z(c[109]) );
  XOR U531 ( .A(b[10]), .B(n402), .Z(n403) );
  XNOR U532 ( .A(a[10]), .B(n403), .Z(c[10]) );
  XOR U533 ( .A(a[110]), .B(n406), .Z(n405) );
  XNOR U534 ( .A(b[110]), .B(n405), .Z(c[110]) );
  XOR U535 ( .A(a[111]), .B(n408), .Z(n407) );
  XNOR U536 ( .A(b[111]), .B(n407), .Z(c[111]) );
  XOR U537 ( .A(a[112]), .B(n410), .Z(n409) );
  XNOR U538 ( .A(b[112]), .B(n409), .Z(c[112]) );
  XOR U539 ( .A(a[113]), .B(n412), .Z(n411) );
  XNOR U540 ( .A(b[113]), .B(n411), .Z(c[113]) );
  XOR U541 ( .A(a[114]), .B(n414), .Z(n413) );
  XNOR U542 ( .A(b[114]), .B(n413), .Z(c[114]) );
  XOR U543 ( .A(a[115]), .B(n416), .Z(n415) );
  XNOR U544 ( .A(b[115]), .B(n415), .Z(c[115]) );
  XOR U545 ( .A(a[116]), .B(n418), .Z(n417) );
  XNOR U546 ( .A(b[116]), .B(n417), .Z(c[116]) );
  XOR U547 ( .A(a[117]), .B(n420), .Z(n419) );
  XNOR U548 ( .A(b[117]), .B(n419), .Z(c[117]) );
  XOR U549 ( .A(a[118]), .B(n422), .Z(n421) );
  XNOR U550 ( .A(b[118]), .B(n421), .Z(c[118]) );
  XOR U551 ( .A(a[119]), .B(n426), .Z(n423) );
  XNOR U552 ( .A(b[119]), .B(n423), .Z(c[119]) );
  XOR U553 ( .A(b[11]), .B(n424), .Z(n425) );
  XNOR U554 ( .A(a[11]), .B(n425), .Z(c[11]) );
  XOR U555 ( .A(a[120]), .B(n428), .Z(n427) );
  XNOR U556 ( .A(b[120]), .B(n427), .Z(c[120]) );
  XOR U557 ( .A(a[121]), .B(n430), .Z(n429) );
  XNOR U558 ( .A(b[121]), .B(n429), .Z(c[121]) );
  XOR U559 ( .A(a[122]), .B(n432), .Z(n431) );
  XNOR U560 ( .A(b[122]), .B(n431), .Z(c[122]) );
  XOR U561 ( .A(a[123]), .B(n434), .Z(n433) );
  XNOR U562 ( .A(b[123]), .B(n433), .Z(c[123]) );
  XOR U563 ( .A(a[124]), .B(n436), .Z(n435) );
  XNOR U564 ( .A(b[124]), .B(n435), .Z(c[124]) );
  XOR U565 ( .A(a[125]), .B(n438), .Z(n437) );
  XNOR U566 ( .A(b[125]), .B(n437), .Z(c[125]) );
  XOR U567 ( .A(a[126]), .B(n440), .Z(n439) );
  XNOR U568 ( .A(b[126]), .B(n439), .Z(c[126]) );
  XOR U569 ( .A(b[12]), .B(n441), .Z(n442) );
  XNOR U570 ( .A(a[12]), .B(n442), .Z(c[12]) );
  XOR U571 ( .A(b[13]), .B(n443), .Z(n444) );
  XNOR U572 ( .A(a[13]), .B(n444), .Z(c[13]) );
  XOR U573 ( .A(b[14]), .B(n445), .Z(n446) );
  XNOR U574 ( .A(a[14]), .B(n446), .Z(c[14]) );
  XOR U575 ( .A(b[15]), .B(n447), .Z(n448) );
  XNOR U576 ( .A(a[15]), .B(n448), .Z(c[15]) );
  XOR U577 ( .A(b[16]), .B(n449), .Z(n450) );
  XNOR U578 ( .A(a[16]), .B(n450), .Z(c[16]) );
  XOR U579 ( .A(b[17]), .B(n451), .Z(n452) );
  XNOR U580 ( .A(a[17]), .B(n452), .Z(c[17]) );
  XOR U581 ( .A(b[18]), .B(n453), .Z(n454) );
  XNOR U582 ( .A(a[18]), .B(n454), .Z(c[18]) );
  XOR U583 ( .A(b[19]), .B(n455), .Z(n456) );
  XNOR U584 ( .A(a[19]), .B(n456), .Z(c[19]) );
  XOR U585 ( .A(a[1]), .B(b[1]), .Z(n457) );
  XNOR U586 ( .A(n458), .B(n457), .Z(c[1]) );
  XOR U587 ( .A(b[20]), .B(n459), .Z(n460) );
  XNOR U588 ( .A(a[20]), .B(n460), .Z(c[20]) );
  XOR U589 ( .A(b[21]), .B(n461), .Z(n462) );
  XNOR U590 ( .A(a[21]), .B(n462), .Z(c[21]) );
  XOR U591 ( .A(b[22]), .B(n463), .Z(n464) );
  XNOR U592 ( .A(a[22]), .B(n464), .Z(c[22]) );
  XOR U593 ( .A(b[23]), .B(n465), .Z(n466) );
  XNOR U594 ( .A(a[23]), .B(n466), .Z(c[23]) );
  XOR U595 ( .A(b[24]), .B(n467), .Z(n468) );
  XNOR U596 ( .A(a[24]), .B(n468), .Z(c[24]) );
  XNOR U597 ( .A(b[25]), .B(a[25]), .Z(n469) );
  XNOR U598 ( .A(n470), .B(n469), .Z(c[25]) );
  XOR U599 ( .A(b[26]), .B(n471), .Z(n472) );
  XNOR U600 ( .A(a[26]), .B(n472), .Z(c[26]) );
  XOR U601 ( .A(b[27]), .B(n473), .Z(n474) );
  XNOR U602 ( .A(a[27]), .B(n474), .Z(c[27]) );
  XOR U603 ( .A(b[28]), .B(n475), .Z(n476) );
  XNOR U604 ( .A(a[28]), .B(n476), .Z(c[28]) );
  XOR U605 ( .A(b[29]), .B(n477), .Z(n478) );
  XNOR U606 ( .A(a[29]), .B(n478), .Z(c[29]) );
  XOR U607 ( .A(b[2]), .B(n479), .Z(n480) );
  XNOR U608 ( .A(a[2]), .B(n480), .Z(c[2]) );
  XOR U609 ( .A(b[30]), .B(n481), .Z(n482) );
  XNOR U610 ( .A(a[30]), .B(n482), .Z(c[30]) );
  XOR U611 ( .A(b[31]), .B(n483), .Z(n484) );
  XNOR U612 ( .A(a[31]), .B(n484), .Z(c[31]) );
  XOR U613 ( .A(b[32]), .B(n485), .Z(n486) );
  XNOR U614 ( .A(a[32]), .B(n486), .Z(c[32]) );
  XOR U615 ( .A(b[33]), .B(n487), .Z(n488) );
  XNOR U616 ( .A(a[33]), .B(n488), .Z(c[33]) );
  XOR U617 ( .A(b[34]), .B(n489), .Z(n490) );
  XNOR U618 ( .A(a[34]), .B(n490), .Z(c[34]) );
  XOR U619 ( .A(b[35]), .B(n491), .Z(n492) );
  XNOR U620 ( .A(a[35]), .B(n492), .Z(c[35]) );
  XOR U621 ( .A(b[36]), .B(n493), .Z(n494) );
  XNOR U622 ( .A(a[36]), .B(n494), .Z(c[36]) );
  XOR U623 ( .A(b[37]), .B(n495), .Z(n496) );
  XNOR U624 ( .A(a[37]), .B(n496), .Z(c[37]) );
  XOR U625 ( .A(b[38]), .B(n497), .Z(n498) );
  XNOR U626 ( .A(a[38]), .B(n498), .Z(c[38]) );
  XOR U627 ( .A(b[39]), .B(n499), .Z(n500) );
  XNOR U628 ( .A(a[39]), .B(n500), .Z(c[39]) );
  XOR U629 ( .A(b[3]), .B(n501), .Z(n502) );
  XNOR U630 ( .A(a[3]), .B(n502), .Z(c[3]) );
  XOR U631 ( .A(b[40]), .B(n503), .Z(n504) );
  XNOR U632 ( .A(a[40]), .B(n504), .Z(c[40]) );
  XOR U633 ( .A(b[41]), .B(n505), .Z(n506) );
  XNOR U634 ( .A(a[41]), .B(n506), .Z(c[41]) );
  XOR U635 ( .A(b[42]), .B(n507), .Z(n508) );
  XNOR U636 ( .A(a[42]), .B(n508), .Z(c[42]) );
  XOR U637 ( .A(b[43]), .B(n509), .Z(n510) );
  XNOR U638 ( .A(a[43]), .B(n510), .Z(c[43]) );
  XOR U639 ( .A(b[44]), .B(n511), .Z(n512) );
  XNOR U640 ( .A(a[44]), .B(n512), .Z(c[44]) );
  XOR U641 ( .A(b[45]), .B(n513), .Z(n514) );
  XNOR U642 ( .A(a[45]), .B(n514), .Z(c[45]) );
  XOR U643 ( .A(b[46]), .B(n515), .Z(n516) );
  XNOR U644 ( .A(a[46]), .B(n516), .Z(c[46]) );
  XOR U645 ( .A(b[47]), .B(n517), .Z(n518) );
  XNOR U646 ( .A(a[47]), .B(n518), .Z(c[47]) );
  XOR U647 ( .A(b[48]), .B(n519), .Z(n520) );
  XNOR U648 ( .A(a[48]), .B(n520), .Z(c[48]) );
  XOR U649 ( .A(b[49]), .B(n521), .Z(n522) );
  XNOR U650 ( .A(a[49]), .B(n522), .Z(c[49]) );
  XOR U651 ( .A(b[4]), .B(n523), .Z(n524) );
  XNOR U652 ( .A(a[4]), .B(n524), .Z(c[4]) );
  XOR U653 ( .A(b[50]), .B(n525), .Z(n526) );
  XNOR U654 ( .A(a[50]), .B(n526), .Z(c[50]) );
  XOR U655 ( .A(b[51]), .B(n527), .Z(n528) );
  XNOR U656 ( .A(a[51]), .B(n528), .Z(c[51]) );
  XOR U657 ( .A(b[52]), .B(n529), .Z(n530) );
  XNOR U658 ( .A(a[52]), .B(n530), .Z(c[52]) );
  XOR U659 ( .A(b[53]), .B(n531), .Z(n532) );
  XNOR U660 ( .A(a[53]), .B(n532), .Z(c[53]) );
  XOR U661 ( .A(b[54]), .B(n533), .Z(n534) );
  XNOR U662 ( .A(a[54]), .B(n534), .Z(c[54]) );
  XOR U663 ( .A(b[55]), .B(n535), .Z(n536) );
  XNOR U664 ( .A(a[55]), .B(n536), .Z(c[55]) );
  XOR U665 ( .A(b[56]), .B(n537), .Z(n538) );
  XNOR U666 ( .A(a[56]), .B(n538), .Z(c[56]) );
  XOR U667 ( .A(b[57]), .B(n539), .Z(n540) );
  XNOR U668 ( .A(a[57]), .B(n540), .Z(c[57]) );
  XOR U669 ( .A(b[58]), .B(n541), .Z(n542) );
  XNOR U670 ( .A(a[58]), .B(n542), .Z(c[58]) );
  XOR U671 ( .A(b[59]), .B(n543), .Z(n544) );
  XNOR U672 ( .A(a[59]), .B(n544), .Z(c[59]) );
  XOR U673 ( .A(b[5]), .B(n545), .Z(n546) );
  XNOR U674 ( .A(a[5]), .B(n546), .Z(c[5]) );
  XOR U675 ( .A(b[60]), .B(n547), .Z(n548) );
  XNOR U676 ( .A(a[60]), .B(n548), .Z(c[60]) );
  XOR U677 ( .A(b[61]), .B(n549), .Z(n550) );
  XNOR U678 ( .A(a[61]), .B(n550), .Z(c[61]) );
  XOR U679 ( .A(b[62]), .B(n551), .Z(n552) );
  XNOR U680 ( .A(a[62]), .B(n552), .Z(c[62]) );
  XOR U681 ( .A(b[63]), .B(n553), .Z(n554) );
  XNOR U682 ( .A(a[63]), .B(n554), .Z(c[63]) );
  XOR U683 ( .A(b[64]), .B(n555), .Z(n556) );
  XNOR U684 ( .A(a[64]), .B(n556), .Z(c[64]) );
  XOR U685 ( .A(b[65]), .B(n557), .Z(n558) );
  XNOR U686 ( .A(a[65]), .B(n558), .Z(c[65]) );
  XOR U687 ( .A(b[66]), .B(n559), .Z(n560) );
  XNOR U688 ( .A(a[66]), .B(n560), .Z(c[66]) );
  XOR U689 ( .A(b[67]), .B(n561), .Z(n562) );
  XNOR U690 ( .A(a[67]), .B(n562), .Z(c[67]) );
  XOR U691 ( .A(b[68]), .B(n563), .Z(n564) );
  XNOR U692 ( .A(a[68]), .B(n564), .Z(c[68]) );
  XOR U693 ( .A(b[69]), .B(n565), .Z(n566) );
  XNOR U694 ( .A(a[69]), .B(n566), .Z(c[69]) );
  XOR U695 ( .A(b[6]), .B(n567), .Z(n568) );
  XNOR U696 ( .A(a[6]), .B(n568), .Z(c[6]) );
  XOR U697 ( .A(b[70]), .B(n569), .Z(n570) );
  XNOR U698 ( .A(a[70]), .B(n570), .Z(c[70]) );
  XOR U699 ( .A(b[71]), .B(n571), .Z(n572) );
  XNOR U700 ( .A(a[71]), .B(n572), .Z(c[71]) );
  XOR U701 ( .A(b[72]), .B(n573), .Z(n574) );
  XNOR U702 ( .A(a[72]), .B(n574), .Z(c[72]) );
  XOR U703 ( .A(b[73]), .B(n575), .Z(n576) );
  XNOR U704 ( .A(a[73]), .B(n576), .Z(c[73]) );
  XOR U705 ( .A(b[74]), .B(n577), .Z(n578) );
  XNOR U706 ( .A(a[74]), .B(n578), .Z(c[74]) );
  XOR U707 ( .A(b[75]), .B(n579), .Z(n580) );
  XNOR U708 ( .A(a[75]), .B(n580), .Z(c[75]) );
  XOR U709 ( .A(b[76]), .B(n581), .Z(n582) );
  XNOR U710 ( .A(a[76]), .B(n582), .Z(c[76]) );
  XOR U711 ( .A(b[77]), .B(n583), .Z(n584) );
  XNOR U712 ( .A(a[77]), .B(n584), .Z(c[77]) );
  XOR U713 ( .A(b[78]), .B(n585), .Z(n586) );
  XNOR U714 ( .A(a[78]), .B(n586), .Z(c[78]) );
  XOR U715 ( .A(b[79]), .B(n587), .Z(n588) );
  XNOR U716 ( .A(a[79]), .B(n588), .Z(c[79]) );
  XOR U717 ( .A(b[7]), .B(n589), .Z(n590) );
  XNOR U718 ( .A(a[7]), .B(n590), .Z(c[7]) );
  XOR U719 ( .A(b[80]), .B(n591), .Z(n592) );
  XNOR U720 ( .A(a[80]), .B(n592), .Z(c[80]) );
  XOR U721 ( .A(b[81]), .B(n593), .Z(n594) );
  XNOR U722 ( .A(a[81]), .B(n594), .Z(c[81]) );
  XOR U723 ( .A(b[82]), .B(n595), .Z(n596) );
  XNOR U724 ( .A(a[82]), .B(n596), .Z(c[82]) );
  XOR U725 ( .A(b[83]), .B(n597), .Z(n598) );
  XNOR U726 ( .A(a[83]), .B(n598), .Z(c[83]) );
  XOR U727 ( .A(b[84]), .B(n599), .Z(n600) );
  XNOR U728 ( .A(a[84]), .B(n600), .Z(c[84]) );
  XOR U729 ( .A(b[85]), .B(n601), .Z(n602) );
  XNOR U730 ( .A(a[85]), .B(n602), .Z(c[85]) );
  XOR U731 ( .A(b[86]), .B(n603), .Z(n604) );
  XNOR U732 ( .A(a[86]), .B(n604), .Z(c[86]) );
  XOR U733 ( .A(b[87]), .B(n605), .Z(n606) );
  XNOR U734 ( .A(a[87]), .B(n606), .Z(c[87]) );
  XOR U735 ( .A(b[88]), .B(n607), .Z(n608) );
  XNOR U736 ( .A(a[88]), .B(n608), .Z(c[88]) );
  XOR U737 ( .A(b[89]), .B(n609), .Z(n610) );
  XNOR U738 ( .A(a[89]), .B(n610), .Z(c[89]) );
  XOR U739 ( .A(b[8]), .B(n611), .Z(n612) );
  XNOR U740 ( .A(a[8]), .B(n612), .Z(c[8]) );
  XOR U741 ( .A(b[90]), .B(n613), .Z(n614) );
  XNOR U742 ( .A(a[90]), .B(n614), .Z(c[90]) );
  XOR U743 ( .A(b[91]), .B(n615), .Z(n616) );
  XNOR U744 ( .A(a[91]), .B(n616), .Z(c[91]) );
  XOR U745 ( .A(b[92]), .B(n617), .Z(n618) );
  XNOR U746 ( .A(a[92]), .B(n618), .Z(c[92]) );
  XOR U747 ( .A(b[93]), .B(n619), .Z(n620) );
  XNOR U748 ( .A(a[93]), .B(n620), .Z(c[93]) );
  XOR U749 ( .A(b[94]), .B(n621), .Z(n622) );
  XNOR U750 ( .A(a[94]), .B(n622), .Z(c[94]) );
  XOR U751 ( .A(b[95]), .B(n623), .Z(n624) );
  XNOR U752 ( .A(a[95]), .B(n624), .Z(c[95]) );
  XOR U753 ( .A(b[96]), .B(n625), .Z(n626) );
  XNOR U754 ( .A(a[96]), .B(n626), .Z(c[96]) );
  XOR U755 ( .A(b[97]), .B(n627), .Z(n628) );
  XNOR U756 ( .A(a[97]), .B(n628), .Z(c[97]) );
  XOR U757 ( .A(b[98]), .B(n629), .Z(n630) );
  XNOR U758 ( .A(a[98]), .B(n630), .Z(c[98]) );
  XOR U759 ( .A(a[99]), .B(n631), .Z(n632) );
  XNOR U760 ( .A(b[99]), .B(n632), .Z(c[99]) );
  XOR U761 ( .A(a[9]), .B(n633), .Z(n634) );
  XNOR U762 ( .A(b[9]), .B(n634), .Z(c[9]) );
endmodule

