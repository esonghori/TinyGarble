
module matrixMult_N_M_1_N3_M32 ( clk, rst, x, y, o );
  input [95:0] x;
  input [287:0] y;
  output [95:0] o;
  input clk, rst;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042;

  DFF \oi_reg[0][31]  ( .D(N64), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \oi_reg[0][30]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \oi_reg[0][29]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \oi_reg[0][28]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \oi_reg[0][27]  ( .D(N60), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \oi_reg[0][26]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \oi_reg[0][25]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \oi_reg[0][24]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \oi_reg[0][23]  ( .D(N56), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \oi_reg[0][22]  ( .D(N55), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \oi_reg[0][21]  ( .D(N54), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \oi_reg[0][20]  ( .D(N53), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \oi_reg[0][19]  ( .D(N52), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \oi_reg[0][18]  ( .D(N51), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \oi_reg[0][17]  ( .D(N50), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \oi_reg[0][16]  ( .D(N49), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \oi_reg[0][15]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \oi_reg[0][14]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \oi_reg[0][13]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \oi_reg[0][12]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \oi_reg[0][11]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \oi_reg[0][10]  ( .D(N43), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \oi_reg[0][9]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \oi_reg[0][8]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \oi_reg[0][7]  ( .D(N40), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \oi_reg[0][6]  ( .D(N39), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \oi_reg[0][5]  ( .D(N38), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \oi_reg[0][4]  ( .D(N37), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \oi_reg[0][3]  ( .D(N36), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \oi_reg[0][2]  ( .D(N35), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \oi_reg[0][1]  ( .D(N34), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \oi_reg[0][0]  ( .D(N33), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \oi_reg[1][31]  ( .D(N128), .CLK(clk), .RST(rst), .Q(o[63]) );
  DFF \oi_reg[1][30]  ( .D(N127), .CLK(clk), .RST(rst), .Q(o[62]) );
  DFF \oi_reg[1][29]  ( .D(N126), .CLK(clk), .RST(rst), .Q(o[61]) );
  DFF \oi_reg[1][28]  ( .D(N125), .CLK(clk), .RST(rst), .Q(o[60]) );
  DFF \oi_reg[1][27]  ( .D(N124), .CLK(clk), .RST(rst), .Q(o[59]) );
  DFF \oi_reg[1][26]  ( .D(N123), .CLK(clk), .RST(rst), .Q(o[58]) );
  DFF \oi_reg[1][25]  ( .D(N122), .CLK(clk), .RST(rst), .Q(o[57]) );
  DFF \oi_reg[1][24]  ( .D(N121), .CLK(clk), .RST(rst), .Q(o[56]) );
  DFF \oi_reg[1][23]  ( .D(N120), .CLK(clk), .RST(rst), .Q(o[55]) );
  DFF \oi_reg[1][22]  ( .D(N119), .CLK(clk), .RST(rst), .Q(o[54]) );
  DFF \oi_reg[1][21]  ( .D(N118), .CLK(clk), .RST(rst), .Q(o[53]) );
  DFF \oi_reg[1][20]  ( .D(N117), .CLK(clk), .RST(rst), .Q(o[52]) );
  DFF \oi_reg[1][19]  ( .D(N116), .CLK(clk), .RST(rst), .Q(o[51]) );
  DFF \oi_reg[1][18]  ( .D(N115), .CLK(clk), .RST(rst), .Q(o[50]) );
  DFF \oi_reg[1][17]  ( .D(N114), .CLK(clk), .RST(rst), .Q(o[49]) );
  DFF \oi_reg[1][16]  ( .D(N113), .CLK(clk), .RST(rst), .Q(o[48]) );
  DFF \oi_reg[1][15]  ( .D(N112), .CLK(clk), .RST(rst), .Q(o[47]) );
  DFF \oi_reg[1][14]  ( .D(N111), .CLK(clk), .RST(rst), .Q(o[46]) );
  DFF \oi_reg[1][13]  ( .D(N110), .CLK(clk), .RST(rst), .Q(o[45]) );
  DFF \oi_reg[1][12]  ( .D(N109), .CLK(clk), .RST(rst), .Q(o[44]) );
  DFF \oi_reg[1][11]  ( .D(N108), .CLK(clk), .RST(rst), .Q(o[43]) );
  DFF \oi_reg[1][10]  ( .D(N107), .CLK(clk), .RST(rst), .Q(o[42]) );
  DFF \oi_reg[1][9]  ( .D(N106), .CLK(clk), .RST(rst), .Q(o[41]) );
  DFF \oi_reg[1][8]  ( .D(N105), .CLK(clk), .RST(rst), .Q(o[40]) );
  DFF \oi_reg[1][7]  ( .D(N104), .CLK(clk), .RST(rst), .Q(o[39]) );
  DFF \oi_reg[1][6]  ( .D(N103), .CLK(clk), .RST(rst), .Q(o[38]) );
  DFF \oi_reg[1][5]  ( .D(N102), .CLK(clk), .RST(rst), .Q(o[37]) );
  DFF \oi_reg[1][4]  ( .D(N101), .CLK(clk), .RST(rst), .Q(o[36]) );
  DFF \oi_reg[1][3]  ( .D(N100), .CLK(clk), .RST(rst), .Q(o[35]) );
  DFF \oi_reg[1][2]  ( .D(N99), .CLK(clk), .RST(rst), .Q(o[34]) );
  DFF \oi_reg[1][1]  ( .D(N98), .CLK(clk), .RST(rst), .Q(o[33]) );
  DFF \oi_reg[1][0]  ( .D(N97), .CLK(clk), .RST(rst), .Q(o[32]) );
  DFF \oi_reg[2][31]  ( .D(N192), .CLK(clk), .RST(rst), .Q(o[95]) );
  DFF \oi_reg[2][30]  ( .D(N191), .CLK(clk), .RST(rst), .Q(o[94]) );
  DFF \oi_reg[2][29]  ( .D(N190), .CLK(clk), .RST(rst), .Q(o[93]) );
  DFF \oi_reg[2][28]  ( .D(N189), .CLK(clk), .RST(rst), .Q(o[92]) );
  DFF \oi_reg[2][27]  ( .D(N188), .CLK(clk), .RST(rst), .Q(o[91]) );
  DFF \oi_reg[2][26]  ( .D(N187), .CLK(clk), .RST(rst), .Q(o[90]) );
  DFF \oi_reg[2][25]  ( .D(N186), .CLK(clk), .RST(rst), .Q(o[89]) );
  DFF \oi_reg[2][24]  ( .D(N185), .CLK(clk), .RST(rst), .Q(o[88]) );
  DFF \oi_reg[2][23]  ( .D(N184), .CLK(clk), .RST(rst), .Q(o[87]) );
  DFF \oi_reg[2][22]  ( .D(N183), .CLK(clk), .RST(rst), .Q(o[86]) );
  DFF \oi_reg[2][21]  ( .D(N182), .CLK(clk), .RST(rst), .Q(o[85]) );
  DFF \oi_reg[2][20]  ( .D(N181), .CLK(clk), .RST(rst), .Q(o[84]) );
  DFF \oi_reg[2][19]  ( .D(N180), .CLK(clk), .RST(rst), .Q(o[83]) );
  DFF \oi_reg[2][18]  ( .D(N179), .CLK(clk), .RST(rst), .Q(o[82]) );
  DFF \oi_reg[2][17]  ( .D(N178), .CLK(clk), .RST(rst), .Q(o[81]) );
  DFF \oi_reg[2][16]  ( .D(N177), .CLK(clk), .RST(rst), .Q(o[80]) );
  DFF \oi_reg[2][15]  ( .D(N176), .CLK(clk), .RST(rst), .Q(o[79]) );
  DFF \oi_reg[2][14]  ( .D(N175), .CLK(clk), .RST(rst), .Q(o[78]) );
  DFF \oi_reg[2][13]  ( .D(N174), .CLK(clk), .RST(rst), .Q(o[77]) );
  DFF \oi_reg[2][12]  ( .D(N173), .CLK(clk), .RST(rst), .Q(o[76]) );
  DFF \oi_reg[2][11]  ( .D(N172), .CLK(clk), .RST(rst), .Q(o[75]) );
  DFF \oi_reg[2][10]  ( .D(N171), .CLK(clk), .RST(rst), .Q(o[74]) );
  DFF \oi_reg[2][9]  ( .D(N170), .CLK(clk), .RST(rst), .Q(o[73]) );
  DFF \oi_reg[2][8]  ( .D(N169), .CLK(clk), .RST(rst), .Q(o[72]) );
  DFF \oi_reg[2][7]  ( .D(N168), .CLK(clk), .RST(rst), .Q(o[71]) );
  DFF \oi_reg[2][6]  ( .D(N167), .CLK(clk), .RST(rst), .Q(o[70]) );
  DFF \oi_reg[2][5]  ( .D(N166), .CLK(clk), .RST(rst), .Q(o[69]) );
  DFF \oi_reg[2][4]  ( .D(N165), .CLK(clk), .RST(rst), .Q(o[68]) );
  DFF \oi_reg[2][3]  ( .D(N164), .CLK(clk), .RST(rst), .Q(o[67]) );
  DFF \oi_reg[2][2]  ( .D(N163), .CLK(clk), .RST(rst), .Q(o[66]) );
  DFF \oi_reg[2][1]  ( .D(N162), .CLK(clk), .RST(rst), .Q(o[65]) );
  DFF \oi_reg[2][0]  ( .D(N161), .CLK(clk), .RST(rst), .Q(o[64]) );
  XNOR U3 ( .A(n7527), .B(n7526), .Z(n7548) );
  XNOR U4 ( .A(n6421), .B(n6422), .Z(n6405) );
  XNOR U5 ( .A(n652), .B(n651), .Z(n643) );
  XNOR U6 ( .A(n1221), .B(n1220), .Z(n1227) );
  XNOR U7 ( .A(n5578), .B(n5579), .Z(n5571) );
  XOR U8 ( .A(n7807), .B(n7808), .Z(n7868) );
  XNOR U9 ( .A(n4296), .B(n4295), .Z(n4297) );
  XNOR U10 ( .A(n1068), .B(n1069), .Z(n1056) );
  XNOR U11 ( .A(n6405), .B(n6404), .Z(n6406) );
  XOR U12 ( .A(n6567), .B(n6568), .Z(n6559) );
  XNOR U13 ( .A(n7698), .B(n7699), .Z(n7631) );
  XOR U14 ( .A(n3441), .B(n3442), .Z(n3411) );
  XOR U15 ( .A(n3574), .B(n3575), .Z(n3562) );
  XOR U16 ( .A(n3663), .B(n3664), .Z(n3665) );
  XOR U17 ( .A(n587), .B(n588), .Z(n575) );
  XNOR U18 ( .A(n649), .B(n650), .Z(n652) );
  XNOR U19 ( .A(n757), .B(n758), .Z(n760) );
  XNOR U20 ( .A(n833), .B(n834), .Z(n835) );
  XNOR U21 ( .A(n1218), .B(n1219), .Z(n1221) );
  XNOR U22 ( .A(n2066), .B(n2067), .Z(n2069) );
  XNOR U23 ( .A(n7084), .B(n7085), .Z(n7012) );
  NAND U24 ( .A(n4436), .B(n3410), .Z(n1) );
  XOR U25 ( .A(n3410), .B(n4436), .Z(n2) );
  NANDN U26 ( .A(n3409), .B(n2), .Z(n3) );
  NAND U27 ( .A(n1), .B(n3), .Z(n3533) );
  XNOR U28 ( .A(n4660), .B(n4661), .Z(n4637) );
  XNOR U29 ( .A(n5323), .B(n5322), .Z(n5252) );
  XNOR U30 ( .A(n5329), .B(n5328), .Z(n5246) );
  XOR U31 ( .A(n2433), .B(n2434), .Z(n2535) );
  XNOR U32 ( .A(n5570), .B(n5571), .Z(n5573) );
  XOR U33 ( .A(n7439), .B(n7440), .Z(n7441) );
  XNOR U34 ( .A(n1458), .B(n1459), .Z(n1461) );
  XNOR U35 ( .A(n6343), .B(n6344), .Z(n6345) );
  XNOR U36 ( .A(n6919), .B(n6920), .Z(n6921) );
  XNOR U37 ( .A(n7262), .B(n7263), .Z(n7265) );
  XNOR U38 ( .A(n7316), .B(n7317), .Z(n7319) );
  XNOR U39 ( .A(n7516), .B(n7515), .Z(n7549) );
  XNOR U40 ( .A(n7848), .B(n7849), .Z(n7851) );
  XOR U41 ( .A(n7842), .B(n7843), .Z(n7844) );
  XOR U42 ( .A(n7880), .B(n7881), .Z(n7882) );
  XNOR U43 ( .A(n3348), .B(n3349), .Z(n3350) );
  XOR U44 ( .A(n3738), .B(n3739), .Z(n3776) );
  XNOR U45 ( .A(n3835), .B(n3834), .Z(n3836) );
  XOR U46 ( .A(n4289), .B(n4290), .Z(n4291) );
  XOR U47 ( .A(n4385), .B(n4386), .Z(n4387) );
  XNOR U48 ( .A(n4739), .B(n4738), .Z(n4696) );
  XNOR U49 ( .A(n4857), .B(n4858), .Z(n4860) );
  XNOR U50 ( .A(n947), .B(n946), .Z(n948) );
  XOR U51 ( .A(n996), .B(n997), .Z(n952) );
  XOR U52 ( .A(n1873), .B(n1874), .Z(n1875) );
  XOR U53 ( .A(n6368), .B(n6369), .Z(n6370) );
  XOR U54 ( .A(n7372), .B(n7373), .Z(n7364) );
  XNOR U55 ( .A(n7824), .B(n7825), .Z(n7827) );
  XNOR U56 ( .A(n8031), .B(n8032), .Z(n8034) );
  XNOR U57 ( .A(n3356), .B(n3590), .Z(n3373) );
  XOR U58 ( .A(n3453), .B(n3454), .Z(n3455) );
  XNOR U59 ( .A(n3556), .B(n3557), .Z(n3559) );
  XOR U60 ( .A(n3789), .B(n3790), .Z(n3791) );
  XOR U61 ( .A(n3647), .B(n3648), .Z(n3689) );
  XNOR U62 ( .A(n4283), .B(n4284), .Z(n4286) );
  XOR U63 ( .A(n4237), .B(n4238), .Z(n4240) );
  XNOR U64 ( .A(n4606), .B(n4607), .Z(n4598) );
  XNOR U65 ( .A(n427), .B(n1482), .Z(n428) );
  XNOR U66 ( .A(n515), .B(n516), .Z(n499) );
  XNOR U67 ( .A(n531), .B(n532), .Z(n526) );
  XOR U68 ( .A(n660), .B(n661), .Z(n697) );
  XOR U69 ( .A(n751), .B(n752), .Z(n753) );
  XNOR U70 ( .A(n760), .B(n759), .Z(n775) );
  XOR U71 ( .A(n1224), .B(n1225), .Z(n1226) );
  XNOR U72 ( .A(n1188), .B(n1189), .Z(n1220) );
  XNOR U73 ( .A(n1230), .B(n1231), .Z(n1233) );
  XNOR U74 ( .A(n1312), .B(n1313), .Z(n1315) );
  XNOR U75 ( .A(n1410), .B(n1411), .Z(n1403) );
  XNOR U76 ( .A(n6529), .B(n6530), .Z(n6532) );
  XNOR U77 ( .A(n6560), .B(n6559), .Z(n6561) );
  XNOR U78 ( .A(n7630), .B(n7631), .Z(n7641) );
  XNOR U79 ( .A(n7636), .B(n7637), .Z(n7646) );
  XOR U80 ( .A(n7836), .B(n7837), .Z(n7838) );
  XNOR U81 ( .A(n8200), .B(n8201), .Z(n8114) );
  NANDN U82 ( .A(n8080), .B(n8079), .Z(n4) );
  NANDN U83 ( .A(n8082), .B(n8081), .Z(n5) );
  NAND U84 ( .A(n4), .B(n5), .Z(n8326) );
  XOR U85 ( .A(n3502), .B(n3503), .Z(n3526) );
  XNOR U86 ( .A(n3636), .B(n3637), .Z(n3639) );
  XNOR U87 ( .A(n3796), .B(n3795), .Z(n3797) );
  XNOR U88 ( .A(n4118), .B(n4119), .Z(n4122) );
  XOR U89 ( .A(n4339), .B(n4340), .Z(n4331) );
  XOR U90 ( .A(n4481), .B(n4482), .Z(n4483) );
  XNOR U91 ( .A(n4642), .B(n4643), .Z(n4652) );
  XNOR U92 ( .A(n4636), .B(n4637), .Z(n4646) );
  XNOR U93 ( .A(n5314), .B(n5315), .Z(n5317) );
  XNOR U94 ( .A(n5320), .B(n5321), .Z(n5323) );
  XNOR U95 ( .A(n5326), .B(n5327), .Z(n5329) );
  XNOR U96 ( .A(n810), .B(n809), .Z(n811) );
  XOR U97 ( .A(n898), .B(n899), .Z(n900) );
  XNOR U98 ( .A(n830), .B(n829), .Z(n869) );
  XOR U99 ( .A(n1628), .B(n1629), .Z(n1514) );
  XNOR U100 ( .A(n1948), .B(n1949), .Z(n1951) );
  XOR U101 ( .A(n1855), .B(n1856), .Z(n1857) );
  XOR U102 ( .A(n2215), .B(n2216), .Z(n2217) );
  XNOR U103 ( .A(n2211), .B(n2212), .Z(n2125) );
  XOR U104 ( .A(n6157), .B(n6158), .Z(n6169) );
  XOR U105 ( .A(n6523), .B(n6524), .Z(n6525) );
  XNOR U106 ( .A(n7013), .B(n7012), .Z(n7108) );
  XNOR U107 ( .A(n8050), .B(n8049), .Z(n8051) );
  XOR U108 ( .A(n8442), .B(n8443), .Z(n8482) );
  NANDN U109 ( .A(n8276), .B(n8275), .Z(n6) );
  NANDN U110 ( .A(n8278), .B(n8277), .Z(n7) );
  NAND U111 ( .A(n6), .B(n7), .Z(n8507) );
  XNOR U112 ( .A(n3532), .B(n3533), .Z(n3535) );
  XOR U113 ( .A(n4104), .B(n4105), .Z(n4106) );
  XNOR U114 ( .A(n5534), .B(n5535), .Z(n5537) );
  XNOR U115 ( .A(n645), .B(n646), .Z(n715) );
  NANDN U116 ( .A(n2333), .B(n2332), .Z(n8) );
  NANDN U117 ( .A(n2331), .B(n2330), .Z(n9) );
  AND U118 ( .A(n8), .B(n9), .Z(n2526) );
  NANDN U119 ( .A(n2323), .B(n2322), .Z(n10) );
  NANDN U120 ( .A(n2325), .B(n2324), .Z(n11) );
  NAND U121 ( .A(n10), .B(n11), .Z(n2426) );
  XNOR U122 ( .A(n2656), .B(n2657), .Z(n2668) );
  XNOR U123 ( .A(n5572), .B(n5573), .Z(n5582) );
  XNOR U124 ( .A(n5784), .B(n5783), .Z(n5764) );
  XNOR U125 ( .A(n2680), .B(n2681), .Z(n2660) );
  NANDN U126 ( .A(n2532), .B(n2531), .Z(n12) );
  NANDN U127 ( .A(n2534), .B(n2533), .Z(n13) );
  NAND U128 ( .A(n12), .B(n13), .Z(n2565) );
  XNOR U129 ( .A(n3042), .B(n3043), .Z(n3039) );
  XNOR U130 ( .A(n1846), .B(n1845), .Z(n1902) );
  XNOR U131 ( .A(n7130), .B(n7131), .Z(n7133) );
  XNOR U132 ( .A(n7198), .B(n7199), .Z(n7201) );
  XOR U133 ( .A(n7447), .B(n7448), .Z(n7378) );
  XOR U134 ( .A(n7505), .B(n7506), .Z(n7507) );
  XOR U135 ( .A(n7562), .B(n7563), .Z(n7606) );
  XNOR U136 ( .A(n7566), .B(n7567), .Z(n7568) );
  XOR U137 ( .A(n7702), .B(n7703), .Z(n7704) );
  XOR U138 ( .A(n3819), .B(n3820), .Z(n3821) );
  XOR U139 ( .A(n3912), .B(n3913), .Z(n3914) );
  XOR U140 ( .A(n4175), .B(n4176), .Z(n4177) );
  XOR U141 ( .A(n4190), .B(n4313), .Z(n4157) );
  XNOR U142 ( .A(n4145), .B(n4146), .Z(n4164) );
  XOR U143 ( .A(n4393), .B(n4394), .Z(n4411) );
  XNOR U144 ( .A(n4554), .B(n4555), .Z(n4557) );
  XOR U145 ( .A(n4562), .B(n4563), .Z(n4575) );
  XNOR U146 ( .A(n4798), .B(n4797), .Z(n4891) );
  XOR U147 ( .A(n4865), .B(n4866), .Z(n4883) );
  XNOR U148 ( .A(n4937), .B(n4938), .Z(n4940) );
  XNOR U149 ( .A(n1081), .B(n1154), .Z(n1061) );
  XNOR U150 ( .A(n1461), .B(n1460), .Z(n1416) );
  XNOR U151 ( .A(n1605), .B(n1606), .Z(n1607) );
  XOR U152 ( .A(n1662), .B(n1663), .Z(n1664) );
  XNOR U153 ( .A(n1863), .B(n1864), .Z(n1801) );
  XNOR U154 ( .A(n1849), .B(n1850), .Z(n1852) );
  XOR U155 ( .A(n1867), .B(n1868), .Z(n1870) );
  XOR U156 ( .A(n2042), .B(n2043), .Z(n2044) );
  XOR U157 ( .A(n1980), .B(n1981), .Z(n2004) );
  XOR U158 ( .A(n2054), .B(n2055), .Z(n2056) );
  XOR U159 ( .A(n6415), .B(n6416), .Z(n6417) );
  XOR U160 ( .A(n6553), .B(n6554), .Z(n6555) );
  XNOR U161 ( .A(n6595), .B(n6596), .Z(n6598) );
  XOR U162 ( .A(n6668), .B(n6669), .Z(n6651) );
  XNOR U163 ( .A(n7235), .B(n7234), .Z(n7236) );
  XNOR U164 ( .A(n7463), .B(n7464), .Z(n7466) );
  XOR U165 ( .A(n7744), .B(n7745), .Z(n7746) );
  XNOR U166 ( .A(n7845), .B(n7844), .Z(n7774) );
  XOR U167 ( .A(n8109), .B(n8110), .Z(n8149) );
  XNOR U168 ( .A(n3374), .B(n3373), .Z(n3375) );
  XOR U169 ( .A(n3506), .B(n3507), .Z(n3500) );
  XNOR U170 ( .A(n3601), .B(n3600), .Z(n3602) );
  XOR U171 ( .A(n3768), .B(n3769), .Z(n3770) );
  XNOR U172 ( .A(n3660), .B(n3659), .Z(n3666) );
  XNOR U173 ( .A(n3690), .B(n3689), .Z(n3691) );
  XOR U174 ( .A(n4045), .B(n4046), .Z(n4034) );
  XNOR U175 ( .A(n4170), .B(n4169), .Z(n4171) );
  XNOR U176 ( .A(n4251), .B(n4252), .Z(n4243) );
  XNOR U177 ( .A(n4286), .B(n4285), .Z(n4239) );
  XNOR U178 ( .A(n4381), .B(n4382), .Z(n4374) );
  XOR U179 ( .A(n4403), .B(n4404), .Z(n4405) );
  XOR U180 ( .A(n4578), .B(n4579), .Z(n4580) );
  XNOR U181 ( .A(n4702), .B(n4703), .Z(n4673) );
  XOR U182 ( .A(n4810), .B(n4811), .Z(n4834) );
  XNOR U183 ( .A(n5345), .B(n5346), .Z(n5347) );
  XNOR U184 ( .A(n5198), .B(n5199), .Z(n5201) );
  XNOR U185 ( .A(n5167), .B(n5168), .Z(n5114) );
  XNOR U186 ( .A(n569), .B(n570), .Z(n572) );
  XNOR U187 ( .A(n614), .B(n613), .Z(n615) );
  XOR U188 ( .A(n673), .B(n672), .Z(n651) );
  XNOR U189 ( .A(n698), .B(n697), .Z(n699) );
  XOR U190 ( .A(n779), .B(n780), .Z(n759) );
  XOR U191 ( .A(n772), .B(n773), .Z(n774) );
  XNOR U192 ( .A(n827), .B(n828), .Z(n830) );
  XOR U193 ( .A(n985), .B(n986), .Z(n987) );
  XOR U194 ( .A(n940), .B(n941), .Z(n942) );
  XNOR U195 ( .A(n1056), .B(n1055), .Z(n1057) );
  XOR U196 ( .A(n1103), .B(n1104), .Z(n1105) );
  XOR U197 ( .A(n1266), .B(n1267), .Z(n1268) );
  XOR U198 ( .A(n1320), .B(n1321), .Z(n1354) );
  XNOR U199 ( .A(n1753), .B(n1754), .Z(n1756) );
  XNOR U200 ( .A(n1658), .B(n1659), .Z(n1768) );
  XNOR U201 ( .A(n1748), .B(n1979), .Z(n1700) );
  XOR U202 ( .A(n1705), .B(n1706), .Z(n1707) );
  XNOR U203 ( .A(n2016), .B(n2017), .Z(n2060) );
  OR U204 ( .A(n2038), .B(n2039), .Z(n14) );
  NAND U205 ( .A(n2040), .B(n2041), .Z(n15) );
  AND U206 ( .A(n14), .B(n15), .Z(n2132) );
  XOR U207 ( .A(n2120), .B(n2121), .Z(n2160) );
  XOR U208 ( .A(n6398), .B(n6399), .Z(n6400) );
  XNOR U209 ( .A(n6690), .B(n6691), .Z(n6693) );
  XOR U210 ( .A(n6765), .B(n6766), .Z(n6720) );
  XOR U211 ( .A(n6928), .B(n6927), .Z(n6901) );
  XNOR U212 ( .A(n7330), .B(n7331), .Z(n7335) );
  XNOR U213 ( .A(n7588), .B(n7589), .Z(n7499) );
  XNOR U214 ( .A(n7768), .B(n7769), .Z(n7771) );
  XOR U215 ( .A(n7886), .B(n7887), .Z(n7889) );
  XOR U216 ( .A(n8448), .B(n8449), .Z(n8496) );
  XNOR U217 ( .A(n3340), .B(n3339), .Z(n3380) );
  XOR U218 ( .A(n3403), .B(n3404), .Z(n3405) );
  XNOR U219 ( .A(n3563), .B(n3562), .Z(n3564) );
  XNOR U220 ( .A(n3815), .B(n3816), .Z(n3843) );
  XNOR U221 ( .A(n3727), .B(n3728), .Z(n3720) );
  XNOR U222 ( .A(n4841), .B(n4842), .Z(n4898) );
  XOR U223 ( .A(n5043), .B(n5044), .Z(n4913) );
  XNOR U224 ( .A(n4981), .B(n4982), .Z(n5036) );
  NAND U225 ( .A(n5110), .B(n5109), .Z(n16) );
  NANDN U226 ( .A(n5108), .B(n5107), .Z(n17) );
  AND U227 ( .A(n16), .B(n17), .Z(n5255) );
  XNOR U228 ( .A(n5317), .B(n5316), .Z(n5322) );
  XNOR U229 ( .A(n5298), .B(n5299), .Z(n5328) );
  XOR U230 ( .A(n429), .B(n428), .Z(n440) );
  XNOR U231 ( .A(n576), .B(n575), .Z(n577) );
  XNOR U232 ( .A(n741), .B(n742), .Z(n734) );
  XOR U233 ( .A(n1013), .B(n1014), .Z(n1015) );
  XOR U234 ( .A(n1037), .B(n1038), .Z(n1109) );
  XNOR U235 ( .A(n1362), .B(n1363), .Z(n1367) );
  XOR U236 ( .A(n1496), .B(n1497), .Z(n1498) );
  XOR U237 ( .A(n1906), .B(n1907), .Z(n1908) );
  XNOR U238 ( .A(n2445), .B(n2446), .Z(n2452) );
  XOR U239 ( .A(n2496), .B(n2497), .Z(n2415) );
  NANDN U240 ( .A(n2115), .B(n2114), .Z(n18) );
  NANDN U241 ( .A(n2117), .B(n2116), .Z(n19) );
  NAND U242 ( .A(n18), .B(n19), .Z(n2265) );
  XNOR U243 ( .A(n7469), .B(n7470), .Z(n7472) );
  XOR U244 ( .A(n7960), .B(n7961), .Z(n7916) );
  XNOR U245 ( .A(n8360), .B(n8361), .Z(n8363) );
  XNOR U246 ( .A(n8472), .B(n8473), .Z(n8485) );
  NANDN U247 ( .A(n8280), .B(n8279), .Z(n20) );
  NANDN U248 ( .A(n8282), .B(n8281), .Z(n21) );
  NAND U249 ( .A(n20), .B(n21), .Z(n8509) );
  NAND U250 ( .A(n8255), .B(n8256), .Z(n22) );
  NANDN U251 ( .A(n8254), .B(n8253), .Z(n23) );
  NAND U252 ( .A(n22), .B(n23), .Z(n8515) );
  NANDN U253 ( .A(n8286), .B(n8285), .Z(n24) );
  NANDN U254 ( .A(n8284), .B(n8283), .Z(n25) );
  AND U255 ( .A(n24), .B(n25), .Z(n8518) );
  XOR U256 ( .A(n8578), .B(n8579), .Z(n8661) );
  XNOR U257 ( .A(n8714), .B(n8715), .Z(n8719) );
  XNOR U258 ( .A(n8798), .B(n8799), .Z(n8796) );
  XNOR U259 ( .A(n8764), .B(n8765), .Z(n8763) );
  XNOR U260 ( .A(n3702), .B(n3701), .Z(n3703) );
  XOR U261 ( .A(n4957), .B(n4958), .Z(n4907) );
  XOR U262 ( .A(n5510), .B(n5511), .Z(n5512) );
  XOR U263 ( .A(n5516), .B(n5517), .Z(n5518) );
  XOR U264 ( .A(n5486), .B(n5487), .Z(n5488) );
  XOR U265 ( .A(n5480), .B(n5481), .Z(n5482) );
  XOR U266 ( .A(n5590), .B(n5591), .Z(n5668) );
  XNOR U267 ( .A(n5791), .B(n5792), .Z(n5789) );
  XOR U268 ( .A(n393), .B(n394), .Z(n344) );
  XNOR U269 ( .A(n487), .B(n488), .Z(n480) );
  XNOR U270 ( .A(n716), .B(n715), .Z(n717) );
  XOR U271 ( .A(n922), .B(n923), .Z(n924) );
  XOR U272 ( .A(n1384), .B(n1385), .Z(n1386) );
  XNOR U273 ( .A(n1951), .B(n1950), .Z(n1936) );
  XNOR U274 ( .A(n2377), .B(n2378), .Z(n2380) );
  XNOR U275 ( .A(n2525), .B(n2526), .Z(n2528) );
  NAND U276 ( .A(n2302), .B(n2303), .Z(n26) );
  NANDN U277 ( .A(n2301), .B(n2300), .Z(n27) );
  NAND U278 ( .A(n26), .B(n27), .Z(n2434) );
  NAND U279 ( .A(n2328), .B(n2329), .Z(n28) );
  NANDN U280 ( .A(n2327), .B(n2326), .Z(n29) );
  NAND U281 ( .A(n28), .B(n29), .Z(n2428) );
  XOR U282 ( .A(n2577), .B(n2578), .Z(n2657) );
  XNOR U283 ( .A(n2692), .B(n2693), .Z(n2715) );
  XNOR U284 ( .A(n2792), .B(n2793), .Z(n2790) );
  XOR U285 ( .A(n2647), .B(n2646), .Z(n2673) );
  XNOR U286 ( .A(n2778), .B(n2779), .Z(n2777) );
  NAND U287 ( .A(n6103), .B(n6073), .Z(n30) );
  XOR U288 ( .A(n6073), .B(n6103), .Z(n31) );
  NANDN U289 ( .A(n6074), .B(n31), .Z(n32) );
  NAND U290 ( .A(n30), .B(n32), .Z(n6085) );
  XOR U291 ( .A(n6090), .B(n6091), .Z(n6093) );
  XNOR U292 ( .A(n6224), .B(n6225), .Z(n6266) );
  XNOR U293 ( .A(n6326), .B(n6327), .Z(n6329) );
  XOR U294 ( .A(n6607), .B(n6608), .Z(n6609) );
  XNOR U295 ( .A(n6708), .B(n6709), .Z(n6711) );
  XNOR U296 ( .A(n7649), .B(n7648), .Z(n7624) );
  XNOR U297 ( .A(n7894), .B(n7895), .Z(n7765) );
  XNOR U298 ( .A(n8685), .B(n8686), .Z(n8668) );
  XNOR U299 ( .A(n8771), .B(n8770), .Z(n8745) );
  NANDN U300 ( .A(n8525), .B(n8524), .Z(n33) );
  NANDN U301 ( .A(n8527), .B(n8526), .Z(n34) );
  NAND U302 ( .A(n33), .B(n34), .Z(n8546) );
  NAND U303 ( .A(n3111), .B(n3081), .Z(n35) );
  XOR U304 ( .A(n3081), .B(n3111), .Z(n36) );
  NANDN U305 ( .A(n3082), .B(n36), .Z(n37) );
  NAND U306 ( .A(n35), .B(n37), .Z(n3093) );
  XOR U307 ( .A(n3098), .B(n3099), .Z(n3101) );
  XNOR U308 ( .A(n3305), .B(n3306), .Z(n3283) );
  XOR U309 ( .A(n3465), .B(n3466), .Z(n3467) );
  XOR U310 ( .A(n3612), .B(n3613), .Z(n3614) );
  XOR U311 ( .A(n4231), .B(n4232), .Z(n4233) );
  XNOR U312 ( .A(n4349), .B(n4350), .Z(n4352) );
  XOR U313 ( .A(n4493), .B(n4494), .Z(n4495) );
  XNOR U314 ( .A(n4655), .B(n4654), .Z(n4630) );
  XNOR U315 ( .A(n4903), .B(n4904), .Z(n4768) );
  XNOR U316 ( .A(n5692), .B(n5693), .Z(n5675) );
  XNOR U317 ( .A(n5777), .B(n5778), .Z(n5776) );
  NAND U318 ( .A(n121), .B(n91), .Z(n38) );
  XOR U319 ( .A(n91), .B(n121), .Z(n39) );
  NANDN U320 ( .A(n92), .B(n39), .Z(n40) );
  NAND U321 ( .A(n38), .B(n40), .Z(n103) );
  XNOR U322 ( .A(n316), .B(n317), .Z(n294) );
  XNOR U323 ( .A(n559), .B(n560), .Z(n628) );
  XOR U324 ( .A(n727), .B(n728), .Z(n729) );
  XOR U325 ( .A(n821), .B(n822), .Z(n823) );
  XOR U326 ( .A(n2078), .B(n2079), .Z(n2080) );
  XOR U327 ( .A(n2233), .B(n2234), .Z(n2235) );
  XNOR U328 ( .A(n3020), .B(n3021), .Z(n3019) );
  XNOR U329 ( .A(n2785), .B(n2784), .Z(n3005) );
  XNOR U330 ( .A(n6147), .B(n6148), .Z(n6142) );
  XNOR U331 ( .A(n7230), .B(n7231), .Z(n7225) );
  XNOR U332 ( .A(n8218), .B(n8219), .Z(n8213) );
  XNOR U333 ( .A(n3155), .B(n3156), .Z(n3150) );
  XNOR U334 ( .A(n5055), .B(n5056), .Z(n5050) );
  XNOR U335 ( .A(n5224), .B(n5225), .Z(n5219) );
  XOR U336 ( .A(n6032), .B(n6033), .Z(n5739) );
  XNOR U337 ( .A(n165), .B(n166), .Z(n160) );
  XNOR U338 ( .A(n1141), .B(n1142), .Z(n1136) );
  XNOR U339 ( .A(n1646), .B(n1647), .Z(n1641) );
  NAND U340 ( .A(n2568), .B(n2567), .Z(n41) );
  NANDN U341 ( .A(n2566), .B(n2565), .Z(n42) );
  AND U342 ( .A(n41), .B(n42), .Z(n3036) );
  IV U343 ( .A(y[195]), .Z(n43) );
  IV U344 ( .A(y[231]), .Z(n44) );
  IV U345 ( .A(x[64]), .Z(n45) );
  IV U346 ( .A(x[65]), .Z(n46) );
  IV U347 ( .A(x[66]), .Z(n47) );
  IV U348 ( .A(x[67]), .Z(n48) );
  IV U349 ( .A(x[68]), .Z(n49) );
  IV U350 ( .A(x[69]), .Z(n50) );
  IV U351 ( .A(x[70]), .Z(n51) );
  IV U352 ( .A(x[71]), .Z(n52) );
  IV U353 ( .A(x[72]), .Z(n53) );
  IV U354 ( .A(x[73]), .Z(n54) );
  IV U355 ( .A(x[74]), .Z(n55) );
  IV U356 ( .A(x[75]), .Z(n56) );
  IV U357 ( .A(x[76]), .Z(n57) );
  IV U358 ( .A(x[77]), .Z(n58) );
  IV U359 ( .A(x[78]), .Z(n59) );
  IV U360 ( .A(x[79]), .Z(n60) );
  IV U361 ( .A(x[82]), .Z(n61) );
  ANDN U362 ( .B(y[192]), .A(n45), .Z(n794) );
  XOR U363 ( .A(n794), .B(o[0]), .Z(N33) );
  ANDN U364 ( .B(y[192]), .A(n46), .Z(n62) );
  IV U365 ( .A(y[193]), .Z(n2857) );
  NANDN U366 ( .A(n2857), .B(x[64]), .Z(n68) );
  XNOR U367 ( .A(n68), .B(o[1]), .Z(n63) );
  XOR U368 ( .A(n62), .B(n63), .Z(n64) );
  AND U369 ( .A(o[0]), .B(n794), .Z(n65) );
  XOR U370 ( .A(n64), .B(n65), .Z(N34) );
  OR U371 ( .A(n63), .B(n62), .Z(n67) );
  NANDN U372 ( .A(n65), .B(n64), .Z(n66) );
  NAND U373 ( .A(n67), .B(n66), .Z(n70) );
  NANDN U374 ( .A(n45), .B(y[194]), .Z(n81) );
  XOR U375 ( .A(n81), .B(o[2]), .Z(n69) );
  XNOR U376 ( .A(n70), .B(n69), .Z(n72) );
  ANDN U377 ( .B(o[1]), .A(n68), .Z(n75) );
  AND U378 ( .A(x[66]), .B(y[192]), .Z(n76) );
  XNOR U379 ( .A(n75), .B(n76), .Z(n78) );
  AND U380 ( .A(x[65]), .B(y[193]), .Z(n77) );
  XNOR U381 ( .A(n78), .B(n77), .Z(n71) );
  XNOR U382 ( .A(n72), .B(n71), .Z(N35) );
  NAND U383 ( .A(n70), .B(n69), .Z(n74) );
  OR U384 ( .A(n72), .B(n71), .Z(n73) );
  NAND U385 ( .A(n74), .B(n73), .Z(n85) );
  OR U386 ( .A(n76), .B(n75), .Z(n80) );
  OR U387 ( .A(n78), .B(n77), .Z(n79) );
  AND U388 ( .A(n80), .B(n79), .Z(n86) );
  XNOR U389 ( .A(n85), .B(n86), .Z(n87) );
  NANDN U390 ( .A(n2857), .B(x[66]), .Z(n97) );
  XNOR U391 ( .A(n97), .B(o[3]), .Z(n91) );
  NANDN U392 ( .A(n81), .B(o[2]), .Z(n94) );
  ANDN U393 ( .B(x[64]), .A(n43), .Z(n83) );
  IV U394 ( .A(y[192]), .Z(n2902) );
  NANDN U395 ( .A(n2902), .B(x[67]), .Z(n82) );
  XOR U396 ( .A(n83), .B(n82), .Z(n93) );
  XNOR U397 ( .A(n94), .B(n93), .Z(n92) );
  AND U398 ( .A(x[65]), .B(y[194]), .Z(n121) );
  XOR U399 ( .A(n92), .B(n121), .Z(n84) );
  XOR U400 ( .A(n91), .B(n84), .Z(n88) );
  XNOR U401 ( .A(n87), .B(n88), .Z(N36) );
  NANDN U402 ( .A(n86), .B(n85), .Z(n90) );
  NAND U403 ( .A(n88), .B(n87), .Z(n89) );
  NAND U404 ( .A(n90), .B(n89), .Z(n102) );
  XNOR U405 ( .A(n102), .B(n103), .Z(n104) );
  AND U406 ( .A(y[195]), .B(x[67]), .Z(n169) );
  NAND U407 ( .A(n794), .B(n169), .Z(n96) );
  OR U408 ( .A(n94), .B(n93), .Z(n95) );
  NAND U409 ( .A(n96), .B(n95), .Z(n109) );
  NANDN U410 ( .A(n97), .B(o[3]), .Z(n118) );
  IV U411 ( .A(y[196]), .Z(n2897) );
  ANDN U412 ( .B(x[64]), .A(n2897), .Z(n99) );
  ANDN U413 ( .B(y[192]), .A(n49), .Z(n98) );
  XNOR U414 ( .A(n99), .B(n98), .Z(n117) );
  XOR U415 ( .A(n118), .B(n117), .Z(n108) );
  XNOR U416 ( .A(n109), .B(n108), .Z(n111) );
  ANDN U417 ( .B(y[195]), .A(n46), .Z(n101) );
  IV U418 ( .A(y[194]), .Z(n2602) );
  NANDN U419 ( .A(n2602), .B(x[66]), .Z(n100) );
  XOR U420 ( .A(n101), .B(n100), .Z(n123) );
  NANDN U421 ( .A(n2857), .B(x[67]), .Z(n114) );
  XNOR U422 ( .A(n114), .B(o[4]), .Z(n122) );
  XOR U423 ( .A(n123), .B(n122), .Z(n110) );
  XOR U424 ( .A(n111), .B(n110), .Z(n105) );
  XOR U425 ( .A(n104), .B(n105), .Z(N37) );
  NANDN U426 ( .A(n103), .B(n102), .Z(n107) );
  NANDN U427 ( .A(n105), .B(n104), .Z(n106) );
  NAND U428 ( .A(n107), .B(n106), .Z(n126) );
  NAND U429 ( .A(n109), .B(n108), .Z(n113) );
  OR U430 ( .A(n111), .B(n110), .Z(n112) );
  NAND U431 ( .A(n113), .B(n112), .Z(n127) );
  XNOR U432 ( .A(n126), .B(n127), .Z(n128) );
  NANDN U433 ( .A(n114), .B(o[4]), .Z(n145) );
  IV U434 ( .A(y[197]), .Z(n1746) );
  ANDN U435 ( .B(x[64]), .A(n1746), .Z(n116) );
  ANDN U436 ( .B(y[192]), .A(n50), .Z(n115) );
  XNOR U437 ( .A(n116), .B(n115), .Z(n144) );
  XOR U438 ( .A(n145), .B(n144), .Z(n140) );
  AND U439 ( .A(y[195]), .B(x[66]), .Z(n138) );
  AND U440 ( .A(x[65]), .B(y[196]), .Z(n153) );
  AND U441 ( .A(x[68]), .B(y[193]), .Z(n148) );
  XOR U442 ( .A(o[5]), .B(n148), .Z(n151) );
  AND U443 ( .A(x[67]), .B(y[194]), .Z(n152) );
  XNOR U444 ( .A(n151), .B(n152), .Z(n154) );
  XNOR U445 ( .A(n153), .B(n154), .Z(n139) );
  XNOR U446 ( .A(n138), .B(n139), .Z(n141) );
  XNOR U447 ( .A(n140), .B(n141), .Z(n135) );
  AND U448 ( .A(y[196]), .B(x[68]), .Z(n234) );
  NAND U449 ( .A(n794), .B(n234), .Z(n120) );
  OR U450 ( .A(n118), .B(n117), .Z(n119) );
  NAND U451 ( .A(n120), .B(n119), .Z(n133) );
  NAND U452 ( .A(n121), .B(n138), .Z(n125) );
  NANDN U453 ( .A(n123), .B(n122), .Z(n124) );
  NAND U454 ( .A(n125), .B(n124), .Z(n132) );
  XNOR U455 ( .A(n133), .B(n132), .Z(n134) );
  XNOR U456 ( .A(n135), .B(n134), .Z(n129) );
  XOR U457 ( .A(n128), .B(n129), .Z(N38) );
  NANDN U458 ( .A(n127), .B(n126), .Z(n131) );
  NANDN U459 ( .A(n129), .B(n128), .Z(n130) );
  NAND U460 ( .A(n131), .B(n130), .Z(n157) );
  OR U461 ( .A(n133), .B(n132), .Z(n137) );
  OR U462 ( .A(n135), .B(n134), .Z(n136) );
  AND U463 ( .A(n137), .B(n136), .Z(n158) );
  XNOR U464 ( .A(n157), .B(n158), .Z(n159) );
  OR U465 ( .A(n139), .B(n138), .Z(n143) );
  OR U466 ( .A(n141), .B(n140), .Z(n142) );
  AND U467 ( .A(n143), .B(n142), .Z(n163) );
  NANDN U468 ( .A(n50), .B(y[197]), .Z(n520) );
  NANDN U469 ( .A(n520), .B(n794), .Z(n147) );
  OR U470 ( .A(n145), .B(n144), .Z(n146) );
  NAND U471 ( .A(n147), .B(n146), .Z(n186) );
  NAND U472 ( .A(n148), .B(o[5]), .Z(n176) );
  ANDN U473 ( .B(y[198]), .A(n45), .Z(n150) );
  ANDN U474 ( .B(y[192]), .A(n51), .Z(n149) );
  XNOR U475 ( .A(n150), .B(n149), .Z(n175) );
  XOR U476 ( .A(n176), .B(n175), .Z(n185) );
  XNOR U477 ( .A(n186), .B(n185), .Z(n188) );
  ANDN U478 ( .B(y[193]), .A(n50), .Z(n179) );
  XNOR U479 ( .A(o[6]), .B(n179), .Z(n180) );
  ANDN U480 ( .B(y[197]), .A(n46), .Z(n456) );
  XOR U481 ( .A(n180), .B(n456), .Z(n182) );
  ANDN U482 ( .B(x[68]), .A(n2602), .Z(n181) );
  XOR U483 ( .A(n182), .B(n181), .Z(n170) );
  ANDN U484 ( .B(x[66]), .A(n2897), .Z(n503) );
  XNOR U485 ( .A(n169), .B(n503), .Z(n171) );
  XOR U486 ( .A(n170), .B(n171), .Z(n187) );
  XNOR U487 ( .A(n188), .B(n187), .Z(n164) );
  XNOR U488 ( .A(n163), .B(n164), .Z(n165) );
  OR U489 ( .A(n152), .B(n151), .Z(n156) );
  OR U490 ( .A(n154), .B(n153), .Z(n155) );
  AND U491 ( .A(n156), .B(n155), .Z(n166) );
  XOR U492 ( .A(n159), .B(n160), .Z(N39) );
  NANDN U493 ( .A(n158), .B(n157), .Z(n162) );
  NANDN U494 ( .A(n160), .B(n159), .Z(n161) );
  NAND U495 ( .A(n162), .B(n161), .Z(n222) );
  OR U496 ( .A(n164), .B(n163), .Z(n168) );
  OR U497 ( .A(n166), .B(n165), .Z(n167) );
  AND U498 ( .A(n168), .B(n167), .Z(n223) );
  XNOR U499 ( .A(n222), .B(n223), .Z(n224) );
  OR U500 ( .A(n169), .B(n503), .Z(n173) );
  NANDN U501 ( .A(n171), .B(n170), .Z(n172) );
  NAND U502 ( .A(n173), .B(n172), .Z(n219) );
  IV U503 ( .A(y[198]), .Z(n2651) );
  ANDN U504 ( .B(x[70]), .A(n2651), .Z(n174) );
  NAND U505 ( .A(n794), .B(n174), .Z(n178) );
  OR U506 ( .A(n176), .B(n175), .Z(n177) );
  AND U507 ( .A(n178), .B(n177), .Z(n217) );
  ANDN U508 ( .B(x[65]), .A(n2651), .Z(n585) );
  NANDN U509 ( .A(n2857), .B(x[70]), .Z(n203) );
  XNOR U510 ( .A(o[7]), .B(n203), .Z(n206) );
  XNOR U511 ( .A(n585), .B(n206), .Z(n207) );
  AND U512 ( .A(y[194]), .B(x[69]), .Z(n364) );
  XNOR U513 ( .A(n207), .B(n364), .Z(n216) );
  XOR U514 ( .A(n217), .B(n216), .Z(n218) );
  XNOR U515 ( .A(n219), .B(n218), .Z(n228) );
  AND U516 ( .A(x[66]), .B(y[197]), .Z(n676) );
  AND U517 ( .A(y[196]), .B(x[67]), .Z(n199) );
  AND U518 ( .A(y[195]), .B(x[68]), .Z(n375) );
  XNOR U519 ( .A(n199), .B(n375), .Z(n200) );
  XOR U520 ( .A(n676), .B(n200), .Z(n210) );
  IV U521 ( .A(y[199]), .Z(n2878) );
  NANDN U522 ( .A(n2878), .B(x[64]), .Z(n196) );
  AND U523 ( .A(n179), .B(o[6]), .Z(n194) );
  NANDN U524 ( .A(n52), .B(y[192]), .Z(n193) );
  XNOR U525 ( .A(n194), .B(n193), .Z(n195) );
  XOR U526 ( .A(n196), .B(n195), .Z(n211) );
  XNOR U527 ( .A(n210), .B(n211), .Z(n213) );
  NANDN U528 ( .A(n180), .B(n456), .Z(n184) );
  NANDN U529 ( .A(n182), .B(n181), .Z(n183) );
  AND U530 ( .A(n184), .B(n183), .Z(n212) );
  XOR U531 ( .A(n213), .B(n212), .Z(n229) );
  XOR U532 ( .A(n228), .B(n229), .Z(n231) );
  OR U533 ( .A(n186), .B(n185), .Z(n190) );
  OR U534 ( .A(n188), .B(n187), .Z(n189) );
  AND U535 ( .A(n190), .B(n189), .Z(n230) );
  XOR U536 ( .A(n231), .B(n230), .Z(n225) );
  XNOR U537 ( .A(n224), .B(n225), .Z(N40) );
  IV U538 ( .A(y[200]), .Z(n2512) );
  ANDN U539 ( .B(x[64]), .A(n2512), .Z(n192) );
  NANDN U540 ( .A(n2902), .B(x[72]), .Z(n191) );
  XOR U541 ( .A(n192), .B(n191), .Z(n247) );
  NANDN U542 ( .A(n2857), .B(x[71]), .Z(n250) );
  XNOR U543 ( .A(n250), .B(o[8]), .Z(n246) );
  XOR U544 ( .A(n247), .B(n246), .Z(n269) );
  NANDN U545 ( .A(n194), .B(n193), .Z(n198) );
  NAND U546 ( .A(n196), .B(n195), .Z(n197) );
  NAND U547 ( .A(n198), .B(n197), .Z(n268) );
  XOR U548 ( .A(n269), .B(n268), .Z(n270) );
  OR U549 ( .A(n375), .B(n199), .Z(n202) );
  OR U550 ( .A(n200), .B(n676), .Z(n201) );
  NAND U551 ( .A(n202), .B(n201), .Z(n271) );
  XNOR U552 ( .A(n270), .B(n271), .Z(n282) );
  AND U553 ( .A(x[70]), .B(y[194]), .Z(n235) );
  XNOR U554 ( .A(n234), .B(n235), .Z(n237) );
  ANDN U555 ( .B(y[198]), .A(n47), .Z(n236) );
  IV U556 ( .A(n236), .Z(n804) );
  XOR U557 ( .A(n237), .B(n804), .Z(n240) );
  AND U558 ( .A(x[67]), .B(y[197]), .Z(n1080) );
  XNOR U559 ( .A(n240), .B(n1080), .Z(n242) );
  NANDN U560 ( .A(n203), .B(o[7]), .Z(n259) );
  ANDN U561 ( .B(y[199]), .A(n46), .Z(n205) );
  ANDN U562 ( .B(x[69]), .A(n43), .Z(n204) );
  XNOR U563 ( .A(n205), .B(n204), .Z(n258) );
  XOR U564 ( .A(n259), .B(n258), .Z(n241) );
  XNOR U565 ( .A(n242), .B(n241), .Z(n262) );
  NAND U566 ( .A(n585), .B(n206), .Z(n209) );
  NANDN U567 ( .A(n207), .B(n364), .Z(n208) );
  AND U568 ( .A(n209), .B(n208), .Z(n263) );
  XOR U569 ( .A(n262), .B(n263), .Z(n265) );
  OR U570 ( .A(n211), .B(n210), .Z(n215) );
  OR U571 ( .A(n213), .B(n212), .Z(n214) );
  AND U572 ( .A(n215), .B(n214), .Z(n264) );
  XOR U573 ( .A(n265), .B(n264), .Z(n280) );
  NANDN U574 ( .A(n217), .B(n216), .Z(n221) );
  OR U575 ( .A(n219), .B(n218), .Z(n220) );
  NAND U576 ( .A(n221), .B(n220), .Z(n281) );
  XNOR U577 ( .A(n280), .B(n281), .Z(n283) );
  XNOR U578 ( .A(n282), .B(n283), .Z(n277) );
  NANDN U579 ( .A(n223), .B(n222), .Z(n227) );
  NAND U580 ( .A(n225), .B(n224), .Z(n226) );
  NAND U581 ( .A(n227), .B(n226), .Z(n274) );
  NANDN U582 ( .A(n229), .B(n228), .Z(n233) );
  OR U583 ( .A(n231), .B(n230), .Z(n232) );
  AND U584 ( .A(n233), .B(n232), .Z(n275) );
  XNOR U585 ( .A(n274), .B(n275), .Z(n276) );
  XOR U586 ( .A(n277), .B(n276), .Z(N41) );
  OR U587 ( .A(n235), .B(n234), .Z(n239) );
  OR U588 ( .A(n237), .B(n236), .Z(n238) );
  NAND U589 ( .A(n239), .B(n238), .Z(n315) );
  OR U590 ( .A(n240), .B(n1080), .Z(n244) );
  OR U591 ( .A(n242), .B(n241), .Z(n243) );
  NAND U592 ( .A(n244), .B(n243), .Z(n314) );
  XNOR U593 ( .A(n315), .B(n314), .Z(n316) );
  ANDN U594 ( .B(y[200]), .A(n53), .Z(n245) );
  NAND U595 ( .A(n794), .B(n245), .Z(n249) );
  NANDN U596 ( .A(n247), .B(n246), .Z(n248) );
  NAND U597 ( .A(n249), .B(n248), .Z(n301) );
  NANDN U598 ( .A(n250), .B(o[8]), .Z(n335) );
  ANDN U599 ( .B(y[194]), .A(n52), .Z(n252) );
  ANDN U600 ( .B(x[69]), .A(n2897), .Z(n251) );
  XNOR U601 ( .A(n252), .B(n251), .Z(n334) );
  XOR U602 ( .A(n335), .B(n334), .Z(n299) );
  IV U603 ( .A(y[201]), .Z(n2837) );
  ANDN U604 ( .B(x[64]), .A(n2837), .Z(n254) );
  NANDN U605 ( .A(n2902), .B(x[73]), .Z(n253) );
  XOR U606 ( .A(n254), .B(n253), .Z(n327) );
  NANDN U607 ( .A(n2857), .B(x[72]), .Z(n320) );
  XOR U608 ( .A(n320), .B(o[9]), .Z(n326) );
  XNOR U609 ( .A(n327), .B(n326), .Z(n298) );
  XOR U610 ( .A(n299), .B(n298), .Z(n300) );
  XNOR U611 ( .A(n301), .B(n300), .Z(n310) );
  ANDN U612 ( .B(y[197]), .A(n49), .Z(n783) );
  ANDN U613 ( .B(y[195]), .A(n51), .Z(n256) );
  ANDN U614 ( .B(y[200]), .A(n46), .Z(n255) );
  XNOR U615 ( .A(n256), .B(n255), .Z(n322) );
  XNOR U616 ( .A(n783), .B(n322), .Z(n304) );
  AND U617 ( .A(x[66]), .B(y[199]), .Z(n1000) );
  NANDN U618 ( .A(n48), .B(y[198]), .Z(n655) );
  XOR U619 ( .A(n1000), .B(n655), .Z(n305) );
  XNOR U620 ( .A(n304), .B(n305), .Z(n308) );
  NANDN U621 ( .A(n43), .B(x[65]), .Z(n321) );
  ANDN U622 ( .B(y[199]), .A(n50), .Z(n257) );
  NANDN U623 ( .A(n321), .B(n257), .Z(n261) );
  OR U624 ( .A(n259), .B(n258), .Z(n260) );
  AND U625 ( .A(n261), .B(n260), .Z(n309) );
  XOR U626 ( .A(n308), .B(n309), .Z(n311) );
  XOR U627 ( .A(n310), .B(n311), .Z(n317) );
  NANDN U628 ( .A(n263), .B(n262), .Z(n267) );
  OR U629 ( .A(n265), .B(n264), .Z(n266) );
  NAND U630 ( .A(n267), .B(n266), .Z(n293) );
  OR U631 ( .A(n269), .B(n268), .Z(n273) );
  NANDN U632 ( .A(n271), .B(n270), .Z(n272) );
  NAND U633 ( .A(n273), .B(n272), .Z(n292) );
  XOR U634 ( .A(n293), .B(n292), .Z(n295) );
  XNOR U635 ( .A(n294), .B(n295), .Z(n289) );
  NANDN U636 ( .A(n275), .B(n274), .Z(n279) );
  NANDN U637 ( .A(n277), .B(n276), .Z(n278) );
  NAND U638 ( .A(n279), .B(n278), .Z(n286) );
  OR U639 ( .A(n281), .B(n280), .Z(n285) );
  OR U640 ( .A(n283), .B(n282), .Z(n284) );
  AND U641 ( .A(n285), .B(n284), .Z(n287) );
  XNOR U642 ( .A(n286), .B(n287), .Z(n288) );
  XOR U643 ( .A(n289), .B(n288), .Z(N42) );
  NANDN U644 ( .A(n287), .B(n286), .Z(n291) );
  NANDN U645 ( .A(n289), .B(n288), .Z(n290) );
  NAND U646 ( .A(n291), .B(n290), .Z(n338) );
  OR U647 ( .A(n293), .B(n292), .Z(n297) );
  NAND U648 ( .A(n295), .B(n294), .Z(n296) );
  AND U649 ( .A(n297), .B(n296), .Z(n339) );
  XNOR U650 ( .A(n338), .B(n339), .Z(n340) );
  NANDN U651 ( .A(n299), .B(n298), .Z(n303) );
  OR U652 ( .A(n301), .B(n300), .Z(n302) );
  NAND U653 ( .A(n303), .B(n302), .Z(n398) );
  NANDN U654 ( .A(n1000), .B(n655), .Z(n307) );
  OR U655 ( .A(n305), .B(n304), .Z(n306) );
  NAND U656 ( .A(n307), .B(n306), .Z(n397) );
  XOR U657 ( .A(n398), .B(n397), .Z(n399) );
  NANDN U658 ( .A(n309), .B(n308), .Z(n313) );
  NANDN U659 ( .A(n311), .B(n310), .Z(n312) );
  AND U660 ( .A(n313), .B(n312), .Z(n400) );
  XNOR U661 ( .A(n399), .B(n400), .Z(n346) );
  OR U662 ( .A(n315), .B(n314), .Z(n319) );
  OR U663 ( .A(n317), .B(n316), .Z(n318) );
  NAND U664 ( .A(n319), .B(n318), .Z(n345) );
  AND U665 ( .A(y[202]), .B(x[64]), .Z(n382) );
  ANDN U666 ( .B(o[9]), .A(n320), .Z(n380) );
  AND U667 ( .A(x[74]), .B(y[192]), .Z(n381) );
  XNOR U668 ( .A(n380), .B(n381), .Z(n383) );
  XOR U669 ( .A(n382), .B(n383), .Z(n371) );
  AND U670 ( .A(x[67]), .B(y[199]), .Z(n1331) );
  AND U671 ( .A(x[66]), .B(y[200]), .Z(n360) );
  XNOR U672 ( .A(n1331), .B(n360), .Z(n361) );
  AND U673 ( .A(x[65]), .B(y[201]), .Z(n1283) );
  XOR U674 ( .A(n361), .B(n1283), .Z(n369) );
  AND U675 ( .A(x[70]), .B(y[200]), .Z(n694) );
  NANDN U676 ( .A(n321), .B(n694), .Z(n324) );
  NANDN U677 ( .A(n322), .B(n783), .Z(n323) );
  AND U678 ( .A(n324), .B(n323), .Z(n370) );
  XNOR U679 ( .A(n369), .B(n370), .Z(n372) );
  XNOR U680 ( .A(n371), .B(n372), .Z(n391) );
  ANDN U681 ( .B(x[73]), .A(n2837), .Z(n325) );
  NAND U682 ( .A(n794), .B(n325), .Z(n329) );
  OR U683 ( .A(n327), .B(n326), .Z(n328) );
  NAND U684 ( .A(n329), .B(n328), .Z(n392) );
  XOR U685 ( .A(n391), .B(n392), .Z(n394) );
  ANDN U686 ( .B(x[72]), .A(n2602), .Z(n330) );
  XOR U687 ( .A(n330), .B(n520), .Z(n366) );
  NANDN U688 ( .A(n2857), .B(x[73]), .Z(n388) );
  XOR U689 ( .A(n388), .B(o[10]), .Z(n365) );
  XNOR U690 ( .A(n366), .B(n365), .Z(n350) );
  ANDN U691 ( .B(y[196]), .A(n51), .Z(n602) );
  ANDN U692 ( .B(y[195]), .A(n52), .Z(n332) );
  NANDN U693 ( .A(n49), .B(y[198]), .Z(n331) );
  XOR U694 ( .A(n332), .B(n331), .Z(n377) );
  XNOR U695 ( .A(n602), .B(n377), .Z(n351) );
  XOR U696 ( .A(n350), .B(n351), .Z(n353) );
  ANDN U697 ( .B(x[71]), .A(n2897), .Z(n333) );
  NAND U698 ( .A(n333), .B(n364), .Z(n337) );
  OR U699 ( .A(n335), .B(n334), .Z(n336) );
  NAND U700 ( .A(n337), .B(n336), .Z(n352) );
  XNOR U701 ( .A(n353), .B(n352), .Z(n393) );
  XOR U702 ( .A(n345), .B(n344), .Z(n347) );
  XNOR U703 ( .A(n346), .B(n347), .Z(n341) );
  XOR U704 ( .A(n340), .B(n341), .Z(N43) );
  NANDN U705 ( .A(n339), .B(n338), .Z(n343) );
  NANDN U706 ( .A(n341), .B(n340), .Z(n342) );
  NAND U707 ( .A(n343), .B(n342), .Z(n403) );
  NANDN U708 ( .A(n345), .B(n344), .Z(n349) );
  OR U709 ( .A(n347), .B(n346), .Z(n348) );
  AND U710 ( .A(n349), .B(n348), .Z(n404) );
  XNOR U711 ( .A(n403), .B(n404), .Z(n405) );
  NANDN U712 ( .A(n351), .B(n350), .Z(n355) );
  OR U713 ( .A(n353), .B(n352), .Z(n354) );
  NAND U714 ( .A(n355), .B(n354), .Z(n435) );
  ANDN U715 ( .B(y[196]), .A(n52), .Z(n357) );
  NANDN U716 ( .A(n54), .B(y[194]), .Z(n356) );
  XOR U717 ( .A(n357), .B(n356), .Z(n467) );
  NANDN U718 ( .A(n43), .B(x[72]), .Z(n466) );
  XNOR U719 ( .A(n467), .B(n466), .Z(n429) );
  AND U720 ( .A(x[67]), .B(y[200]), .Z(n1482) );
  NANDN U721 ( .A(n49), .B(y[199]), .Z(n453) );
  ANDN U722 ( .B(y[201]), .A(n47), .Z(n359) );
  ANDN U723 ( .B(x[69]), .A(n2651), .Z(n358) );
  XNOR U724 ( .A(n359), .B(n358), .Z(n452) );
  XNOR U725 ( .A(n453), .B(n452), .Z(n427) );
  OR U726 ( .A(n360), .B(n1331), .Z(n363) );
  OR U727 ( .A(n361), .B(n1283), .Z(n362) );
  AND U728 ( .A(n363), .B(n362), .Z(n438) );
  AND U729 ( .A(y[197]), .B(x[72]), .Z(n1208) );
  NAND U730 ( .A(n364), .B(n1208), .Z(n368) );
  OR U731 ( .A(n366), .B(n365), .Z(n367) );
  NAND U732 ( .A(n368), .B(n367), .Z(n439) );
  XNOR U733 ( .A(n438), .B(n439), .Z(n441) );
  XOR U734 ( .A(n440), .B(n441), .Z(n432) );
  OR U735 ( .A(n370), .B(n369), .Z(n374) );
  OR U736 ( .A(n372), .B(n371), .Z(n373) );
  NAND U737 ( .A(n374), .B(n373), .Z(n418) );
  ANDN U738 ( .B(x[71]), .A(n2651), .Z(n376) );
  NAND U739 ( .A(n376), .B(n375), .Z(n379) );
  NANDN U740 ( .A(n377), .B(n602), .Z(n378) );
  NAND U741 ( .A(n379), .B(n378), .Z(n416) );
  OR U742 ( .A(n381), .B(n380), .Z(n385) );
  OR U743 ( .A(n383), .B(n382), .Z(n384) );
  NAND U744 ( .A(n385), .B(n384), .Z(n424) );
  ANDN U745 ( .B(x[70]), .A(n1746), .Z(n387) );
  IV U746 ( .A(y[202]), .Z(n2906) );
  NANDN U747 ( .A(n2906), .B(x[65]), .Z(n386) );
  XOR U748 ( .A(n387), .B(n386), .Z(n459) );
  NANDN U749 ( .A(n2857), .B(x[74]), .Z(n470) );
  XOR U750 ( .A(n470), .B(o[11]), .Z(n458) );
  XNOR U751 ( .A(n459), .B(n458), .Z(n422) );
  NANDN U752 ( .A(n388), .B(o[10]), .Z(n463) );
  ANDN U753 ( .B(y[203]), .A(n45), .Z(n390) );
  NANDN U754 ( .A(n2902), .B(x[75]), .Z(n389) );
  XOR U755 ( .A(n390), .B(n389), .Z(n462) );
  XNOR U756 ( .A(n463), .B(n462), .Z(n421) );
  XOR U757 ( .A(n422), .B(n421), .Z(n423) );
  XNOR U758 ( .A(n424), .B(n423), .Z(n415) );
  XNOR U759 ( .A(n416), .B(n415), .Z(n417) );
  XNOR U760 ( .A(n418), .B(n417), .Z(n433) );
  XNOR U761 ( .A(n432), .B(n433), .Z(n434) );
  XNOR U762 ( .A(n435), .B(n434), .Z(n409) );
  NANDN U763 ( .A(n392), .B(n391), .Z(n396) );
  OR U764 ( .A(n394), .B(n393), .Z(n395) );
  AND U765 ( .A(n396), .B(n395), .Z(n410) );
  XOR U766 ( .A(n409), .B(n410), .Z(n412) );
  OR U767 ( .A(n398), .B(n397), .Z(n402) );
  NANDN U768 ( .A(n400), .B(n399), .Z(n401) );
  NAND U769 ( .A(n402), .B(n401), .Z(n411) );
  XOR U770 ( .A(n412), .B(n411), .Z(n406) );
  XNOR U771 ( .A(n405), .B(n406), .Z(N44) );
  NANDN U772 ( .A(n404), .B(n403), .Z(n408) );
  NAND U773 ( .A(n406), .B(n405), .Z(n407) );
  NAND U774 ( .A(n408), .B(n407), .Z(n473) );
  NANDN U775 ( .A(n410), .B(n409), .Z(n414) );
  OR U776 ( .A(n412), .B(n411), .Z(n413) );
  AND U777 ( .A(n414), .B(n413), .Z(n474) );
  XNOR U778 ( .A(n473), .B(n474), .Z(n475) );
  OR U779 ( .A(n416), .B(n415), .Z(n420) );
  OR U780 ( .A(n418), .B(n417), .Z(n419) );
  AND U781 ( .A(n420), .B(n419), .Z(n488) );
  OR U782 ( .A(n422), .B(n421), .Z(n426) );
  NANDN U783 ( .A(n424), .B(n423), .Z(n425) );
  NAND U784 ( .A(n426), .B(n425), .Z(n486) );
  NANDN U785 ( .A(n427), .B(n1482), .Z(n431) );
  NANDN U786 ( .A(n429), .B(n428), .Z(n430) );
  NAND U787 ( .A(n431), .B(n430), .Z(n485) );
  XNOR U788 ( .A(n486), .B(n485), .Z(n487) );
  NAND U789 ( .A(n433), .B(n432), .Z(n437) );
  OR U790 ( .A(n435), .B(n434), .Z(n436) );
  NAND U791 ( .A(n437), .B(n436), .Z(n479) );
  XNOR U792 ( .A(n480), .B(n479), .Z(n482) );
  OR U793 ( .A(n439), .B(n438), .Z(n443) );
  NANDN U794 ( .A(n441), .B(n440), .Z(n442) );
  NAND U795 ( .A(n443), .B(n442), .Z(n494) );
  ANDN U796 ( .B(y[197]), .A(n52), .Z(n445) );
  NANDN U797 ( .A(n50), .B(y[199]), .Z(n444) );
  XOR U798 ( .A(n445), .B(n444), .Z(n522) );
  ANDN U799 ( .B(x[74]), .A(n2602), .Z(n447) );
  NANDN U800 ( .A(n54), .B(y[195]), .Z(n446) );
  XOR U801 ( .A(n447), .B(n446), .Z(n544) );
  NANDN U802 ( .A(n49), .B(y[200]), .Z(n543) );
  XNOR U803 ( .A(n544), .B(n543), .Z(n521) );
  XNOR U804 ( .A(n522), .B(n521), .Z(n515) );
  IV U805 ( .A(y[204]), .Z(n2905) );
  ANDN U806 ( .B(x[64]), .A(n2905), .Z(n449) );
  NANDN U807 ( .A(n2902), .B(x[76]), .Z(n448) );
  XOR U808 ( .A(n449), .B(n448), .Z(n536) );
  NANDN U809 ( .A(n56), .B(y[193]), .Z(n510) );
  XOR U810 ( .A(o[12]), .B(n510), .Z(n535) );
  XOR U811 ( .A(n536), .B(n535), .Z(n513) );
  ANDN U812 ( .B(x[72]), .A(n2897), .Z(n451) );
  NANDN U813 ( .A(n2906), .B(x[66]), .Z(n450) );
  XOR U814 ( .A(n451), .B(n450), .Z(n506) );
  NANDN U815 ( .A(n48), .B(y[201]), .Z(n505) );
  XNOR U816 ( .A(n506), .B(n505), .Z(n514) );
  XOR U817 ( .A(n513), .B(n514), .Z(n516) );
  AND U818 ( .A(y[201]), .B(x[69]), .Z(n656) );
  NANDN U819 ( .A(n804), .B(n656), .Z(n455) );
  OR U820 ( .A(n453), .B(n452), .Z(n454) );
  NAND U821 ( .A(n455), .B(n454), .Z(n498) );
  ANDN U822 ( .B(x[70]), .A(n2906), .Z(n457) );
  NAND U823 ( .A(n457), .B(n456), .Z(n461) );
  OR U824 ( .A(n459), .B(n458), .Z(n460) );
  NAND U825 ( .A(n461), .B(n460), .Z(n497) );
  XOR U826 ( .A(n498), .B(n497), .Z(n500) );
  XNOR U827 ( .A(n499), .B(n500), .Z(n491) );
  AND U828 ( .A(y[203]), .B(x[75]), .Z(n1614) );
  NAND U829 ( .A(n794), .B(n1614), .Z(n465) );
  OR U830 ( .A(n463), .B(n462), .Z(n464) );
  NAND U831 ( .A(n465), .B(n464), .Z(n527) );
  NANDN U832 ( .A(n2602), .B(x[71]), .Z(n681) );
  NANDN U833 ( .A(n54), .B(y[196]), .Z(n1042) );
  OR U834 ( .A(n681), .B(n1042), .Z(n469) );
  OR U835 ( .A(n467), .B(n466), .Z(n468) );
  NAND U836 ( .A(n469), .B(n468), .Z(n525) );
  NANDN U837 ( .A(n470), .B(o[11]), .Z(n532) );
  ANDN U838 ( .B(y[203]), .A(n46), .Z(n472) );
  NANDN U839 ( .A(n2651), .B(x[70]), .Z(n471) );
  XOR U840 ( .A(n472), .B(n471), .Z(n531) );
  XOR U841 ( .A(n525), .B(n526), .Z(n528) );
  XOR U842 ( .A(n527), .B(n528), .Z(n492) );
  XNOR U843 ( .A(n491), .B(n492), .Z(n493) );
  XNOR U844 ( .A(n494), .B(n493), .Z(n481) );
  XNOR U845 ( .A(n482), .B(n481), .Z(n476) );
  XOR U846 ( .A(n475), .B(n476), .Z(N45) );
  NANDN U847 ( .A(n474), .B(n473), .Z(n478) );
  NANDN U848 ( .A(n476), .B(n475), .Z(n477) );
  NAND U849 ( .A(n478), .B(n477), .Z(n619) );
  OR U850 ( .A(n480), .B(n479), .Z(n484) );
  OR U851 ( .A(n482), .B(n481), .Z(n483) );
  AND U852 ( .A(n484), .B(n483), .Z(n620) );
  XNOR U853 ( .A(n619), .B(n620), .Z(n621) );
  OR U854 ( .A(n486), .B(n485), .Z(n490) );
  OR U855 ( .A(n488), .B(n487), .Z(n489) );
  AND U856 ( .A(n490), .B(n489), .Z(n625) );
  NANDN U857 ( .A(n492), .B(n491), .Z(n496) );
  NANDN U858 ( .A(n494), .B(n493), .Z(n495) );
  NAND U859 ( .A(n496), .B(n495), .Z(n626) );
  XOR U860 ( .A(n625), .B(n626), .Z(n627) );
  OR U861 ( .A(n498), .B(n497), .Z(n502) );
  NAND U862 ( .A(n500), .B(n499), .Z(n501) );
  AND U863 ( .A(n502), .B(n501), .Z(n557) );
  ANDN U864 ( .B(x[72]), .A(n2906), .Z(n504) );
  NAND U865 ( .A(n504), .B(n503), .Z(n508) );
  OR U866 ( .A(n506), .B(n505), .Z(n507) );
  NAND U867 ( .A(n508), .B(n507), .Z(n578) );
  ANDN U868 ( .B(y[199]), .A(n51), .Z(n509) );
  XOR U869 ( .A(n509), .B(n1042), .Z(n605) );
  NANDN U870 ( .A(n47), .B(y[203]), .Z(n604) );
  XNOR U871 ( .A(n605), .B(n604), .Z(n576) );
  NANDN U872 ( .A(n510), .B(o[12]), .Z(n588) );
  ANDN U873 ( .B(y[204]), .A(n46), .Z(n512) );
  NANDN U874 ( .A(n2651), .B(x[71]), .Z(n511) );
  XOR U875 ( .A(n512), .B(n511), .Z(n587) );
  XNOR U876 ( .A(n578), .B(n577), .Z(n554) );
  NANDN U877 ( .A(n514), .B(n513), .Z(n518) );
  OR U878 ( .A(n516), .B(n515), .Z(n517) );
  AND U879 ( .A(n518), .B(n517), .Z(n551) );
  ANDN U880 ( .B(x[71]), .A(n2878), .Z(n519) );
  NANDN U881 ( .A(n520), .B(n519), .Z(n524) );
  OR U882 ( .A(n522), .B(n521), .Z(n523) );
  AND U883 ( .A(n524), .B(n523), .Z(n552) );
  XOR U884 ( .A(n551), .B(n552), .Z(n553) );
  XNOR U885 ( .A(n554), .B(n553), .Z(n558) );
  XNOR U886 ( .A(n557), .B(n558), .Z(n559) );
  NANDN U887 ( .A(n526), .B(n525), .Z(n530) );
  NANDN U888 ( .A(n528), .B(n527), .Z(n529) );
  NAND U889 ( .A(n530), .B(n529), .Z(n566) );
  AND U890 ( .A(y[203]), .B(x[70]), .Z(n1008) );
  NAND U891 ( .A(n585), .B(n1008), .Z(n534) );
  OR U892 ( .A(n532), .B(n531), .Z(n533) );
  NAND U893 ( .A(n534), .B(n533), .Z(n571) );
  AND U894 ( .A(x[76]), .B(y[204]), .Z(n1827) );
  NAND U895 ( .A(n794), .B(n1827), .Z(n538) );
  OR U896 ( .A(n536), .B(n535), .Z(n537) );
  AND U897 ( .A(n538), .B(n537), .Z(n569) );
  ANDN U898 ( .B(y[194]), .A(n56), .Z(n540) );
  NANDN U899 ( .A(n55), .B(y[195]), .Z(n539) );
  XNOR U900 ( .A(n540), .B(n539), .Z(n591) );
  XNOR U901 ( .A(n1208), .B(n591), .Z(n570) );
  XOR U902 ( .A(n571), .B(n572), .Z(n563) );
  ANDN U903 ( .B(y[194]), .A(n54), .Z(n542) );
  ANDN U904 ( .B(y[195]), .A(n55), .Z(n541) );
  NAND U905 ( .A(n542), .B(n541), .Z(n546) );
  OR U906 ( .A(n544), .B(n543), .Z(n545) );
  NAND U907 ( .A(n546), .B(n545), .Z(n616) );
  IV U908 ( .A(y[205]), .Z(n1613) );
  ANDN U909 ( .B(x[64]), .A(n1613), .Z(n548) );
  NANDN U910 ( .A(n2902), .B(x[77]), .Z(n547) );
  XOR U911 ( .A(n548), .B(n547), .Z(n599) );
  NANDN U912 ( .A(n57), .B(y[193]), .Z(n610) );
  XOR U913 ( .A(o[13]), .B(n610), .Z(n598) );
  XNOR U914 ( .A(n599), .B(n598), .Z(n614) );
  ANDN U915 ( .B(x[69]), .A(n2512), .Z(n550) );
  NANDN U916 ( .A(n2906), .B(x[67]), .Z(n549) );
  XOR U917 ( .A(n550), .B(n549), .Z(n595) );
  NANDN U918 ( .A(n2837), .B(x[68]), .Z(n594) );
  XOR U919 ( .A(n595), .B(n594), .Z(n613) );
  XOR U920 ( .A(n616), .B(n615), .Z(n564) );
  XNOR U921 ( .A(n563), .B(n564), .Z(n565) );
  XOR U922 ( .A(n566), .B(n565), .Z(n560) );
  XOR U923 ( .A(n627), .B(n628), .Z(n622) );
  XOR U924 ( .A(n621), .B(n622), .Z(N46) );
  OR U925 ( .A(n552), .B(n551), .Z(n556) );
  NANDN U926 ( .A(n554), .B(n553), .Z(n555) );
  NAND U927 ( .A(n556), .B(n555), .Z(n640) );
  OR U928 ( .A(n558), .B(n557), .Z(n562) );
  OR U929 ( .A(n560), .B(n559), .Z(n561) );
  AND U930 ( .A(n562), .B(n561), .Z(n637) );
  NANDN U931 ( .A(n564), .B(n563), .Z(n568) );
  NANDN U932 ( .A(n566), .B(n565), .Z(n567) );
  AND U933 ( .A(n568), .B(n567), .Z(n718) );
  OR U934 ( .A(n570), .B(n569), .Z(n574) );
  NANDN U935 ( .A(n572), .B(n571), .Z(n573) );
  AND U936 ( .A(n574), .B(n573), .Z(n645) );
  NANDN U937 ( .A(n576), .B(n575), .Z(n580) );
  NAND U938 ( .A(n578), .B(n577), .Z(n579) );
  AND U939 ( .A(n580), .B(n579), .Z(n644) );
  ANDN U940 ( .B(y[203]), .A(n48), .Z(n582) );
  NANDN U941 ( .A(n2651), .B(x[72]), .Z(n581) );
  XNOR U942 ( .A(n582), .B(n581), .Z(n657) );
  XNOR U943 ( .A(n656), .B(n657), .Z(n672) );
  AND U944 ( .A(x[68]), .B(y[202]), .Z(n671) );
  AND U945 ( .A(y[196]), .B(x[74]), .Z(n1337) );
  ANDN U946 ( .B(y[204]), .A(n47), .Z(n584) );
  ANDN U947 ( .B(x[73]), .A(n1746), .Z(n583) );
  XNOR U948 ( .A(n584), .B(n583), .Z(n677) );
  XOR U949 ( .A(n1337), .B(n677), .Z(n670) );
  XOR U950 ( .A(n671), .B(n670), .Z(n673) );
  ANDN U951 ( .B(x[71]), .A(n2905), .Z(n586) );
  NAND U952 ( .A(n586), .B(n585), .Z(n590) );
  OR U953 ( .A(n588), .B(n587), .Z(n589) );
  AND U954 ( .A(n590), .B(n589), .Z(n649) );
  NANDN U955 ( .A(n55), .B(y[194]), .Z(n1213) );
  ANDN U956 ( .B(y[195]), .A(n56), .Z(n692) );
  IV U957 ( .A(n692), .Z(n763) );
  OR U958 ( .A(n1213), .B(n763), .Z(n593) );
  NAND U959 ( .A(n591), .B(n1208), .Z(n592) );
  AND U960 ( .A(n593), .B(n592), .Z(n650) );
  XOR U961 ( .A(n644), .B(n643), .Z(n646) );
  AND U962 ( .A(x[69]), .B(y[202]), .Z(n778) );
  NAND U963 ( .A(n1482), .B(n778), .Z(n597) );
  OR U964 ( .A(n595), .B(n594), .Z(n596) );
  NAND U965 ( .A(n597), .B(n596), .Z(n705) );
  NAND U966 ( .A(y[205]), .B(x[65]), .Z(n691) );
  XOR U967 ( .A(n692), .B(n691), .Z(n693) );
  XOR U968 ( .A(n694), .B(n693), .Z(n704) );
  ANDN U969 ( .B(x[77]), .A(n1613), .Z(n2191) );
  NAND U970 ( .A(n794), .B(n2191), .Z(n601) );
  OR U971 ( .A(n599), .B(n598), .Z(n600) );
  AND U972 ( .A(n601), .B(n600), .Z(n703) );
  XNOR U973 ( .A(n704), .B(n703), .Z(n706) );
  XOR U974 ( .A(n705), .B(n706), .Z(n711) );
  ANDN U975 ( .B(y[199]), .A(n54), .Z(n603) );
  NAND U976 ( .A(n603), .B(n602), .Z(n607) );
  OR U977 ( .A(n605), .B(n604), .Z(n606) );
  AND U978 ( .A(n607), .B(n606), .Z(n700) );
  ANDN U979 ( .B(y[194]), .A(n57), .Z(n609) );
  NANDN U980 ( .A(n2878), .B(x[71]), .Z(n608) );
  XOR U981 ( .A(n609), .B(n608), .Z(n683) );
  NANDN U982 ( .A(n58), .B(y[193]), .Z(n686) );
  XOR U983 ( .A(o[14]), .B(n686), .Z(n682) );
  XNOR U984 ( .A(n683), .B(n682), .Z(n698) );
  NANDN U985 ( .A(n610), .B(o[13]), .Z(n661) );
  IV U986 ( .A(y[206]), .Z(n2876) );
  ANDN U987 ( .B(x[64]), .A(n2876), .Z(n612) );
  NANDN U988 ( .A(n2902), .B(x[78]), .Z(n611) );
  XOR U989 ( .A(n612), .B(n611), .Z(n660) );
  XOR U990 ( .A(n700), .B(n699), .Z(n709) );
  NANDN U991 ( .A(n614), .B(n613), .Z(n618) );
  NAND U992 ( .A(n616), .B(n615), .Z(n617) );
  NAND U993 ( .A(n618), .B(n617), .Z(n710) );
  XOR U994 ( .A(n709), .B(n710), .Z(n712) );
  XOR U995 ( .A(n711), .B(n712), .Z(n716) );
  XOR U996 ( .A(n718), .B(n717), .Z(n638) );
  XNOR U997 ( .A(n637), .B(n638), .Z(n639) );
  XNOR U998 ( .A(n640), .B(n639), .Z(n634) );
  NANDN U999 ( .A(n620), .B(n619), .Z(n624) );
  NANDN U1000 ( .A(n622), .B(n621), .Z(n623) );
  NAND U1001 ( .A(n624), .B(n623), .Z(n631) );
  OR U1002 ( .A(n626), .B(n625), .Z(n630) );
  NANDN U1003 ( .A(n628), .B(n627), .Z(n629) );
  AND U1004 ( .A(n630), .B(n629), .Z(n632) );
  XNOR U1005 ( .A(n631), .B(n632), .Z(n633) );
  XOR U1006 ( .A(n634), .B(n633), .Z(N47) );
  NANDN U1007 ( .A(n632), .B(n631), .Z(n636) );
  NANDN U1008 ( .A(n634), .B(n633), .Z(n635) );
  NAND U1009 ( .A(n636), .B(n635), .Z(n721) );
  OR U1010 ( .A(n638), .B(n637), .Z(n642) );
  OR U1011 ( .A(n640), .B(n639), .Z(n641) );
  AND U1012 ( .A(n642), .B(n641), .Z(n722) );
  XNOR U1013 ( .A(n721), .B(n722), .Z(n723) );
  NANDN U1014 ( .A(n644), .B(n643), .Z(n648) );
  OR U1015 ( .A(n646), .B(n645), .Z(n647) );
  NAND U1016 ( .A(n648), .B(n647), .Z(n812) );
  OR U1017 ( .A(n650), .B(n649), .Z(n654) );
  NANDN U1018 ( .A(n652), .B(n651), .Z(n653) );
  AND U1019 ( .A(n654), .B(n653), .Z(n747) );
  NANDN U1020 ( .A(n53), .B(y[203]), .Z(n1089) );
  OR U1021 ( .A(n1089), .B(n655), .Z(n659) );
  NAND U1022 ( .A(n657), .B(n656), .Z(n658) );
  NAND U1023 ( .A(n659), .B(n658), .Z(n773) );
  ANDN U1024 ( .B(x[78]), .A(n2876), .Z(n2472) );
  NAND U1025 ( .A(n794), .B(n2472), .Z(n663) );
  OR U1026 ( .A(n661), .B(n660), .Z(n662) );
  NAND U1027 ( .A(n663), .B(n662), .Z(n772) );
  NANDN U1028 ( .A(n59), .B(y[193]), .Z(n799) );
  XOR U1029 ( .A(o[15]), .B(n799), .Z(n791) );
  ANDN U1030 ( .B(y[206]), .A(n46), .Z(n665) );
  NANDN U1031 ( .A(n53), .B(y[199]), .Z(n664) );
  XOR U1032 ( .A(n665), .B(n664), .Z(n790) );
  XOR U1033 ( .A(n791), .B(n790), .Z(n757) );
  ANDN U1034 ( .B(x[66]), .A(n1613), .Z(n667) );
  NANDN U1035 ( .A(n2651), .B(x[73]), .Z(n666) );
  XOR U1036 ( .A(n667), .B(n666), .Z(n806) );
  NANDN U1037 ( .A(n48), .B(y[204]), .Z(n805) );
  XOR U1038 ( .A(n806), .B(n805), .Z(n758) );
  AND U1039 ( .A(x[71]), .B(y[200]), .Z(n1160) );
  ANDN U1040 ( .B(x[74]), .A(n1746), .Z(n669) );
  NANDN U1041 ( .A(n49), .B(y[203]), .Z(n668) );
  XOR U1042 ( .A(n669), .B(n668), .Z(n784) );
  XNOR U1043 ( .A(n1160), .B(n784), .Z(n779) );
  ANDN U1044 ( .B(y[201]), .A(n51), .Z(n851) );
  XNOR U1045 ( .A(n778), .B(n851), .Z(n780) );
  XOR U1046 ( .A(n774), .B(n775), .Z(n745) );
  NANDN U1047 ( .A(n671), .B(n670), .Z(n675) );
  NANDN U1048 ( .A(n673), .B(n672), .Z(n674) );
  NAND U1049 ( .A(n675), .B(n674), .Z(n746) );
  XNOR U1050 ( .A(n745), .B(n746), .Z(n748) );
  XNOR U1051 ( .A(n747), .B(n748), .Z(n810) );
  AND U1052 ( .A(y[204]), .B(x[73]), .Z(n1433) );
  NAND U1053 ( .A(n676), .B(n1433), .Z(n679) );
  NANDN U1054 ( .A(n677), .B(n1337), .Z(n678) );
  AND U1055 ( .A(n679), .B(n678), .Z(n739) );
  ANDN U1056 ( .B(x[76]), .A(n2878), .Z(n680) );
  NANDN U1057 ( .A(n681), .B(n680), .Z(n685) );
  OR U1058 ( .A(n683), .B(n682), .Z(n684) );
  NAND U1059 ( .A(n685), .B(n684), .Z(n754) );
  NANDN U1060 ( .A(n686), .B(o[14]), .Z(n796) );
  IV U1061 ( .A(y[207]), .Z(n2852) );
  ANDN U1062 ( .B(x[64]), .A(n2852), .Z(n688) );
  NANDN U1063 ( .A(n2902), .B(x[79]), .Z(n687) );
  XOR U1064 ( .A(n688), .B(n687), .Z(n795) );
  XOR U1065 ( .A(n796), .B(n795), .Z(n751) );
  ANDN U1066 ( .B(y[195]), .A(n57), .Z(n690) );
  NANDN U1067 ( .A(n2897), .B(x[75]), .Z(n689) );
  XOR U1068 ( .A(n690), .B(n689), .Z(n765) );
  NANDN U1069 ( .A(n2602), .B(x[77]), .Z(n764) );
  XOR U1070 ( .A(n765), .B(n764), .Z(n752) );
  XNOR U1071 ( .A(n754), .B(n753), .Z(n740) );
  XNOR U1072 ( .A(n739), .B(n740), .Z(n741) );
  NANDN U1073 ( .A(n692), .B(n691), .Z(n696) );
  OR U1074 ( .A(n694), .B(n693), .Z(n695) );
  NAND U1075 ( .A(n696), .B(n695), .Z(n742) );
  NANDN U1076 ( .A(n698), .B(n697), .Z(n702) );
  NANDN U1077 ( .A(n700), .B(n699), .Z(n701) );
  AND U1078 ( .A(n702), .B(n701), .Z(n733) );
  XNOR U1079 ( .A(n734), .B(n733), .Z(n736) );
  OR U1080 ( .A(n704), .B(n703), .Z(n708) );
  NANDN U1081 ( .A(n706), .B(n705), .Z(n707) );
  AND U1082 ( .A(n708), .B(n707), .Z(n735) );
  XOR U1083 ( .A(n736), .B(n735), .Z(n809) );
  XNOR U1084 ( .A(n812), .B(n811), .Z(n728) );
  NANDN U1085 ( .A(n710), .B(n709), .Z(n714) );
  NANDN U1086 ( .A(n712), .B(n711), .Z(n713) );
  NAND U1087 ( .A(n714), .B(n713), .Z(n727) );
  NANDN U1088 ( .A(n716), .B(n715), .Z(n720) );
  NANDN U1089 ( .A(n718), .B(n717), .Z(n719) );
  NAND U1090 ( .A(n720), .B(n719), .Z(n730) );
  XNOR U1091 ( .A(n729), .B(n730), .Z(n724) );
  XOR U1092 ( .A(n723), .B(n724), .Z(N48) );
  NANDN U1093 ( .A(n722), .B(n721), .Z(n726) );
  NANDN U1094 ( .A(n724), .B(n723), .Z(n725) );
  NAND U1095 ( .A(n726), .B(n725), .Z(n815) );
  OR U1096 ( .A(n728), .B(n727), .Z(n732) );
  NANDN U1097 ( .A(n730), .B(n729), .Z(n731) );
  NAND U1098 ( .A(n732), .B(n731), .Z(n816) );
  XNOR U1099 ( .A(n815), .B(n816), .Z(n817) );
  OR U1100 ( .A(n734), .B(n733), .Z(n738) );
  OR U1101 ( .A(n736), .B(n735), .Z(n737) );
  NAND U1102 ( .A(n738), .B(n737), .Z(n907) );
  OR U1103 ( .A(n740), .B(n739), .Z(n744) );
  OR U1104 ( .A(n742), .B(n741), .Z(n743) );
  NAND U1105 ( .A(n744), .B(n743), .Z(n905) );
  OR U1106 ( .A(n746), .B(n745), .Z(n750) );
  OR U1107 ( .A(n748), .B(n747), .Z(n749) );
  NAND U1108 ( .A(n750), .B(n749), .Z(n904) );
  XOR U1109 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U1110 ( .A(n907), .B(n906), .Z(n824) );
  OR U1111 ( .A(n752), .B(n751), .Z(n756) );
  NANDN U1112 ( .A(n754), .B(n753), .Z(n755) );
  NAND U1113 ( .A(n756), .B(n755), .Z(n901) );
  OR U1114 ( .A(n758), .B(n757), .Z(n762) );
  NANDN U1115 ( .A(n760), .B(n759), .Z(n761) );
  AND U1116 ( .A(n762), .B(n761), .Z(n898) );
  AND U1117 ( .A(x[76]), .B(y[196]), .Z(n1576) );
  NANDN U1118 ( .A(n763), .B(n1576), .Z(n767) );
  OR U1119 ( .A(n765), .B(n764), .Z(n766) );
  NAND U1120 ( .A(n767), .B(n766), .Z(n894) );
  ANDN U1121 ( .B(x[66]), .A(n2876), .Z(n769) );
  NANDN U1122 ( .A(n54), .B(y[199]), .Z(n768) );
  XOR U1123 ( .A(n769), .B(n768), .Z(n884) );
  NANDN U1124 ( .A(n1613), .B(x[67]), .Z(n883) );
  XOR U1125 ( .A(n884), .B(n883), .Z(n892) );
  ANDN U1126 ( .B(x[77]), .A(n43), .Z(n771) );
  NANDN U1127 ( .A(n50), .B(y[203]), .Z(n770) );
  XNOR U1128 ( .A(n771), .B(n770), .Z(n857) );
  XNOR U1129 ( .A(n1576), .B(n857), .Z(n893) );
  XOR U1130 ( .A(n892), .B(n893), .Z(n895) );
  XNOR U1131 ( .A(n894), .B(n895), .Z(n899) );
  XNOR U1132 ( .A(n901), .B(n900), .Z(n872) );
  OR U1133 ( .A(n773), .B(n772), .Z(n777) );
  NAND U1134 ( .A(n775), .B(n774), .Z(n776) );
  NAND U1135 ( .A(n777), .B(n776), .Z(n870) );
  OR U1136 ( .A(n778), .B(n851), .Z(n782) );
  OR U1137 ( .A(n780), .B(n779), .Z(n781) );
  AND U1138 ( .A(n782), .B(n781), .Z(n827) );
  AND U1139 ( .A(y[203]), .B(x[74]), .Z(n1478) );
  NAND U1140 ( .A(n783), .B(n1478), .Z(n786) );
  NANDN U1141 ( .A(n784), .B(n1160), .Z(n785) );
  NAND U1142 ( .A(n786), .B(n785), .Z(n866) );
  NANDN U1143 ( .A(n45), .B(y[208]), .Z(n840) );
  IV U1144 ( .A(x[80]), .Z(n8890) );
  NANDN U1145 ( .A(n8890), .B(y[192]), .Z(n839) );
  XOR U1146 ( .A(n840), .B(n839), .Z(n841) );
  NANDN U1147 ( .A(n60), .B(y[193]), .Z(n860) );
  XOR U1148 ( .A(o[16]), .B(n860), .Z(n842) );
  XOR U1149 ( .A(n841), .B(n842), .Z(n864) );
  ANDN U1150 ( .B(y[201]), .A(n52), .Z(n788) );
  NANDN U1151 ( .A(n2906), .B(x[70]), .Z(n787) );
  XOR U1152 ( .A(n788), .B(n787), .Z(n853) );
  NANDN U1153 ( .A(n55), .B(y[198]), .Z(n852) );
  XOR U1154 ( .A(n853), .B(n852), .Z(n863) );
  XNOR U1155 ( .A(n864), .B(n863), .Z(n865) );
  XNOR U1156 ( .A(n866), .B(n865), .Z(n878) );
  NANDN U1157 ( .A(n53), .B(y[206]), .Z(n1735) );
  ANDN U1158 ( .B(x[65]), .A(n2878), .Z(n789) );
  NANDN U1159 ( .A(n1735), .B(n789), .Z(n793) );
  OR U1160 ( .A(n791), .B(n790), .Z(n792) );
  AND U1161 ( .A(n793), .B(n792), .Z(n875) );
  NANDN U1162 ( .A(n60), .B(y[207]), .Z(n2830) );
  NANDN U1163 ( .A(n2830), .B(n794), .Z(n798) );
  OR U1164 ( .A(n796), .B(n795), .Z(n797) );
  AND U1165 ( .A(n798), .B(n797), .Z(n876) );
  XOR U1166 ( .A(n875), .B(n876), .Z(n877) );
  XNOR U1167 ( .A(n878), .B(n877), .Z(n828) );
  NANDN U1168 ( .A(n799), .B(o[15]), .Z(n848) );
  ANDN U1169 ( .B(y[207]), .A(n46), .Z(n801) );
  NANDN U1170 ( .A(n53), .B(y[200]), .Z(n800) );
  XOR U1171 ( .A(n801), .B(n800), .Z(n847) );
  XOR U1172 ( .A(n848), .B(n847), .Z(n836) );
  ANDN U1173 ( .B(y[197]), .A(n56), .Z(n803) );
  NANDN U1174 ( .A(n2602), .B(x[78]), .Z(n802) );
  XOR U1175 ( .A(n803), .B(n802), .Z(n889) );
  NANDN U1176 ( .A(n49), .B(y[204]), .Z(n888) );
  XOR U1177 ( .A(n889), .B(n888), .Z(n833) );
  AND U1178 ( .A(y[205]), .B(x[73]), .Z(n1572) );
  NANDN U1179 ( .A(n804), .B(n1572), .Z(n808) );
  OR U1180 ( .A(n806), .B(n805), .Z(n807) );
  NAND U1181 ( .A(n808), .B(n807), .Z(n834) );
  XOR U1182 ( .A(n836), .B(n835), .Z(n829) );
  XNOR U1183 ( .A(n870), .B(n869), .Z(n871) );
  XOR U1184 ( .A(n872), .B(n871), .Z(n821) );
  NANDN U1185 ( .A(n810), .B(n809), .Z(n814) );
  NAND U1186 ( .A(n812), .B(n811), .Z(n813) );
  AND U1187 ( .A(n814), .B(n813), .Z(n822) );
  XNOR U1188 ( .A(n824), .B(n823), .Z(n818) );
  XOR U1189 ( .A(n817), .B(n818), .Z(N49) );
  NANDN U1190 ( .A(n816), .B(n815), .Z(n820) );
  NANDN U1191 ( .A(n818), .B(n817), .Z(n819) );
  NAND U1192 ( .A(n820), .B(n819), .Z(n910) );
  OR U1193 ( .A(n822), .B(n821), .Z(n826) );
  NANDN U1194 ( .A(n824), .B(n823), .Z(n825) );
  NAND U1195 ( .A(n826), .B(n825), .Z(n911) );
  XNOR U1196 ( .A(n910), .B(n911), .Z(n912) );
  OR U1197 ( .A(n828), .B(n827), .Z(n832) );
  NANDN U1198 ( .A(n830), .B(n829), .Z(n831) );
  NAND U1199 ( .A(n832), .B(n831), .Z(n1016) );
  OR U1200 ( .A(n834), .B(n833), .Z(n838) );
  OR U1201 ( .A(n836), .B(n835), .Z(n837) );
  AND U1202 ( .A(n838), .B(n837), .Z(n1013) );
  OR U1203 ( .A(n840), .B(n839), .Z(n844) );
  NANDN U1204 ( .A(n842), .B(n841), .Z(n843) );
  AND U1205 ( .A(n844), .B(n843), .Z(n949) );
  ANDN U1206 ( .B(y[207]), .A(n47), .Z(n846) );
  NANDN U1207 ( .A(n55), .B(y[199]), .Z(n845) );
  XOR U1208 ( .A(n846), .B(n845), .Z(n1002) );
  NANDN U1209 ( .A(n2876), .B(x[67]), .Z(n1001) );
  XNOR U1210 ( .A(n1002), .B(n1001), .Z(n947) );
  NANDN U1211 ( .A(n8890), .B(y[193]), .Z(n974) );
  XOR U1212 ( .A(o[17]), .B(n974), .Z(n959) );
  IV U1213 ( .A(x[81]), .Z(n8626) );
  ANDN U1214 ( .B(y[192]), .A(n8626), .Z(n958) );
  XOR U1215 ( .A(n959), .B(n958), .Z(n961) );
  IV U1216 ( .A(y[209]), .Z(n2851) );
  ANDN U1217 ( .B(x[64]), .A(n2851), .Z(n960) );
  XNOR U1218 ( .A(n961), .B(n960), .Z(n946) );
  XOR U1219 ( .A(n949), .B(n948), .Z(n943) );
  NANDN U1220 ( .A(n53), .B(y[207]), .Z(n1571) );
  AND U1221 ( .A(x[65]), .B(y[200]), .Z(n1067) );
  NANDN U1222 ( .A(n1571), .B(n1067), .Z(n850) );
  OR U1223 ( .A(n848), .B(n847), .Z(n849) );
  NAND U1224 ( .A(n850), .B(n849), .Z(n941) );
  NOR U1225 ( .A(n52), .B(n2906), .Z(n881) );
  IV U1226 ( .A(n881), .Z(n1088) );
  NANDN U1227 ( .A(n1088), .B(n851), .Z(n855) );
  OR U1228 ( .A(n853), .B(n852), .Z(n854) );
  NAND U1229 ( .A(n855), .B(n854), .Z(n940) );
  XOR U1230 ( .A(n943), .B(n942), .Z(n928) );
  AND U1231 ( .A(y[203]), .B(x[77]), .Z(n1752) );
  IV U1232 ( .A(n1752), .Z(n1819) );
  ANDN U1233 ( .B(y[195]), .A(n50), .Z(n856) );
  NANDN U1234 ( .A(n1819), .B(n856), .Z(n859) );
  NAND U1235 ( .A(n857), .B(n1576), .Z(n858) );
  NAND U1236 ( .A(n859), .B(n858), .Z(n954) );
  NANDN U1237 ( .A(n57), .B(y[197]), .Z(n981) );
  AND U1238 ( .A(x[78]), .B(y[195]), .Z(n980) );
  NANDN U1239 ( .A(n60), .B(y[194]), .Z(n979) );
  XOR U1240 ( .A(n980), .B(n979), .Z(n982) );
  XNOR U1241 ( .A(n981), .B(n982), .Z(n953) );
  NANDN U1242 ( .A(n860), .B(o[16]), .Z(n997) );
  ANDN U1243 ( .B(y[208]), .A(n46), .Z(n862) );
  NANDN U1244 ( .A(n54), .B(y[200]), .Z(n861) );
  XOR U1245 ( .A(n862), .B(n861), .Z(n996) );
  XOR U1246 ( .A(n953), .B(n952), .Z(n955) );
  XOR U1247 ( .A(n954), .B(n955), .Z(n929) );
  XNOR U1248 ( .A(n928), .B(n929), .Z(n931) );
  NANDN U1249 ( .A(n864), .B(n863), .Z(n868) );
  NAND U1250 ( .A(n866), .B(n865), .Z(n867) );
  AND U1251 ( .A(n868), .B(n867), .Z(n930) );
  XOR U1252 ( .A(n931), .B(n930), .Z(n1014) );
  XNOR U1253 ( .A(n1016), .B(n1015), .Z(n917) );
  NAND U1254 ( .A(n870), .B(n869), .Z(n874) );
  OR U1255 ( .A(n872), .B(n871), .Z(n873) );
  NAND U1256 ( .A(n874), .B(n873), .Z(n925) );
  OR U1257 ( .A(n876), .B(n875), .Z(n880) );
  NANDN U1258 ( .A(n878), .B(n877), .Z(n879) );
  NAND U1259 ( .A(n880), .B(n879), .Z(n937) );
  AND U1260 ( .A(y[205]), .B(x[68]), .Z(n971) );
  AND U1261 ( .A(x[75]), .B(y[198]), .Z(n969) );
  AND U1262 ( .A(y[196]), .B(x[77]), .Z(n968) );
  XNOR U1263 ( .A(n969), .B(n968), .Z(n970) );
  XNOR U1264 ( .A(n971), .B(n970), .Z(n991) );
  NANDN U1265 ( .A(n2905), .B(x[69]), .Z(n1010) );
  NANDN U1266 ( .A(n53), .B(y[201]), .Z(n1007) );
  XNOR U1267 ( .A(n1008), .B(n1007), .Z(n1009) );
  XOR U1268 ( .A(n1010), .B(n1009), .Z(n992) );
  XNOR U1269 ( .A(n991), .B(n992), .Z(n993) );
  XOR U1270 ( .A(n881), .B(n993), .Z(n988) );
  ANDN U1271 ( .B(y[206]), .A(n54), .Z(n882) );
  NAND U1272 ( .A(n882), .B(n1000), .Z(n886) );
  OR U1273 ( .A(n884), .B(n883), .Z(n885) );
  NAND U1274 ( .A(n886), .B(n885), .Z(n986) );
  NANDN U1275 ( .A(n2602), .B(x[75]), .Z(n1050) );
  ANDN U1276 ( .B(x[78]), .A(n1746), .Z(n887) );
  NANDN U1277 ( .A(n1050), .B(n887), .Z(n891) );
  OR U1278 ( .A(n889), .B(n888), .Z(n890) );
  NAND U1279 ( .A(n891), .B(n890), .Z(n985) );
  XNOR U1280 ( .A(n988), .B(n987), .Z(n935) );
  NANDN U1281 ( .A(n893), .B(n892), .Z(n897) );
  NANDN U1282 ( .A(n895), .B(n894), .Z(n896) );
  AND U1283 ( .A(n897), .B(n896), .Z(n934) );
  XOR U1284 ( .A(n935), .B(n934), .Z(n936) );
  XNOR U1285 ( .A(n937), .B(n936), .Z(n923) );
  OR U1286 ( .A(n899), .B(n898), .Z(n903) );
  NAND U1287 ( .A(n901), .B(n900), .Z(n902) );
  NAND U1288 ( .A(n903), .B(n902), .Z(n922) );
  XNOR U1289 ( .A(n925), .B(n924), .Z(n916) );
  XNOR U1290 ( .A(n917), .B(n916), .Z(n919) );
  OR U1291 ( .A(n905), .B(n904), .Z(n909) );
  NANDN U1292 ( .A(n907), .B(n906), .Z(n908) );
  AND U1293 ( .A(n909), .B(n908), .Z(n918) );
  XOR U1294 ( .A(n919), .B(n918), .Z(n913) );
  XNOR U1295 ( .A(n912), .B(n913), .Z(N50) );
  NANDN U1296 ( .A(n911), .B(n910), .Z(n915) );
  NAND U1297 ( .A(n913), .B(n912), .Z(n914) );
  NAND U1298 ( .A(n915), .B(n914), .Z(n1019) );
  OR U1299 ( .A(n917), .B(n916), .Z(n921) );
  OR U1300 ( .A(n919), .B(n918), .Z(n920) );
  AND U1301 ( .A(n921), .B(n920), .Z(n1020) );
  XNOR U1302 ( .A(n1019), .B(n1020), .Z(n1021) );
  OR U1303 ( .A(n923), .B(n922), .Z(n927) );
  NANDN U1304 ( .A(n925), .B(n924), .Z(n926) );
  NAND U1305 ( .A(n927), .B(n926), .Z(n1028) );
  OR U1306 ( .A(n929), .B(n928), .Z(n933) );
  OR U1307 ( .A(n931), .B(n930), .Z(n932) );
  NAND U1308 ( .A(n933), .B(n932), .Z(n1128) );
  OR U1309 ( .A(n935), .B(n934), .Z(n939) );
  NAND U1310 ( .A(n937), .B(n936), .Z(n938) );
  NAND U1311 ( .A(n939), .B(n938), .Z(n1127) );
  XOR U1312 ( .A(n1128), .B(n1127), .Z(n1129) );
  OR U1313 ( .A(n941), .B(n940), .Z(n945) );
  NAND U1314 ( .A(n943), .B(n942), .Z(n944) );
  NAND U1315 ( .A(n945), .B(n944), .Z(n1106) );
  NANDN U1316 ( .A(n947), .B(n946), .Z(n951) );
  NANDN U1317 ( .A(n949), .B(n948), .Z(n950) );
  AND U1318 ( .A(n951), .B(n950), .Z(n1103) );
  NANDN U1319 ( .A(n953), .B(n952), .Z(n957) );
  NANDN U1320 ( .A(n955), .B(n954), .Z(n956) );
  AND U1321 ( .A(n957), .B(n956), .Z(n1104) );
  XNOR U1322 ( .A(n1106), .B(n1105), .Z(n1033) );
  NANDN U1323 ( .A(n959), .B(n958), .Z(n963) );
  NANDN U1324 ( .A(n961), .B(n960), .Z(n962) );
  NAND U1325 ( .A(n963), .B(n962), .Z(n1110) );
  ANDN U1326 ( .B(y[203]), .A(n52), .Z(n965) );
  NANDN U1327 ( .A(n2906), .B(x[72]), .Z(n964) );
  XOR U1328 ( .A(n965), .B(n964), .Z(n1091) );
  NANDN U1329 ( .A(n49), .B(y[206]), .Z(n1090) );
  XOR U1330 ( .A(n1091), .B(n1090), .Z(n1037) );
  AND U1331 ( .A(y[204]), .B(x[70]), .Z(n1551) );
  NANDN U1332 ( .A(n1613), .B(x[69]), .Z(n1192) );
  XOR U1333 ( .A(n1551), .B(n1192), .Z(n1038) );
  XNOR U1334 ( .A(n1110), .B(n1109), .Z(n1111) );
  NANDN U1335 ( .A(n47), .B(y[208]), .Z(n1052) );
  ANDN U1336 ( .B(y[194]), .A(n8890), .Z(n967) );
  NANDN U1337 ( .A(n2878), .B(x[75]), .Z(n966) );
  XOR U1338 ( .A(n967), .B(n966), .Z(n1051) );
  XOR U1339 ( .A(n1052), .B(n1051), .Z(n1112) );
  XOR U1340 ( .A(n1111), .B(n1112), .Z(n1123) );
  OR U1341 ( .A(n969), .B(n968), .Z(n973) );
  OR U1342 ( .A(n971), .B(n970), .Z(n972) );
  NAND U1343 ( .A(n973), .B(n972), .Z(n1058) );
  NANDN U1344 ( .A(n974), .B(o[17]), .Z(n1069) );
  ANDN U1345 ( .B(x[65]), .A(n2851), .Z(n976) );
  NANDN U1346 ( .A(n55), .B(y[200]), .Z(n975) );
  XOR U1347 ( .A(n976), .B(n975), .Z(n1068) );
  ANDN U1348 ( .B(y[196]), .A(n59), .Z(n978) );
  NANDN U1349 ( .A(n2837), .B(x[73]), .Z(n977) );
  XOR U1350 ( .A(n978), .B(n977), .Z(n1044) );
  NANDN U1351 ( .A(n60), .B(y[195]), .Z(n1043) );
  XOR U1352 ( .A(n1044), .B(n1043), .Z(n1055) );
  XOR U1353 ( .A(n1058), .B(n1057), .Z(n1122) );
  NANDN U1354 ( .A(n980), .B(n979), .Z(n984) );
  NANDN U1355 ( .A(n982), .B(n981), .Z(n983) );
  AND U1356 ( .A(n984), .B(n983), .Z(n1121) );
  XOR U1357 ( .A(n1122), .B(n1121), .Z(n1124) );
  XNOR U1358 ( .A(n1123), .B(n1124), .Z(n1031) );
  OR U1359 ( .A(n986), .B(n985), .Z(n990) );
  NANDN U1360 ( .A(n988), .B(n987), .Z(n989) );
  NAND U1361 ( .A(n990), .B(n989), .Z(n1100) );
  NANDN U1362 ( .A(n992), .B(n991), .Z(n995) );
  NANDN U1363 ( .A(n1088), .B(n993), .Z(n994) );
  NAND U1364 ( .A(n995), .B(n994), .Z(n1098) );
  AND U1365 ( .A(y[208]), .B(x[73]), .Z(n2039) );
  NAND U1366 ( .A(n2039), .B(n1067), .Z(n999) );
  OR U1367 ( .A(n997), .B(n996), .Z(n998) );
  NAND U1368 ( .A(n999), .B(n998), .Z(n1118) );
  ANDN U1369 ( .B(x[74]), .A(n2852), .Z(n2038) );
  NAND U1370 ( .A(n1000), .B(n2038), .Z(n1004) );
  OR U1371 ( .A(n1002), .B(n1001), .Z(n1003) );
  NAND U1372 ( .A(n1004), .B(n1003), .Z(n1063) );
  NANDN U1373 ( .A(n45), .B(y[210]), .Z(n1073) );
  NANDN U1374 ( .A(n61), .B(y[192]), .Z(n1072) );
  XOR U1375 ( .A(n1073), .B(n1072), .Z(n1074) );
  NANDN U1376 ( .A(n8626), .B(y[193]), .Z(n1094) );
  XOR U1377 ( .A(o[18]), .B(n1094), .Z(n1075) );
  XOR U1378 ( .A(n1074), .B(n1075), .Z(n1062) );
  AND U1379 ( .A(x[76]), .B(y[198]), .Z(n1154) );
  ANDN U1380 ( .B(y[207]), .A(n48), .Z(n1006) );
  NANDN U1381 ( .A(n58), .B(y[197]), .Z(n1005) );
  XOR U1382 ( .A(n1006), .B(n1005), .Z(n1081) );
  XOR U1383 ( .A(n1062), .B(n1061), .Z(n1064) );
  XOR U1384 ( .A(n1063), .B(n1064), .Z(n1115) );
  NANDN U1385 ( .A(n1008), .B(n1007), .Z(n1012) );
  NAND U1386 ( .A(n1010), .B(n1009), .Z(n1011) );
  AND U1387 ( .A(n1012), .B(n1011), .Z(n1116) );
  XOR U1388 ( .A(n1115), .B(n1116), .Z(n1117) );
  XNOR U1389 ( .A(n1118), .B(n1117), .Z(n1097) );
  XOR U1390 ( .A(n1098), .B(n1097), .Z(n1099) );
  XNOR U1391 ( .A(n1100), .B(n1099), .Z(n1032) );
  XNOR U1392 ( .A(n1031), .B(n1032), .Z(n1034) );
  XNOR U1393 ( .A(n1033), .B(n1034), .Z(n1130) );
  XNOR U1394 ( .A(n1129), .B(n1130), .Z(n1025) );
  OR U1395 ( .A(n1014), .B(n1013), .Z(n1018) );
  NAND U1396 ( .A(n1016), .B(n1015), .Z(n1017) );
  NAND U1397 ( .A(n1018), .B(n1017), .Z(n1026) );
  XOR U1398 ( .A(n1025), .B(n1026), .Z(n1027) );
  XOR U1399 ( .A(n1028), .B(n1027), .Z(n1022) );
  XOR U1400 ( .A(n1021), .B(n1022), .Z(N51) );
  NANDN U1401 ( .A(n1020), .B(n1019), .Z(n1024) );
  NANDN U1402 ( .A(n1022), .B(n1021), .Z(n1023) );
  NAND U1403 ( .A(n1024), .B(n1023), .Z(n1133) );
  OR U1404 ( .A(n1026), .B(n1025), .Z(n1030) );
  NAND U1405 ( .A(n1028), .B(n1027), .Z(n1029) );
  NAND U1406 ( .A(n1030), .B(n1029), .Z(n1134) );
  XNOR U1407 ( .A(n1133), .B(n1134), .Z(n1135) );
  OR U1408 ( .A(n1032), .B(n1031), .Z(n1036) );
  OR U1409 ( .A(n1034), .B(n1033), .Z(n1035) );
  AND U1410 ( .A(n1036), .B(n1035), .Z(n1139) );
  NANDN U1411 ( .A(n1551), .B(n1192), .Z(n1040) );
  OR U1412 ( .A(n1038), .B(n1037), .Z(n1039) );
  NAND U1413 ( .A(n1040), .B(n1039), .Z(n1232) );
  ANDN U1414 ( .B(y[197]), .A(n59), .Z(n1041) );
  XOR U1415 ( .A(n1041), .B(n1089), .Z(n1210) );
  NANDN U1416 ( .A(n46), .B(y[210]), .Z(n1209) );
  XOR U1417 ( .A(n1210), .B(n1209), .Z(n1176) );
  AND U1418 ( .A(x[78]), .B(y[201]), .Z(n1681) );
  NANDN U1419 ( .A(n1042), .B(n1681), .Z(n1046) );
  OR U1420 ( .A(n1044), .B(n1043), .Z(n1045) );
  NAND U1421 ( .A(n1046), .B(n1045), .Z(n1175) );
  NANDN U1422 ( .A(n47), .B(y[209]), .Z(n1157) );
  ANDN U1423 ( .B(y[199]), .A(n57), .Z(n1048) );
  ANDN U1424 ( .B(y[198]), .A(n58), .Z(n1047) );
  XNOR U1425 ( .A(n1048), .B(n1047), .Z(n1156) );
  XOR U1426 ( .A(n1157), .B(n1156), .Z(n1174) );
  XNOR U1427 ( .A(n1175), .B(n1174), .Z(n1177) );
  XNOR U1428 ( .A(n1176), .B(n1177), .Z(n1230) );
  ANDN U1429 ( .B(x[80]), .A(n2878), .Z(n1049) );
  NANDN U1430 ( .A(n1050), .B(n1049), .Z(n1054) );
  OR U1431 ( .A(n1052), .B(n1051), .Z(n1053) );
  NAND U1432 ( .A(n1054), .B(n1053), .Z(n1231) );
  XOR U1433 ( .A(n1232), .B(n1233), .Z(n1236) );
  NANDN U1434 ( .A(n1056), .B(n1055), .Z(n1060) );
  NANDN U1435 ( .A(n1058), .B(n1057), .Z(n1059) );
  NAND U1436 ( .A(n1060), .B(n1059), .Z(n1225) );
  NANDN U1437 ( .A(n1062), .B(n1061), .Z(n1066) );
  NANDN U1438 ( .A(n1064), .B(n1063), .Z(n1065) );
  NAND U1439 ( .A(n1066), .B(n1065), .Z(n1224) );
  ANDN U1440 ( .B(x[74]), .A(n2851), .Z(n2335) );
  NAND U1441 ( .A(n1067), .B(n2335), .Z(n1071) );
  OR U1442 ( .A(n1069), .B(n1068), .Z(n1070) );
  AND U1443 ( .A(n1071), .B(n1070), .Z(n1188) );
  OR U1444 ( .A(n1073), .B(n1072), .Z(n1077) );
  NANDN U1445 ( .A(n1075), .B(n1074), .Z(n1076) );
  NAND U1446 ( .A(n1077), .B(n1076), .Z(n1186) );
  ANDN U1447 ( .B(x[80]), .A(n43), .Z(n1079) );
  NANDN U1448 ( .A(n2906), .B(x[73]), .Z(n1078) );
  XOR U1449 ( .A(n1079), .B(n1078), .Z(n1147) );
  ANDN U1450 ( .B(y[196]), .A(n60), .Z(n1146) );
  XOR U1451 ( .A(n1147), .B(n1146), .Z(n1187) );
  XOR U1452 ( .A(n1186), .B(n1187), .Z(n1189) );
  ANDN U1453 ( .B(x[77]), .A(n2852), .Z(n2439) );
  NAND U1454 ( .A(n1080), .B(n2439), .Z(n1083) );
  NANDN U1455 ( .A(n1081), .B(n1154), .Z(n1082) );
  NAND U1456 ( .A(n1083), .B(n1082), .Z(n1181) );
  ANDN U1457 ( .B(y[204]), .A(n52), .Z(n1085) );
  NANDN U1458 ( .A(n2512), .B(x[75]), .Z(n1084) );
  XOR U1459 ( .A(n1085), .B(n1084), .Z(n1162) );
  NANDN U1460 ( .A(n48), .B(y[208]), .Z(n1161) );
  XOR U1461 ( .A(n1162), .B(n1161), .Z(n1180) );
  XNOR U1462 ( .A(n1181), .B(n1180), .Z(n1183) );
  ANDN U1463 ( .B(y[193]), .A(n61), .Z(n1167) );
  XNOR U1464 ( .A(o[19]), .B(n1167), .Z(n1215) );
  ANDN U1465 ( .B(y[201]), .A(n55), .Z(n1087) );
  NANDN U1466 ( .A(n8626), .B(y[194]), .Z(n1086) );
  XNOR U1467 ( .A(n1087), .B(n1086), .Z(n1214) );
  XOR U1468 ( .A(n1215), .B(n1214), .Z(n1182) );
  XOR U1469 ( .A(n1183), .B(n1182), .Z(n1218) );
  OR U1470 ( .A(n1089), .B(n1088), .Z(n1093) );
  OR U1471 ( .A(n1091), .B(n1090), .Z(n1092) );
  NAND U1472 ( .A(n1093), .B(n1092), .Z(n1170) );
  NANDN U1473 ( .A(n1094), .B(o[18]), .Z(n1201) );
  NANDN U1474 ( .A(n45), .B(y[211]), .Z(n1199) );
  IV U1475 ( .A(x[83]), .Z(n8824) );
  NANDN U1476 ( .A(n8824), .B(y[192]), .Z(n1198) );
  XOR U1477 ( .A(n1199), .B(n1198), .Z(n1200) );
  XNOR U1478 ( .A(n1201), .B(n1200), .Z(n1168) );
  AND U1479 ( .A(y[207]), .B(x[68]), .Z(n1324) );
  ANDN U1480 ( .B(x[70]), .A(n1613), .Z(n1096) );
  NANDN U1481 ( .A(n50), .B(y[206]), .Z(n1095) );
  XNOR U1482 ( .A(n1096), .B(n1095), .Z(n1193) );
  XNOR U1483 ( .A(n1324), .B(n1193), .Z(n1169) );
  XOR U1484 ( .A(n1168), .B(n1169), .Z(n1171) );
  XNOR U1485 ( .A(n1170), .B(n1171), .Z(n1219) );
  XOR U1486 ( .A(n1226), .B(n1227), .Z(n1237) );
  XNOR U1487 ( .A(n1236), .B(n1237), .Z(n1238) );
  OR U1488 ( .A(n1098), .B(n1097), .Z(n1102) );
  NAND U1489 ( .A(n1100), .B(n1099), .Z(n1101) );
  NAND U1490 ( .A(n1102), .B(n1101), .Z(n1239) );
  XOR U1491 ( .A(n1238), .B(n1239), .Z(n1244) );
  OR U1492 ( .A(n1104), .B(n1103), .Z(n1108) );
  NANDN U1493 ( .A(n1106), .B(n1105), .Z(n1107) );
  NAND U1494 ( .A(n1108), .B(n1107), .Z(n1243) );
  NANDN U1495 ( .A(n1110), .B(n1109), .Z(n1114) );
  NANDN U1496 ( .A(n1112), .B(n1111), .Z(n1113) );
  AND U1497 ( .A(n1114), .B(n1113), .Z(n1251) );
  NANDN U1498 ( .A(n1116), .B(n1115), .Z(n1120) );
  OR U1499 ( .A(n1118), .B(n1117), .Z(n1119) );
  AND U1500 ( .A(n1120), .B(n1119), .Z(n1248) );
  NANDN U1501 ( .A(n1122), .B(n1121), .Z(n1126) );
  NANDN U1502 ( .A(n1124), .B(n1123), .Z(n1125) );
  NAND U1503 ( .A(n1126), .B(n1125), .Z(n1249) );
  XNOR U1504 ( .A(n1248), .B(n1249), .Z(n1250) );
  XOR U1505 ( .A(n1251), .B(n1250), .Z(n1242) );
  XOR U1506 ( .A(n1243), .B(n1242), .Z(n1245) );
  XOR U1507 ( .A(n1244), .B(n1245), .Z(n1140) );
  XNOR U1508 ( .A(n1139), .B(n1140), .Z(n1141) );
  OR U1509 ( .A(n1128), .B(n1127), .Z(n1132) );
  NANDN U1510 ( .A(n1130), .B(n1129), .Z(n1131) );
  AND U1511 ( .A(n1132), .B(n1131), .Z(n1142) );
  XOR U1512 ( .A(n1135), .B(n1136), .Z(N52) );
  NANDN U1513 ( .A(n1134), .B(n1133), .Z(n1138) );
  NANDN U1514 ( .A(n1136), .B(n1135), .Z(n1137) );
  NAND U1515 ( .A(n1138), .B(n1137), .Z(n1254) );
  OR U1516 ( .A(n1140), .B(n1139), .Z(n1144) );
  OR U1517 ( .A(n1142), .B(n1141), .Z(n1143) );
  AND U1518 ( .A(n1144), .B(n1143), .Z(n1255) );
  XNOR U1519 ( .A(n1254), .B(n1255), .Z(n1256) );
  ANDN U1520 ( .B(y[195]), .A(n54), .Z(n1145) );
  ANDN U1521 ( .B(y[202]), .A(n8890), .Z(n2091) );
  NAND U1522 ( .A(n1145), .B(n2091), .Z(n1149) );
  NANDN U1523 ( .A(n1147), .B(n1146), .Z(n1148) );
  AND U1524 ( .A(n1149), .B(n1148), .Z(n1313) );
  ANDN U1525 ( .B(y[197]), .A(n60), .Z(n1151) );
  NANDN U1526 ( .A(n54), .B(y[203]), .Z(n1150) );
  XOR U1527 ( .A(n1151), .B(n1150), .Z(n1290) );
  NANDN U1528 ( .A(n59), .B(y[198]), .Z(n1289) );
  XOR U1529 ( .A(n1290), .B(n1289), .Z(n1348) );
  IV U1530 ( .A(y[210]), .Z(n2702) );
  NANDN U1531 ( .A(n2702), .B(x[66]), .Z(n1339) );
  ANDN U1532 ( .B(x[80]), .A(n2897), .Z(n1153) );
  NANDN U1533 ( .A(n2906), .B(x[74]), .Z(n1152) );
  XOR U1534 ( .A(n1153), .B(n1152), .Z(n1338) );
  XNOR U1535 ( .A(n1339), .B(n1338), .Z(n1349) );
  XOR U1536 ( .A(n1348), .B(n1349), .Z(n1351) );
  ANDN U1537 ( .B(x[77]), .A(n2878), .Z(n1155) );
  NAND U1538 ( .A(n1155), .B(n1154), .Z(n1159) );
  OR U1539 ( .A(n1157), .B(n1156), .Z(n1158) );
  AND U1540 ( .A(n1159), .B(n1158), .Z(n1350) );
  XNOR U1541 ( .A(n1351), .B(n1350), .Z(n1312) );
  AND U1542 ( .A(x[75]), .B(y[204]), .Z(n1742) );
  NAND U1543 ( .A(n1742), .B(n1160), .Z(n1164) );
  OR U1544 ( .A(n1162), .B(n1161), .Z(n1163) );
  AND U1545 ( .A(n1164), .B(n1163), .Z(n1356) );
  ANDN U1546 ( .B(y[211]), .A(n46), .Z(n1166) );
  NANDN U1547 ( .A(n2837), .B(x[75]), .Z(n1165) );
  XOR U1548 ( .A(n1166), .B(n1165), .Z(n1285) );
  ANDN U1549 ( .B(y[193]), .A(n8824), .Z(n1293) );
  XOR U1550 ( .A(o[20]), .B(n1293), .Z(n1284) );
  XOR U1551 ( .A(n1285), .B(n1284), .Z(n1355) );
  NAND U1552 ( .A(o[19]), .B(n1167), .Z(n1321) );
  NANDN U1553 ( .A(n2902), .B(x[84]), .Z(n1319) );
  IV U1554 ( .A(y[212]), .Z(n2449) );
  ANDN U1555 ( .B(x[64]), .A(n2449), .Z(n1318) );
  XOR U1556 ( .A(n1319), .B(n1318), .Z(n1320) );
  XOR U1557 ( .A(n1355), .B(n1354), .Z(n1357) );
  XOR U1558 ( .A(n1356), .B(n1357), .Z(n1314) );
  XNOR U1559 ( .A(n1315), .B(n1314), .Z(n1269) );
  NANDN U1560 ( .A(n1169), .B(n1168), .Z(n1173) );
  NANDN U1561 ( .A(n1171), .B(n1170), .Z(n1172) );
  NAND U1562 ( .A(n1173), .B(n1172), .Z(n1267) );
  NAND U1563 ( .A(n1175), .B(n1174), .Z(n1179) );
  NANDN U1564 ( .A(n1177), .B(n1176), .Z(n1178) );
  NAND U1565 ( .A(n1179), .B(n1178), .Z(n1266) );
  XOR U1566 ( .A(n1269), .B(n1268), .Z(n1308) );
  NAND U1567 ( .A(n1181), .B(n1180), .Z(n1185) );
  OR U1568 ( .A(n1183), .B(n1182), .Z(n1184) );
  NAND U1569 ( .A(n1185), .B(n1184), .Z(n1307) );
  NANDN U1570 ( .A(n1187), .B(n1186), .Z(n1191) );
  OR U1571 ( .A(n1189), .B(n1188), .Z(n1190) );
  NAND U1572 ( .A(n1191), .B(n1190), .Z(n1275) );
  AND U1573 ( .A(y[206]), .B(x[70]), .Z(n1294) );
  NANDN U1574 ( .A(n1192), .B(n1294), .Z(n1195) );
  NAND U1575 ( .A(n1193), .B(n1324), .Z(n1194) );
  AND U1576 ( .A(n1195), .B(n1194), .Z(n1303) );
  NANDN U1577 ( .A(n8626), .B(y[195]), .Z(n1280) );
  ANDN U1578 ( .B(y[200]), .A(n57), .Z(n1197) );
  ANDN U1579 ( .B(x[82]), .A(n2602), .Z(n1196) );
  XNOR U1580 ( .A(n1197), .B(n1196), .Z(n1279) );
  XOR U1581 ( .A(n1280), .B(n1279), .Z(n1300) );
  OR U1582 ( .A(n1199), .B(n1198), .Z(n1203) );
  NANDN U1583 ( .A(n1201), .B(n1200), .Z(n1202) );
  AND U1584 ( .A(n1203), .B(n1202), .Z(n1301) );
  XNOR U1585 ( .A(n1300), .B(n1301), .Z(n1302) );
  XOR U1586 ( .A(n1303), .B(n1302), .Z(n1272) );
  NANDN U1587 ( .A(n52), .B(y[205]), .Z(n1326) );
  ANDN U1588 ( .B(x[69]), .A(n2852), .Z(n1205) );
  NANDN U1589 ( .A(n49), .B(y[208]), .Z(n1204) );
  XOR U1590 ( .A(n1205), .B(n1204), .Z(n1325) );
  XNOR U1591 ( .A(n1326), .B(n1325), .Z(n1295) );
  XOR U1592 ( .A(n1294), .B(n1295), .Z(n1297) );
  NANDN U1593 ( .A(n53), .B(y[204]), .Z(n1334) );
  ANDN U1594 ( .B(x[67]), .A(n2851), .Z(n1207) );
  NANDN U1595 ( .A(n2878), .B(x[77]), .Z(n1206) );
  XOR U1596 ( .A(n1207), .B(n1206), .Z(n1333) );
  XNOR U1597 ( .A(n1334), .B(n1333), .Z(n1296) );
  XNOR U1598 ( .A(n1297), .B(n1296), .Z(n1344) );
  AND U1599 ( .A(y[203]), .B(x[78]), .Z(n1984) );
  NAND U1600 ( .A(n1984), .B(n1208), .Z(n1212) );
  OR U1601 ( .A(n1210), .B(n1209), .Z(n1211) );
  NAND U1602 ( .A(n1212), .B(n1211), .Z(n1343) );
  ANDN U1603 ( .B(x[81]), .A(n2837), .Z(n2104) );
  NANDN U1604 ( .A(n1213), .B(n2104), .Z(n1217) );
  NANDN U1605 ( .A(n1215), .B(n1214), .Z(n1216) );
  NAND U1606 ( .A(n1217), .B(n1216), .Z(n1342) );
  XOR U1607 ( .A(n1343), .B(n1342), .Z(n1345) );
  XNOR U1608 ( .A(n1344), .B(n1345), .Z(n1273) );
  XNOR U1609 ( .A(n1272), .B(n1273), .Z(n1274) );
  XNOR U1610 ( .A(n1275), .B(n1274), .Z(n1306) );
  XOR U1611 ( .A(n1307), .B(n1306), .Z(n1309) );
  XOR U1612 ( .A(n1308), .B(n1309), .Z(n1366) );
  OR U1613 ( .A(n1219), .B(n1218), .Z(n1223) );
  NANDN U1614 ( .A(n1221), .B(n1220), .Z(n1222) );
  NAND U1615 ( .A(n1223), .B(n1222), .Z(n1361) );
  OR U1616 ( .A(n1225), .B(n1224), .Z(n1229) );
  NAND U1617 ( .A(n1227), .B(n1226), .Z(n1228) );
  NAND U1618 ( .A(n1229), .B(n1228), .Z(n1360) );
  XNOR U1619 ( .A(n1361), .B(n1360), .Z(n1362) );
  OR U1620 ( .A(n1231), .B(n1230), .Z(n1235) );
  NANDN U1621 ( .A(n1233), .B(n1232), .Z(n1234) );
  NAND U1622 ( .A(n1235), .B(n1234), .Z(n1363) );
  XNOR U1623 ( .A(n1366), .B(n1367), .Z(n1369) );
  NANDN U1624 ( .A(n1237), .B(n1236), .Z(n1241) );
  NANDN U1625 ( .A(n1239), .B(n1238), .Z(n1240) );
  AND U1626 ( .A(n1241), .B(n1240), .Z(n1368) );
  XOR U1627 ( .A(n1369), .B(n1368), .Z(n1260) );
  NANDN U1628 ( .A(n1243), .B(n1242), .Z(n1247) );
  NANDN U1629 ( .A(n1245), .B(n1244), .Z(n1246) );
  AND U1630 ( .A(n1247), .B(n1246), .Z(n1261) );
  XNOR U1631 ( .A(n1260), .B(n1261), .Z(n1263) );
  OR U1632 ( .A(n1249), .B(n1248), .Z(n1253) );
  OR U1633 ( .A(n1251), .B(n1250), .Z(n1252) );
  NAND U1634 ( .A(n1253), .B(n1252), .Z(n1262) );
  XOR U1635 ( .A(n1263), .B(n1262), .Z(n1257) );
  XOR U1636 ( .A(n1256), .B(n1257), .Z(N53) );
  NANDN U1637 ( .A(n1255), .B(n1254), .Z(n1259) );
  NANDN U1638 ( .A(n1257), .B(n1256), .Z(n1258) );
  NAND U1639 ( .A(n1259), .B(n1258), .Z(n1372) );
  NAND U1640 ( .A(n1261), .B(n1260), .Z(n1265) );
  OR U1641 ( .A(n1263), .B(n1262), .Z(n1264) );
  NAND U1642 ( .A(n1265), .B(n1264), .Z(n1373) );
  XNOR U1643 ( .A(n1372), .B(n1373), .Z(n1374) );
  OR U1644 ( .A(n1267), .B(n1266), .Z(n1271) );
  NANDN U1645 ( .A(n1269), .B(n1268), .Z(n1270) );
  NAND U1646 ( .A(n1271), .B(n1270), .Z(n1499) );
  NANDN U1647 ( .A(n1273), .B(n1272), .Z(n1277) );
  NANDN U1648 ( .A(n1275), .B(n1274), .Z(n1276) );
  AND U1649 ( .A(n1277), .B(n1276), .Z(n1496) );
  ANDN U1650 ( .B(x[76]), .A(n2602), .Z(n1278) );
  ANDN U1651 ( .B(x[82]), .A(n2512), .Z(n2103) );
  NAND U1652 ( .A(n1278), .B(n2103), .Z(n1282) );
  OR U1653 ( .A(n1280), .B(n1279), .Z(n1281) );
  AND U1654 ( .A(n1282), .B(n1281), .Z(n1411) );
  NANDN U1655 ( .A(n56), .B(y[211]), .Z(n2921) );
  NANDN U1656 ( .A(n2921), .B(n1283), .Z(n1287) );
  NANDN U1657 ( .A(n1285), .B(n1284), .Z(n1286) );
  AND U1658 ( .A(n1287), .B(n1286), .Z(n1408) );
  ANDN U1659 ( .B(y[208]), .A(n50), .Z(n1488) );
  NANDN U1660 ( .A(n8890), .B(y[197]), .Z(n1489) );
  XOR U1661 ( .A(n1488), .B(n1489), .Z(n1491) );
  NANDN U1662 ( .A(n60), .B(y[198]), .Z(n1490) );
  XOR U1663 ( .A(n1491), .B(n1490), .Z(n1452) );
  ANDN U1664 ( .B(y[197]), .A(n54), .Z(n1288) );
  AND U1665 ( .A(y[203]), .B(x[79]), .Z(n2096) );
  NAND U1666 ( .A(n1288), .B(n2096), .Z(n1292) );
  OR U1667 ( .A(n1290), .B(n1289), .Z(n1291) );
  NAND U1668 ( .A(n1292), .B(n1291), .Z(n1453) );
  XNOR U1669 ( .A(n1452), .B(n1453), .Z(n1455) );
  AND U1670 ( .A(y[213]), .B(x[64]), .Z(n1472) );
  AND U1671 ( .A(n1293), .B(o[20]), .Z(n1470) );
  AND U1672 ( .A(x[85]), .B(y[192]), .Z(n1471) );
  XNOR U1673 ( .A(n1470), .B(n1471), .Z(n1473) );
  XNOR U1674 ( .A(n1472), .B(n1473), .Z(n1454) );
  XOR U1675 ( .A(n1455), .B(n1454), .Z(n1409) );
  XNOR U1676 ( .A(n1408), .B(n1409), .Z(n1410) );
  NANDN U1677 ( .A(n1295), .B(n1294), .Z(n1299) );
  OR U1678 ( .A(n1297), .B(n1296), .Z(n1298) );
  AND U1679 ( .A(n1299), .B(n1298), .Z(n1402) );
  XNOR U1680 ( .A(n1403), .B(n1402), .Z(n1405) );
  NANDN U1681 ( .A(n1301), .B(n1300), .Z(n1305) );
  NANDN U1682 ( .A(n1303), .B(n1302), .Z(n1304) );
  AND U1683 ( .A(n1305), .B(n1304), .Z(n1404) );
  XOR U1684 ( .A(n1405), .B(n1404), .Z(n1497) );
  XNOR U1685 ( .A(n1499), .B(n1498), .Z(n1387) );
  NANDN U1686 ( .A(n1307), .B(n1306), .Z(n1311) );
  OR U1687 ( .A(n1309), .B(n1308), .Z(n1310) );
  AND U1688 ( .A(n1311), .B(n1310), .Z(n1384) );
  OR U1689 ( .A(n1313), .B(n1312), .Z(n1317) );
  NANDN U1690 ( .A(n1315), .B(n1314), .Z(n1316) );
  NAND U1691 ( .A(n1317), .B(n1316), .Z(n1393) );
  NANDN U1692 ( .A(n1319), .B(n1318), .Z(n1323) );
  OR U1693 ( .A(n1321), .B(n1320), .Z(n1322) );
  AND U1694 ( .A(n1323), .B(n1322), .Z(n1414) );
  NAND U1695 ( .A(n1324), .B(n1488), .Z(n1328) );
  OR U1696 ( .A(n1326), .B(n1325), .Z(n1327) );
  AND U1697 ( .A(n1328), .B(n1327), .Z(n1415) );
  XOR U1698 ( .A(n1414), .B(n1415), .Z(n1417) );
  AND U1699 ( .A(y[207]), .B(x[70]), .Z(n1465) );
  AND U1700 ( .A(y[206]), .B(x[71]), .Z(n1570) );
  AND U1701 ( .A(x[78]), .B(y[199]), .Z(n1464) );
  XNOR U1702 ( .A(n1570), .B(n1464), .Z(n1466) );
  XNOR U1703 ( .A(n1465), .B(n1466), .Z(n1435) );
  NANDN U1704 ( .A(n1613), .B(x[72]), .Z(n1432) );
  XOR U1705 ( .A(n1433), .B(n1432), .Z(n1434) );
  XNOR U1706 ( .A(n1435), .B(n1434), .Z(n1460) );
  NANDN U1707 ( .A(n49), .B(y[209]), .Z(n1484) );
  ANDN U1708 ( .B(x[77]), .A(n2512), .Z(n1330) );
  ANDN U1709 ( .B(y[210]), .A(n48), .Z(n1329) );
  XNOR U1710 ( .A(n1330), .B(n1329), .Z(n1483) );
  XNOR U1711 ( .A(n1484), .B(n1483), .Z(n1458) );
  NANDN U1712 ( .A(n57), .B(y[201]), .Z(n1440) );
  AND U1713 ( .A(x[66]), .B(y[211]), .Z(n1439) );
  NANDN U1714 ( .A(n2897), .B(x[81]), .Z(n1438) );
  XOR U1715 ( .A(n1439), .B(n1438), .Z(n1441) );
  XNOR U1716 ( .A(n1440), .B(n1441), .Z(n1459) );
  XNOR U1717 ( .A(n1417), .B(n1416), .Z(n1428) );
  NANDN U1718 ( .A(n2906), .B(x[75]), .Z(n1449) );
  IV U1719 ( .A(x[84]), .Z(n8885) );
  NANDN U1720 ( .A(n8885), .B(y[193]), .Z(n1487) );
  XOR U1721 ( .A(o[21]), .B(n1487), .Z(n1447) );
  NANDN U1722 ( .A(n2602), .B(x[83]), .Z(n1446) );
  XNOR U1723 ( .A(n1447), .B(n1446), .Z(n1448) );
  XNOR U1724 ( .A(n1449), .B(n1448), .Z(n1421) );
  AND U1725 ( .A(x[65]), .B(y[212]), .Z(n1476) );
  AND U1726 ( .A(y[195]), .B(x[82]), .Z(n1477) );
  XNOR U1727 ( .A(n1476), .B(n1477), .Z(n1479) );
  XNOR U1728 ( .A(n1478), .B(n1479), .Z(n1420) );
  XOR U1729 ( .A(n1421), .B(n1420), .Z(n1423) );
  ANDN U1730 ( .B(y[209]), .A(n58), .Z(n1332) );
  NAND U1731 ( .A(n1332), .B(n1331), .Z(n1336) );
  OR U1732 ( .A(n1334), .B(n1333), .Z(n1335) );
  AND U1733 ( .A(n1336), .B(n1335), .Z(n1422) );
  XOR U1734 ( .A(n1423), .B(n1422), .Z(n1427) );
  NAND U1735 ( .A(n1337), .B(n2091), .Z(n1341) );
  OR U1736 ( .A(n1339), .B(n1338), .Z(n1340) );
  NAND U1737 ( .A(n1341), .B(n1340), .Z(n1426) );
  XNOR U1738 ( .A(n1427), .B(n1426), .Z(n1429) );
  XNOR U1739 ( .A(n1428), .B(n1429), .Z(n1391) );
  OR U1740 ( .A(n1343), .B(n1342), .Z(n1347) );
  NAND U1741 ( .A(n1345), .B(n1344), .Z(n1346) );
  AND U1742 ( .A(n1347), .B(n1346), .Z(n1396) );
  NANDN U1743 ( .A(n1349), .B(n1348), .Z(n1353) );
  OR U1744 ( .A(n1351), .B(n1350), .Z(n1352) );
  NAND U1745 ( .A(n1353), .B(n1352), .Z(n1397) );
  XOR U1746 ( .A(n1396), .B(n1397), .Z(n1398) );
  NANDN U1747 ( .A(n1355), .B(n1354), .Z(n1359) );
  OR U1748 ( .A(n1357), .B(n1356), .Z(n1358) );
  NAND U1749 ( .A(n1359), .B(n1358), .Z(n1399) );
  XNOR U1750 ( .A(n1398), .B(n1399), .Z(n1390) );
  XOR U1751 ( .A(n1391), .B(n1390), .Z(n1392) );
  XOR U1752 ( .A(n1393), .B(n1392), .Z(n1385) );
  XOR U1753 ( .A(n1387), .B(n1386), .Z(n1381) );
  OR U1754 ( .A(n1361), .B(n1360), .Z(n1365) );
  OR U1755 ( .A(n1363), .B(n1362), .Z(n1364) );
  NAND U1756 ( .A(n1365), .B(n1364), .Z(n1379) );
  OR U1757 ( .A(n1367), .B(n1366), .Z(n1371) );
  OR U1758 ( .A(n1369), .B(n1368), .Z(n1370) );
  NAND U1759 ( .A(n1371), .B(n1370), .Z(n1378) );
  XNOR U1760 ( .A(n1379), .B(n1378), .Z(n1380) );
  XNOR U1761 ( .A(n1381), .B(n1380), .Z(n1375) );
  XOR U1762 ( .A(n1374), .B(n1375), .Z(N54) );
  NANDN U1763 ( .A(n1373), .B(n1372), .Z(n1377) );
  NANDN U1764 ( .A(n1375), .B(n1374), .Z(n1376) );
  NAND U1765 ( .A(n1377), .B(n1376), .Z(n1502) );
  OR U1766 ( .A(n1379), .B(n1378), .Z(n1383) );
  OR U1767 ( .A(n1381), .B(n1380), .Z(n1382) );
  AND U1768 ( .A(n1383), .B(n1382), .Z(n1503) );
  XNOR U1769 ( .A(n1502), .B(n1503), .Z(n1504) );
  OR U1770 ( .A(n1385), .B(n1384), .Z(n1389) );
  NANDN U1771 ( .A(n1387), .B(n1386), .Z(n1388) );
  NAND U1772 ( .A(n1389), .B(n1388), .Z(n1511) );
  OR U1773 ( .A(n1391), .B(n1390), .Z(n1395) );
  NAND U1774 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U1775 ( .A(n1395), .B(n1394), .Z(n1633) );
  OR U1776 ( .A(n1397), .B(n1396), .Z(n1401) );
  NANDN U1777 ( .A(n1399), .B(n1398), .Z(n1400) );
  AND U1778 ( .A(n1401), .B(n1400), .Z(n1632) );
  XOR U1779 ( .A(n1633), .B(n1632), .Z(n1634) );
  OR U1780 ( .A(n1403), .B(n1402), .Z(n1407) );
  OR U1781 ( .A(n1405), .B(n1404), .Z(n1406) );
  NAND U1782 ( .A(n1407), .B(n1406), .Z(n1515) );
  OR U1783 ( .A(n1409), .B(n1408), .Z(n1413) );
  OR U1784 ( .A(n1411), .B(n1410), .Z(n1412) );
  NAND U1785 ( .A(n1413), .B(n1412), .Z(n1629) );
  OR U1786 ( .A(n1415), .B(n1414), .Z(n1419) );
  NAND U1787 ( .A(n1417), .B(n1416), .Z(n1418) );
  NAND U1788 ( .A(n1419), .B(n1418), .Z(n1627) );
  NANDN U1789 ( .A(n1421), .B(n1420), .Z(n1425) );
  OR U1790 ( .A(n1423), .B(n1422), .Z(n1424) );
  NAND U1791 ( .A(n1425), .B(n1424), .Z(n1626) );
  XNOR U1792 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U1793 ( .A(n1515), .B(n1514), .Z(n1517) );
  OR U1794 ( .A(n1427), .B(n1426), .Z(n1431) );
  NANDN U1795 ( .A(n1429), .B(n1428), .Z(n1430) );
  NAND U1796 ( .A(n1431), .B(n1430), .Z(n1523) );
  NANDN U1797 ( .A(n1433), .B(n1432), .Z(n1437) );
  OR U1798 ( .A(n1435), .B(n1434), .Z(n1436) );
  AND U1799 ( .A(n1437), .B(n1436), .Z(n1540) );
  NANDN U1800 ( .A(n1439), .B(n1438), .Z(n1443) );
  NANDN U1801 ( .A(n1441), .B(n1440), .Z(n1442) );
  NAND U1802 ( .A(n1443), .B(n1442), .Z(n1608) );
  ANDN U1803 ( .B(x[82]), .A(n2897), .Z(n1445) );
  NANDN U1804 ( .A(n2906), .B(x[76]), .Z(n1444) );
  XOR U1805 ( .A(n1445), .B(n1444), .Z(n1578) );
  NANDN U1806 ( .A(n2702), .B(x[68]), .Z(n1577) );
  XNOR U1807 ( .A(n1578), .B(n1577), .Z(n1605) );
  NANDN U1808 ( .A(n50), .B(y[209]), .Z(n1545) );
  NANDN U1809 ( .A(n1746), .B(x[81]), .Z(n1544) );
  XOR U1810 ( .A(n1545), .B(n1544), .Z(n1546) );
  NANDN U1811 ( .A(n8890), .B(y[198]), .Z(n1547) );
  XOR U1812 ( .A(n1546), .B(n1547), .Z(n1606) );
  XOR U1813 ( .A(n1608), .B(n1607), .Z(n1538) );
  OR U1814 ( .A(n1447), .B(n1446), .Z(n1451) );
  OR U1815 ( .A(n1449), .B(n1448), .Z(n1450) );
  NAND U1816 ( .A(n1451), .B(n1450), .Z(n1539) );
  XNOR U1817 ( .A(n1538), .B(n1539), .Z(n1541) );
  XOR U1818 ( .A(n1540), .B(n1541), .Z(n1521) );
  OR U1819 ( .A(n1453), .B(n1452), .Z(n1457) );
  OR U1820 ( .A(n1455), .B(n1454), .Z(n1456) );
  AND U1821 ( .A(n1457), .B(n1456), .Z(n1526) );
  OR U1822 ( .A(n1459), .B(n1458), .Z(n1463) );
  NANDN U1823 ( .A(n1461), .B(n1460), .Z(n1462) );
  NAND U1824 ( .A(n1463), .B(n1462), .Z(n1527) );
  XOR U1825 ( .A(n1526), .B(n1527), .Z(n1528) );
  OR U1826 ( .A(n1464), .B(n1570), .Z(n1468) );
  OR U1827 ( .A(n1466), .B(n1465), .Z(n1467) );
  NAND U1828 ( .A(n1468), .B(n1467), .Z(n1596) );
  ANDN U1829 ( .B(y[207]), .A(n52), .Z(n1469) );
  XNOR U1830 ( .A(n1469), .B(n1735), .Z(n1573) );
  XNOR U1831 ( .A(n1572), .B(n1573), .Z(n1594) );
  NANDN U1832 ( .A(n45), .B(y[214]), .Z(n1582) );
  IV U1833 ( .A(x[86]), .Z(n8864) );
  NANDN U1834 ( .A(n8864), .B(y[192]), .Z(n1581) );
  XOR U1835 ( .A(n1582), .B(n1581), .Z(n1583) );
  IV U1836 ( .A(x[85]), .Z(n8827) );
  NANDN U1837 ( .A(n8827), .B(y[193]), .Z(n1550) );
  XOR U1838 ( .A(o[22]), .B(n1550), .Z(n1584) );
  XOR U1839 ( .A(n1583), .B(n1584), .Z(n1593) );
  XOR U1840 ( .A(n1594), .B(n1593), .Z(n1595) );
  XNOR U1841 ( .A(n1596), .B(n1595), .Z(n1602) );
  OR U1842 ( .A(n1471), .B(n1470), .Z(n1475) );
  OR U1843 ( .A(n1473), .B(n1472), .Z(n1474) );
  AND U1844 ( .A(n1475), .B(n1474), .Z(n1599) );
  OR U1845 ( .A(n1477), .B(n1476), .Z(n1481) );
  OR U1846 ( .A(n1479), .B(n1478), .Z(n1480) );
  AND U1847 ( .A(n1481), .B(n1480), .Z(n1600) );
  XOR U1848 ( .A(n1599), .B(n1600), .Z(n1601) );
  XOR U1849 ( .A(n1602), .B(n1601), .Z(n1535) );
  AND U1850 ( .A(x[77]), .B(y[210]), .Z(n2923) );
  NAND U1851 ( .A(n1482), .B(n2923), .Z(n1486) );
  OR U1852 ( .A(n1484), .B(n1483), .Z(n1485) );
  AND U1853 ( .A(n1486), .B(n1485), .Z(n1587) );
  NANDN U1854 ( .A(n2512), .B(x[78]), .Z(n1621) );
  NANDN U1855 ( .A(n48), .B(y[211]), .Z(n1620) );
  XOR U1856 ( .A(n1621), .B(n1620), .Z(n1622) );
  NANDN U1857 ( .A(n43), .B(x[83]), .Z(n1623) );
  XOR U1858 ( .A(n1622), .B(n1623), .Z(n1588) );
  XNOR U1859 ( .A(n1587), .B(n1588), .Z(n1590) );
  NANDN U1860 ( .A(n1487), .B(o[21]), .Z(n1617) );
  NANDN U1861 ( .A(n46), .B(y[213]), .Z(n1615) );
  XOR U1862 ( .A(n1614), .B(n1615), .Z(n1616) );
  XNOR U1863 ( .A(n1617), .B(n1616), .Z(n1589) );
  XOR U1864 ( .A(n1590), .B(n1589), .Z(n1532) );
  NANDN U1865 ( .A(n2449), .B(x[66]), .Z(n1557) );
  NANDN U1866 ( .A(n2602), .B(x[84]), .Z(n1556) );
  XOR U1867 ( .A(n1557), .B(n1556), .Z(n1558) );
  NANDN U1868 ( .A(n58), .B(y[201]), .Z(n1559) );
  XOR U1869 ( .A(n1558), .B(n1559), .Z(n1565) );
  NANDN U1870 ( .A(n1489), .B(n1488), .Z(n1493) );
  OR U1871 ( .A(n1491), .B(n1490), .Z(n1492) );
  NAND U1872 ( .A(n1493), .B(n1492), .Z(n1563) );
  ANDN U1873 ( .B(y[208]), .A(n51), .Z(n1495) );
  NANDN U1874 ( .A(n55), .B(y[204]), .Z(n1494) );
  XOR U1875 ( .A(n1495), .B(n1494), .Z(n1553) );
  NANDN U1876 ( .A(n60), .B(y[199]), .Z(n1552) );
  XOR U1877 ( .A(n1553), .B(n1552), .Z(n1562) );
  XNOR U1878 ( .A(n1563), .B(n1562), .Z(n1564) );
  XOR U1879 ( .A(n1565), .B(n1564), .Z(n1533) );
  XNOR U1880 ( .A(n1532), .B(n1533), .Z(n1534) );
  XNOR U1881 ( .A(n1535), .B(n1534), .Z(n1529) );
  XOR U1882 ( .A(n1528), .B(n1529), .Z(n1520) );
  XNOR U1883 ( .A(n1521), .B(n1520), .Z(n1522) );
  XNOR U1884 ( .A(n1523), .B(n1522), .Z(n1516) );
  XNOR U1885 ( .A(n1517), .B(n1516), .Z(n1635) );
  XNOR U1886 ( .A(n1634), .B(n1635), .Z(n1508) );
  OR U1887 ( .A(n1497), .B(n1496), .Z(n1501) );
  NAND U1888 ( .A(n1499), .B(n1498), .Z(n1500) );
  NAND U1889 ( .A(n1501), .B(n1500), .Z(n1509) );
  XOR U1890 ( .A(n1508), .B(n1509), .Z(n1510) );
  XNOR U1891 ( .A(n1511), .B(n1510), .Z(n1505) );
  XOR U1892 ( .A(n1504), .B(n1505), .Z(N55) );
  NANDN U1893 ( .A(n1503), .B(n1502), .Z(n1507) );
  NANDN U1894 ( .A(n1505), .B(n1504), .Z(n1506) );
  NAND U1895 ( .A(n1507), .B(n1506), .Z(n1638) );
  OR U1896 ( .A(n1509), .B(n1508), .Z(n1513) );
  NANDN U1897 ( .A(n1511), .B(n1510), .Z(n1512) );
  NAND U1898 ( .A(n1513), .B(n1512), .Z(n1639) );
  XNOR U1899 ( .A(n1638), .B(n1639), .Z(n1640) );
  NANDN U1900 ( .A(n1515), .B(n1514), .Z(n1519) );
  OR U1901 ( .A(n1517), .B(n1516), .Z(n1518) );
  AND U1902 ( .A(n1519), .B(n1518), .Z(n1644) );
  NANDN U1903 ( .A(n1521), .B(n1520), .Z(n1525) );
  NANDN U1904 ( .A(n1523), .B(n1522), .Z(n1524) );
  NAND U1905 ( .A(n1525), .B(n1524), .Z(n1651) );
  OR U1906 ( .A(n1527), .B(n1526), .Z(n1531) );
  NANDN U1907 ( .A(n1529), .B(n1528), .Z(n1530) );
  AND U1908 ( .A(n1531), .B(n1530), .Z(n1773) );
  OR U1909 ( .A(n1533), .B(n1532), .Z(n1537) );
  OR U1910 ( .A(n1535), .B(n1534), .Z(n1536) );
  AND U1911 ( .A(n1537), .B(n1536), .Z(n1772) );
  OR U1912 ( .A(n1539), .B(n1538), .Z(n1543) );
  OR U1913 ( .A(n1541), .B(n1540), .Z(n1542) );
  AND U1914 ( .A(n1543), .B(n1542), .Z(n1771) );
  XNOR U1915 ( .A(n1772), .B(n1771), .Z(n1774) );
  XNOR U1916 ( .A(n1773), .B(n1774), .Z(n1650) );
  XOR U1917 ( .A(n1651), .B(n1650), .Z(n1652) );
  NANDN U1918 ( .A(n2906), .B(x[77]), .Z(n1676) );
  NANDN U1919 ( .A(n47), .B(y[213]), .Z(n1675) );
  XOR U1920 ( .A(n1676), .B(n1675), .Z(n1677) );
  NANDN U1921 ( .A(n2602), .B(x[85]), .Z(n1678) );
  XNOR U1922 ( .A(n1677), .B(n1678), .Z(n1713) );
  OR U1923 ( .A(n1545), .B(n1544), .Z(n1549) );
  NANDN U1924 ( .A(n1547), .B(n1546), .Z(n1548) );
  NAND U1925 ( .A(n1549), .B(n1548), .Z(n1711) );
  NANDN U1926 ( .A(n1550), .B(o[22]), .Z(n1732) );
  NANDN U1927 ( .A(n57), .B(y[203]), .Z(n1730) );
  NANDN U1928 ( .A(n46), .B(y[214]), .Z(n1729) );
  XOR U1929 ( .A(n1730), .B(n1729), .Z(n1731) );
  XOR U1930 ( .A(n1732), .B(n1731), .Z(n1712) );
  XOR U1931 ( .A(n1711), .B(n1712), .Z(n1714) );
  XOR U1932 ( .A(n1713), .B(n1714), .Z(n1755) );
  NANDN U1933 ( .A(n48), .B(y[212]), .Z(n1682) );
  XOR U1934 ( .A(n1681), .B(n1682), .Z(n1684) );
  IV U1935 ( .A(y[211]), .Z(n2937) );
  NANDN U1936 ( .A(n2937), .B(x[68]), .Z(n1683) );
  XOR U1937 ( .A(n1684), .B(n1683), .Z(n1695) );
  ANDN U1938 ( .B(y[208]), .A(n55), .Z(n2144) );
  NAND U1939 ( .A(n1551), .B(n2144), .Z(n1555) );
  OR U1940 ( .A(n1553), .B(n1552), .Z(n1554) );
  NAND U1941 ( .A(n1555), .B(n1554), .Z(n1693) );
  AND U1942 ( .A(y[198]), .B(x[81]), .Z(n1832) );
  NANDN U1943 ( .A(n50), .B(y[210]), .Z(n1669) );
  NANDN U1944 ( .A(n1746), .B(x[82]), .Z(n1668) );
  XOR U1945 ( .A(n1669), .B(n1668), .Z(n1670) );
  XNOR U1946 ( .A(n1832), .B(n1670), .Z(n1694) );
  XOR U1947 ( .A(n1693), .B(n1694), .Z(n1696) );
  XNOR U1948 ( .A(n1695), .B(n1696), .Z(n1753) );
  OR U1949 ( .A(n1557), .B(n1556), .Z(n1561) );
  NANDN U1950 ( .A(n1559), .B(n1558), .Z(n1560) );
  NAND U1951 ( .A(n1561), .B(n1560), .Z(n1754) );
  XOR U1952 ( .A(n1755), .B(n1756), .Z(n1717) );
  NAND U1953 ( .A(n1563), .B(n1562), .Z(n1567) );
  OR U1954 ( .A(n1565), .B(n1564), .Z(n1566) );
  AND U1955 ( .A(n1567), .B(n1566), .Z(n1718) );
  XOR U1956 ( .A(n1717), .B(n1718), .Z(n1719) );
  NANDN U1957 ( .A(n45), .B(y[215]), .Z(n1724) );
  IV U1958 ( .A(x[87]), .Z(n8656) );
  NANDN U1959 ( .A(n8656), .B(y[192]), .Z(n1723) );
  XOR U1960 ( .A(n1724), .B(n1723), .Z(n1725) );
  NANDN U1961 ( .A(n8864), .B(y[193]), .Z(n1751) );
  XOR U1962 ( .A(o[23]), .B(n1751), .Z(n1726) );
  XOR U1963 ( .A(n1725), .B(n1726), .Z(n1701) );
  AND U1964 ( .A(y[196]), .B(x[83]), .Z(n1979) );
  ANDN U1965 ( .B(y[199]), .A(n8890), .Z(n1569) );
  NANDN U1966 ( .A(n8885), .B(y[195]), .Z(n1568) );
  XOR U1967 ( .A(n1569), .B(n1568), .Z(n1748) );
  NANDN U1968 ( .A(n1571), .B(n1570), .Z(n1575) );
  NAND U1969 ( .A(n1573), .B(n1572), .Z(n1574) );
  NAND U1970 ( .A(n1575), .B(n1574), .Z(n1699) );
  XNOR U1971 ( .A(n1700), .B(n1699), .Z(n1702) );
  XNOR U1972 ( .A(n1701), .B(n1702), .Z(n1708) );
  ANDN U1973 ( .B(y[202]), .A(n61), .Z(n2456) );
  IV U1974 ( .A(n2456), .Z(n2346) );
  NANDN U1975 ( .A(n2346), .B(n1576), .Z(n1580) );
  OR U1976 ( .A(n1578), .B(n1577), .Z(n1579) );
  AND U1977 ( .A(n1580), .B(n1579), .Z(n1705) );
  OR U1978 ( .A(n1582), .B(n1581), .Z(n1586) );
  NANDN U1979 ( .A(n1584), .B(n1583), .Z(n1585) );
  AND U1980 ( .A(n1586), .B(n1585), .Z(n1706) );
  XOR U1981 ( .A(n1708), .B(n1707), .Z(n1720) );
  XOR U1982 ( .A(n1719), .B(n1720), .Z(n1759) );
  OR U1983 ( .A(n1588), .B(n1587), .Z(n1592) );
  OR U1984 ( .A(n1590), .B(n1589), .Z(n1591) );
  AND U1985 ( .A(n1592), .B(n1591), .Z(n1656) );
  OR U1986 ( .A(n1594), .B(n1593), .Z(n1598) );
  NANDN U1987 ( .A(n1596), .B(n1595), .Z(n1597) );
  AND U1988 ( .A(n1598), .B(n1597), .Z(n1657) );
  XNOR U1989 ( .A(n1656), .B(n1657), .Z(n1658) );
  OR U1990 ( .A(n1600), .B(n1599), .Z(n1604) );
  NANDN U1991 ( .A(n1602), .B(n1601), .Z(n1603) );
  NAND U1992 ( .A(n1604), .B(n1603), .Z(n1659) );
  OR U1993 ( .A(n1606), .B(n1605), .Z(n1610) );
  OR U1994 ( .A(n1608), .B(n1607), .Z(n1609) );
  AND U1995 ( .A(n1610), .B(n1609), .Z(n1765) );
  ANDN U1996 ( .B(x[72]), .A(n2852), .Z(n1612) );
  NANDN U1997 ( .A(n54), .B(y[206]), .Z(n1611) );
  XOR U1998 ( .A(n1612), .B(n1611), .Z(n1737) );
  NANDN U1999 ( .A(n52), .B(y[208]), .Z(n1736) );
  XOR U2000 ( .A(n1737), .B(n1736), .Z(n1687) );
  NANDN U2001 ( .A(n1613), .B(x[74]), .Z(n1688) );
  XNOR U2002 ( .A(n1687), .B(n1688), .Z(n1689) );
  NANDN U2003 ( .A(n51), .B(y[209]), .Z(n1741) );
  NANDN U2004 ( .A(n60), .B(y[200]), .Z(n1740) );
  XOR U2005 ( .A(n1741), .B(n1740), .Z(n1743) );
  XNOR U2006 ( .A(n1742), .B(n1743), .Z(n1690) );
  XOR U2007 ( .A(n1689), .B(n1690), .Z(n1665) );
  NANDN U2008 ( .A(n1615), .B(n1614), .Z(n1619) );
  OR U2009 ( .A(n1617), .B(n1616), .Z(n1618) );
  NAND U2010 ( .A(n1619), .B(n1618), .Z(n1663) );
  OR U2011 ( .A(n1621), .B(n1620), .Z(n1625) );
  NANDN U2012 ( .A(n1623), .B(n1622), .Z(n1624) );
  NAND U2013 ( .A(n1625), .B(n1624), .Z(n1662) );
  XOR U2014 ( .A(n1665), .B(n1664), .Z(n1766) );
  XOR U2015 ( .A(n1765), .B(n1766), .Z(n1767) );
  XNOR U2016 ( .A(n1768), .B(n1767), .Z(n1760) );
  XNOR U2017 ( .A(n1759), .B(n1760), .Z(n1762) );
  OR U2018 ( .A(n1627), .B(n1626), .Z(n1631) );
  OR U2019 ( .A(n1629), .B(n1628), .Z(n1630) );
  AND U2020 ( .A(n1631), .B(n1630), .Z(n1761) );
  XNOR U2021 ( .A(n1762), .B(n1761), .Z(n1653) );
  XOR U2022 ( .A(n1652), .B(n1653), .Z(n1645) );
  XNOR U2023 ( .A(n1644), .B(n1645), .Z(n1646) );
  OR U2024 ( .A(n1633), .B(n1632), .Z(n1637) );
  NANDN U2025 ( .A(n1635), .B(n1634), .Z(n1636) );
  AND U2026 ( .A(n1637), .B(n1636), .Z(n1647) );
  XOR U2027 ( .A(n1640), .B(n1641), .Z(N56) );
  NANDN U2028 ( .A(n1639), .B(n1638), .Z(n1643) );
  NANDN U2029 ( .A(n1641), .B(n1640), .Z(n1642) );
  NAND U2030 ( .A(n1643), .B(n1642), .Z(n1777) );
  OR U2031 ( .A(n1645), .B(n1644), .Z(n1649) );
  OR U2032 ( .A(n1647), .B(n1646), .Z(n1648) );
  AND U2033 ( .A(n1649), .B(n1648), .Z(n1778) );
  XNOR U2034 ( .A(n1777), .B(n1778), .Z(n1779) );
  OR U2035 ( .A(n1651), .B(n1650), .Z(n1655) );
  NANDN U2036 ( .A(n1653), .B(n1652), .Z(n1654) );
  AND U2037 ( .A(n1655), .B(n1654), .Z(n1783) );
  OR U2038 ( .A(n1657), .B(n1656), .Z(n1661) );
  OR U2039 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U2040 ( .A(n1661), .B(n1660), .Z(n1913) );
  OR U2041 ( .A(n1663), .B(n1662), .Z(n1667) );
  NAND U2042 ( .A(n1665), .B(n1664), .Z(n1666) );
  NAND U2043 ( .A(n1667), .B(n1666), .Z(n1797) );
  AND U2044 ( .A(x[87]), .B(y[193]), .Z(n1831) );
  XNOR U2045 ( .A(o[24]), .B(n1831), .Z(n1846) );
  NANDN U2046 ( .A(n45), .B(y[216]), .Z(n1844) );
  IV U2047 ( .A(x[88]), .Z(n8865) );
  NANDN U2048 ( .A(n8865), .B(y[192]), .Z(n1843) );
  XOR U2049 ( .A(n1844), .B(n1843), .Z(n1845) );
  OR U2050 ( .A(n1669), .B(n1668), .Z(n1672) );
  NAND U2051 ( .A(n1670), .B(n1832), .Z(n1671) );
  AND U2052 ( .A(n1672), .B(n1671), .Z(n1901) );
  NANDN U2053 ( .A(n52), .B(y[209]), .Z(n1834) );
  ANDN U2054 ( .B(x[82]), .A(n2651), .Z(n1674) );
  ANDN U2055 ( .B(x[81]), .A(n2878), .Z(n1673) );
  XNOR U2056 ( .A(n1674), .B(n1673), .Z(n1833) );
  XNOR U2057 ( .A(n1834), .B(n1833), .Z(n1900) );
  XOR U2058 ( .A(n1901), .B(n1900), .Z(n1903) );
  XOR U2059 ( .A(n1902), .B(n1903), .Z(n1869) );
  OR U2060 ( .A(n1676), .B(n1675), .Z(n1680) );
  NANDN U2061 ( .A(n1678), .B(n1677), .Z(n1679) );
  AND U2062 ( .A(n1680), .B(n1679), .Z(n1867) );
  NANDN U2063 ( .A(n1682), .B(n1681), .Z(n1686) );
  OR U2064 ( .A(n1684), .B(n1683), .Z(n1685) );
  AND U2065 ( .A(n1686), .B(n1685), .Z(n1868) );
  XOR U2066 ( .A(n1869), .B(n1870), .Z(n1796) );
  NANDN U2067 ( .A(n1688), .B(n1687), .Z(n1692) );
  NANDN U2068 ( .A(n1690), .B(n1689), .Z(n1691) );
  NAND U2069 ( .A(n1692), .B(n1691), .Z(n1795) );
  XNOR U2070 ( .A(n1796), .B(n1795), .Z(n1798) );
  XOR U2071 ( .A(n1797), .B(n1798), .Z(n1909) );
  NANDN U2072 ( .A(n1694), .B(n1693), .Z(n1698) );
  NANDN U2073 ( .A(n1696), .B(n1695), .Z(n1697) );
  NAND U2074 ( .A(n1698), .B(n1697), .Z(n1858) );
  OR U2075 ( .A(n1700), .B(n1699), .Z(n1704) );
  NANDN U2076 ( .A(n1702), .B(n1701), .Z(n1703) );
  AND U2077 ( .A(n1704), .B(n1703), .Z(n1855) );
  OR U2078 ( .A(n1706), .B(n1705), .Z(n1710) );
  NANDN U2079 ( .A(n1708), .B(n1707), .Z(n1709) );
  NAND U2080 ( .A(n1710), .B(n1709), .Z(n1856) );
  XNOR U2081 ( .A(n1858), .B(n1857), .Z(n1906) );
  NANDN U2082 ( .A(n1712), .B(n1711), .Z(n1716) );
  NANDN U2083 ( .A(n1714), .B(n1713), .Z(n1715) );
  AND U2084 ( .A(n1716), .B(n1715), .Z(n1907) );
  XOR U2085 ( .A(n1909), .B(n1908), .Z(n1912) );
  XNOR U2086 ( .A(n1913), .B(n1912), .Z(n1915) );
  NANDN U2087 ( .A(n1718), .B(n1717), .Z(n1722) );
  OR U2088 ( .A(n1720), .B(n1719), .Z(n1721) );
  NAND U2089 ( .A(n1722), .B(n1721), .Z(n1792) );
  NANDN U2090 ( .A(n53), .B(y[208]), .Z(n1808) );
  NANDN U2091 ( .A(n56), .B(y[205]), .Z(n1807) );
  XOR U2092 ( .A(n1808), .B(n1807), .Z(n1809) );
  NANDN U2093 ( .A(n2906), .B(x[78]), .Z(n1810) );
  XOR U2094 ( .A(n1809), .B(n1810), .Z(n1815) );
  AND U2095 ( .A(y[207]), .B(x[73]), .Z(n1814) );
  NAND U2096 ( .A(y[206]), .B(x[74]), .Z(n1813) );
  XOR U2097 ( .A(n1814), .B(n1813), .Z(n1816) );
  XOR U2098 ( .A(n1815), .B(n1816), .Z(n1851) );
  OR U2099 ( .A(n1724), .B(n1723), .Z(n1728) );
  NANDN U2100 ( .A(n1726), .B(n1725), .Z(n1727) );
  AND U2101 ( .A(n1728), .B(n1727), .Z(n1849) );
  NANDN U2102 ( .A(n2837), .B(x[79]), .Z(n1838) );
  NANDN U2103 ( .A(n48), .B(y[213]), .Z(n1837) );
  XOR U2104 ( .A(n1838), .B(n1837), .Z(n1839) );
  NANDN U2105 ( .A(n2449), .B(x[68]), .Z(n1840) );
  XOR U2106 ( .A(n1839), .B(n1840), .Z(n1850) );
  XNOR U2107 ( .A(n1851), .B(n1852), .Z(n1803) );
  OR U2108 ( .A(n1730), .B(n1729), .Z(n1734) );
  NANDN U2109 ( .A(n1732), .B(n1731), .Z(n1733) );
  AND U2110 ( .A(n1734), .B(n1733), .Z(n1863) );
  NANDN U2111 ( .A(n1735), .B(n1814), .Z(n1739) );
  OR U2112 ( .A(n1737), .B(n1736), .Z(n1738) );
  NAND U2113 ( .A(n1739), .B(n1738), .Z(n1861) );
  NANDN U2114 ( .A(n50), .B(y[211]), .Z(n1893) );
  NANDN U2115 ( .A(n43), .B(x[85]), .Z(n1892) );
  XOR U2116 ( .A(n1893), .B(n1892), .Z(n1894) );
  NANDN U2117 ( .A(n8890), .B(y[200]), .Z(n1895) );
  XOR U2118 ( .A(n1894), .B(n1895), .Z(n1882) );
  OR U2119 ( .A(n1741), .B(n1740), .Z(n1745) );
  NAND U2120 ( .A(n1743), .B(n1742), .Z(n1744) );
  AND U2121 ( .A(n1745), .B(n1744), .Z(n1879) );
  NANDN U2122 ( .A(n2702), .B(x[70]), .Z(n1887) );
  NANDN U2123 ( .A(n1746), .B(x[83]), .Z(n1886) );
  XOR U2124 ( .A(n1887), .B(n1886), .Z(n1888) );
  NANDN U2125 ( .A(n2897), .B(x[84]), .Z(n1889) );
  XOR U2126 ( .A(n1888), .B(n1889), .Z(n1880) );
  XOR U2127 ( .A(n1879), .B(n1880), .Z(n1881) );
  XOR U2128 ( .A(n1882), .B(n1881), .Z(n1862) );
  XOR U2129 ( .A(n1861), .B(n1862), .Z(n1864) );
  NANDN U2130 ( .A(n47), .B(y[214]), .Z(n1826) );
  NANDN U2131 ( .A(n2602), .B(x[86]), .Z(n1825) );
  XNOR U2132 ( .A(n1826), .B(n1825), .Z(n1828) );
  XOR U2133 ( .A(n1827), .B(n1828), .Z(n1876) );
  ANDN U2134 ( .B(y[195]), .A(n8890), .Z(n1747) );
  ANDN U2135 ( .B(x[84]), .A(n2878), .Z(n2289) );
  NAND U2136 ( .A(n1747), .B(n2289), .Z(n1750) );
  NANDN U2137 ( .A(n1748), .B(n1979), .Z(n1749) );
  AND U2138 ( .A(n1750), .B(n1749), .Z(n1873) );
  NANDN U2139 ( .A(n1751), .B(o[23]), .Z(n1822) );
  IV U2140 ( .A(y[215]), .Z(n2894) );
  NANDN U2141 ( .A(n2894), .B(x[65]), .Z(n1820) );
  XNOR U2142 ( .A(n1752), .B(n1820), .Z(n1821) );
  XOR U2143 ( .A(n1822), .B(n1821), .Z(n1874) );
  XNOR U2144 ( .A(n1876), .B(n1875), .Z(n1802) );
  XOR U2145 ( .A(n1801), .B(n1802), .Z(n1804) );
  XOR U2146 ( .A(n1803), .B(n1804), .Z(n1789) );
  OR U2147 ( .A(n1754), .B(n1753), .Z(n1758) );
  NANDN U2148 ( .A(n1756), .B(n1755), .Z(n1757) );
  NAND U2149 ( .A(n1758), .B(n1757), .Z(n1790) );
  XOR U2150 ( .A(n1789), .B(n1790), .Z(n1791) );
  XOR U2151 ( .A(n1792), .B(n1791), .Z(n1914) );
  XNOR U2152 ( .A(n1915), .B(n1914), .Z(n1784) );
  XOR U2153 ( .A(n1783), .B(n1784), .Z(n1785) );
  OR U2154 ( .A(n1760), .B(n1759), .Z(n1764) );
  OR U2155 ( .A(n1762), .B(n1761), .Z(n1763) );
  NAND U2156 ( .A(n1764), .B(n1763), .Z(n1921) );
  OR U2157 ( .A(n1766), .B(n1765), .Z(n1770) );
  NANDN U2158 ( .A(n1768), .B(n1767), .Z(n1769) );
  AND U2159 ( .A(n1770), .B(n1769), .Z(n1918) );
  OR U2160 ( .A(n1772), .B(n1771), .Z(n1776) );
  OR U2161 ( .A(n1774), .B(n1773), .Z(n1775) );
  NAND U2162 ( .A(n1776), .B(n1775), .Z(n1919) );
  XNOR U2163 ( .A(n1918), .B(n1919), .Z(n1920) );
  XOR U2164 ( .A(n1921), .B(n1920), .Z(n1786) );
  XOR U2165 ( .A(n1785), .B(n1786), .Z(n1780) );
  XOR U2166 ( .A(n1779), .B(n1780), .Z(N57) );
  NANDN U2167 ( .A(n1778), .B(n1777), .Z(n1782) );
  NANDN U2168 ( .A(n1780), .B(n1779), .Z(n1781) );
  NAND U2169 ( .A(n1782), .B(n1781), .Z(n1924) );
  OR U2170 ( .A(n1784), .B(n1783), .Z(n1788) );
  NANDN U2171 ( .A(n1786), .B(n1785), .Z(n1787) );
  AND U2172 ( .A(n1788), .B(n1787), .Z(n1925) );
  XNOR U2173 ( .A(n1924), .B(n1925), .Z(n1926) );
  OR U2174 ( .A(n1790), .B(n1789), .Z(n1794) );
  NAND U2175 ( .A(n1792), .B(n1791), .Z(n1793) );
  NAND U2176 ( .A(n1794), .B(n1793), .Z(n1944) );
  OR U2177 ( .A(n1796), .B(n1795), .Z(n1800) );
  NANDN U2178 ( .A(n1798), .B(n1797), .Z(n1799) );
  NAND U2179 ( .A(n1800), .B(n1799), .Z(n2068) );
  NANDN U2180 ( .A(n1802), .B(n1801), .Z(n1806) );
  OR U2181 ( .A(n1804), .B(n1803), .Z(n1805) );
  AND U2182 ( .A(n1806), .B(n1805), .Z(n2066) );
  OR U2183 ( .A(n1808), .B(n1807), .Z(n1812) );
  NANDN U2184 ( .A(n1810), .B(n1809), .Z(n1811) );
  NAND U2185 ( .A(n1812), .B(n1811), .Z(n1999) );
  ANDN U2186 ( .B(y[206]), .A(n56), .Z(n1958) );
  ANDN U2187 ( .B(y[205]), .A(n57), .Z(n1956) );
  ANDN U2188 ( .B(y[210]), .A(n52), .Z(n1955) );
  XOR U2189 ( .A(n1956), .B(n1955), .Z(n1957) );
  XOR U2190 ( .A(n1958), .B(n1957), .Z(n1996) );
  NANDN U2191 ( .A(n58), .B(y[204]), .Z(n1991) );
  NANDN U2192 ( .A(n46), .B(y[216]), .Z(n1990) );
  XOR U2193 ( .A(n1991), .B(n1990), .Z(n1992) );
  NANDN U2194 ( .A(n8865), .B(y[193]), .Z(n1954) );
  XOR U2195 ( .A(o[25]), .B(n1954), .Z(n1993) );
  XOR U2196 ( .A(n1992), .B(n1993), .Z(n1997) );
  XNOR U2197 ( .A(n1996), .B(n1997), .Z(n1998) );
  XNOR U2198 ( .A(n1999), .B(n1998), .Z(n2055) );
  NANDN U2199 ( .A(n1814), .B(n1813), .Z(n1818) );
  NANDN U2200 ( .A(n1816), .B(n1815), .Z(n1817) );
  NAND U2201 ( .A(n1818), .B(n1817), .Z(n2054) );
  OR U2202 ( .A(n1820), .B(n1819), .Z(n1824) );
  NANDN U2203 ( .A(n1822), .B(n1821), .Z(n1823) );
  NAND U2204 ( .A(n1824), .B(n1823), .Z(n2045) );
  OR U2205 ( .A(n1826), .B(n1825), .Z(n1830) );
  NANDN U2206 ( .A(n1828), .B(n1827), .Z(n1829) );
  AND U2207 ( .A(n1830), .B(n1829), .Z(n2042) );
  NANDN U2208 ( .A(n2851), .B(x[72]), .Z(n2041) );
  XOR U2209 ( .A(n2038), .B(n2039), .Z(n2040) );
  XNOR U2210 ( .A(n2041), .B(n2040), .Z(n2026) );
  AND U2211 ( .A(n1831), .B(o[24]), .Z(n2035) );
  NAND U2212 ( .A(x[89]), .B(y[192]), .Z(n2032) );
  NANDN U2213 ( .A(n45), .B(y[217]), .Z(n2033) );
  XNOR U2214 ( .A(n2032), .B(n2033), .Z(n2034) );
  XOR U2215 ( .A(n2035), .B(n2034), .Z(n2027) );
  XOR U2216 ( .A(n2026), .B(n2027), .Z(n2029) );
  ANDN U2217 ( .B(x[82]), .A(n2878), .Z(n1885) );
  IV U2218 ( .A(n1885), .Z(n1973) );
  NANDN U2219 ( .A(n1973), .B(n1832), .Z(n1836) );
  OR U2220 ( .A(n1834), .B(n1833), .Z(n1835) );
  NAND U2221 ( .A(n1836), .B(n1835), .Z(n2028) );
  XOR U2222 ( .A(n2029), .B(n2028), .Z(n2043) );
  XNOR U2223 ( .A(n2045), .B(n2044), .Z(n2057) );
  XOR U2224 ( .A(n2056), .B(n2057), .Z(n2062) );
  OR U2225 ( .A(n1838), .B(n1837), .Z(n1842) );
  NANDN U2226 ( .A(n1840), .B(n1839), .Z(n1841) );
  AND U2227 ( .A(n1842), .B(n1841), .Z(n2016) );
  OR U2228 ( .A(n1844), .B(n1843), .Z(n1848) );
  NANDN U2229 ( .A(n1846), .B(n1845), .Z(n1847) );
  NAND U2230 ( .A(n1848), .B(n1847), .Z(n2014) );
  NANDN U2231 ( .A(n48), .B(y[214]), .Z(n1987) );
  NANDN U2232 ( .A(n47), .B(y[215]), .Z(n1985) );
  XOR U2233 ( .A(n1984), .B(n1985), .Z(n1986) );
  XNOR U2234 ( .A(n1987), .B(n1986), .Z(n2015) );
  XOR U2235 ( .A(n2014), .B(n2015), .Z(n2017) );
  OR U2236 ( .A(n1850), .B(n1849), .Z(n1854) );
  NANDN U2237 ( .A(n1852), .B(n1851), .Z(n1853) );
  NAND U2238 ( .A(n1854), .B(n1853), .Z(n2061) );
  XOR U2239 ( .A(n2060), .B(n2061), .Z(n2063) );
  XOR U2240 ( .A(n2062), .B(n2063), .Z(n2067) );
  XOR U2241 ( .A(n2068), .B(n2069), .Z(n1942) );
  OR U2242 ( .A(n1856), .B(n1855), .Z(n1860) );
  NANDN U2243 ( .A(n1858), .B(n1857), .Z(n1859) );
  AND U2244 ( .A(n1860), .B(n1859), .Z(n1937) );
  NANDN U2245 ( .A(n1862), .B(n1861), .Z(n1866) );
  OR U2246 ( .A(n1864), .B(n1863), .Z(n1865) );
  NAND U2247 ( .A(n1866), .B(n1865), .Z(n1949) );
  OR U2248 ( .A(n1868), .B(n1867), .Z(n1872) );
  NAND U2249 ( .A(n1870), .B(n1869), .Z(n1871) );
  NAND U2250 ( .A(n1872), .B(n1871), .Z(n1948) );
  OR U2251 ( .A(n1874), .B(n1873), .Z(n1878) );
  NANDN U2252 ( .A(n1876), .B(n1875), .Z(n1877) );
  NAND U2253 ( .A(n1878), .B(n1877), .Z(n2023) );
  OR U2254 ( .A(n1880), .B(n1879), .Z(n1884) );
  NANDN U2255 ( .A(n1882), .B(n1881), .Z(n1883) );
  NAND U2256 ( .A(n1884), .B(n1883), .Z(n2021) );
  ANDN U2257 ( .B(y[194]), .A(n8656), .Z(n1970) );
  IV U2258 ( .A(y[213]), .Z(n2705) );
  ANDN U2259 ( .B(x[68]), .A(n2705), .Z(n1968) );
  ANDN U2260 ( .B(y[201]), .A(n8890), .Z(n1967) );
  XOR U2261 ( .A(n1968), .B(n1967), .Z(n1969) );
  XOR U2262 ( .A(n1970), .B(n1969), .Z(n2010) );
  ANDN U2263 ( .B(y[202]), .A(n60), .Z(n1976) );
  ANDN U2264 ( .B(y[211]), .A(n51), .Z(n1974) );
  XOR U2265 ( .A(n1885), .B(n1974), .Z(n1975) );
  XOR U2266 ( .A(n1976), .B(n1975), .Z(n2008) );
  OR U2267 ( .A(n1887), .B(n1886), .Z(n1891) );
  NANDN U2268 ( .A(n1889), .B(n1888), .Z(n1890) );
  AND U2269 ( .A(n1891), .B(n1890), .Z(n2009) );
  XOR U2270 ( .A(n2008), .B(n2009), .Z(n2011) );
  XNOR U2271 ( .A(n2010), .B(n2011), .Z(n2048) );
  ANDN U2272 ( .B(y[195]), .A(n8864), .Z(n1964) );
  ANDN U2273 ( .B(x[69]), .A(n2449), .Z(n1962) );
  ANDN U2274 ( .B(x[81]), .A(n2512), .Z(n1961) );
  XOR U2275 ( .A(n1962), .B(n1961), .Z(n1963) );
  XOR U2276 ( .A(n1964), .B(n1963), .Z(n2002) );
  OR U2277 ( .A(n1893), .B(n1892), .Z(n1897) );
  NANDN U2278 ( .A(n1895), .B(n1894), .Z(n1896) );
  AND U2279 ( .A(n1897), .B(n1896), .Z(n2003) );
  XOR U2280 ( .A(n2002), .B(n2003), .Z(n2005) );
  NANDN U2281 ( .A(n8885), .B(y[197]), .Z(n1981) );
  ANDN U2282 ( .B(y[198]), .A(n8824), .Z(n1899) );
  NANDN U2283 ( .A(n8827), .B(y[196]), .Z(n1898) );
  XOR U2284 ( .A(n1899), .B(n1898), .Z(n1980) );
  XNOR U2285 ( .A(n2005), .B(n2004), .Z(n2049) );
  XNOR U2286 ( .A(n2048), .B(n2049), .Z(n2051) );
  OR U2287 ( .A(n1901), .B(n1900), .Z(n1905) );
  NAND U2288 ( .A(n1903), .B(n1902), .Z(n1904) );
  NAND U2289 ( .A(n1905), .B(n1904), .Z(n2050) );
  XOR U2290 ( .A(n2051), .B(n2050), .Z(n2020) );
  XNOR U2291 ( .A(n2021), .B(n2020), .Z(n2022) );
  XNOR U2292 ( .A(n2023), .B(n2022), .Z(n1950) );
  XOR U2293 ( .A(n1937), .B(n1936), .Z(n1939) );
  OR U2294 ( .A(n1907), .B(n1906), .Z(n1911) );
  NAND U2295 ( .A(n1909), .B(n1908), .Z(n1910) );
  NAND U2296 ( .A(n1911), .B(n1910), .Z(n1938) );
  XOR U2297 ( .A(n1939), .B(n1938), .Z(n1943) );
  XOR U2298 ( .A(n1942), .B(n1943), .Z(n1945) );
  XNOR U2299 ( .A(n1944), .B(n1945), .Z(n1933) );
  OR U2300 ( .A(n1913), .B(n1912), .Z(n1917) );
  OR U2301 ( .A(n1915), .B(n1914), .Z(n1916) );
  AND U2302 ( .A(n1917), .B(n1916), .Z(n1930) );
  OR U2303 ( .A(n1919), .B(n1918), .Z(n1923) );
  OR U2304 ( .A(n1921), .B(n1920), .Z(n1922) );
  NAND U2305 ( .A(n1923), .B(n1922), .Z(n1931) );
  XOR U2306 ( .A(n1930), .B(n1931), .Z(n1932) );
  XOR U2307 ( .A(n1933), .B(n1932), .Z(n1927) );
  XOR U2308 ( .A(n1926), .B(n1927), .Z(N58) );
  NANDN U2309 ( .A(n1925), .B(n1924), .Z(n1929) );
  NANDN U2310 ( .A(n1927), .B(n1926), .Z(n1928) );
  NAND U2311 ( .A(n1929), .B(n1928), .Z(n2072) );
  OR U2312 ( .A(n1931), .B(n1930), .Z(n1935) );
  NANDN U2313 ( .A(n1933), .B(n1932), .Z(n1934) );
  AND U2314 ( .A(n1935), .B(n1934), .Z(n2073) );
  XNOR U2315 ( .A(n2072), .B(n2073), .Z(n2074) );
  NANDN U2316 ( .A(n1937), .B(n1936), .Z(n1941) );
  OR U2317 ( .A(n1939), .B(n1938), .Z(n1940) );
  NAND U2318 ( .A(n1941), .B(n1940), .Z(n2081) );
  NANDN U2319 ( .A(n1943), .B(n1942), .Z(n1947) );
  NANDN U2320 ( .A(n1945), .B(n1944), .Z(n1946) );
  AND U2321 ( .A(n1947), .B(n1946), .Z(n2078) );
  OR U2322 ( .A(n1949), .B(n1948), .Z(n1953) );
  NANDN U2323 ( .A(n1951), .B(n1950), .Z(n1952) );
  NAND U2324 ( .A(n1953), .B(n1952), .Z(n2222) );
  NANDN U2325 ( .A(n1954), .B(o[25]), .Z(n2186) );
  NAND U2326 ( .A(x[78]), .B(y[204]), .Z(n2184) );
  NAND U2327 ( .A(x[65]), .B(y[217]), .Z(n2185) );
  XNOR U2328 ( .A(n2184), .B(n2185), .Z(n2187) );
  XNOR U2329 ( .A(n2186), .B(n2187), .Z(n2136) );
  NANDN U2330 ( .A(n45), .B(y[218]), .Z(n2149) );
  AND U2331 ( .A(y[192]), .B(x[90]), .Z(n2148) );
  XNOR U2332 ( .A(n2149), .B(n2148), .Z(n2151) );
  NANDN U2333 ( .A(n2857), .B(x[89]), .Z(n2196) );
  XNOR U2334 ( .A(n2196), .B(o[26]), .Z(n2150) );
  XNOR U2335 ( .A(n2151), .B(n2150), .Z(n2137) );
  XNOR U2336 ( .A(n2136), .B(n2137), .Z(n2139) );
  OR U2337 ( .A(n1956), .B(n1955), .Z(n1960) );
  NANDN U2338 ( .A(n1958), .B(n1957), .Z(n1959) );
  NAND U2339 ( .A(n1960), .B(n1959), .Z(n2138) );
  XOR U2340 ( .A(n2139), .B(n2138), .Z(n2117) );
  OR U2341 ( .A(n1962), .B(n1961), .Z(n1966) );
  NANDN U2342 ( .A(n1964), .B(n1963), .Z(n1965) );
  NAND U2343 ( .A(n1966), .B(n1965), .Z(n2114) );
  OR U2344 ( .A(n1968), .B(n1967), .Z(n1972) );
  NANDN U2345 ( .A(n1970), .B(n1969), .Z(n1971) );
  AND U2346 ( .A(n1972), .B(n1971), .Z(n2115) );
  XNOR U2347 ( .A(n2114), .B(n2115), .Z(n2116) );
  XOR U2348 ( .A(n2117), .B(n2116), .Z(n2157) );
  NAND U2349 ( .A(x[68]), .B(y[214]), .Z(n2102) );
  XOR U2350 ( .A(n2103), .B(n2102), .Z(n2105) );
  XNOR U2351 ( .A(n2104), .B(n2105), .Z(n2108) );
  NANDN U2352 ( .A(n1974), .B(n1973), .Z(n1978) );
  NANDN U2353 ( .A(n1976), .B(n1975), .Z(n1977) );
  NAND U2354 ( .A(n1978), .B(n1977), .Z(n2109) );
  XOR U2355 ( .A(n2108), .B(n2109), .Z(n2111) );
  NANDN U2356 ( .A(n2878), .B(x[83]), .Z(n2179) );
  AND U2357 ( .A(x[75]), .B(y[207]), .Z(n2178) );
  XNOR U2358 ( .A(n2179), .B(n2178), .Z(n2180) );
  NANDN U2359 ( .A(n2894), .B(x[67]), .Z(n2181) );
  XNOR U2360 ( .A(n2180), .B(n2181), .Z(n2110) );
  XOR U2361 ( .A(n2111), .B(n2110), .Z(n2154) );
  ANDN U2362 ( .B(x[85]), .A(n2651), .Z(n2282) );
  NAND U2363 ( .A(n1979), .B(n2282), .Z(n1983) );
  OR U2364 ( .A(n1981), .B(n1980), .Z(n1982) );
  NAND U2365 ( .A(n1983), .B(n1982), .Z(n2085) );
  NANDN U2366 ( .A(n8864), .B(y[196]), .Z(n2093) );
  NANDN U2367 ( .A(n43), .B(x[87]), .Z(n2090) );
  XNOR U2368 ( .A(n2091), .B(n2090), .Z(n2092) );
  XNOR U2369 ( .A(n2093), .B(n2092), .Z(n2084) );
  XNOR U2370 ( .A(n2085), .B(n2084), .Z(n2087) );
  NAND U2371 ( .A(x[84]), .B(y[198]), .Z(n2192) );
  NAND U2372 ( .A(y[197]), .B(x[85]), .Z(n2190) );
  XOR U2373 ( .A(n2191), .B(n2190), .Z(n2193) );
  XOR U2374 ( .A(n2192), .B(n2193), .Z(n2086) );
  XNOR U2375 ( .A(n2087), .B(n2086), .Z(n2155) );
  XOR U2376 ( .A(n2154), .B(n2155), .Z(n2156) );
  XOR U2377 ( .A(n2157), .B(n2156), .Z(n2162) );
  NANDN U2378 ( .A(n1985), .B(n1984), .Z(n1989) );
  OR U2379 ( .A(n1987), .B(n1986), .Z(n1988) );
  NAND U2380 ( .A(n1989), .B(n1988), .Z(n2119) );
  OR U2381 ( .A(n1991), .B(n1990), .Z(n1995) );
  NANDN U2382 ( .A(n1993), .B(n1992), .Z(n1994) );
  NAND U2383 ( .A(n1995), .B(n1994), .Z(n2118) );
  XNOR U2384 ( .A(n2119), .B(n2118), .Z(n2120) );
  NAND U2385 ( .A(y[209]), .B(x[73]), .Z(n2199) );
  NAND U2386 ( .A(x[70]), .B(y[212]), .Z(n2197) );
  NAND U2387 ( .A(x[72]), .B(y[210]), .Z(n2198) );
  XNOR U2388 ( .A(n2197), .B(n2198), .Z(n2200) );
  XOR U2389 ( .A(n2199), .B(n2200), .Z(n2175) );
  AND U2390 ( .A(x[71]), .B(y[211]), .Z(n2172) );
  NAND U2391 ( .A(x[76]), .B(y[206]), .Z(n2142) );
  NAND U2392 ( .A(y[213]), .B(x[69]), .Z(n2143) );
  XNOR U2393 ( .A(n2142), .B(n2143), .Z(n2145) );
  XNOR U2394 ( .A(n2144), .B(n2145), .Z(n2173) );
  XNOR U2395 ( .A(n2172), .B(n2173), .Z(n2174) );
  XNOR U2396 ( .A(n2175), .B(n2174), .Z(n2121) );
  NANDN U2397 ( .A(n1997), .B(n1996), .Z(n2001) );
  NAND U2398 ( .A(n1999), .B(n1998), .Z(n2000) );
  AND U2399 ( .A(n2001), .B(n2000), .Z(n2161) );
  XNOR U2400 ( .A(n2160), .B(n2161), .Z(n2163) );
  XNOR U2401 ( .A(n2162), .B(n2163), .Z(n2124) );
  NANDN U2402 ( .A(n2003), .B(n2002), .Z(n2007) );
  NANDN U2403 ( .A(n2005), .B(n2004), .Z(n2006) );
  NAND U2404 ( .A(n2007), .B(n2006), .Z(n2210) );
  NANDN U2405 ( .A(n2009), .B(n2008), .Z(n2013) );
  NANDN U2406 ( .A(n2011), .B(n2010), .Z(n2012) );
  NAND U2407 ( .A(n2013), .B(n2012), .Z(n2209) );
  XNOR U2408 ( .A(n2210), .B(n2209), .Z(n2211) );
  NANDN U2409 ( .A(n2015), .B(n2014), .Z(n2019) );
  OR U2410 ( .A(n2017), .B(n2016), .Z(n2018) );
  NAND U2411 ( .A(n2019), .B(n2018), .Z(n2212) );
  XOR U2412 ( .A(n2124), .B(n2125), .Z(n2127) );
  NANDN U2413 ( .A(n2021), .B(n2020), .Z(n2025) );
  NANDN U2414 ( .A(n2023), .B(n2022), .Z(n2024) );
  AND U2415 ( .A(n2025), .B(n2024), .Z(n2126) );
  XOR U2416 ( .A(n2127), .B(n2126), .Z(n2221) );
  XNOR U2417 ( .A(n2222), .B(n2221), .Z(n2224) );
  NANDN U2418 ( .A(n2027), .B(n2026), .Z(n2031) );
  NANDN U2419 ( .A(n2029), .B(n2028), .Z(n2030) );
  AND U2420 ( .A(n2031), .B(n2030), .Z(n2203) );
  NANDN U2421 ( .A(n47), .B(y[216]), .Z(n2097) );
  XNOR U2422 ( .A(n2097), .B(n2096), .Z(n2099) );
  AND U2423 ( .A(x[88]), .B(y[194]), .Z(n2098) );
  XOR U2424 ( .A(n2099), .B(n2098), .Z(n2130) );
  NAND U2425 ( .A(n2033), .B(n2032), .Z(n2037) );
  OR U2426 ( .A(n2035), .B(n2034), .Z(n2036) );
  AND U2427 ( .A(n2037), .B(n2036), .Z(n2131) );
  XNOR U2428 ( .A(n2130), .B(n2131), .Z(n2133) );
  XOR U2429 ( .A(n2133), .B(n2132), .Z(n2204) );
  XNOR U2430 ( .A(n2203), .B(n2204), .Z(n2206) );
  OR U2431 ( .A(n2043), .B(n2042), .Z(n2047) );
  NAND U2432 ( .A(n2045), .B(n2044), .Z(n2046) );
  AND U2433 ( .A(n2047), .B(n2046), .Z(n2205) );
  XOR U2434 ( .A(n2206), .B(n2205), .Z(n2169) );
  OR U2435 ( .A(n2049), .B(n2048), .Z(n2053) );
  OR U2436 ( .A(n2051), .B(n2050), .Z(n2052) );
  AND U2437 ( .A(n2053), .B(n2052), .Z(n2166) );
  OR U2438 ( .A(n2055), .B(n2054), .Z(n2059) );
  NANDN U2439 ( .A(n2057), .B(n2056), .Z(n2058) );
  NAND U2440 ( .A(n2059), .B(n2058), .Z(n2167) );
  XOR U2441 ( .A(n2166), .B(n2167), .Z(n2168) );
  XOR U2442 ( .A(n2169), .B(n2168), .Z(n2223) );
  XNOR U2443 ( .A(n2224), .B(n2223), .Z(n2218) );
  NANDN U2444 ( .A(n2061), .B(n2060), .Z(n2065) );
  NANDN U2445 ( .A(n2063), .B(n2062), .Z(n2064) );
  NAND U2446 ( .A(n2065), .B(n2064), .Z(n2216) );
  OR U2447 ( .A(n2067), .B(n2066), .Z(n2071) );
  NANDN U2448 ( .A(n2069), .B(n2068), .Z(n2070) );
  NAND U2449 ( .A(n2071), .B(n2070), .Z(n2215) );
  XNOR U2450 ( .A(n2218), .B(n2217), .Z(n2079) );
  XNOR U2451 ( .A(n2081), .B(n2080), .Z(n2075) );
  XOR U2452 ( .A(n2074), .B(n2075), .Z(N59) );
  NANDN U2453 ( .A(n2073), .B(n2072), .Z(n2077) );
  NANDN U2454 ( .A(n2075), .B(n2074), .Z(n2076) );
  NAND U2455 ( .A(n2077), .B(n2076), .Z(n2227) );
  OR U2456 ( .A(n2079), .B(n2078), .Z(n2083) );
  NANDN U2457 ( .A(n2081), .B(n2080), .Z(n2082) );
  NAND U2458 ( .A(n2083), .B(n2082), .Z(n2228) );
  XNOR U2459 ( .A(n2227), .B(n2228), .Z(n2229) );
  OR U2460 ( .A(n2085), .B(n2084), .Z(n2089) );
  OR U2461 ( .A(n2087), .B(n2086), .Z(n2088) );
  NAND U2462 ( .A(n2089), .B(n2088), .Z(n2252) );
  NANDN U2463 ( .A(n2091), .B(n2090), .Z(n2095) );
  NAND U2464 ( .A(n2093), .B(n2092), .Z(n2094) );
  NAND U2465 ( .A(n2095), .B(n2094), .Z(n2326) );
  NANDN U2466 ( .A(n2097), .B(n2096), .Z(n2101) );
  NAND U2467 ( .A(n2099), .B(n2098), .Z(n2100) );
  NAND U2468 ( .A(n2101), .B(n2100), .Z(n2327) );
  XNOR U2469 ( .A(n2326), .B(n2327), .Z(n2329) );
  NANDN U2470 ( .A(n2103), .B(n2102), .Z(n2107) );
  OR U2471 ( .A(n2105), .B(n2104), .Z(n2106) );
  NAND U2472 ( .A(n2107), .B(n2106), .Z(n2322) );
  NAND U2473 ( .A(y[210]), .B(x[73]), .Z(n2283) );
  NAND U2474 ( .A(y[201]), .B(x[82]), .Z(n2281) );
  XOR U2475 ( .A(n2282), .B(n2281), .Z(n2284) );
  XOR U2476 ( .A(n2283), .B(n2284), .Z(n2323) );
  XNOR U2477 ( .A(n2322), .B(n2323), .Z(n2324) );
  NAND U2478 ( .A(x[64]), .B(y[219]), .Z(n2271) );
  AND U2479 ( .A(y[193]), .B(x[90]), .Z(n2287) );
  XOR U2480 ( .A(o[27]), .B(n2287), .Z(n2270) );
  NAND U2481 ( .A(y[192]), .B(x[91]), .Z(n2269) );
  XOR U2482 ( .A(n2270), .B(n2269), .Z(n2272) );
  XOR U2483 ( .A(n2271), .B(n2272), .Z(n2325) );
  XNOR U2484 ( .A(n2324), .B(n2325), .Z(n2328) );
  XNOR U2485 ( .A(n2329), .B(n2328), .Z(n2263) );
  NANDN U2486 ( .A(n2109), .B(n2108), .Z(n2113) );
  NANDN U2487 ( .A(n2111), .B(n2110), .Z(n2112) );
  AND U2488 ( .A(n2113), .B(n2112), .Z(n2264) );
  XOR U2489 ( .A(n2263), .B(n2264), .Z(n2266) );
  XNOR U2490 ( .A(n2266), .B(n2265), .Z(n2251) );
  XNOR U2491 ( .A(n2252), .B(n2251), .Z(n2254) );
  OR U2492 ( .A(n2119), .B(n2118), .Z(n2123) );
  OR U2493 ( .A(n2121), .B(n2120), .Z(n2122) );
  NAND U2494 ( .A(n2123), .B(n2122), .Z(n2253) );
  XNOR U2495 ( .A(n2254), .B(n2253), .Z(n2377) );
  NANDN U2496 ( .A(n2125), .B(n2124), .Z(n2129) );
  OR U2497 ( .A(n2127), .B(n2126), .Z(n2128) );
  NAND U2498 ( .A(n2129), .B(n2128), .Z(n2378) );
  NAND U2499 ( .A(n2131), .B(n2130), .Z(n2135) );
  NANDN U2500 ( .A(n2133), .B(n2132), .Z(n2134) );
  NAND U2501 ( .A(n2135), .B(n2134), .Z(n2260) );
  OR U2502 ( .A(n2137), .B(n2136), .Z(n2141) );
  OR U2503 ( .A(n2139), .B(n2138), .Z(n2140) );
  NAND U2504 ( .A(n2141), .B(n2140), .Z(n2258) );
  AND U2505 ( .A(x[76]), .B(y[207]), .Z(n2353) );
  AND U2506 ( .A(y[206]), .B(x[77]), .Z(n2354) );
  XNOR U2507 ( .A(n2353), .B(n2354), .Z(n2356) );
  NANDN U2508 ( .A(n56), .B(y[208]), .Z(n2337) );
  NANDN U2509 ( .A(n8890), .B(y[203]), .Z(n2334) );
  XNOR U2510 ( .A(n2335), .B(n2334), .Z(n2336) );
  XNOR U2511 ( .A(n2337), .B(n2336), .Z(n2355) );
  XNOR U2512 ( .A(n2356), .B(n2355), .Z(n2306) );
  AND U2513 ( .A(y[216]), .B(x[67]), .Z(n2361) );
  AND U2514 ( .A(y[217]), .B(x[66]), .Z(n2359) );
  AND U2515 ( .A(x[79]), .B(y[204]), .Z(n2360) );
  XNOR U2516 ( .A(n2359), .B(n2360), .Z(n2362) );
  XOR U2517 ( .A(n2361), .B(n2362), .Z(n2304) );
  NANDN U2518 ( .A(n2705), .B(x[70]), .Z(n2296) );
  NAND U2519 ( .A(y[194]), .B(x[89]), .Z(n2294) );
  NANDN U2520 ( .A(n8824), .B(y[200]), .Z(n2295) );
  XNOR U2521 ( .A(n2294), .B(n2295), .Z(n2297) );
  XNOR U2522 ( .A(n2296), .B(n2297), .Z(n2305) );
  XNOR U2523 ( .A(n2304), .B(n2305), .Z(n2307) );
  XNOR U2524 ( .A(n2306), .B(n2307), .Z(n2333) );
  NAND U2525 ( .A(n2143), .B(n2142), .Z(n2147) );
  OR U2526 ( .A(n2145), .B(n2144), .Z(n2146) );
  NAND U2527 ( .A(n2147), .B(n2146), .Z(n2330) );
  NANDN U2528 ( .A(n2149), .B(n2148), .Z(n2153) );
  NAND U2529 ( .A(n2151), .B(n2150), .Z(n2152) );
  NAND U2530 ( .A(n2153), .B(n2152), .Z(n2331) );
  XNOR U2531 ( .A(n2330), .B(n2331), .Z(n2332) );
  XOR U2532 ( .A(n2333), .B(n2332), .Z(n2257) );
  XNOR U2533 ( .A(n2258), .B(n2257), .Z(n2259) );
  XNOR U2534 ( .A(n2260), .B(n2259), .Z(n2245) );
  NANDN U2535 ( .A(n2155), .B(n2154), .Z(n2159) );
  OR U2536 ( .A(n2157), .B(n2156), .Z(n2158) );
  NAND U2537 ( .A(n2159), .B(n2158), .Z(n2246) );
  XOR U2538 ( .A(n2245), .B(n2246), .Z(n2248) );
  OR U2539 ( .A(n2161), .B(n2160), .Z(n2165) );
  OR U2540 ( .A(n2163), .B(n2162), .Z(n2164) );
  AND U2541 ( .A(n2165), .B(n2164), .Z(n2247) );
  XNOR U2542 ( .A(n2248), .B(n2247), .Z(n2379) );
  XNOR U2543 ( .A(n2380), .B(n2379), .Z(n2373) );
  OR U2544 ( .A(n2167), .B(n2166), .Z(n2171) );
  NANDN U2545 ( .A(n2169), .B(n2168), .Z(n2170) );
  AND U2546 ( .A(n2171), .B(n2170), .Z(n2371) );
  OR U2547 ( .A(n2173), .B(n2172), .Z(n2177) );
  OR U2548 ( .A(n2175), .B(n2174), .Z(n2176) );
  AND U2549 ( .A(n2177), .B(n2176), .Z(n2241) );
  NANDN U2550 ( .A(n2179), .B(n2178), .Z(n2183) );
  NANDN U2551 ( .A(n2181), .B(n2180), .Z(n2182) );
  NAND U2552 ( .A(n2183), .B(n2182), .Z(n2312) );
  AND U2553 ( .A(x[86]), .B(y[197]), .Z(n2342) );
  AND U2554 ( .A(y[196]), .B(x[87]), .Z(n2340) );
  AND U2555 ( .A(x[72]), .B(y[211]), .Z(n2341) );
  XNOR U2556 ( .A(n2340), .B(n2341), .Z(n2343) );
  XOR U2557 ( .A(n2342), .B(n2343), .Z(n2310) );
  NANDN U2558 ( .A(n52), .B(y[212]), .Z(n2290) );
  NANDN U2559 ( .A(n43), .B(x[88]), .Z(n2288) );
  XOR U2560 ( .A(n2289), .B(n2288), .Z(n2291) );
  XNOR U2561 ( .A(n2290), .B(n2291), .Z(n2311) );
  XNOR U2562 ( .A(n2310), .B(n2311), .Z(n2313) );
  XNOR U2563 ( .A(n2312), .B(n2313), .Z(n2239) );
  NAND U2564 ( .A(n2185), .B(n2184), .Z(n2189) );
  NANDN U2565 ( .A(n2187), .B(n2186), .Z(n2188) );
  NAND U2566 ( .A(n2189), .B(n2188), .Z(n2301) );
  NANDN U2567 ( .A(n2191), .B(n2190), .Z(n2195) );
  NANDN U2568 ( .A(n2193), .B(n2192), .Z(n2194) );
  AND U2569 ( .A(n2195), .B(n2194), .Z(n2300) );
  XNOR U2570 ( .A(n2301), .B(n2300), .Z(n2303) );
  AND U2571 ( .A(y[205]), .B(x[78]), .Z(n2349) );
  ANDN U2572 ( .B(o[26]), .A(n2196), .Z(n2347) );
  AND U2573 ( .A(y[218]), .B(x[65]), .Z(n2348) );
  XNOR U2574 ( .A(n2347), .B(n2348), .Z(n2350) );
  XOR U2575 ( .A(n2349), .B(n2350), .Z(n2317) );
  NANDN U2576 ( .A(n8626), .B(y[202]), .Z(n2276) );
  AND U2577 ( .A(y[215]), .B(x[68]), .Z(n2275) );
  XNOR U2578 ( .A(n2276), .B(n2275), .Z(n2278) );
  AND U2579 ( .A(y[214]), .B(x[69]), .Z(n2277) );
  XOR U2580 ( .A(n2278), .B(n2277), .Z(n2316) );
  XOR U2581 ( .A(n2317), .B(n2316), .Z(n2319) );
  NAND U2582 ( .A(n2198), .B(n2197), .Z(n2202) );
  NANDN U2583 ( .A(n2200), .B(n2199), .Z(n2201) );
  NAND U2584 ( .A(n2202), .B(n2201), .Z(n2318) );
  XOR U2585 ( .A(n2319), .B(n2318), .Z(n2302) );
  XOR U2586 ( .A(n2303), .B(n2302), .Z(n2240) );
  XNOR U2587 ( .A(n2239), .B(n2240), .Z(n2242) );
  XOR U2588 ( .A(n2241), .B(n2242), .Z(n2365) );
  OR U2589 ( .A(n2204), .B(n2203), .Z(n2208) );
  OR U2590 ( .A(n2206), .B(n2205), .Z(n2207) );
  AND U2591 ( .A(n2208), .B(n2207), .Z(n2366) );
  XNOR U2592 ( .A(n2365), .B(n2366), .Z(n2368) );
  OR U2593 ( .A(n2210), .B(n2209), .Z(n2214) );
  OR U2594 ( .A(n2212), .B(n2211), .Z(n2213) );
  NAND U2595 ( .A(n2214), .B(n2213), .Z(n2367) );
  XOR U2596 ( .A(n2368), .B(n2367), .Z(n2372) );
  XNOR U2597 ( .A(n2371), .B(n2372), .Z(n2374) );
  XNOR U2598 ( .A(n2373), .B(n2374), .Z(n2236) );
  OR U2599 ( .A(n2216), .B(n2215), .Z(n2220) );
  NAND U2600 ( .A(n2218), .B(n2217), .Z(n2219) );
  AND U2601 ( .A(n2220), .B(n2219), .Z(n2233) );
  NAND U2602 ( .A(n2222), .B(n2221), .Z(n2226) );
  OR U2603 ( .A(n2224), .B(n2223), .Z(n2225) );
  NAND U2604 ( .A(n2226), .B(n2225), .Z(n2234) );
  XNOR U2605 ( .A(n2236), .B(n2235), .Z(n2230) );
  XOR U2606 ( .A(n2229), .B(n2230), .Z(N60) );
  NANDN U2607 ( .A(n2228), .B(n2227), .Z(n2232) );
  NANDN U2608 ( .A(n2230), .B(n2229), .Z(n2231) );
  NAND U2609 ( .A(n2232), .B(n2231), .Z(n2383) );
  OR U2610 ( .A(n2234), .B(n2233), .Z(n2238) );
  NANDN U2611 ( .A(n2236), .B(n2235), .Z(n2237) );
  NAND U2612 ( .A(n2238), .B(n2237), .Z(n2384) );
  XNOR U2613 ( .A(n2383), .B(n2384), .Z(n2385) );
  OR U2614 ( .A(n2240), .B(n2239), .Z(n2244) );
  OR U2615 ( .A(n2242), .B(n2241), .Z(n2243) );
  AND U2616 ( .A(n2244), .B(n2243), .Z(n2544) );
  NANDN U2617 ( .A(n2246), .B(n2245), .Z(n2250) );
  OR U2618 ( .A(n2248), .B(n2247), .Z(n2249) );
  NAND U2619 ( .A(n2250), .B(n2249), .Z(n2542) );
  OR U2620 ( .A(n2252), .B(n2251), .Z(n2256) );
  OR U2621 ( .A(n2254), .B(n2253), .Z(n2255) );
  NAND U2622 ( .A(n2256), .B(n2255), .Z(n2541) );
  XOR U2623 ( .A(n2542), .B(n2541), .Z(n2543) );
  XNOR U2624 ( .A(n2544), .B(n2543), .Z(n2549) );
  OR U2625 ( .A(n2258), .B(n2257), .Z(n2262) );
  OR U2626 ( .A(n2260), .B(n2259), .Z(n2261) );
  NAND U2627 ( .A(n2262), .B(n2261), .Z(n2531) );
  NANDN U2628 ( .A(n2264), .B(n2263), .Z(n2268) );
  OR U2629 ( .A(n2266), .B(n2265), .Z(n2267) );
  NAND U2630 ( .A(n2268), .B(n2267), .Z(n2532) );
  XNOR U2631 ( .A(n2531), .B(n2532), .Z(n2533) );
  NANDN U2632 ( .A(n2270), .B(n2269), .Z(n2274) );
  NANDN U2633 ( .A(n2272), .B(n2271), .Z(n2273) );
  AND U2634 ( .A(n2274), .B(n2273), .Z(n2413) );
  NANDN U2635 ( .A(n2276), .B(n2275), .Z(n2280) );
  NAND U2636 ( .A(n2278), .B(n2277), .Z(n2279) );
  NAND U2637 ( .A(n2280), .B(n2279), .Z(n2414) );
  XOR U2638 ( .A(n2413), .B(n2414), .Z(n2416) );
  NANDN U2639 ( .A(n2282), .B(n2281), .Z(n2286) );
  NANDN U2640 ( .A(n2284), .B(n2283), .Z(n2285) );
  AND U2641 ( .A(n2286), .B(n2285), .Z(n2494) );
  AND U2642 ( .A(x[74]), .B(y[210]), .Z(n2508) );
  AND U2643 ( .A(y[211]), .B(x[73]), .Z(n2506) );
  AND U2644 ( .A(y[212]), .B(x[72]), .Z(n2507) );
  XNOR U2645 ( .A(n2506), .B(n2507), .Z(n2509) );
  XNOR U2646 ( .A(n2508), .B(n2509), .Z(n2495) );
  XNOR U2647 ( .A(n2494), .B(n2495), .Z(n2496) );
  AND U2648 ( .A(y[220]), .B(x[64]), .Z(n2515) );
  AND U2649 ( .A(n2287), .B(o[27]), .Z(n2513) );
  AND U2650 ( .A(x[92]), .B(y[192]), .Z(n2514) );
  XNOR U2651 ( .A(n2513), .B(n2514), .Z(n2516) );
  XNOR U2652 ( .A(n2515), .B(n2516), .Z(n2497) );
  XNOR U2653 ( .A(n2416), .B(n2415), .Z(n2398) );
  AND U2654 ( .A(y[219]), .B(x[65]), .Z(n2470) );
  AND U2655 ( .A(y[195]), .B(x[89]), .Z(n2471) );
  XNOR U2656 ( .A(n2470), .B(n2471), .Z(n2473) );
  XNOR U2657 ( .A(n2472), .B(n2473), .Z(n2409) );
  AND U2658 ( .A(y[204]), .B(x[80]), .Z(n2478) );
  AND U2659 ( .A(y[218]), .B(x[66]), .Z(n2476) );
  AND U2660 ( .A(y[196]), .B(x[88]), .Z(n2477) );
  XNOR U2661 ( .A(n2476), .B(n2477), .Z(n2479) );
  XOR U2662 ( .A(n2478), .B(n2479), .Z(n2407) );
  NANDN U2663 ( .A(n2289), .B(n2288), .Z(n2293) );
  NANDN U2664 ( .A(n2291), .B(n2290), .Z(n2292) );
  NAND U2665 ( .A(n2293), .B(n2292), .Z(n2408) );
  XNOR U2666 ( .A(n2407), .B(n2408), .Z(n2410) );
  XNOR U2667 ( .A(n2409), .B(n2410), .Z(n2396) );
  AND U2668 ( .A(y[197]), .B(x[87]), .Z(n2437) );
  AND U2669 ( .A(y[217]), .B(x[67]), .Z(n2438) );
  XNOR U2670 ( .A(n2437), .B(n2438), .Z(n2440) );
  XOR U2671 ( .A(n2439), .B(n2440), .Z(n2421) );
  AND U2672 ( .A(x[69]), .B(y[215]), .Z(n2464) );
  AND U2673 ( .A(y[200]), .B(x[84]), .Z(n2462) );
  AND U2674 ( .A(y[199]), .B(x[85]), .Z(n2463) );
  XNOR U2675 ( .A(n2462), .B(n2463), .Z(n2465) );
  XOR U2676 ( .A(n2464), .B(n2465), .Z(n2419) );
  NAND U2677 ( .A(n2295), .B(n2294), .Z(n2299) );
  NANDN U2678 ( .A(n2297), .B(n2296), .Z(n2298) );
  NAND U2679 ( .A(n2299), .B(n2298), .Z(n2420) );
  XNOR U2680 ( .A(n2419), .B(n2420), .Z(n2422) );
  XNOR U2681 ( .A(n2421), .B(n2422), .Z(n2395) );
  XOR U2682 ( .A(n2396), .B(n2395), .Z(n2397) );
  XNOR U2683 ( .A(n2398), .B(n2397), .Z(n2536) );
  OR U2684 ( .A(n2305), .B(n2304), .Z(n2309) );
  NANDN U2685 ( .A(n2307), .B(n2306), .Z(n2308) );
  NAND U2686 ( .A(n2309), .B(n2308), .Z(n2432) );
  OR U2687 ( .A(n2311), .B(n2310), .Z(n2315) );
  NANDN U2688 ( .A(n2313), .B(n2312), .Z(n2314) );
  NAND U2689 ( .A(n2315), .B(n2314), .Z(n2431) );
  XNOR U2690 ( .A(n2432), .B(n2431), .Z(n2433) );
  XOR U2691 ( .A(n2536), .B(n2535), .Z(n2538) );
  NANDN U2692 ( .A(n2317), .B(n2316), .Z(n2321) );
  OR U2693 ( .A(n2319), .B(n2318), .Z(n2320) );
  AND U2694 ( .A(n2321), .B(n2320), .Z(n2425) );
  XOR U2695 ( .A(n2425), .B(n2426), .Z(n2427) );
  XNOR U2696 ( .A(n2427), .B(n2428), .Z(n2527) );
  AND U2697 ( .A(x[71]), .B(y[213]), .Z(n2484) );
  AND U2698 ( .A(y[209]), .B(x[75]), .Z(n2482) );
  AND U2699 ( .A(y[208]), .B(x[76]), .Z(n2483) );
  XNOR U2700 ( .A(n2482), .B(n2483), .Z(n2485) );
  XOR U2701 ( .A(n2484), .B(n2485), .Z(n2450) );
  NANDN U2702 ( .A(n2335), .B(n2334), .Z(n2339) );
  NAND U2703 ( .A(n2337), .B(n2336), .Z(n2338) );
  NAND U2704 ( .A(n2339), .B(n2338), .Z(n2451) );
  XNOR U2705 ( .A(n2450), .B(n2451), .Z(n2453) );
  NANDN U2706 ( .A(n60), .B(y[205]), .Z(n2444) );
  ANDN U2707 ( .B(x[90]), .A(n2602), .Z(n2443) );
  XOR U2708 ( .A(n2444), .B(n2443), .Z(n2445) );
  ANDN U2709 ( .B(x[91]), .A(n2857), .Z(n2601) );
  XNOR U2710 ( .A(o[28]), .B(n2601), .Z(n2446) );
  XOR U2711 ( .A(n2453), .B(n2452), .Z(n2401) );
  OR U2712 ( .A(n2341), .B(n2340), .Z(n2345) );
  OR U2713 ( .A(n2343), .B(n2342), .Z(n2344) );
  AND U2714 ( .A(n2345), .B(n2344), .Z(n2488) );
  AND U2715 ( .A(y[214]), .B(x[70]), .Z(n2458) );
  AND U2716 ( .A(x[83]), .B(y[201]), .Z(n2457) );
  XOR U2717 ( .A(n2346), .B(n2457), .Z(n2459) );
  XNOR U2718 ( .A(n2458), .B(n2459), .Z(n2489) );
  XOR U2719 ( .A(n2488), .B(n2489), .Z(n2491) );
  NANDN U2720 ( .A(n8626), .B(y[203]), .Z(n2502) );
  AND U2721 ( .A(y[216]), .B(x[68]), .Z(n2501) );
  NANDN U2722 ( .A(n8864), .B(y[198]), .Z(n2500) );
  XOR U2723 ( .A(n2501), .B(n2500), .Z(n2503) );
  XNOR U2724 ( .A(n2502), .B(n2503), .Z(n2490) );
  XNOR U2725 ( .A(n2491), .B(n2490), .Z(n2402) );
  XNOR U2726 ( .A(n2401), .B(n2402), .Z(n2404) );
  OR U2727 ( .A(n2348), .B(n2347), .Z(n2352) );
  OR U2728 ( .A(n2350), .B(n2349), .Z(n2351) );
  AND U2729 ( .A(n2352), .B(n2351), .Z(n2521) );
  OR U2730 ( .A(n2354), .B(n2353), .Z(n2358) );
  OR U2731 ( .A(n2356), .B(n2355), .Z(n2357) );
  AND U2732 ( .A(n2358), .B(n2357), .Z(n2520) );
  OR U2733 ( .A(n2360), .B(n2359), .Z(n2364) );
  OR U2734 ( .A(n2362), .B(n2361), .Z(n2363) );
  AND U2735 ( .A(n2364), .B(n2363), .Z(n2519) );
  XNOR U2736 ( .A(n2520), .B(n2519), .Z(n2522) );
  XNOR U2737 ( .A(n2521), .B(n2522), .Z(n2403) );
  XNOR U2738 ( .A(n2404), .B(n2403), .Z(n2525) );
  XNOR U2739 ( .A(n2527), .B(n2528), .Z(n2537) );
  XNOR U2740 ( .A(n2538), .B(n2537), .Z(n2534) );
  XOR U2741 ( .A(n2533), .B(n2534), .Z(n2547) );
  OR U2742 ( .A(n2366), .B(n2365), .Z(n2370) );
  OR U2743 ( .A(n2368), .B(n2367), .Z(n2369) );
  AND U2744 ( .A(n2370), .B(n2369), .Z(n2548) );
  XOR U2745 ( .A(n2547), .B(n2548), .Z(n2550) );
  XNOR U2746 ( .A(n2549), .B(n2550), .Z(n2389) );
  OR U2747 ( .A(n2372), .B(n2371), .Z(n2376) );
  NANDN U2748 ( .A(n2374), .B(n2373), .Z(n2375) );
  AND U2749 ( .A(n2376), .B(n2375), .Z(n2390) );
  XOR U2750 ( .A(n2389), .B(n2390), .Z(n2392) );
  OR U2751 ( .A(n2378), .B(n2377), .Z(n2382) );
  OR U2752 ( .A(n2380), .B(n2379), .Z(n2381) );
  NAND U2753 ( .A(n2382), .B(n2381), .Z(n2391) );
  XOR U2754 ( .A(n2392), .B(n2391), .Z(n2386) );
  XNOR U2755 ( .A(n2385), .B(n2386), .Z(N61) );
  NANDN U2756 ( .A(n2384), .B(n2383), .Z(n2388) );
  NAND U2757 ( .A(n2386), .B(n2385), .Z(n2387) );
  NAND U2758 ( .A(n2388), .B(n2387), .Z(n2553) );
  NANDN U2759 ( .A(n2390), .B(n2389), .Z(n2394) );
  OR U2760 ( .A(n2392), .B(n2391), .Z(n2393) );
  AND U2761 ( .A(n2394), .B(n2393), .Z(n2554) );
  XNOR U2762 ( .A(n2553), .B(n2554), .Z(n2555) );
  NANDN U2763 ( .A(n2396), .B(n2395), .Z(n2400) );
  OR U2764 ( .A(n2398), .B(n2397), .Z(n2399) );
  AND U2765 ( .A(n2400), .B(n2399), .Z(n2722) );
  OR U2766 ( .A(n2402), .B(n2401), .Z(n2406) );
  OR U2767 ( .A(n2404), .B(n2403), .Z(n2405) );
  NAND U2768 ( .A(n2406), .B(n2405), .Z(n2733) );
  OR U2769 ( .A(n2408), .B(n2407), .Z(n2412) );
  NANDN U2770 ( .A(n2410), .B(n2409), .Z(n2411) );
  NAND U2771 ( .A(n2412), .B(n2411), .Z(n2572) );
  OR U2772 ( .A(n2414), .B(n2413), .Z(n2418) );
  NAND U2773 ( .A(n2416), .B(n2415), .Z(n2417) );
  AND U2774 ( .A(n2418), .B(n2417), .Z(n2569) );
  OR U2775 ( .A(n2420), .B(n2419), .Z(n2424) );
  OR U2776 ( .A(n2422), .B(n2421), .Z(n2423) );
  NAND U2777 ( .A(n2424), .B(n2423), .Z(n2570) );
  XNOR U2778 ( .A(n2569), .B(n2570), .Z(n2571) );
  XOR U2779 ( .A(n2572), .B(n2571), .Z(n2732) );
  XNOR U2780 ( .A(n2733), .B(n2732), .Z(n2735) );
  OR U2781 ( .A(n2426), .B(n2425), .Z(n2430) );
  NANDN U2782 ( .A(n2428), .B(n2427), .Z(n2429) );
  AND U2783 ( .A(n2430), .B(n2429), .Z(n2734) );
  XOR U2784 ( .A(n2735), .B(n2734), .Z(n2720) );
  OR U2785 ( .A(n2432), .B(n2431), .Z(n2436) );
  OR U2786 ( .A(n2434), .B(n2433), .Z(n2435) );
  AND U2787 ( .A(n2436), .B(n2435), .Z(n2721) );
  XNOR U2788 ( .A(n2720), .B(n2721), .Z(n2723) );
  XOR U2789 ( .A(n2722), .B(n2723), .Z(n2728) );
  OR U2790 ( .A(n2438), .B(n2437), .Z(n2442) );
  OR U2791 ( .A(n2440), .B(n2439), .Z(n2441) );
  AND U2792 ( .A(n2442), .B(n2441), .Z(n2575) );
  NANDN U2793 ( .A(n2444), .B(n2443), .Z(n2448) );
  OR U2794 ( .A(n2446), .B(n2445), .Z(n2447) );
  NAND U2795 ( .A(n2448), .B(n2447), .Z(n2576) );
  XNOR U2796 ( .A(n2575), .B(n2576), .Z(n2577) );
  ANDN U2797 ( .B(x[73]), .A(n2449), .Z(n2696) );
  IV U2798 ( .A(n2696), .Z(n2818) );
  AND U2799 ( .A(y[216]), .B(x[69]), .Z(n2587) );
  AND U2800 ( .A(y[211]), .B(x[74]), .Z(n2588) );
  XNOR U2801 ( .A(n2587), .B(n2588), .Z(n2590) );
  AND U2802 ( .A(y[217]), .B(x[68]), .Z(n2589) );
  XNOR U2803 ( .A(n2590), .B(n2589), .Z(n2697) );
  XOR U2804 ( .A(n2818), .B(n2697), .Z(n2699) );
  AND U2805 ( .A(y[213]), .B(x[72]), .Z(n2619) );
  AND U2806 ( .A(y[214]), .B(x[71]), .Z(n2620) );
  XNOR U2807 ( .A(n2619), .B(n2620), .Z(n2622) );
  AND U2808 ( .A(x[70]), .B(y[215]), .Z(n2621) );
  XNOR U2809 ( .A(n2622), .B(n2621), .Z(n2698) );
  XNOR U2810 ( .A(n2699), .B(n2698), .Z(n2578) );
  OR U2811 ( .A(n2451), .B(n2450), .Z(n2455) );
  OR U2812 ( .A(n2453), .B(n2452), .Z(n2454) );
  AND U2813 ( .A(n2455), .B(n2454), .Z(n2654) );
  OR U2814 ( .A(n2457), .B(n2456), .Z(n2461) );
  OR U2815 ( .A(n2459), .B(n2458), .Z(n2460) );
  NAND U2816 ( .A(n2461), .B(n2460), .Z(n2687) );
  AND U2817 ( .A(x[78]), .B(y[207]), .Z(n2635) );
  AND U2818 ( .A(y[196]), .B(x[89]), .Z(n2633) );
  AND U2819 ( .A(y[195]), .B(x[90]), .Z(n2634) );
  XNOR U2820 ( .A(n2633), .B(n2634), .Z(n2636) );
  XOR U2821 ( .A(n2635), .B(n2636), .Z(n2685) );
  AND U2822 ( .A(y[221]), .B(x[64]), .Z(n2710) );
  AND U2823 ( .A(x[92]), .B(y[193]), .Z(n2650) );
  XOR U2824 ( .A(o[29]), .B(n2650), .Z(n2708) );
  AND U2825 ( .A(x[93]), .B(y[192]), .Z(n2709) );
  XNOR U2826 ( .A(n2708), .B(n2709), .Z(n2711) );
  XNOR U2827 ( .A(n2710), .B(n2711), .Z(n2684) );
  XOR U2828 ( .A(n2685), .B(n2684), .Z(n2686) );
  XOR U2829 ( .A(n2687), .B(n2686), .Z(n2663) );
  OR U2830 ( .A(n2463), .B(n2462), .Z(n2467) );
  OR U2831 ( .A(n2465), .B(n2464), .Z(n2466) );
  AND U2832 ( .A(n2467), .B(n2466), .Z(n2627) );
  AND U2833 ( .A(y[205]), .B(x[80]), .Z(n2599) );
  NANDN U2834 ( .A(n2857), .B(o[28]), .Z(n2468) );
  XOR U2835 ( .A(n2602), .B(n2468), .Z(n2469) );
  NAND U2836 ( .A(x[91]), .B(n2469), .Z(n2600) );
  XNOR U2837 ( .A(n2599), .B(n2600), .Z(n2628) );
  XOR U2838 ( .A(n2627), .B(n2628), .Z(n2630) );
  NANDN U2839 ( .A(n47), .B(y[219]), .Z(n2595) );
  AND U2840 ( .A(y[203]), .B(x[82]), .Z(n2594) );
  NANDN U2841 ( .A(n8824), .B(y[202]), .Z(n2593) );
  XOR U2842 ( .A(n2594), .B(n2593), .Z(n2596) );
  XNOR U2843 ( .A(n2595), .B(n2596), .Z(n2629) );
  XNOR U2844 ( .A(n2630), .B(n2629), .Z(n2661) );
  OR U2845 ( .A(n2471), .B(n2470), .Z(n2475) );
  OR U2846 ( .A(n2473), .B(n2472), .Z(n2474) );
  AND U2847 ( .A(n2475), .B(n2474), .Z(n2681) );
  OR U2848 ( .A(n2477), .B(n2476), .Z(n2481) );
  OR U2849 ( .A(n2479), .B(n2478), .Z(n2480) );
  AND U2850 ( .A(n2481), .B(n2480), .Z(n2678) );
  OR U2851 ( .A(n2483), .B(n2482), .Z(n2487) );
  OR U2852 ( .A(n2485), .B(n2484), .Z(n2486) );
  AND U2853 ( .A(n2487), .B(n2486), .Z(n2581) );
  AND U2854 ( .A(x[75]), .B(y[210]), .Z(n2607) );
  AND U2855 ( .A(y[204]), .B(x[81]), .Z(n2608) );
  XNOR U2856 ( .A(n2607), .B(n2608), .Z(n2610) );
  AND U2857 ( .A(y[218]), .B(x[67]), .Z(n2609) );
  XNOR U2858 ( .A(n2610), .B(n2609), .Z(n2582) );
  XOR U2859 ( .A(n2581), .B(n2582), .Z(n2584) );
  ANDN U2860 ( .B(y[198]), .A(n8656), .Z(n2613) );
  IV U2861 ( .A(n2613), .Z(n2968) );
  AND U2862 ( .A(x[88]), .B(y[197]), .Z(n2614) );
  XOR U2863 ( .A(n2968), .B(n2614), .Z(n2616) );
  AND U2864 ( .A(y[208]), .B(x[77]), .Z(n2615) );
  XOR U2865 ( .A(n2616), .B(n2615), .Z(n2583) );
  XNOR U2866 ( .A(n2584), .B(n2583), .Z(n2679) );
  XNOR U2867 ( .A(n2678), .B(n2679), .Z(n2680) );
  XOR U2868 ( .A(n2661), .B(n2660), .Z(n2662) );
  XNOR U2869 ( .A(n2663), .B(n2662), .Z(n2655) );
  XNOR U2870 ( .A(n2654), .B(n2655), .Z(n2656) );
  OR U2871 ( .A(n2489), .B(n2488), .Z(n2493) );
  NAND U2872 ( .A(n2491), .B(n2490), .Z(n2492) );
  AND U2873 ( .A(n2493), .B(n2492), .Z(n2666) );
  OR U2874 ( .A(n2495), .B(n2494), .Z(n2499) );
  OR U2875 ( .A(n2497), .B(n2496), .Z(n2498) );
  AND U2876 ( .A(n2499), .B(n2498), .Z(n2714) );
  NANDN U2877 ( .A(n2501), .B(n2500), .Z(n2505) );
  NANDN U2878 ( .A(n2503), .B(n2502), .Z(n2504) );
  AND U2879 ( .A(n2505), .B(n2504), .Z(n2690) );
  ANDN U2880 ( .B(y[209]), .A(n57), .Z(n2641) );
  IV U2881 ( .A(n2641), .Z(n2924) );
  AND U2882 ( .A(x[86]), .B(y[199]), .Z(n2639) );
  AND U2883 ( .A(y[220]), .B(x[65]), .Z(n2640) );
  XNOR U2884 ( .A(n2639), .B(n2640), .Z(n2642) );
  XOR U2885 ( .A(n2924), .B(n2642), .Z(n2675) );
  OR U2886 ( .A(n2507), .B(n2506), .Z(n2511) );
  OR U2887 ( .A(n2509), .B(n2508), .Z(n2510) );
  AND U2888 ( .A(n2511), .B(n2510), .Z(n2672) );
  NANDN U2889 ( .A(n60), .B(y[206]), .Z(n2646) );
  ANDN U2890 ( .B(x[85]), .A(n2512), .Z(n2838) );
  NANDN U2891 ( .A(n8885), .B(y[201]), .Z(n2645) );
  XOR U2892 ( .A(n2838), .B(n2645), .Z(n2647) );
  XNOR U2893 ( .A(n2672), .B(n2673), .Z(n2674) );
  XNOR U2894 ( .A(n2675), .B(n2674), .Z(n2691) );
  XNOR U2895 ( .A(n2690), .B(n2691), .Z(n2692) );
  OR U2896 ( .A(n2514), .B(n2513), .Z(n2518) );
  OR U2897 ( .A(n2516), .B(n2515), .Z(n2517) );
  AND U2898 ( .A(n2518), .B(n2517), .Z(n2693) );
  XNOR U2899 ( .A(n2714), .B(n2715), .Z(n2717) );
  OR U2900 ( .A(n2520), .B(n2519), .Z(n2524) );
  OR U2901 ( .A(n2522), .B(n2521), .Z(n2523) );
  AND U2902 ( .A(n2524), .B(n2523), .Z(n2716) );
  XNOR U2903 ( .A(n2717), .B(n2716), .Z(n2667) );
  XNOR U2904 ( .A(n2666), .B(n2667), .Z(n2669) );
  XOR U2905 ( .A(n2668), .B(n2669), .Z(n2726) );
  OR U2906 ( .A(n2526), .B(n2525), .Z(n2530) );
  OR U2907 ( .A(n2528), .B(n2527), .Z(n2529) );
  NAND U2908 ( .A(n2530), .B(n2529), .Z(n2727) );
  XOR U2909 ( .A(n2726), .B(n2727), .Z(n2729) );
  XNOR U2910 ( .A(n2728), .B(n2729), .Z(n2567) );
  NANDN U2911 ( .A(n2536), .B(n2535), .Z(n2540) );
  OR U2912 ( .A(n2538), .B(n2537), .Z(n2539) );
  AND U2913 ( .A(n2540), .B(n2539), .Z(n2566) );
  XNOR U2914 ( .A(n2565), .B(n2566), .Z(n2568) );
  XNOR U2915 ( .A(n2567), .B(n2568), .Z(n2562) );
  OR U2916 ( .A(n2542), .B(n2541), .Z(n2546) );
  NANDN U2917 ( .A(n2544), .B(n2543), .Z(n2545) );
  AND U2918 ( .A(n2546), .B(n2545), .Z(n2559) );
  NANDN U2919 ( .A(n2548), .B(n2547), .Z(n2552) );
  OR U2920 ( .A(n2550), .B(n2549), .Z(n2551) );
  NAND U2921 ( .A(n2552), .B(n2551), .Z(n2560) );
  XNOR U2922 ( .A(n2559), .B(n2560), .Z(n2561) );
  XOR U2923 ( .A(n2562), .B(n2561), .Z(n2556) );
  XNOR U2924 ( .A(n2555), .B(n2556), .Z(N62) );
  NANDN U2925 ( .A(n2554), .B(n2553), .Z(n2558) );
  NAND U2926 ( .A(n2556), .B(n2555), .Z(n2557) );
  AND U2927 ( .A(n2558), .B(n2557), .Z(n2740) );
  OR U2928 ( .A(n2560), .B(n2559), .Z(n2564) );
  OR U2929 ( .A(n2562), .B(n2561), .Z(n2563) );
  AND U2930 ( .A(n2564), .B(n2563), .Z(n2741) );
  XNOR U2931 ( .A(n2740), .B(n2741), .Z(n2739) );
  OR U2932 ( .A(n2570), .B(n2569), .Z(n2574) );
  OR U2933 ( .A(n2572), .B(n2571), .Z(n2573) );
  NAND U2934 ( .A(n2574), .B(n2573), .Z(n2747) );
  OR U2935 ( .A(n2576), .B(n2575), .Z(n2580) );
  OR U2936 ( .A(n2578), .B(n2577), .Z(n2579) );
  AND U2937 ( .A(n2580), .B(n2579), .Z(n3002) );
  OR U2938 ( .A(n2582), .B(n2581), .Z(n2586) );
  NAND U2939 ( .A(n2584), .B(n2583), .Z(n2585) );
  AND U2940 ( .A(n2586), .B(n2585), .Z(n3004) );
  OR U2941 ( .A(n2588), .B(n2587), .Z(n2592) );
  OR U2942 ( .A(n2590), .B(n2589), .Z(n2591) );
  AND U2943 ( .A(n2592), .B(n2591), .Z(n2783) );
  NANDN U2944 ( .A(n51), .B(y[216]), .Z(n2973) );
  NANDN U2945 ( .A(n50), .B(y[217]), .Z(n2975) );
  NANDN U2946 ( .A(n8824), .B(y[203]), .Z(n2974) );
  XNOR U2947 ( .A(n2975), .B(n2974), .Z(n2972) );
  XNOR U2948 ( .A(n2973), .B(n2972), .Z(n2870) );
  NANDN U2949 ( .A(n2594), .B(n2593), .Z(n2598) );
  NANDN U2950 ( .A(n2596), .B(n2595), .Z(n2597) );
  AND U2951 ( .A(n2598), .B(n2597), .Z(n2872) );
  NANDN U2952 ( .A(n49), .B(y[218]), .Z(n2842) );
  NANDN U2953 ( .A(n48), .B(y[219]), .Z(n2844) );
  ANDN U2954 ( .B(x[82]), .A(n2905), .Z(n2843) );
  XNOR U2955 ( .A(n2844), .B(n2843), .Z(n2841) );
  XNOR U2956 ( .A(n2842), .B(n2841), .Z(n2873) );
  XOR U2957 ( .A(n2872), .B(n2873), .Z(n2871) );
  XNOR U2958 ( .A(n2870), .B(n2871), .Z(n2782) );
  XNOR U2959 ( .A(n2783), .B(n2782), .Z(n2785) );
  OR U2960 ( .A(n2600), .B(n2599), .Z(n2606) );
  NAND U2961 ( .A(o[28]), .B(n2601), .Z(n2604) );
  NANDN U2962 ( .A(n2602), .B(x[91]), .Z(n2603) );
  AND U2963 ( .A(n2604), .B(n2603), .Z(n2605) );
  ANDN U2964 ( .B(n2606), .A(n2605), .Z(n2784) );
  XNOR U2965 ( .A(n3004), .B(n3005), .Z(n3003) );
  XNOR U2966 ( .A(n3002), .B(n3003), .Z(n3027) );
  OR U2967 ( .A(n2608), .B(n2607), .Z(n2612) );
  OR U2968 ( .A(n2610), .B(n2609), .Z(n2611) );
  NAND U2969 ( .A(n2612), .B(n2611), .Z(n2791) );
  NANDN U2970 ( .A(n2906), .B(x[84]), .Z(n2961) );
  ANDN U2971 ( .B(y[208]), .A(n59), .Z(n2960) );
  XOR U2972 ( .A(n2961), .B(n2960), .Z(n2959) );
  ANDN U2973 ( .B(y[214]), .A(n53), .Z(n2958) );
  XOR U2974 ( .A(n2959), .B(n2958), .Z(n2793) );
  NANDN U2975 ( .A(n2902), .B(x[94]), .Z(n2824) );
  NANDN U2976 ( .A(n2857), .B(x[93]), .Z(n2877) );
  XNOR U2977 ( .A(o[30]), .B(n2877), .Z(n2823) );
  XOR U2978 ( .A(n2824), .B(n2823), .Z(n2822) );
  ANDN U2979 ( .B(y[222]), .A(n45), .Z(n2821) );
  XOR U2980 ( .A(n2822), .B(n2821), .Z(n2792) );
  XOR U2981 ( .A(n2791), .B(n2790), .Z(n2766) );
  OR U2982 ( .A(n2614), .B(n2613), .Z(n2618) );
  OR U2983 ( .A(n2616), .B(n2615), .Z(n2617) );
  AND U2984 ( .A(n2618), .B(n2617), .Z(n2767) );
  XNOR U2985 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2986 ( .A(n2620), .B(n2619), .Z(n2624) );
  OR U2987 ( .A(n2622), .B(n2621), .Z(n2623) );
  AND U2988 ( .A(n2624), .B(n2623), .Z(n2803) );
  NANDN U2989 ( .A(n8626), .B(y[205]), .Z(n2928) );
  NANDN U2990 ( .A(n47), .B(y[220]), .Z(n2930) );
  IV U2991 ( .A(x[90]), .Z(n8901) );
  NANDN U2992 ( .A(n8901), .B(y[196]), .Z(n2929) );
  XNOR U2993 ( .A(n2930), .B(n2929), .Z(n2927) );
  XNOR U2994 ( .A(n2928), .B(n2927), .Z(n2804) );
  NANDN U2995 ( .A(n2894), .B(x[71]), .Z(n2836) );
  ANDN U2996 ( .B(y[200]), .A(n8864), .Z(n2626) );
  ANDN U2997 ( .B(x[85]), .A(n2837), .Z(n2625) );
  XNOR U2998 ( .A(n2626), .B(n2625), .Z(n2835) );
  XOR U2999 ( .A(n2836), .B(n2835), .Z(n2805) );
  XNOR U3000 ( .A(n2804), .B(n2805), .Z(n2802) );
  XOR U3001 ( .A(n2803), .B(n2802), .Z(n2764) );
  XNOR U3002 ( .A(n2765), .B(n2764), .Z(n2759) );
  OR U3003 ( .A(n2628), .B(n2627), .Z(n2632) );
  NAND U3004 ( .A(n2630), .B(n2629), .Z(n2631) );
  NAND U3005 ( .A(n2632), .B(n2631), .Z(n2756) );
  OR U3006 ( .A(n2634), .B(n2633), .Z(n2638) );
  OR U3007 ( .A(n2636), .B(n2635), .Z(n2637) );
  AND U3008 ( .A(n2638), .B(n2637), .Z(n2776) );
  OR U3009 ( .A(n2640), .B(n2639), .Z(n2644) );
  OR U3010 ( .A(n2642), .B(n2641), .Z(n2643) );
  AND U3011 ( .A(n2644), .B(n2643), .Z(n2779) );
  NANDN U3012 ( .A(n2838), .B(n2645), .Z(n2649) );
  NANDN U3013 ( .A(n2647), .B(n2646), .Z(n2648) );
  AND U3014 ( .A(n2649), .B(n2648), .Z(n2796) );
  NAND U3015 ( .A(n2650), .B(o[29]), .Z(n2953) );
  IV U3016 ( .A(x[92]), .Z(n8654) );
  NANDN U3017 ( .A(n8654), .B(y[194]), .Z(n2955) );
  NANDN U3018 ( .A(n8890), .B(y[206]), .Z(n2954) );
  XNOR U3019 ( .A(n2955), .B(n2954), .Z(n2952) );
  XNOR U3020 ( .A(n2953), .B(n2952), .Z(n2798) );
  IV U3021 ( .A(x[89]), .Z(n8928) );
  NANDN U3022 ( .A(n8928), .B(y[197]), .Z(n2967) );
  ANDN U3023 ( .B(y[199]), .A(n8656), .Z(n2653) );
  NANDN U3024 ( .A(n2651), .B(x[88]), .Z(n2652) );
  XOR U3025 ( .A(n2653), .B(n2652), .Z(n2966) );
  XOR U3026 ( .A(n2967), .B(n2966), .Z(n2799) );
  XOR U3027 ( .A(n2798), .B(n2799), .Z(n2797) );
  XNOR U3028 ( .A(n2796), .B(n2797), .Z(n2778) );
  XOR U3029 ( .A(n2776), .B(n2777), .Z(n2757) );
  XNOR U3030 ( .A(n2756), .B(n2757), .Z(n2758) );
  XNOR U3031 ( .A(n2759), .B(n2758), .Z(n3026) );
  XNOR U3032 ( .A(n3027), .B(n3026), .Z(n3025) );
  OR U3033 ( .A(n2655), .B(n2654), .Z(n2659) );
  OR U3034 ( .A(n2657), .B(n2656), .Z(n2658) );
  NAND U3035 ( .A(n2659), .B(n2658), .Z(n3024) );
  XOR U3036 ( .A(n3025), .B(n3024), .Z(n2746) );
  XNOR U3037 ( .A(n2747), .B(n2746), .Z(n2745) );
  OR U3038 ( .A(n2661), .B(n2660), .Z(n2665) );
  NANDN U3039 ( .A(n2663), .B(n2662), .Z(n2664) );
  NAND U3040 ( .A(n2665), .B(n2664), .Z(n2744) );
  XNOR U3041 ( .A(n2745), .B(n2744), .Z(n3020) );
  OR U3042 ( .A(n2667), .B(n2666), .Z(n2671) );
  NANDN U3043 ( .A(n2669), .B(n2668), .Z(n2670) );
  NAND U3044 ( .A(n2671), .B(n2670), .Z(n3021) );
  OR U3045 ( .A(n2673), .B(n2672), .Z(n2677) );
  OR U3046 ( .A(n2675), .B(n2674), .Z(n2676) );
  AND U3047 ( .A(n2677), .B(n2676), .Z(n2753) );
  OR U3048 ( .A(n2679), .B(n2678), .Z(n2683) );
  OR U3049 ( .A(n2681), .B(n2680), .Z(n2682) );
  AND U3050 ( .A(n2683), .B(n2682), .Z(n2752) );
  XOR U3051 ( .A(n2753), .B(n2752), .Z(n2750) );
  NANDN U3052 ( .A(n2685), .B(n2684), .Z(n2689) );
  OR U3053 ( .A(n2687), .B(n2686), .Z(n2688) );
  NAND U3054 ( .A(n2689), .B(n2688), .Z(n2751) );
  XNOR U3055 ( .A(n2750), .B(n2751), .Z(n2998) );
  OR U3056 ( .A(n2691), .B(n2690), .Z(n2695) );
  OR U3057 ( .A(n2693), .B(n2692), .Z(n2694) );
  NAND U3058 ( .A(n2695), .B(n2694), .Z(n2771) );
  OR U3059 ( .A(n2697), .B(n2696), .Z(n2701) );
  OR U3060 ( .A(n2699), .B(n2698), .Z(n2700) );
  NAND U3061 ( .A(n2701), .B(n2700), .Z(n2773) );
  NANDN U3062 ( .A(n43), .B(x[91]), .Z(n2832) );
  ANDN U3063 ( .B(y[221]), .A(n46), .Z(n2831) );
  XNOR U3064 ( .A(n2832), .B(n2831), .Z(n2829) );
  XOR U3065 ( .A(n2829), .B(n2830), .Z(n2810) );
  ANDN U3066 ( .B(x[77]), .A(n2851), .Z(n2704) );
  NANDN U3067 ( .A(n2702), .B(x[76]), .Z(n2703) );
  XOR U3068 ( .A(n2704), .B(n2703), .Z(n2922) );
  XNOR U3069 ( .A(n2922), .B(n2921), .Z(n2817) );
  ANDN U3070 ( .B(y[212]), .A(n55), .Z(n2707) );
  ANDN U3071 ( .B(x[73]), .A(n2705), .Z(n2706) );
  XNOR U3072 ( .A(n2707), .B(n2706), .Z(n2816) );
  XOR U3073 ( .A(n2817), .B(n2816), .Z(n2813) );
  OR U3074 ( .A(n2709), .B(n2708), .Z(n2713) );
  OR U3075 ( .A(n2711), .B(n2710), .Z(n2712) );
  AND U3076 ( .A(n2713), .B(n2712), .Z(n2812) );
  XNOR U3077 ( .A(n2813), .B(n2812), .Z(n2811) );
  XNOR U3078 ( .A(n2810), .B(n2811), .Z(n2772) );
  XNOR U3079 ( .A(n2773), .B(n2772), .Z(n2770) );
  XNOR U3080 ( .A(n2771), .B(n2770), .Z(n2999) );
  XNOR U3081 ( .A(n2998), .B(n2999), .Z(n2997) );
  OR U3082 ( .A(n2715), .B(n2714), .Z(n2719) );
  OR U3083 ( .A(n2717), .B(n2716), .Z(n2718) );
  NAND U3084 ( .A(n2719), .B(n2718), .Z(n2996) );
  XNOR U3085 ( .A(n2997), .B(n2996), .Z(n3018) );
  XOR U3086 ( .A(n3019), .B(n3018), .Z(n3038) );
  OR U3087 ( .A(n2721), .B(n2720), .Z(n2725) );
  OR U3088 ( .A(n2723), .B(n2722), .Z(n2724) );
  AND U3089 ( .A(n2725), .B(n2724), .Z(n3044) );
  NANDN U3090 ( .A(n2727), .B(n2726), .Z(n2731) );
  OR U3091 ( .A(n2729), .B(n2728), .Z(n2730) );
  NAND U3092 ( .A(n2731), .B(n2730), .Z(n3045) );
  XNOR U3093 ( .A(n3044), .B(n3045), .Z(n3042) );
  OR U3094 ( .A(n2733), .B(n2732), .Z(n2737) );
  OR U3095 ( .A(n2735), .B(n2734), .Z(n2736) );
  NAND U3096 ( .A(n2737), .B(n2736), .Z(n3043) );
  XNOR U3097 ( .A(n3038), .B(n3039), .Z(n3037) );
  XOR U3098 ( .A(n3036), .B(n3037), .Z(n2738) );
  XOR U3099 ( .A(n2739), .B(n2738), .Z(N63) );
  NANDN U3100 ( .A(n2739), .B(n2738), .Z(n2743) );
  OR U3101 ( .A(n2741), .B(n2740), .Z(n2742) );
  AND U3102 ( .A(n2743), .B(n2742), .Z(n3035) );
  OR U3103 ( .A(n2745), .B(n2744), .Z(n2749) );
  OR U3104 ( .A(n2747), .B(n2746), .Z(n2748) );
  AND U3105 ( .A(n2749), .B(n2748), .Z(n3017) );
  NANDN U3106 ( .A(n2751), .B(n2750), .Z(n2755) );
  NOR U3107 ( .A(n2753), .B(n2752), .Z(n2754) );
  ANDN U3108 ( .B(n2755), .A(n2754), .Z(n2763) );
  NOR U3109 ( .A(n2757), .B(n2756), .Z(n2761) );
  ANDN U3110 ( .B(n2759), .A(n2758), .Z(n2760) );
  OR U3111 ( .A(n2761), .B(n2760), .Z(n2762) );
  XNOR U3112 ( .A(n2763), .B(n2762), .Z(n3015) );
  OR U3113 ( .A(n2765), .B(n2764), .Z(n2769) );
  OR U3114 ( .A(n2767), .B(n2766), .Z(n2768) );
  AND U3115 ( .A(n2769), .B(n2768), .Z(n3013) );
  OR U3116 ( .A(n2771), .B(n2770), .Z(n2775) );
  OR U3117 ( .A(n2773), .B(n2772), .Z(n2774) );
  AND U3118 ( .A(n2775), .B(n2774), .Z(n2995) );
  OR U3119 ( .A(n2777), .B(n2776), .Z(n2781) );
  OR U3120 ( .A(n2779), .B(n2778), .Z(n2780) );
  AND U3121 ( .A(n2781), .B(n2780), .Z(n2789) );
  NOR U3122 ( .A(n2783), .B(n2782), .Z(n2787) );
  NOR U3123 ( .A(n2785), .B(n2784), .Z(n2786) );
  OR U3124 ( .A(n2787), .B(n2786), .Z(n2788) );
  XNOR U3125 ( .A(n2789), .B(n2788), .Z(n2993) );
  OR U3126 ( .A(n2791), .B(n2790), .Z(n2795) );
  OR U3127 ( .A(n2793), .B(n2792), .Z(n2794) );
  AND U3128 ( .A(n2795), .B(n2794), .Z(n2991) );
  OR U3129 ( .A(n2797), .B(n2796), .Z(n2801) );
  NANDN U3130 ( .A(n2799), .B(n2798), .Z(n2800) );
  AND U3131 ( .A(n2801), .B(n2800), .Z(n2809) );
  NANDN U3132 ( .A(n2803), .B(n2802), .Z(n2807) );
  NANDN U3133 ( .A(n2805), .B(n2804), .Z(n2806) );
  NAND U3134 ( .A(n2807), .B(n2806), .Z(n2808) );
  XNOR U3135 ( .A(n2809), .B(n2808), .Z(n2989) );
  NANDN U3136 ( .A(n2811), .B(n2810), .Z(n2815) );
  OR U3137 ( .A(n2813), .B(n2812), .Z(n2814) );
  AND U3138 ( .A(n2815), .B(n2814), .Z(n2987) );
  OR U3139 ( .A(n2817), .B(n2816), .Z(n2820) );
  NANDN U3140 ( .A(n55), .B(y[213]), .Z(n2943) );
  OR U3141 ( .A(n2943), .B(n2818), .Z(n2819) );
  AND U3142 ( .A(n2820), .B(n2819), .Z(n2828) );
  NANDN U3143 ( .A(n2822), .B(n2821), .Z(n2826) );
  NANDN U3144 ( .A(n2824), .B(n2823), .Z(n2825) );
  NAND U3145 ( .A(n2826), .B(n2825), .Z(n2827) );
  XNOR U3146 ( .A(n2828), .B(n2827), .Z(n2985) );
  NANDN U3147 ( .A(n2830), .B(n2829), .Z(n2834) );
  NANDN U3148 ( .A(n2832), .B(n2831), .Z(n2833) );
  AND U3149 ( .A(n2834), .B(n2833), .Z(n2869) );
  OR U3150 ( .A(n2836), .B(n2835), .Z(n2840) );
  NANDN U3151 ( .A(n2837), .B(x[86]), .Z(n2879) );
  NANDN U3152 ( .A(n2879), .B(n2838), .Z(n2839) );
  AND U3153 ( .A(n2840), .B(n2839), .Z(n2848) );
  NANDN U3154 ( .A(n2842), .B(n2841), .Z(n2846) );
  NANDN U3155 ( .A(n2844), .B(n2843), .Z(n2845) );
  NAND U3156 ( .A(n2846), .B(n2845), .Z(n2847) );
  XNOR U3157 ( .A(n2848), .B(n2847), .Z(n2867) );
  ANDN U3158 ( .B(y[203]), .A(n8885), .Z(n2850) );
  NANDN U3159 ( .A(n54), .B(y[214]), .Z(n2849) );
  XNOR U3160 ( .A(n2850), .B(n2849), .Z(n2856) );
  ANDN U3161 ( .B(x[78]), .A(n2851), .Z(n2854) );
  NANDN U3162 ( .A(n2852), .B(x[80]), .Z(n2853) );
  XNOR U3163 ( .A(n2854), .B(n2853), .Z(n2855) );
  XOR U3164 ( .A(n2856), .B(n2855), .Z(n2865) );
  IV U3165 ( .A(x[93]), .Z(n8893) );
  ANDN U3166 ( .B(y[194]), .A(n8893), .Z(n2859) );
  NANDN U3167 ( .A(n2857), .B(x[94]), .Z(n2858) );
  XNOR U3168 ( .A(n2859), .B(n2858), .Z(n2863) );
  ANDN U3169 ( .B(y[220]), .A(n48), .Z(n2861) );
  NANDN U3170 ( .A(n61), .B(y[205]), .Z(n2860) );
  XNOR U3171 ( .A(n2861), .B(n2860), .Z(n2862) );
  XNOR U3172 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3173 ( .A(n2865), .B(n2864), .Z(n2866) );
  XNOR U3174 ( .A(n2867), .B(n2866), .Z(n2868) );
  XNOR U3175 ( .A(n2869), .B(n2868), .Z(n2951) );
  NAND U3176 ( .A(n2871), .B(n2870), .Z(n2875) );
  OR U3177 ( .A(n2873), .B(n2872), .Z(n2874) );
  AND U3178 ( .A(n2875), .B(n2874), .Z(n2949) );
  ANDN U3179 ( .B(x[81]), .A(n2876), .Z(n2885) );
  ANDN U3180 ( .B(o[30]), .A(n2877), .Z(n2883) );
  XOR U3181 ( .A(n2923), .B(o[31]), .Z(n2881) );
  NANDN U3182 ( .A(n2878), .B(x[88]), .Z(n2969) );
  XNOR U3183 ( .A(n2879), .B(n2969), .Z(n2880) );
  XNOR U3184 ( .A(n2881), .B(n2880), .Z(n2882) );
  XNOR U3185 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3186 ( .A(n2885), .B(n2884), .Z(n2893) );
  ANDN U3187 ( .B(y[216]), .A(n52), .Z(n2887) );
  NANDN U3188 ( .A(n51), .B(y[217]), .Z(n2886) );
  XNOR U3189 ( .A(n2887), .B(n2886), .Z(n2891) );
  ANDN U3190 ( .B(y[221]), .A(n47), .Z(n2889) );
  NANDN U3191 ( .A(n50), .B(y[218]), .Z(n2888) );
  XNOR U3192 ( .A(n2889), .B(n2888), .Z(n2890) );
  XNOR U3193 ( .A(n2891), .B(n2890), .Z(n2892) );
  XNOR U3194 ( .A(n2893), .B(n2892), .Z(n2947) );
  ANDN U3195 ( .B(y[198]), .A(n8928), .Z(n2896) );
  NANDN U3196 ( .A(n2894), .B(x[72]), .Z(n2895) );
  XNOR U3197 ( .A(n2896), .B(n2895), .Z(n2901) );
  ANDN U3198 ( .B(y[200]), .A(n8656), .Z(n2899) );
  NANDN U3199 ( .A(n2897), .B(x[91]), .Z(n2898) );
  XNOR U3200 ( .A(n2899), .B(n2898), .Z(n2900) );
  XOR U3201 ( .A(n2901), .B(n2900), .Z(n2912) );
  ANDN U3202 ( .B(y[219]), .A(n49), .Z(n2904) );
  NANDN U3203 ( .A(n2902), .B(x[95]), .Z(n2903) );
  XNOR U3204 ( .A(n2904), .B(n2903), .Z(n2910) );
  ANDN U3205 ( .B(x[83]), .A(n2905), .Z(n2908) );
  NANDN U3206 ( .A(n2906), .B(x[85]), .Z(n2907) );
  XNOR U3207 ( .A(n2908), .B(n2907), .Z(n2909) );
  XNOR U3208 ( .A(n2910), .B(n2909), .Z(n2911) );
  XNOR U3209 ( .A(n2912), .B(n2911), .Z(n2920) );
  ANDN U3210 ( .B(y[222]), .A(n46), .Z(n2914) );
  NANDN U3211 ( .A(n8654), .B(y[195]), .Z(n2913) );
  XNOR U3212 ( .A(n2914), .B(n2913), .Z(n2918) );
  ANDN U3213 ( .B(y[208]), .A(n60), .Z(n2916) );
  NANDN U3214 ( .A(n45), .B(y[223]), .Z(n2915) );
  XNOR U3215 ( .A(n2916), .B(n2915), .Z(n2917) );
  XNOR U3216 ( .A(n2918), .B(n2917), .Z(n2919) );
  XNOR U3217 ( .A(n2920), .B(n2919), .Z(n2936) );
  OR U3218 ( .A(n2922), .B(n2921), .Z(n2926) );
  NANDN U3219 ( .A(n2924), .B(n2923), .Z(n2925) );
  AND U3220 ( .A(n2926), .B(n2925), .Z(n2934) );
  OR U3221 ( .A(n2928), .B(n2927), .Z(n2932) );
  OR U3222 ( .A(n2930), .B(n2929), .Z(n2931) );
  NAND U3223 ( .A(n2932), .B(n2931), .Z(n2933) );
  XNOR U3224 ( .A(n2934), .B(n2933), .Z(n2935) );
  XOR U3225 ( .A(n2936), .B(n2935), .Z(n2945) );
  ANDN U3226 ( .B(y[212]), .A(n56), .Z(n2939) );
  NANDN U3227 ( .A(n2937), .B(x[76]), .Z(n2938) );
  XNOR U3228 ( .A(n2939), .B(n2938), .Z(n2941) );
  NANDN U3229 ( .A(n8901), .B(y[197]), .Z(n2940) );
  XNOR U3230 ( .A(n2941), .B(n2940), .Z(n2942) );
  XOR U3231 ( .A(n2943), .B(n2942), .Z(n2944) );
  XNOR U3232 ( .A(n2945), .B(n2944), .Z(n2946) );
  XNOR U3233 ( .A(n2947), .B(n2946), .Z(n2948) );
  XNOR U3234 ( .A(n2949), .B(n2948), .Z(n2950) );
  XOR U3235 ( .A(n2951), .B(n2950), .Z(n2983) );
  OR U3236 ( .A(n2953), .B(n2952), .Z(n2957) );
  OR U3237 ( .A(n2955), .B(n2954), .Z(n2956) );
  AND U3238 ( .A(n2957), .B(n2956), .Z(n2965) );
  NANDN U3239 ( .A(n2959), .B(n2958), .Z(n2963) );
  NANDN U3240 ( .A(n2961), .B(n2960), .Z(n2962) );
  NAND U3241 ( .A(n2963), .B(n2962), .Z(n2964) );
  XNOR U3242 ( .A(n2965), .B(n2964), .Z(n2981) );
  OR U3243 ( .A(n2967), .B(n2966), .Z(n2971) );
  OR U3244 ( .A(n2969), .B(n2968), .Z(n2970) );
  AND U3245 ( .A(n2971), .B(n2970), .Z(n2979) );
  OR U3246 ( .A(n2973), .B(n2972), .Z(n2977) );
  OR U3247 ( .A(n2975), .B(n2974), .Z(n2976) );
  NAND U3248 ( .A(n2977), .B(n2976), .Z(n2978) );
  XNOR U3249 ( .A(n2979), .B(n2978), .Z(n2980) );
  XNOR U3250 ( .A(n2981), .B(n2980), .Z(n2982) );
  XNOR U3251 ( .A(n2983), .B(n2982), .Z(n2984) );
  XNOR U3252 ( .A(n2985), .B(n2984), .Z(n2986) );
  XNOR U3253 ( .A(n2987), .B(n2986), .Z(n2988) );
  XNOR U3254 ( .A(n2989), .B(n2988), .Z(n2990) );
  XNOR U3255 ( .A(n2991), .B(n2990), .Z(n2992) );
  XNOR U3256 ( .A(n2993), .B(n2992), .Z(n2994) );
  XNOR U3257 ( .A(n2995), .B(n2994), .Z(n3011) );
  OR U3258 ( .A(n2997), .B(n2996), .Z(n3001) );
  OR U3259 ( .A(n2999), .B(n2998), .Z(n3000) );
  AND U3260 ( .A(n3001), .B(n3000), .Z(n3009) );
  OR U3261 ( .A(n3003), .B(n3002), .Z(n3007) );
  OR U3262 ( .A(n3005), .B(n3004), .Z(n3006) );
  NAND U3263 ( .A(n3007), .B(n3006), .Z(n3008) );
  XNOR U3264 ( .A(n3009), .B(n3008), .Z(n3010) );
  XNOR U3265 ( .A(n3011), .B(n3010), .Z(n3012) );
  XNOR U3266 ( .A(n3013), .B(n3012), .Z(n3014) );
  XNOR U3267 ( .A(n3015), .B(n3014), .Z(n3016) );
  XNOR U3268 ( .A(n3017), .B(n3016), .Z(n3033) );
  OR U3269 ( .A(n3019), .B(n3018), .Z(n3023) );
  OR U3270 ( .A(n3021), .B(n3020), .Z(n3022) );
  AND U3271 ( .A(n3023), .B(n3022), .Z(n3031) );
  OR U3272 ( .A(n3025), .B(n3024), .Z(n3029) );
  OR U3273 ( .A(n3027), .B(n3026), .Z(n3028) );
  NAND U3274 ( .A(n3029), .B(n3028), .Z(n3030) );
  XNOR U3275 ( .A(n3031), .B(n3030), .Z(n3032) );
  XNOR U3276 ( .A(n3033), .B(n3032), .Z(n3034) );
  XNOR U3277 ( .A(n3035), .B(n3034), .Z(n3051) );
  OR U3278 ( .A(n3037), .B(n3036), .Z(n3041) );
  OR U3279 ( .A(n3039), .B(n3038), .Z(n3040) );
  AND U3280 ( .A(n3041), .B(n3040), .Z(n3049) );
  OR U3281 ( .A(n3043), .B(n3042), .Z(n3047) );
  OR U3282 ( .A(n3045), .B(n3044), .Z(n3046) );
  NAND U3283 ( .A(n3047), .B(n3046), .Z(n3048) );
  XNOR U3284 ( .A(n3049), .B(n3048), .Z(n3050) );
  XNOR U3285 ( .A(n3051), .B(n3050), .Z(N64) );
  IV U3286 ( .A(y[224]), .Z(n5905) );
  ANDN U3287 ( .B(x[64]), .A(n5905), .Z(n3747) );
  XOR U3288 ( .A(n3747), .B(o[32]), .Z(N97) );
  ANDN U3289 ( .B(x[65]), .A(n5905), .Z(n3052) );
  NANDN U3290 ( .A(n45), .B(y[225]), .Z(n3058) );
  XNOR U3291 ( .A(n3058), .B(o[33]), .Z(n3053) );
  XOR U3292 ( .A(n3052), .B(n3053), .Z(n3054) );
  AND U3293 ( .A(o[32]), .B(n3747), .Z(n3055) );
  XOR U3294 ( .A(n3054), .B(n3055), .Z(N98) );
  OR U3295 ( .A(n3053), .B(n3052), .Z(n3057) );
  NANDN U3296 ( .A(n3055), .B(n3054), .Z(n3056) );
  NAND U3297 ( .A(n3057), .B(n3056), .Z(n3060) );
  NANDN U3298 ( .A(n45), .B(y[226]), .Z(n3071) );
  XOR U3299 ( .A(n3071), .B(o[34]), .Z(n3059) );
  XNOR U3300 ( .A(n3060), .B(n3059), .Z(n3062) );
  ANDN U3301 ( .B(o[33]), .A(n3058), .Z(n3065) );
  AND U3302 ( .A(y[224]), .B(x[66]), .Z(n3066) );
  XNOR U3303 ( .A(n3065), .B(n3066), .Z(n3068) );
  AND U3304 ( .A(y[225]), .B(x[65]), .Z(n3067) );
  XNOR U3305 ( .A(n3068), .B(n3067), .Z(n3061) );
  XNOR U3306 ( .A(n3062), .B(n3061), .Z(N99) );
  NAND U3307 ( .A(n3060), .B(n3059), .Z(n3064) );
  OR U3308 ( .A(n3062), .B(n3061), .Z(n3063) );
  NAND U3309 ( .A(n3064), .B(n3063), .Z(n3075) );
  OR U3310 ( .A(n3066), .B(n3065), .Z(n3070) );
  OR U3311 ( .A(n3068), .B(n3067), .Z(n3069) );
  AND U3312 ( .A(n3070), .B(n3069), .Z(n3076) );
  XNOR U3313 ( .A(n3075), .B(n3076), .Z(n3077) );
  NANDN U3314 ( .A(n47), .B(y[225]), .Z(n3083) );
  XNOR U3315 ( .A(n3083), .B(o[35]), .Z(n3081) );
  NANDN U3316 ( .A(n3071), .B(o[34]), .Z(n3087) );
  ANDN U3317 ( .B(x[67]), .A(n5905), .Z(n3073) );
  NANDN U3318 ( .A(n45), .B(y[227]), .Z(n3072) );
  XOR U3319 ( .A(n3073), .B(n3072), .Z(n3086) );
  XNOR U3320 ( .A(n3087), .B(n3086), .Z(n3082) );
  AND U3321 ( .A(y[226]), .B(x[65]), .Z(n3111) );
  XOR U3322 ( .A(n3082), .B(n3111), .Z(n3074) );
  XOR U3323 ( .A(n3081), .B(n3074), .Z(n3078) );
  XNOR U3324 ( .A(n3077), .B(n3078), .Z(N100) );
  NANDN U3325 ( .A(n3076), .B(n3075), .Z(n3080) );
  NAND U3326 ( .A(n3078), .B(n3077), .Z(n3079) );
  NAND U3327 ( .A(n3080), .B(n3079), .Z(n3092) );
  XNOR U3328 ( .A(n3092), .B(n3093), .Z(n3094) );
  NANDN U3329 ( .A(n3083), .B(o[35]), .Z(n3108) );
  ANDN U3330 ( .B(x[68]), .A(n5905), .Z(n3085) );
  ANDN U3331 ( .B(y[228]), .A(n45), .Z(n3084) );
  XNOR U3332 ( .A(n3085), .B(n3084), .Z(n3107) );
  XOR U3333 ( .A(n3108), .B(n3107), .Z(n3100) );
  AND U3334 ( .A(y[227]), .B(x[67]), .Z(n3159) );
  NAND U3335 ( .A(n3747), .B(n3159), .Z(n3089) );
  OR U3336 ( .A(n3087), .B(n3086), .Z(n3088) );
  AND U3337 ( .A(n3089), .B(n3088), .Z(n3098) );
  IV U3338 ( .A(y[227]), .Z(n5714) );
  ANDN U3339 ( .B(x[65]), .A(n5714), .Z(n3091) );
  NANDN U3340 ( .A(n47), .B(y[226]), .Z(n3090) );
  XOR U3341 ( .A(n3091), .B(n3090), .Z(n3113) );
  NANDN U3342 ( .A(n48), .B(y[225]), .Z(n3104) );
  XNOR U3343 ( .A(n3104), .B(o[36]), .Z(n3112) );
  XOR U3344 ( .A(n3113), .B(n3112), .Z(n3099) );
  XOR U3345 ( .A(n3100), .B(n3101), .Z(n3095) );
  XOR U3346 ( .A(n3094), .B(n3095), .Z(N101) );
  NANDN U3347 ( .A(n3093), .B(n3092), .Z(n3097) );
  NANDN U3348 ( .A(n3095), .B(n3094), .Z(n3096) );
  NAND U3349 ( .A(n3097), .B(n3096), .Z(n3116) );
  OR U3350 ( .A(n3099), .B(n3098), .Z(n3103) );
  NAND U3351 ( .A(n3101), .B(n3100), .Z(n3102) );
  NAND U3352 ( .A(n3103), .B(n3102), .Z(n3117) );
  XNOR U3353 ( .A(n3116), .B(n3117), .Z(n3118) );
  NANDN U3354 ( .A(n3104), .B(o[36]), .Z(n3135) );
  ANDN U3355 ( .B(x[69]), .A(n5905), .Z(n3106) );
  ANDN U3356 ( .B(y[229]), .A(n45), .Z(n3105) );
  XNOR U3357 ( .A(n3106), .B(n3105), .Z(n3134) );
  XOR U3358 ( .A(n3135), .B(n3134), .Z(n3130) );
  AND U3359 ( .A(y[227]), .B(x[66]), .Z(n3128) );
  AND U3360 ( .A(y[228]), .B(x[65]), .Z(n3143) );
  AND U3361 ( .A(y[225]), .B(x[68]), .Z(n3138) );
  XOR U3362 ( .A(o[37]), .B(n3138), .Z(n3141) );
  AND U3363 ( .A(y[226]), .B(x[67]), .Z(n3142) );
  XNOR U3364 ( .A(n3141), .B(n3142), .Z(n3144) );
  XNOR U3365 ( .A(n3143), .B(n3144), .Z(n3129) );
  XNOR U3366 ( .A(n3128), .B(n3129), .Z(n3131) );
  XNOR U3367 ( .A(n3130), .B(n3131), .Z(n3125) );
  AND U3368 ( .A(y[228]), .B(x[68]), .Z(n3223) );
  NAND U3369 ( .A(n3747), .B(n3223), .Z(n3110) );
  OR U3370 ( .A(n3108), .B(n3107), .Z(n3109) );
  NAND U3371 ( .A(n3110), .B(n3109), .Z(n3123) );
  NAND U3372 ( .A(n3111), .B(n3128), .Z(n3115) );
  NANDN U3373 ( .A(n3113), .B(n3112), .Z(n3114) );
  NAND U3374 ( .A(n3115), .B(n3114), .Z(n3122) );
  XNOR U3375 ( .A(n3123), .B(n3122), .Z(n3124) );
  XNOR U3376 ( .A(n3125), .B(n3124), .Z(n3119) );
  XOR U3377 ( .A(n3118), .B(n3119), .Z(N102) );
  NANDN U3378 ( .A(n3117), .B(n3116), .Z(n3121) );
  NANDN U3379 ( .A(n3119), .B(n3118), .Z(n3120) );
  NAND U3380 ( .A(n3121), .B(n3120), .Z(n3147) );
  OR U3381 ( .A(n3123), .B(n3122), .Z(n3127) );
  OR U3382 ( .A(n3125), .B(n3124), .Z(n3126) );
  AND U3383 ( .A(n3127), .B(n3126), .Z(n3148) );
  XNOR U3384 ( .A(n3147), .B(n3148), .Z(n3149) );
  OR U3385 ( .A(n3129), .B(n3128), .Z(n3133) );
  OR U3386 ( .A(n3131), .B(n3130), .Z(n3132) );
  AND U3387 ( .A(n3133), .B(n3132), .Z(n3153) );
  NANDN U3388 ( .A(n50), .B(y[229]), .Z(n3495) );
  NANDN U3389 ( .A(n3495), .B(n3747), .Z(n3137) );
  OR U3390 ( .A(n3135), .B(n3134), .Z(n3136) );
  NAND U3391 ( .A(n3137), .B(n3136), .Z(n3176) );
  NAND U3392 ( .A(n3138), .B(o[37]), .Z(n3166) );
  ANDN U3393 ( .B(x[70]), .A(n5905), .Z(n3140) );
  IV U3394 ( .A(y[230]), .Z(n5663) );
  ANDN U3395 ( .B(x[64]), .A(n5663), .Z(n3139) );
  XNOR U3396 ( .A(n3140), .B(n3139), .Z(n3165) );
  XOR U3397 ( .A(n3166), .B(n3165), .Z(n3175) );
  XNOR U3398 ( .A(n3176), .B(n3175), .Z(n3178) );
  ANDN U3399 ( .B(y[229]), .A(n46), .Z(n3435) );
  NANDN U3400 ( .A(n50), .B(y[225]), .Z(n3169) );
  XNOR U3401 ( .A(n3169), .B(o[38]), .Z(n3170) );
  XNOR U3402 ( .A(n3435), .B(n3170), .Z(n3172) );
  ANDN U3403 ( .B(y[226]), .A(n49), .Z(n3171) );
  XOR U3404 ( .A(n3172), .B(n3171), .Z(n3160) );
  ANDN U3405 ( .B(y[228]), .A(n47), .Z(n3477) );
  XNOR U3406 ( .A(n3159), .B(n3477), .Z(n3161) );
  XOR U3407 ( .A(n3160), .B(n3161), .Z(n3177) );
  XNOR U3408 ( .A(n3178), .B(n3177), .Z(n3154) );
  XNOR U3409 ( .A(n3153), .B(n3154), .Z(n3155) );
  OR U3410 ( .A(n3142), .B(n3141), .Z(n3146) );
  OR U3411 ( .A(n3144), .B(n3143), .Z(n3145) );
  AND U3412 ( .A(n3146), .B(n3145), .Z(n3156) );
  XOR U3413 ( .A(n3149), .B(n3150), .Z(N103) );
  NANDN U3414 ( .A(n3148), .B(n3147), .Z(n3152) );
  NANDN U3415 ( .A(n3150), .B(n3149), .Z(n3151) );
  NAND U3416 ( .A(n3152), .B(n3151), .Z(n3211) );
  OR U3417 ( .A(n3154), .B(n3153), .Z(n3158) );
  OR U3418 ( .A(n3156), .B(n3155), .Z(n3157) );
  AND U3419 ( .A(n3158), .B(n3157), .Z(n3212) );
  XNOR U3420 ( .A(n3211), .B(n3212), .Z(n3213) );
  OR U3421 ( .A(n3159), .B(n3477), .Z(n3163) );
  NANDN U3422 ( .A(n3161), .B(n3160), .Z(n3162) );
  NAND U3423 ( .A(n3163), .B(n3162), .Z(n3196) );
  ANDN U3424 ( .B(y[230]), .A(n51), .Z(n3164) );
  NAND U3425 ( .A(n3747), .B(n3164), .Z(n3168) );
  OR U3426 ( .A(n3166), .B(n3165), .Z(n3167) );
  AND U3427 ( .A(n3168), .B(n3167), .Z(n3194) );
  AND U3428 ( .A(y[226]), .B(x[69]), .Z(n3368) );
  ANDN U3429 ( .B(y[230]), .A(n46), .Z(n3572) );
  NANDN U3430 ( .A(n51), .B(y[225]), .Z(n3181) );
  XNOR U3431 ( .A(o[39]), .B(n3181), .Z(n3183) );
  XNOR U3432 ( .A(n3572), .B(n3183), .Z(n3184) );
  XNOR U3433 ( .A(n3368), .B(n3184), .Z(n3193) );
  XOR U3434 ( .A(n3194), .B(n3193), .Z(n3195) );
  XNOR U3435 ( .A(n3196), .B(n3195), .Z(n3217) );
  AND U3436 ( .A(y[229]), .B(x[66]), .Z(n3669) );
  AND U3437 ( .A(y[227]), .B(x[68]), .Z(n3354) );
  AND U3438 ( .A(y[228]), .B(x[67]), .Z(n3207) );
  XNOR U3439 ( .A(n3354), .B(n3207), .Z(n3208) );
  XOR U3440 ( .A(n3669), .B(n3208), .Z(n3187) );
  NANDN U3441 ( .A(n44), .B(x[64]), .Z(n3203) );
  ANDN U3442 ( .B(o[38]), .A(n3169), .Z(n3202) );
  NANDN U3443 ( .A(n5905), .B(x[71]), .Z(n3201) );
  XOR U3444 ( .A(n3202), .B(n3201), .Z(n3204) );
  XNOR U3445 ( .A(n3203), .B(n3204), .Z(n3188) );
  XNOR U3446 ( .A(n3187), .B(n3188), .Z(n3190) );
  NAND U3447 ( .A(n3435), .B(n3170), .Z(n3174) );
  NANDN U3448 ( .A(n3172), .B(n3171), .Z(n3173) );
  AND U3449 ( .A(n3174), .B(n3173), .Z(n3189) );
  XOR U3450 ( .A(n3190), .B(n3189), .Z(n3218) );
  XOR U3451 ( .A(n3217), .B(n3218), .Z(n3220) );
  OR U3452 ( .A(n3176), .B(n3175), .Z(n3180) );
  OR U3453 ( .A(n3178), .B(n3177), .Z(n3179) );
  AND U3454 ( .A(n3180), .B(n3179), .Z(n3219) );
  XOR U3455 ( .A(n3220), .B(n3219), .Z(n3214) );
  XNOR U3456 ( .A(n3213), .B(n3214), .Z(N104) );
  AND U3457 ( .A(y[226]), .B(x[70]), .Z(n3224) );
  XNOR U3458 ( .A(n3223), .B(n3224), .Z(n3226) );
  ANDN U3459 ( .B(x[66]), .A(n5663), .Z(n3225) );
  IV U3460 ( .A(n3225), .Z(n3763) );
  XOR U3461 ( .A(n3226), .B(n3763), .Z(n3229) );
  AND U3462 ( .A(y[229]), .B(x[67]), .Z(n4057) );
  XNOR U3463 ( .A(n3229), .B(n4057), .Z(n3231) );
  NANDN U3464 ( .A(n3181), .B(o[39]), .Z(n3248) );
  ANDN U3465 ( .B(y[231]), .A(n46), .Z(n3742) );
  ANDN U3466 ( .B(x[69]), .A(n5714), .Z(n3182) );
  XNOR U3467 ( .A(n3742), .B(n3182), .Z(n3247) );
  XOR U3468 ( .A(n3248), .B(n3247), .Z(n3230) );
  XNOR U3469 ( .A(n3231), .B(n3230), .Z(n3251) );
  NAND U3470 ( .A(n3572), .B(n3183), .Z(n3186) );
  NANDN U3471 ( .A(n3184), .B(n3368), .Z(n3185) );
  AND U3472 ( .A(n3186), .B(n3185), .Z(n3252) );
  XOR U3473 ( .A(n3251), .B(n3252), .Z(n3254) );
  OR U3474 ( .A(n3188), .B(n3187), .Z(n3192) );
  OR U3475 ( .A(n3190), .B(n3189), .Z(n3191) );
  AND U3476 ( .A(n3192), .B(n3191), .Z(n3253) );
  XOR U3477 ( .A(n3254), .B(n3253), .Z(n3269) );
  NANDN U3478 ( .A(n3194), .B(n3193), .Z(n3198) );
  OR U3479 ( .A(n3196), .B(n3195), .Z(n3197) );
  NAND U3480 ( .A(n3198), .B(n3197), .Z(n3270) );
  XNOR U3481 ( .A(n3269), .B(n3270), .Z(n3272) );
  ANDN U3482 ( .B(x[72]), .A(n5905), .Z(n3200) );
  NANDN U3483 ( .A(n45), .B(y[232]), .Z(n3199) );
  XOR U3484 ( .A(n3200), .B(n3199), .Z(n3236) );
  NANDN U3485 ( .A(n52), .B(y[225]), .Z(n3239) );
  XOR U3486 ( .A(n3239), .B(o[40]), .Z(n3235) );
  XNOR U3487 ( .A(n3236), .B(n3235), .Z(n3258) );
  NANDN U3488 ( .A(n3202), .B(n3201), .Z(n3206) );
  NANDN U3489 ( .A(n3204), .B(n3203), .Z(n3205) );
  NAND U3490 ( .A(n3206), .B(n3205), .Z(n3257) );
  XOR U3491 ( .A(n3258), .B(n3257), .Z(n3259) );
  OR U3492 ( .A(n3207), .B(n3354), .Z(n3210) );
  OR U3493 ( .A(n3208), .B(n3669), .Z(n3209) );
  NAND U3494 ( .A(n3210), .B(n3209), .Z(n3260) );
  XNOR U3495 ( .A(n3259), .B(n3260), .Z(n3271) );
  XNOR U3496 ( .A(n3272), .B(n3271), .Z(n3266) );
  NANDN U3497 ( .A(n3212), .B(n3211), .Z(n3216) );
  NAND U3498 ( .A(n3214), .B(n3213), .Z(n3215) );
  NAND U3499 ( .A(n3216), .B(n3215), .Z(n3263) );
  NANDN U3500 ( .A(n3218), .B(n3217), .Z(n3222) );
  OR U3501 ( .A(n3220), .B(n3219), .Z(n3221) );
  AND U3502 ( .A(n3222), .B(n3221), .Z(n3264) );
  XNOR U3503 ( .A(n3263), .B(n3264), .Z(n3265) );
  XOR U3504 ( .A(n3266), .B(n3265), .Z(N105) );
  OR U3505 ( .A(n3224), .B(n3223), .Z(n3228) );
  OR U3506 ( .A(n3226), .B(n3225), .Z(n3227) );
  NAND U3507 ( .A(n3228), .B(n3227), .Z(n3304) );
  OR U3508 ( .A(n3229), .B(n4057), .Z(n3233) );
  OR U3509 ( .A(n3231), .B(n3230), .Z(n3232) );
  NAND U3510 ( .A(n3233), .B(n3232), .Z(n3303) );
  XNOR U3511 ( .A(n3304), .B(n3303), .Z(n3305) );
  ANDN U3512 ( .B(y[232]), .A(n53), .Z(n3234) );
  NAND U3513 ( .A(n3747), .B(n3234), .Z(n3238) );
  OR U3514 ( .A(n3236), .B(n3235), .Z(n3237) );
  NAND U3515 ( .A(n3238), .B(n3237), .Z(n3290) );
  NANDN U3516 ( .A(n3239), .B(o[40]), .Z(n3310) );
  ANDN U3517 ( .B(y[226]), .A(n52), .Z(n3241) );
  NANDN U3518 ( .A(n50), .B(y[228]), .Z(n3240) );
  XNOR U3519 ( .A(n3241), .B(n3240), .Z(n3309) );
  XNOR U3520 ( .A(n3310), .B(n3309), .Z(n3288) );
  ANDN U3521 ( .B(x[73]), .A(n5905), .Z(n3243) );
  NANDN U3522 ( .A(n45), .B(y[233]), .Z(n3242) );
  XOR U3523 ( .A(n3243), .B(n3242), .Z(n3322) );
  NANDN U3524 ( .A(n53), .B(y[225]), .Z(n3316) );
  XOR U3525 ( .A(n3316), .B(o[41]), .Z(n3321) );
  XNOR U3526 ( .A(n3322), .B(n3321), .Z(n3287) );
  XOR U3527 ( .A(n3288), .B(n3287), .Z(n3289) );
  XNOR U3528 ( .A(n3290), .B(n3289), .Z(n3299) );
  ANDN U3529 ( .B(y[229]), .A(n49), .Z(n3754) );
  IV U3530 ( .A(y[232]), .Z(n5947) );
  ANDN U3531 ( .B(x[65]), .A(n5947), .Z(n3245) );
  NANDN U3532 ( .A(n51), .B(y[227]), .Z(n3244) );
  XNOR U3533 ( .A(n3245), .B(n3244), .Z(n3318) );
  XOR U3534 ( .A(n3754), .B(n3318), .Z(n3293) );
  AND U3535 ( .A(y[231]), .B(x[66]), .Z(n3962) );
  NANDN U3536 ( .A(n5663), .B(x[67]), .Z(n3642) );
  XOR U3537 ( .A(n3962), .B(n3642), .Z(n3294) );
  XNOR U3538 ( .A(n3293), .B(n3294), .Z(n3297) );
  NANDN U3539 ( .A(n46), .B(y[227]), .Z(n3317) );
  ANDN U3540 ( .B(y[231]), .A(n50), .Z(n3246) );
  NANDN U3541 ( .A(n3317), .B(n3246), .Z(n3250) );
  OR U3542 ( .A(n3248), .B(n3247), .Z(n3249) );
  AND U3543 ( .A(n3250), .B(n3249), .Z(n3298) );
  XOR U3544 ( .A(n3297), .B(n3298), .Z(n3300) );
  XOR U3545 ( .A(n3299), .B(n3300), .Z(n3306) );
  NANDN U3546 ( .A(n3252), .B(n3251), .Z(n3256) );
  OR U3547 ( .A(n3254), .B(n3253), .Z(n3255) );
  NAND U3548 ( .A(n3256), .B(n3255), .Z(n3282) );
  OR U3549 ( .A(n3258), .B(n3257), .Z(n3262) );
  NANDN U3550 ( .A(n3260), .B(n3259), .Z(n3261) );
  NAND U3551 ( .A(n3262), .B(n3261), .Z(n3281) );
  XOR U3552 ( .A(n3282), .B(n3281), .Z(n3284) );
  XNOR U3553 ( .A(n3283), .B(n3284), .Z(n3278) );
  NANDN U3554 ( .A(n3264), .B(n3263), .Z(n3268) );
  NANDN U3555 ( .A(n3266), .B(n3265), .Z(n3267) );
  NAND U3556 ( .A(n3268), .B(n3267), .Z(n3275) );
  OR U3557 ( .A(n3270), .B(n3269), .Z(n3274) );
  OR U3558 ( .A(n3272), .B(n3271), .Z(n3273) );
  AND U3559 ( .A(n3274), .B(n3273), .Z(n3276) );
  XNOR U3560 ( .A(n3275), .B(n3276), .Z(n3277) );
  XOR U3561 ( .A(n3278), .B(n3277), .Z(N106) );
  NANDN U3562 ( .A(n3276), .B(n3275), .Z(n3280) );
  NANDN U3563 ( .A(n3278), .B(n3277), .Z(n3279) );
  NAND U3564 ( .A(n3280), .B(n3279), .Z(n3325) );
  OR U3565 ( .A(n3282), .B(n3281), .Z(n3286) );
  NAND U3566 ( .A(n3284), .B(n3283), .Z(n3285) );
  AND U3567 ( .A(n3286), .B(n3285), .Z(n3326) );
  XNOR U3568 ( .A(n3325), .B(n3326), .Z(n3327) );
  NANDN U3569 ( .A(n3288), .B(n3287), .Z(n3292) );
  OR U3570 ( .A(n3290), .B(n3289), .Z(n3291) );
  NAND U3571 ( .A(n3292), .B(n3291), .Z(n3386) );
  NANDN U3572 ( .A(n3962), .B(n3642), .Z(n3296) );
  OR U3573 ( .A(n3294), .B(n3293), .Z(n3295) );
  NAND U3574 ( .A(n3296), .B(n3295), .Z(n3385) );
  XOR U3575 ( .A(n3386), .B(n3385), .Z(n3387) );
  NANDN U3576 ( .A(n3298), .B(n3297), .Z(n3302) );
  NANDN U3577 ( .A(n3300), .B(n3299), .Z(n3301) );
  AND U3578 ( .A(n3302), .B(n3301), .Z(n3388) );
  XNOR U3579 ( .A(n3387), .B(n3388), .Z(n3333) );
  OR U3580 ( .A(n3304), .B(n3303), .Z(n3308) );
  OR U3581 ( .A(n3306), .B(n3305), .Z(n3307) );
  NAND U3582 ( .A(n3308), .B(n3307), .Z(n3332) );
  ANDN U3583 ( .B(y[228]), .A(n52), .Z(n3360) );
  NAND U3584 ( .A(n3360), .B(n3368), .Z(n3312) );
  NANDN U3585 ( .A(n3310), .B(n3309), .Z(n3311) );
  AND U3586 ( .A(n3312), .B(n3311), .Z(n3376) );
  ANDN U3587 ( .B(y[226]), .A(n53), .Z(n3313) );
  XOR U3588 ( .A(n3313), .B(n3495), .Z(n3370) );
  NANDN U3589 ( .A(n54), .B(y[225]), .Z(n3343) );
  XOR U3590 ( .A(o[42]), .B(n3343), .Z(n3369) );
  XNOR U3591 ( .A(n3370), .B(n3369), .Z(n3374) );
  AND U3592 ( .A(y[228]), .B(x[70]), .Z(n3590) );
  ANDN U3593 ( .B(x[71]), .A(n5714), .Z(n3315) );
  NANDN U3594 ( .A(n49), .B(y[230]), .Z(n3314) );
  XOR U3595 ( .A(n3315), .B(n3314), .Z(n3356) );
  XOR U3596 ( .A(n3376), .B(n3375), .Z(n3381) );
  AND U3597 ( .A(y[234]), .B(x[64]), .Z(n3351) );
  ANDN U3598 ( .B(o[41]), .A(n3316), .Z(n3348) );
  AND U3599 ( .A(y[224]), .B(x[74]), .Z(n3349) );
  XNOR U3600 ( .A(n3351), .B(n3350), .Z(n3339) );
  AND U3601 ( .A(y[231]), .B(x[67]), .Z(n4320) );
  AND U3602 ( .A(y[232]), .B(x[66]), .Z(n3364) );
  XNOR U3603 ( .A(n4320), .B(n3364), .Z(n3365) );
  IV U3604 ( .A(y[233]), .Z(n5637) );
  ANDN U3605 ( .B(x[65]), .A(n5637), .Z(n4266) );
  XOR U3606 ( .A(n3365), .B(n4266), .Z(n3338) );
  AND U3607 ( .A(y[232]), .B(x[70]), .Z(n3686) );
  NANDN U3608 ( .A(n3317), .B(n3686), .Z(n3320) );
  NAND U3609 ( .A(n3318), .B(n3754), .Z(n3319) );
  AND U3610 ( .A(n3320), .B(n3319), .Z(n3337) );
  XNOR U3611 ( .A(n3338), .B(n3337), .Z(n3340) );
  AND U3612 ( .A(y[233]), .B(x[73]), .Z(n4021) );
  NAND U3613 ( .A(n3747), .B(n4021), .Z(n3324) );
  OR U3614 ( .A(n3322), .B(n3321), .Z(n3323) );
  NAND U3615 ( .A(n3324), .B(n3323), .Z(n3379) );
  XNOR U3616 ( .A(n3380), .B(n3379), .Z(n3382) );
  XOR U3617 ( .A(n3381), .B(n3382), .Z(n3331) );
  XNOR U3618 ( .A(n3332), .B(n3331), .Z(n3334) );
  XNOR U3619 ( .A(n3333), .B(n3334), .Z(n3328) );
  XOR U3620 ( .A(n3327), .B(n3328), .Z(N107) );
  NANDN U3621 ( .A(n3326), .B(n3325), .Z(n3330) );
  NANDN U3622 ( .A(n3328), .B(n3327), .Z(n3329) );
  NAND U3623 ( .A(n3330), .B(n3329), .Z(n3391) );
  OR U3624 ( .A(n3332), .B(n3331), .Z(n3336) );
  OR U3625 ( .A(n3334), .B(n3333), .Z(n3335) );
  AND U3626 ( .A(n3336), .B(n3335), .Z(n3392) );
  XNOR U3627 ( .A(n3391), .B(n3392), .Z(n3393) );
  OR U3628 ( .A(n3338), .B(n3337), .Z(n3342) );
  NANDN U3629 ( .A(n3340), .B(n3339), .Z(n3341) );
  NAND U3630 ( .A(n3342), .B(n3341), .Z(n3406) );
  NANDN U3631 ( .A(n3343), .B(o[42]), .Z(n3442) );
  ANDN U3632 ( .B(x[75]), .A(n5905), .Z(n3345) );
  NANDN U3633 ( .A(n45), .B(y[235]), .Z(n3344) );
  XOR U3634 ( .A(n3345), .B(n3344), .Z(n3441) );
  IV U3635 ( .A(y[234]), .Z(n5196) );
  ANDN U3636 ( .B(x[65]), .A(n5196), .Z(n3347) );
  NANDN U3637 ( .A(n51), .B(y[229]), .Z(n3346) );
  XOR U3638 ( .A(n3347), .B(n3346), .Z(n3438) );
  NANDN U3639 ( .A(n55), .B(y[225]), .Z(n3450) );
  XOR U3640 ( .A(n3450), .B(o[43]), .Z(n3437) );
  XNOR U3641 ( .A(n3438), .B(n3437), .Z(n3412) );
  XNOR U3642 ( .A(n3411), .B(n3412), .Z(n3413) );
  OR U3643 ( .A(n3349), .B(n3348), .Z(n3353) );
  OR U3644 ( .A(n3351), .B(n3350), .Z(n3352) );
  NAND U3645 ( .A(n3353), .B(n3352), .Z(n3414) );
  XNOR U3646 ( .A(n3413), .B(n3414), .Z(n3403) );
  ANDN U3647 ( .B(y[230]), .A(n52), .Z(n3355) );
  NAND U3648 ( .A(n3355), .B(n3354), .Z(n3358) );
  NANDN U3649 ( .A(n3356), .B(n3590), .Z(n3357) );
  NAND U3650 ( .A(n3358), .B(n3357), .Z(n3404) );
  XOR U3651 ( .A(n3406), .B(n3405), .Z(n3420) );
  NANDN U3652 ( .A(n54), .B(y[226]), .Z(n3359) );
  XOR U3653 ( .A(n3360), .B(n3359), .Z(n3447) );
  NANDN U3654 ( .A(n53), .B(y[227]), .Z(n3446) );
  XOR U3655 ( .A(n3447), .B(n3446), .Z(n3410) );
  ANDN U3656 ( .B(x[67]), .A(n5947), .Z(n4436) );
  IV U3657 ( .A(n4436), .Z(n3581) );
  NANDN U3658 ( .A(n49), .B(y[231]), .Z(n3432) );
  ANDN U3659 ( .B(x[66]), .A(n5637), .Z(n3362) );
  NANDN U3660 ( .A(n50), .B(y[230]), .Z(n3361) );
  XOR U3661 ( .A(n3362), .B(n3361), .Z(n3431) );
  XNOR U3662 ( .A(n3432), .B(n3431), .Z(n3409) );
  XOR U3663 ( .A(n3581), .B(n3409), .Z(n3363) );
  XOR U3664 ( .A(n3410), .B(n3363), .Z(n3456) );
  OR U3665 ( .A(n3364), .B(n4320), .Z(n3367) );
  OR U3666 ( .A(n3365), .B(n4266), .Z(n3366) );
  AND U3667 ( .A(n3367), .B(n3366), .Z(n3453) );
  AND U3668 ( .A(y[229]), .B(x[72]), .Z(n4197) );
  NAND U3669 ( .A(n4197), .B(n3368), .Z(n3372) );
  OR U3670 ( .A(n3370), .B(n3369), .Z(n3371) );
  NAND U3671 ( .A(n3372), .B(n3371), .Z(n3454) );
  XNOR U3672 ( .A(n3456), .B(n3455), .Z(n3418) );
  NANDN U3673 ( .A(n3374), .B(n3373), .Z(n3378) );
  NANDN U3674 ( .A(n3376), .B(n3375), .Z(n3377) );
  AND U3675 ( .A(n3378), .B(n3377), .Z(n3417) );
  XOR U3676 ( .A(n3418), .B(n3417), .Z(n3419) );
  XOR U3677 ( .A(n3420), .B(n3419), .Z(n3397) );
  OR U3678 ( .A(n3380), .B(n3379), .Z(n3384) );
  NANDN U3679 ( .A(n3382), .B(n3381), .Z(n3383) );
  AND U3680 ( .A(n3384), .B(n3383), .Z(n3398) );
  XNOR U3681 ( .A(n3397), .B(n3398), .Z(n3400) );
  OR U3682 ( .A(n3386), .B(n3385), .Z(n3390) );
  NANDN U3683 ( .A(n3388), .B(n3387), .Z(n3389) );
  NAND U3684 ( .A(n3390), .B(n3389), .Z(n3399) );
  XOR U3685 ( .A(n3400), .B(n3399), .Z(n3394) );
  XNOR U3686 ( .A(n3393), .B(n3394), .Z(N108) );
  NANDN U3687 ( .A(n3392), .B(n3391), .Z(n3396) );
  NAND U3688 ( .A(n3394), .B(n3393), .Z(n3395) );
  NAND U3689 ( .A(n3396), .B(n3395), .Z(n3459) );
  OR U3690 ( .A(n3398), .B(n3397), .Z(n3402) );
  OR U3691 ( .A(n3400), .B(n3399), .Z(n3401) );
  AND U3692 ( .A(n3402), .B(n3401), .Z(n3460) );
  XNOR U3693 ( .A(n3459), .B(n3460), .Z(n3461) );
  OR U3694 ( .A(n3404), .B(n3403), .Z(n3408) );
  NANDN U3695 ( .A(n3406), .B(n3405), .Z(n3407) );
  NAND U3696 ( .A(n3408), .B(n3407), .Z(n3534) );
  NANDN U3697 ( .A(n3412), .B(n3411), .Z(n3416) );
  NANDN U3698 ( .A(n3414), .B(n3413), .Z(n3415) );
  NAND U3699 ( .A(n3416), .B(n3415), .Z(n3532) );
  XOR U3700 ( .A(n3534), .B(n3535), .Z(n3468) );
  OR U3701 ( .A(n3418), .B(n3417), .Z(n3422) );
  NAND U3702 ( .A(n3420), .B(n3419), .Z(n3421) );
  AND U3703 ( .A(n3422), .B(n3421), .Z(n3465) );
  ANDN U3704 ( .B(y[229]), .A(n52), .Z(n3424) );
  NANDN U3705 ( .A(n50), .B(y[231]), .Z(n3423) );
  XOR U3706 ( .A(n3424), .B(n3423), .Z(n3497) );
  ANDN U3707 ( .B(y[226]), .A(n55), .Z(n3426) );
  NANDN U3708 ( .A(n54), .B(y[227]), .Z(n3425) );
  XOR U3709 ( .A(n3426), .B(n3425), .Z(n3519) );
  NANDN U3710 ( .A(n49), .B(y[232]), .Z(n3518) );
  XNOR U3711 ( .A(n3519), .B(n3518), .Z(n3496) );
  XOR U3712 ( .A(n3497), .B(n3496), .Z(n3490) );
  ANDN U3713 ( .B(x[76]), .A(n5905), .Z(n3428) );
  NANDN U3714 ( .A(n45), .B(y[236]), .Z(n3427) );
  XOR U3715 ( .A(n3428), .B(n3427), .Z(n3511) );
  NANDN U3716 ( .A(n56), .B(y[225]), .Z(n3485) );
  XOR U3717 ( .A(o[44]), .B(n3485), .Z(n3510) );
  XOR U3718 ( .A(n3511), .B(n3510), .Z(n3488) );
  ANDN U3719 ( .B(x[66]), .A(n5196), .Z(n3430) );
  NANDN U3720 ( .A(n53), .B(y[228]), .Z(n3429) );
  XOR U3721 ( .A(n3430), .B(n3429), .Z(n3480) );
  NANDN U3722 ( .A(n5637), .B(x[67]), .Z(n3479) );
  XNOR U3723 ( .A(n3480), .B(n3479), .Z(n3489) );
  XOR U3724 ( .A(n3488), .B(n3489), .Z(n3491) );
  XOR U3725 ( .A(n3490), .B(n3491), .Z(n3473) );
  AND U3726 ( .A(y[233]), .B(x[69]), .Z(n3643) );
  NANDN U3727 ( .A(n3763), .B(n3643), .Z(n3434) );
  OR U3728 ( .A(n3432), .B(n3431), .Z(n3433) );
  NAND U3729 ( .A(n3434), .B(n3433), .Z(n3472) );
  ANDN U3730 ( .B(y[234]), .A(n51), .Z(n3436) );
  NAND U3731 ( .A(n3436), .B(n3435), .Z(n3440) );
  OR U3732 ( .A(n3438), .B(n3437), .Z(n3439) );
  NAND U3733 ( .A(n3440), .B(n3439), .Z(n3471) );
  XNOR U3734 ( .A(n3472), .B(n3471), .Z(n3474) );
  XNOR U3735 ( .A(n3473), .B(n3474), .Z(n3527) );
  ANDN U3736 ( .B(y[235]), .A(n56), .Z(n4587) );
  NAND U3737 ( .A(n3747), .B(n4587), .Z(n3444) );
  OR U3738 ( .A(n3442), .B(n3441), .Z(n3443) );
  AND U3739 ( .A(n3444), .B(n3443), .Z(n3502) );
  NANDN U3740 ( .A(n52), .B(y[226]), .Z(n3674) );
  ANDN U3741 ( .B(y[228]), .A(n54), .Z(n3445) );
  NANDN U3742 ( .A(n3674), .B(n3445), .Z(n3449) );
  OR U3743 ( .A(n3447), .B(n3446), .Z(n3448) );
  NAND U3744 ( .A(n3449), .B(n3448), .Z(n3501) );
  NANDN U3745 ( .A(n3450), .B(o[43]), .Z(n3507) );
  ANDN U3746 ( .B(y[235]), .A(n46), .Z(n3452) );
  NANDN U3747 ( .A(n51), .B(y[230]), .Z(n3451) );
  XOR U3748 ( .A(n3452), .B(n3451), .Z(n3506) );
  XNOR U3749 ( .A(n3501), .B(n3500), .Z(n3503) );
  XOR U3750 ( .A(n3527), .B(n3526), .Z(n3529) );
  OR U3751 ( .A(n3454), .B(n3453), .Z(n3458) );
  NANDN U3752 ( .A(n3456), .B(n3455), .Z(n3457) );
  AND U3753 ( .A(n3458), .B(n3457), .Z(n3528) );
  XOR U3754 ( .A(n3529), .B(n3528), .Z(n3466) );
  XOR U3755 ( .A(n3468), .B(n3467), .Z(n3462) );
  XOR U3756 ( .A(n3461), .B(n3462), .Z(N109) );
  NANDN U3757 ( .A(n3460), .B(n3459), .Z(n3464) );
  NANDN U3758 ( .A(n3462), .B(n3461), .Z(n3463) );
  NAND U3759 ( .A(n3464), .B(n3463), .Z(n3606) );
  OR U3760 ( .A(n3466), .B(n3465), .Z(n3470) );
  NAND U3761 ( .A(n3468), .B(n3467), .Z(n3469) );
  NAND U3762 ( .A(n3470), .B(n3469), .Z(n3607) );
  XNOR U3763 ( .A(n3606), .B(n3607), .Z(n3608) );
  OR U3764 ( .A(n3472), .B(n3471), .Z(n3476) );
  NANDN U3765 ( .A(n3474), .B(n3473), .Z(n3475) );
  AND U3766 ( .A(n3476), .B(n3475), .Z(n3544) );
  ANDN U3767 ( .B(y[234]), .A(n53), .Z(n3478) );
  NAND U3768 ( .A(n3478), .B(n3477), .Z(n3482) );
  OR U3769 ( .A(n3480), .B(n3479), .Z(n3481) );
  NAND U3770 ( .A(n3482), .B(n3481), .Z(n3565) );
  ANDN U3771 ( .B(x[70]), .A(n44), .Z(n3484) );
  NANDN U3772 ( .A(n54), .B(y[228]), .Z(n3483) );
  XOR U3773 ( .A(n3484), .B(n3483), .Z(n3593) );
  NANDN U3774 ( .A(n47), .B(y[235]), .Z(n3592) );
  XNOR U3775 ( .A(n3593), .B(n3592), .Z(n3563) );
  NANDN U3776 ( .A(n3485), .B(o[44]), .Z(n3575) );
  ANDN U3777 ( .B(y[236]), .A(n46), .Z(n3487) );
  NANDN U3778 ( .A(n52), .B(y[230]), .Z(n3486) );
  XOR U3779 ( .A(n3487), .B(n3486), .Z(n3574) );
  XNOR U3780 ( .A(n3565), .B(n3564), .Z(n3541) );
  NANDN U3781 ( .A(n3489), .B(n3488), .Z(n3493) );
  NANDN U3782 ( .A(n3491), .B(n3490), .Z(n3492) );
  AND U3783 ( .A(n3493), .B(n3492), .Z(n3538) );
  ANDN U3784 ( .B(y[231]), .A(n52), .Z(n3494) );
  NANDN U3785 ( .A(n3495), .B(n3494), .Z(n3499) );
  OR U3786 ( .A(n3497), .B(n3496), .Z(n3498) );
  AND U3787 ( .A(n3499), .B(n3498), .Z(n3539) );
  XOR U3788 ( .A(n3538), .B(n3539), .Z(n3540) );
  XNOR U3789 ( .A(n3541), .B(n3540), .Z(n3545) );
  XOR U3790 ( .A(n3544), .B(n3545), .Z(n3546) );
  NAND U3791 ( .A(n3501), .B(n3500), .Z(n3505) );
  OR U3792 ( .A(n3503), .B(n3502), .Z(n3504) );
  NAND U3793 ( .A(n3505), .B(n3504), .Z(n3553) );
  AND U3794 ( .A(y[235]), .B(x[70]), .Z(n3969) );
  NAND U3795 ( .A(n3572), .B(n3969), .Z(n3509) );
  OR U3796 ( .A(n3507), .B(n3506), .Z(n3508) );
  NAND U3797 ( .A(n3509), .B(n3508), .Z(n3558) );
  AND U3798 ( .A(y[236]), .B(x[76]), .Z(n4797) );
  NAND U3799 ( .A(n3747), .B(n4797), .Z(n3513) );
  OR U3800 ( .A(n3511), .B(n3510), .Z(n3512) );
  AND U3801 ( .A(n3513), .B(n3512), .Z(n3556) );
  ANDN U3802 ( .B(y[226]), .A(n56), .Z(n3515) );
  NANDN U3803 ( .A(n55), .B(y[227]), .Z(n3514) );
  XNOR U3804 ( .A(n3515), .B(n3514), .Z(n3578) );
  XNOR U3805 ( .A(n4197), .B(n3578), .Z(n3557) );
  XOR U3806 ( .A(n3558), .B(n3559), .Z(n3550) );
  ANDN U3807 ( .B(y[226]), .A(n54), .Z(n3517) );
  ANDN U3808 ( .B(y[227]), .A(n55), .Z(n3516) );
  NAND U3809 ( .A(n3517), .B(n3516), .Z(n3521) );
  OR U3810 ( .A(n3519), .B(n3518), .Z(n3520) );
  NAND U3811 ( .A(n3521), .B(n3520), .Z(n3603) );
  ANDN U3812 ( .B(x[77]), .A(n5905), .Z(n3523) );
  NANDN U3813 ( .A(n45), .B(y[237]), .Z(n3522) );
  XOR U3814 ( .A(n3523), .B(n3522), .Z(n3587) );
  NANDN U3815 ( .A(n57), .B(y[225]), .Z(n3597) );
  XOR U3816 ( .A(o[45]), .B(n3597), .Z(n3586) );
  XNOR U3817 ( .A(n3587), .B(n3586), .Z(n3601) );
  ANDN U3818 ( .B(x[67]), .A(n5196), .Z(n3525) );
  NANDN U3819 ( .A(n50), .B(y[232]), .Z(n3524) );
  XOR U3820 ( .A(n3525), .B(n3524), .Z(n3583) );
  NANDN U3821 ( .A(n5637), .B(x[68]), .Z(n3582) );
  XOR U3822 ( .A(n3583), .B(n3582), .Z(n3600) );
  XOR U3823 ( .A(n3603), .B(n3602), .Z(n3551) );
  XNOR U3824 ( .A(n3550), .B(n3551), .Z(n3552) );
  XOR U3825 ( .A(n3553), .B(n3552), .Z(n3547) );
  XNOR U3826 ( .A(n3546), .B(n3547), .Z(n3615) );
  NANDN U3827 ( .A(n3527), .B(n3526), .Z(n3531) );
  NANDN U3828 ( .A(n3529), .B(n3528), .Z(n3530) );
  AND U3829 ( .A(n3531), .B(n3530), .Z(n3612) );
  OR U3830 ( .A(n3533), .B(n3532), .Z(n3537) );
  NANDN U3831 ( .A(n3535), .B(n3534), .Z(n3536) );
  NAND U3832 ( .A(n3537), .B(n3536), .Z(n3613) );
  XNOR U3833 ( .A(n3615), .B(n3614), .Z(n3609) );
  XOR U3834 ( .A(n3608), .B(n3609), .Z(N110) );
  OR U3835 ( .A(n3539), .B(n3538), .Z(n3543) );
  NANDN U3836 ( .A(n3541), .B(n3540), .Z(n3542) );
  NAND U3837 ( .A(n3543), .B(n3542), .Z(n3627) );
  OR U3838 ( .A(n3545), .B(n3544), .Z(n3549) );
  NANDN U3839 ( .A(n3547), .B(n3546), .Z(n3548) );
  AND U3840 ( .A(n3549), .B(n3548), .Z(n3624) );
  NANDN U3841 ( .A(n3551), .B(n3550), .Z(n3555) );
  NANDN U3842 ( .A(n3553), .B(n3552), .Z(n3554) );
  AND U3843 ( .A(n3555), .B(n3554), .Z(n3704) );
  OR U3844 ( .A(n3557), .B(n3556), .Z(n3561) );
  NANDN U3845 ( .A(n3559), .B(n3558), .Z(n3560) );
  NAND U3846 ( .A(n3561), .B(n3560), .Z(n3638) );
  NANDN U3847 ( .A(n3563), .B(n3562), .Z(n3567) );
  NAND U3848 ( .A(n3565), .B(n3564), .Z(n3566) );
  AND U3849 ( .A(n3567), .B(n3566), .Z(n3636) );
  AND U3850 ( .A(y[234]), .B(x[68]), .Z(n3658) );
  ANDN U3851 ( .B(y[228]), .A(n55), .Z(n4326) );
  ANDN U3852 ( .B(y[236]), .A(n47), .Z(n3569) );
  NANDN U3853 ( .A(n54), .B(y[229]), .Z(n3568) );
  XOR U3854 ( .A(n3569), .B(n3568), .Z(n3670) );
  XNOR U3855 ( .A(n4326), .B(n3670), .Z(n3657) );
  XNOR U3856 ( .A(n3658), .B(n3657), .Z(n3660) );
  ANDN U3857 ( .B(y[235]), .A(n48), .Z(n3571) );
  NANDN U3858 ( .A(n53), .B(y[230]), .Z(n3570) );
  XOR U3859 ( .A(n3571), .B(n3570), .Z(n3644) );
  XOR U3860 ( .A(n3643), .B(n3644), .Z(n3659) );
  ANDN U3861 ( .B(y[236]), .A(n52), .Z(n3573) );
  NAND U3862 ( .A(n3573), .B(n3572), .Z(n3577) );
  OR U3863 ( .A(n3575), .B(n3574), .Z(n3576) );
  AND U3864 ( .A(n3577), .B(n3576), .Z(n3663) );
  NANDN U3865 ( .A(n55), .B(y[226]), .Z(n4202) );
  AND U3866 ( .A(x[75]), .B(y[227]), .Z(n3780) );
  NANDN U3867 ( .A(n4202), .B(n3780), .Z(n3580) );
  NAND U3868 ( .A(n3578), .B(n4197), .Z(n3579) );
  AND U3869 ( .A(n3580), .B(n3579), .Z(n3664) );
  XOR U3870 ( .A(n3666), .B(n3665), .Z(n3637) );
  XOR U3871 ( .A(n3638), .B(n3639), .Z(n3701) );
  AND U3872 ( .A(y[234]), .B(x[69]), .Z(n3737) );
  NANDN U3873 ( .A(n3581), .B(n3737), .Z(n3585) );
  OR U3874 ( .A(n3583), .B(n3582), .Z(n3584) );
  NAND U3875 ( .A(n3585), .B(n3584), .Z(n3697) );
  NAND U3876 ( .A(y[237]), .B(x[65]), .Z(n3684) );
  XOR U3877 ( .A(n3780), .B(n3684), .Z(n3685) );
  XOR U3878 ( .A(n3686), .B(n3685), .Z(n3696) );
  AND U3879 ( .A(x[77]), .B(y[237]), .Z(n5184) );
  NAND U3880 ( .A(n3747), .B(n5184), .Z(n3589) );
  OR U3881 ( .A(n3587), .B(n3586), .Z(n3588) );
  AND U3882 ( .A(n3589), .B(n3588), .Z(n3695) );
  XNOR U3883 ( .A(n3696), .B(n3695), .Z(n3698) );
  XOR U3884 ( .A(n3697), .B(n3698), .Z(n3632) );
  ANDN U3885 ( .B(y[231]), .A(n54), .Z(n3591) );
  NAND U3886 ( .A(n3591), .B(n3590), .Z(n3595) );
  OR U3887 ( .A(n3593), .B(n3592), .Z(n3594) );
  AND U3888 ( .A(n3595), .B(n3594), .Z(n3692) );
  ANDN U3889 ( .B(y[226]), .A(n57), .Z(n4255) );
  NANDN U3890 ( .A(n52), .B(y[231]), .Z(n3596) );
  XOR U3891 ( .A(n4255), .B(n3596), .Z(n3676) );
  NANDN U3892 ( .A(n58), .B(y[225]), .Z(n3679) );
  XOR U3893 ( .A(o[46]), .B(n3679), .Z(n3675) );
  XNOR U3894 ( .A(n3676), .B(n3675), .Z(n3690) );
  NANDN U3895 ( .A(n3597), .B(o[45]), .Z(n3648) );
  ANDN U3896 ( .B(x[78]), .A(n5905), .Z(n3599) );
  NANDN U3897 ( .A(n45), .B(y[238]), .Z(n3598) );
  XOR U3898 ( .A(n3599), .B(n3598), .Z(n3647) );
  XOR U3899 ( .A(n3692), .B(n3691), .Z(n3630) );
  NANDN U3900 ( .A(n3601), .B(n3600), .Z(n3605) );
  NAND U3901 ( .A(n3603), .B(n3602), .Z(n3604) );
  NAND U3902 ( .A(n3605), .B(n3604), .Z(n3631) );
  XOR U3903 ( .A(n3630), .B(n3631), .Z(n3633) );
  XOR U3904 ( .A(n3632), .B(n3633), .Z(n3702) );
  XOR U3905 ( .A(n3704), .B(n3703), .Z(n3625) );
  XNOR U3906 ( .A(n3624), .B(n3625), .Z(n3626) );
  XNOR U3907 ( .A(n3627), .B(n3626), .Z(n3621) );
  NANDN U3908 ( .A(n3607), .B(n3606), .Z(n3611) );
  NANDN U3909 ( .A(n3609), .B(n3608), .Z(n3610) );
  NAND U3910 ( .A(n3611), .B(n3610), .Z(n3618) );
  OR U3911 ( .A(n3613), .B(n3612), .Z(n3617) );
  NANDN U3912 ( .A(n3615), .B(n3614), .Z(n3616) );
  NAND U3913 ( .A(n3617), .B(n3616), .Z(n3619) );
  XNOR U3914 ( .A(n3618), .B(n3619), .Z(n3620) );
  XOR U3915 ( .A(n3621), .B(n3620), .Z(N111) );
  NANDN U3916 ( .A(n3619), .B(n3618), .Z(n3623) );
  NANDN U3917 ( .A(n3621), .B(n3620), .Z(n3622) );
  NAND U3918 ( .A(n3623), .B(n3622), .Z(n3707) );
  OR U3919 ( .A(n3625), .B(n3624), .Z(n3629) );
  OR U3920 ( .A(n3627), .B(n3626), .Z(n3628) );
  AND U3921 ( .A(n3629), .B(n3628), .Z(n3708) );
  XNOR U3922 ( .A(n3707), .B(n3708), .Z(n3709) );
  NANDN U3923 ( .A(n3631), .B(n3630), .Z(n3635) );
  NANDN U3924 ( .A(n3633), .B(n3632), .Z(n3634) );
  NAND U3925 ( .A(n3635), .B(n3634), .Z(n3714) );
  OR U3926 ( .A(n3637), .B(n3636), .Z(n3641) );
  NANDN U3927 ( .A(n3639), .B(n3638), .Z(n3640) );
  AND U3928 ( .A(n3641), .B(n3640), .Z(n3798) );
  NANDN U3929 ( .A(n53), .B(y[235]), .Z(n4066) );
  OR U3930 ( .A(n4066), .B(n3642), .Z(n3646) );
  NANDN U3931 ( .A(n3644), .B(n3643), .Z(n3645) );
  NAND U3932 ( .A(n3646), .B(n3645), .Z(n3769) );
  AND U3933 ( .A(x[78]), .B(y[238]), .Z(n5395) );
  NAND U3934 ( .A(n3747), .B(n5395), .Z(n3650) );
  OR U3935 ( .A(n3648), .B(n3647), .Z(n3649) );
  NAND U3936 ( .A(n3650), .B(n3649), .Z(n3768) );
  AND U3937 ( .A(y[232]), .B(x[71]), .Z(n4149) );
  ANDN U3938 ( .B(y[229]), .A(n55), .Z(n3652) );
  NANDN U3939 ( .A(n49), .B(y[235]), .Z(n3651) );
  XOR U3940 ( .A(n3652), .B(n3651), .Z(n3755) );
  XNOR U3941 ( .A(n4149), .B(n3755), .Z(n3738) );
  ANDN U3942 ( .B(x[70]), .A(n5637), .Z(n3864) );
  XNOR U3943 ( .A(n3737), .B(n3864), .Z(n3739) );
  ANDN U3944 ( .B(y[225]), .A(n59), .Z(n3758) );
  XNOR U3945 ( .A(o[47]), .B(n3758), .Z(n3744) );
  IV U3946 ( .A(y[238]), .Z(n5473) );
  ANDN U3947 ( .B(x[65]), .A(n5473), .Z(n3654) );
  NANDN U3948 ( .A(n53), .B(y[231]), .Z(n3653) );
  XNOR U3949 ( .A(n3654), .B(n3653), .Z(n3743) );
  XNOR U3950 ( .A(n3744), .B(n3743), .Z(n3775) );
  NANDN U3951 ( .A(n48), .B(y[236]), .Z(n3765) );
  IV U3952 ( .A(y[237]), .Z(n5332) );
  ANDN U3953 ( .B(x[66]), .A(n5332), .Z(n3656) );
  NANDN U3954 ( .A(n54), .B(y[230]), .Z(n3655) );
  XOR U3955 ( .A(n3656), .B(n3655), .Z(n3764) );
  XNOR U3956 ( .A(n3765), .B(n3764), .Z(n3774) );
  XOR U3957 ( .A(n3775), .B(n3774), .Z(n3777) );
  XOR U3958 ( .A(n3776), .B(n3777), .Z(n3771) );
  XNOR U3959 ( .A(n3770), .B(n3771), .Z(n3731) );
  OR U3960 ( .A(n3658), .B(n3657), .Z(n3662) );
  NANDN U3961 ( .A(n3660), .B(n3659), .Z(n3661) );
  NAND U3962 ( .A(n3662), .B(n3661), .Z(n3732) );
  XNOR U3963 ( .A(n3731), .B(n3732), .Z(n3734) );
  OR U3964 ( .A(n3664), .B(n3663), .Z(n3668) );
  NANDN U3965 ( .A(n3666), .B(n3665), .Z(n3667) );
  AND U3966 ( .A(n3668), .B(n3667), .Z(n3733) );
  XNOR U3967 ( .A(n3734), .B(n3733), .Z(n3796) );
  AND U3968 ( .A(y[236]), .B(x[73]), .Z(n4415) );
  NAND U3969 ( .A(n3669), .B(n4415), .Z(n3672) );
  NANDN U3970 ( .A(n3670), .B(n4326), .Z(n3671) );
  AND U3971 ( .A(n3672), .B(n3671), .Z(n3725) );
  ANDN U3972 ( .B(y[231]), .A(n57), .Z(n3673) );
  NANDN U3973 ( .A(n3674), .B(n3673), .Z(n3678) );
  OR U3974 ( .A(n3676), .B(n3675), .Z(n3677) );
  NAND U3975 ( .A(n3678), .B(n3677), .Z(n3792) );
  NANDN U3976 ( .A(n3679), .B(o[46]), .Z(n3749) );
  ANDN U3977 ( .B(x[79]), .A(n5905), .Z(n3681) );
  NANDN U3978 ( .A(n45), .B(y[239]), .Z(n3680) );
  XOR U3979 ( .A(n3681), .B(n3680), .Z(n3748) );
  XOR U3980 ( .A(n3749), .B(n3748), .Z(n3789) );
  ANDN U3981 ( .B(x[76]), .A(n5714), .Z(n3683) );
  NANDN U3982 ( .A(n56), .B(y[228]), .Z(n3682) );
  XOR U3983 ( .A(n3683), .B(n3682), .Z(n3782) );
  NANDN U3984 ( .A(n58), .B(y[226]), .Z(n3781) );
  XOR U3985 ( .A(n3782), .B(n3781), .Z(n3790) );
  XNOR U3986 ( .A(n3792), .B(n3791), .Z(n3726) );
  XNOR U3987 ( .A(n3725), .B(n3726), .Z(n3727) );
  NANDN U3988 ( .A(n3780), .B(n3684), .Z(n3688) );
  OR U3989 ( .A(n3686), .B(n3685), .Z(n3687) );
  NAND U3990 ( .A(n3688), .B(n3687), .Z(n3728) );
  NANDN U3991 ( .A(n3690), .B(n3689), .Z(n3694) );
  NANDN U3992 ( .A(n3692), .B(n3691), .Z(n3693) );
  AND U3993 ( .A(n3694), .B(n3693), .Z(n3719) );
  XNOR U3994 ( .A(n3720), .B(n3719), .Z(n3722) );
  OR U3995 ( .A(n3696), .B(n3695), .Z(n3700) );
  NANDN U3996 ( .A(n3698), .B(n3697), .Z(n3699) );
  AND U3997 ( .A(n3700), .B(n3699), .Z(n3721) );
  XOR U3998 ( .A(n3722), .B(n3721), .Z(n3795) );
  XNOR U3999 ( .A(n3798), .B(n3797), .Z(n3713) );
  XOR U4000 ( .A(n3714), .B(n3713), .Z(n3716) );
  NANDN U4001 ( .A(n3702), .B(n3701), .Z(n3706) );
  NANDN U4002 ( .A(n3704), .B(n3703), .Z(n3705) );
  NAND U4003 ( .A(n3706), .B(n3705), .Z(n3715) );
  XOR U4004 ( .A(n3716), .B(n3715), .Z(n3710) );
  XOR U4005 ( .A(n3709), .B(n3710), .Z(N112) );
  NANDN U4006 ( .A(n3708), .B(n3707), .Z(n3712) );
  NANDN U4007 ( .A(n3710), .B(n3709), .Z(n3711) );
  NAND U4008 ( .A(n3712), .B(n3711), .Z(n3801) );
  NANDN U4009 ( .A(n3714), .B(n3713), .Z(n3718) );
  OR U4010 ( .A(n3716), .B(n3715), .Z(n3717) );
  NAND U4011 ( .A(n3718), .B(n3717), .Z(n3802) );
  XNOR U4012 ( .A(n3801), .B(n3802), .Z(n3803) );
  OR U4013 ( .A(n3720), .B(n3719), .Z(n3724) );
  OR U4014 ( .A(n3722), .B(n3721), .Z(n3723) );
  NAND U4015 ( .A(n3724), .B(n3723), .Z(n3891) );
  OR U4016 ( .A(n3726), .B(n3725), .Z(n3730) );
  OR U4017 ( .A(n3728), .B(n3727), .Z(n3729) );
  NAND U4018 ( .A(n3730), .B(n3729), .Z(n3889) );
  OR U4019 ( .A(n3732), .B(n3731), .Z(n3736) );
  OR U4020 ( .A(n3734), .B(n3733), .Z(n3735) );
  NAND U4021 ( .A(n3736), .B(n3735), .Z(n3888) );
  XOR U4022 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U4023 ( .A(n3891), .B(n3890), .Z(n3810) );
  OR U4024 ( .A(n3737), .B(n3864), .Z(n3741) );
  OR U4025 ( .A(n3739), .B(n3738), .Z(n3740) );
  AND U4026 ( .A(n3741), .B(n3740), .Z(n3846) );
  NANDN U4027 ( .A(n53), .B(y[238]), .Z(n4742) );
  NANDN U4028 ( .A(n4742), .B(n3742), .Z(n3746) );
  NANDN U4029 ( .A(n3744), .B(n3743), .Z(n3745) );
  AND U4030 ( .A(n3746), .B(n3745), .Z(n3819) );
  ANDN U4031 ( .B(y[239]), .A(n60), .Z(n5920) );
  NAND U4032 ( .A(n3747), .B(n5920), .Z(n3751) );
  OR U4033 ( .A(n3749), .B(n3748), .Z(n3750) );
  AND U4034 ( .A(n3751), .B(n3750), .Z(n3820) );
  NANDN U4035 ( .A(n45), .B(y[240]), .Z(n3876) );
  ANDN U4036 ( .B(x[80]), .A(n5905), .Z(n3875) );
  XNOR U4037 ( .A(n3876), .B(n3875), .Z(n3878) );
  NANDN U4038 ( .A(n60), .B(y[225]), .Z(n3885) );
  XNOR U4039 ( .A(n3885), .B(o[48]), .Z(n3877) );
  XNOR U4040 ( .A(n3878), .B(n3877), .Z(n3859) );
  ANDN U4041 ( .B(x[71]), .A(n5637), .Z(n3753) );
  NANDN U4042 ( .A(n51), .B(y[234]), .Z(n3752) );
  XOR U4043 ( .A(n3753), .B(n3752), .Z(n3866) );
  NANDN U4044 ( .A(n55), .B(y[230]), .Z(n3865) );
  XNOR U4045 ( .A(n3866), .B(n3865), .Z(n3858) );
  XNOR U4046 ( .A(n3859), .B(n3858), .Z(n3861) );
  AND U4047 ( .A(y[235]), .B(x[74]), .Z(n4465) );
  NAND U4048 ( .A(n3754), .B(n4465), .Z(n3757) );
  NANDN U4049 ( .A(n3755), .B(n4149), .Z(n3756) );
  AND U4050 ( .A(n3757), .B(n3756), .Z(n3860) );
  XOR U4051 ( .A(n3861), .B(n3860), .Z(n3822) );
  XOR U4052 ( .A(n3821), .B(n3822), .Z(n3847) );
  XOR U4053 ( .A(n3846), .B(n3847), .Z(n3848) );
  NAND U4054 ( .A(n3758), .B(o[47]), .Z(n3870) );
  IV U4055 ( .A(y[239]), .Z(n5936) );
  ANDN U4056 ( .B(x[65]), .A(n5936), .Z(n3760) );
  NANDN U4057 ( .A(n53), .B(y[232]), .Z(n3759) );
  XOR U4058 ( .A(n3760), .B(n3759), .Z(n3869) );
  XNOR U4059 ( .A(n3870), .B(n3869), .Z(n3854) );
  ANDN U4060 ( .B(y[229]), .A(n56), .Z(n3762) );
  NANDN U4061 ( .A(n59), .B(y[226]), .Z(n3761) );
  XOR U4062 ( .A(n3762), .B(n3761), .Z(n3831) );
  NANDN U4063 ( .A(n49), .B(y[236]), .Z(n3830) );
  XOR U4064 ( .A(n3831), .B(n3830), .Z(n3853) );
  ANDN U4065 ( .B(y[237]), .A(n54), .Z(n4539) );
  NANDN U4066 ( .A(n3763), .B(n4539), .Z(n3767) );
  OR U4067 ( .A(n3765), .B(n3764), .Z(n3766) );
  NAND U4068 ( .A(n3767), .B(n3766), .Z(n3852) );
  XNOR U4069 ( .A(n3853), .B(n3852), .Z(n3855) );
  XOR U4070 ( .A(n3854), .B(n3855), .Z(n3849) );
  XOR U4071 ( .A(n3848), .B(n3849), .Z(n3841) );
  OR U4072 ( .A(n3769), .B(n3768), .Z(n3773) );
  NANDN U4073 ( .A(n3771), .B(n3770), .Z(n3772) );
  AND U4074 ( .A(n3773), .B(n3772), .Z(n3840) );
  XOR U4075 ( .A(n3841), .B(n3840), .Z(n3842) );
  NANDN U4076 ( .A(n3775), .B(n3774), .Z(n3779) );
  NANDN U4077 ( .A(n3777), .B(n3776), .Z(n3778) );
  AND U4078 ( .A(n3779), .B(n3778), .Z(n3813) );
  NANDN U4079 ( .A(n57), .B(y[228]), .Z(n4543) );
  NANDN U4080 ( .A(n4543), .B(n3780), .Z(n3784) );
  OR U4081 ( .A(n3782), .B(n3781), .Z(n3783) );
  NAND U4082 ( .A(n3784), .B(n3783), .Z(n3837) );
  ANDN U4083 ( .B(x[66]), .A(n5473), .Z(n3786) );
  NANDN U4084 ( .A(n54), .B(y[231]), .Z(n3785) );
  XOR U4085 ( .A(n3786), .B(n3785), .Z(n3827) );
  NANDN U4086 ( .A(n5332), .B(x[67]), .Z(n3826) );
  XNOR U4087 ( .A(n3827), .B(n3826), .Z(n3835) );
  ANDN U4088 ( .B(x[77]), .A(n5714), .Z(n3788) );
  ANDN U4089 ( .B(y[235]), .A(n50), .Z(n3787) );
  XNOR U4090 ( .A(n3788), .B(n3787), .Z(n3882) );
  XOR U4091 ( .A(n4543), .B(n3882), .Z(n3834) );
  XOR U4092 ( .A(n3837), .B(n3836), .Z(n3814) );
  XNOR U4093 ( .A(n3813), .B(n3814), .Z(n3815) );
  OR U4094 ( .A(n3790), .B(n3789), .Z(n3794) );
  NANDN U4095 ( .A(n3792), .B(n3791), .Z(n3793) );
  AND U4096 ( .A(n3794), .B(n3793), .Z(n3816) );
  XNOR U4097 ( .A(n3842), .B(n3843), .Z(n3808) );
  NANDN U4098 ( .A(n3796), .B(n3795), .Z(n3800) );
  NANDN U4099 ( .A(n3798), .B(n3797), .Z(n3799) );
  AND U4100 ( .A(n3800), .B(n3799), .Z(n3807) );
  XOR U4101 ( .A(n3808), .B(n3807), .Z(n3809) );
  XNOR U4102 ( .A(n3810), .B(n3809), .Z(n3804) );
  XOR U4103 ( .A(n3803), .B(n3804), .Z(N113) );
  NANDN U4104 ( .A(n3802), .B(n3801), .Z(n3806) );
  NANDN U4105 ( .A(n3804), .B(n3803), .Z(n3805) );
  NAND U4106 ( .A(n3806), .B(n3805), .Z(n3894) );
  OR U4107 ( .A(n3808), .B(n3807), .Z(n3812) );
  NANDN U4108 ( .A(n3810), .B(n3809), .Z(n3811) );
  NAND U4109 ( .A(n3812), .B(n3811), .Z(n3895) );
  XNOR U4110 ( .A(n3894), .B(n3895), .Z(n3896) );
  OR U4111 ( .A(n3814), .B(n3813), .Z(n3818) );
  OR U4112 ( .A(n3816), .B(n3815), .Z(n3817) );
  NAND U4113 ( .A(n3818), .B(n3817), .Z(n3992) );
  OR U4114 ( .A(n3820), .B(n3819), .Z(n3824) );
  NAND U4115 ( .A(n3822), .B(n3821), .Z(n3823) );
  NAND U4116 ( .A(n3824), .B(n3823), .Z(n3988) );
  AND U4117 ( .A(y[234]), .B(x[71]), .Z(n4065) );
  AND U4118 ( .A(y[237]), .B(x[68]), .Z(n3931) );
  AND U4119 ( .A(y[230]), .B(x[75]), .Z(n3929) );
  AND U4120 ( .A(y[228]), .B(x[77]), .Z(n3930) );
  XNOR U4121 ( .A(n3929), .B(n3930), .Z(n3932) );
  XOR U4122 ( .A(n3931), .B(n3932), .Z(n3958) );
  AND U4123 ( .A(y[236]), .B(x[69]), .Z(n3971) );
  AND U4124 ( .A(y[233]), .B(x[72]), .Z(n3970) );
  XNOR U4125 ( .A(n3969), .B(n3970), .Z(n3972) );
  XNOR U4126 ( .A(n3971), .B(n3972), .Z(n3957) );
  XOR U4127 ( .A(n3958), .B(n3957), .Z(n3959) );
  XOR U4128 ( .A(n4065), .B(n3959), .Z(n3953) );
  ANDN U4129 ( .B(y[238]), .A(n54), .Z(n3825) );
  NAND U4130 ( .A(n3825), .B(n3962), .Z(n3829) );
  OR U4131 ( .A(n3827), .B(n3826), .Z(n3828) );
  NAND U4132 ( .A(n3829), .B(n3828), .Z(n3952) );
  NANDN U4133 ( .A(n56), .B(y[226]), .Z(n4027) );
  ANDN U4134 ( .B(y[229]), .A(n59), .Z(n4019) );
  NANDN U4135 ( .A(n4027), .B(n4019), .Z(n3833) );
  OR U4136 ( .A(n3831), .B(n3830), .Z(n3832) );
  NAND U4137 ( .A(n3833), .B(n3832), .Z(n3951) );
  XNOR U4138 ( .A(n3952), .B(n3951), .Z(n3954) );
  XNOR U4139 ( .A(n3953), .B(n3954), .Z(n3986) );
  NANDN U4140 ( .A(n3835), .B(n3834), .Z(n3839) );
  NAND U4141 ( .A(n3837), .B(n3836), .Z(n3838) );
  AND U4142 ( .A(n3839), .B(n3838), .Z(n3985) );
  XOR U4143 ( .A(n3986), .B(n3985), .Z(n3987) );
  XNOR U4144 ( .A(n3988), .B(n3987), .Z(n3991) );
  XNOR U4145 ( .A(n3992), .B(n3991), .Z(n3994) );
  OR U4146 ( .A(n3841), .B(n3840), .Z(n3845) );
  NANDN U4147 ( .A(n3843), .B(n3842), .Z(n3844) );
  NAND U4148 ( .A(n3845), .B(n3844), .Z(n3993) );
  XOR U4149 ( .A(n3994), .B(n3993), .Z(n3900) );
  OR U4150 ( .A(n3847), .B(n3846), .Z(n3851) );
  NANDN U4151 ( .A(n3849), .B(n3848), .Z(n3850) );
  NAND U4152 ( .A(n3851), .B(n3850), .Z(n4000) );
  OR U4153 ( .A(n3853), .B(n3852), .Z(n3857) );
  NANDN U4154 ( .A(n3855), .B(n3854), .Z(n3856) );
  NAND U4155 ( .A(n3857), .B(n3856), .Z(n3998) );
  OR U4156 ( .A(n3859), .B(n3858), .Z(n3863) );
  OR U4157 ( .A(n3861), .B(n3860), .Z(n3862) );
  NAND U4158 ( .A(n3863), .B(n3862), .Z(n3981) );
  NAND U4159 ( .A(n3864), .B(n4065), .Z(n3868) );
  OR U4160 ( .A(n3866), .B(n3865), .Z(n3867) );
  AND U4161 ( .A(n3868), .B(n3867), .Z(n3918) );
  NANDN U4162 ( .A(n53), .B(y[239]), .Z(n4538) );
  AND U4163 ( .A(y[232]), .B(x[65]), .Z(n4044) );
  NANDN U4164 ( .A(n4538), .B(n4044), .Z(n3872) );
  OR U4165 ( .A(n3870), .B(n3869), .Z(n3871) );
  AND U4166 ( .A(n3872), .B(n3871), .Z(n3919) );
  XOR U4167 ( .A(n3918), .B(n3919), .Z(n3920) );
  NANDN U4168 ( .A(n8890), .B(y[225]), .Z(n3924) );
  XOR U4169 ( .A(o[49]), .B(n3924), .Z(n3936) );
  ANDN U4170 ( .B(x[81]), .A(n5905), .Z(n3935) );
  XOR U4171 ( .A(n3936), .B(n3935), .Z(n3938) );
  IV U4172 ( .A(y[241]), .Z(n5874) );
  ANDN U4173 ( .B(x[64]), .A(n5874), .Z(n3937) );
  XOR U4174 ( .A(n3938), .B(n3937), .Z(n3915) );
  ANDN U4175 ( .B(x[66]), .A(n5936), .Z(n3874) );
  NANDN U4176 ( .A(n55), .B(y[231]), .Z(n3873) );
  XOR U4177 ( .A(n3874), .B(n3873), .Z(n3964) );
  ANDN U4178 ( .B(x[67]), .A(n5473), .Z(n3963) );
  XOR U4179 ( .A(n3964), .B(n3963), .Z(n3912) );
  NANDN U4180 ( .A(n3876), .B(n3875), .Z(n3880) );
  NAND U4181 ( .A(n3878), .B(n3877), .Z(n3879) );
  AND U4182 ( .A(n3880), .B(n3879), .Z(n3913) );
  XOR U4183 ( .A(n3915), .B(n3914), .Z(n3921) );
  XNOR U4184 ( .A(n3920), .B(n3921), .Z(n3980) );
  AND U4185 ( .A(y[235]), .B(x[77]), .Z(n4735) );
  IV U4186 ( .A(n4735), .Z(n4789) );
  ANDN U4187 ( .B(y[227]), .A(n50), .Z(n3881) );
  NANDN U4188 ( .A(n4789), .B(n3881), .Z(n3884) );
  OR U4189 ( .A(n3882), .B(n4543), .Z(n3883) );
  AND U4190 ( .A(n3884), .B(n3883), .Z(n3909) );
  AND U4191 ( .A(y[229]), .B(x[76]), .Z(n3947) );
  ANDN U4192 ( .B(x[78]), .A(n5714), .Z(n3945) );
  IV U4193 ( .A(n3945), .Z(n4020) );
  AND U4194 ( .A(y[226]), .B(x[79]), .Z(n3946) );
  XOR U4195 ( .A(n4020), .B(n3946), .Z(n3948) );
  XOR U4196 ( .A(n3947), .B(n3948), .Z(n3907) );
  NANDN U4197 ( .A(n3885), .B(o[48]), .Z(n3976) );
  ANDN U4198 ( .B(y[240]), .A(n46), .Z(n3887) );
  NANDN U4199 ( .A(n54), .B(y[232]), .Z(n3886) );
  XOR U4200 ( .A(n3887), .B(n3886), .Z(n3975) );
  XNOR U4201 ( .A(n3976), .B(n3975), .Z(n3906) );
  XOR U4202 ( .A(n3907), .B(n3906), .Z(n3908) );
  XOR U4203 ( .A(n3909), .B(n3908), .Z(n3979) );
  XOR U4204 ( .A(n3980), .B(n3979), .Z(n3982) );
  XOR U4205 ( .A(n3981), .B(n3982), .Z(n3997) );
  XNOR U4206 ( .A(n3998), .B(n3997), .Z(n3999) );
  XOR U4207 ( .A(n4000), .B(n3999), .Z(n3901) );
  XNOR U4208 ( .A(n3900), .B(n3901), .Z(n3903) );
  OR U4209 ( .A(n3889), .B(n3888), .Z(n3893) );
  NANDN U4210 ( .A(n3891), .B(n3890), .Z(n3892) );
  AND U4211 ( .A(n3893), .B(n3892), .Z(n3902) );
  XOR U4212 ( .A(n3903), .B(n3902), .Z(n3897) );
  XNOR U4213 ( .A(n3896), .B(n3897), .Z(N114) );
  NANDN U4214 ( .A(n3895), .B(n3894), .Z(n3899) );
  NAND U4215 ( .A(n3897), .B(n3896), .Z(n3898) );
  NAND U4216 ( .A(n3899), .B(n3898), .Z(n4003) );
  OR U4217 ( .A(n3901), .B(n3900), .Z(n3905) );
  OR U4218 ( .A(n3903), .B(n3902), .Z(n3904) );
  AND U4219 ( .A(n3905), .B(n3904), .Z(n4004) );
  XNOR U4220 ( .A(n4003), .B(n4004), .Z(n4005) );
  OR U4221 ( .A(n3907), .B(n3906), .Z(n3911) );
  NANDN U4222 ( .A(n3909), .B(n3908), .Z(n3910) );
  AND U4223 ( .A(n3911), .B(n3910), .Z(n4080) );
  OR U4224 ( .A(n3913), .B(n3912), .Z(n3917) );
  NANDN U4225 ( .A(n3915), .B(n3914), .Z(n3916) );
  AND U4226 ( .A(n3917), .B(n3916), .Z(n4081) );
  XOR U4227 ( .A(n4080), .B(n4081), .Z(n4082) );
  OR U4228 ( .A(n3919), .B(n3918), .Z(n3923) );
  NANDN U4229 ( .A(n3921), .B(n3920), .Z(n3922) );
  AND U4230 ( .A(n3923), .B(n3922), .Z(n4083) );
  XNOR U4231 ( .A(n4082), .B(n4083), .Z(n4112) );
  NANDN U4232 ( .A(n3924), .B(o[49]), .Z(n4046) );
  ANDN U4233 ( .B(x[65]), .A(n5874), .Z(n3926) );
  NANDN U4234 ( .A(n55), .B(y[232]), .Z(n3925) );
  XOR U4235 ( .A(n3926), .B(n3925), .Z(n4045) );
  ANDN U4236 ( .B(x[79]), .A(n5714), .Z(n3928) );
  NANDN U4237 ( .A(n59), .B(y[228]), .Z(n3927) );
  XNOR U4238 ( .A(n3928), .B(n3927), .Z(n4022) );
  XNOR U4239 ( .A(n4021), .B(n4022), .Z(n4033) );
  OR U4240 ( .A(n3930), .B(n3929), .Z(n3934) );
  OR U4241 ( .A(n3932), .B(n3931), .Z(n3933) );
  NAND U4242 ( .A(n3934), .B(n3933), .Z(n4032) );
  XNOR U4243 ( .A(n4033), .B(n4032), .Z(n4035) );
  XOR U4244 ( .A(n4034), .B(n4035), .Z(n4099) );
  NANDN U4245 ( .A(n3936), .B(n3935), .Z(n3940) );
  NANDN U4246 ( .A(n3938), .B(n3937), .Z(n3939) );
  NAND U4247 ( .A(n3940), .B(n3939), .Z(n4087) );
  ANDN U4248 ( .B(y[235]), .A(n52), .Z(n3942) );
  NANDN U4249 ( .A(n53), .B(y[234]), .Z(n3941) );
  XOR U4250 ( .A(n3942), .B(n3941), .Z(n4068) );
  NANDN U4251 ( .A(n5473), .B(x[68]), .Z(n4067) );
  XNOR U4252 ( .A(n4068), .B(n4067), .Z(n4015) );
  ANDN U4253 ( .B(x[69]), .A(n5332), .Z(n4189) );
  NANDN U4254 ( .A(n51), .B(y[236]), .Z(n4524) );
  XOR U4255 ( .A(n4189), .B(n4524), .Z(n4016) );
  XNOR U4256 ( .A(n4015), .B(n4016), .Z(n4086) );
  XOR U4257 ( .A(n4087), .B(n4086), .Z(n4089) );
  NANDN U4258 ( .A(n47), .B(y[240]), .Z(n4029) );
  ANDN U4259 ( .B(x[75]), .A(n44), .Z(n3944) );
  ANDN U4260 ( .B(y[226]), .A(n8890), .Z(n3943) );
  XNOR U4261 ( .A(n3944), .B(n3943), .Z(n4028) );
  XOR U4262 ( .A(n4029), .B(n4028), .Z(n4088) );
  XNOR U4263 ( .A(n4089), .B(n4088), .Z(n4098) );
  XOR U4264 ( .A(n4099), .B(n4098), .Z(n4101) );
  OR U4265 ( .A(n3946), .B(n3945), .Z(n3950) );
  OR U4266 ( .A(n3948), .B(n3947), .Z(n3949) );
  NAND U4267 ( .A(n3950), .B(n3949), .Z(n4100) );
  XOR U4268 ( .A(n4101), .B(n4100), .Z(n4111) );
  OR U4269 ( .A(n3952), .B(n3951), .Z(n3956) );
  NANDN U4270 ( .A(n3954), .B(n3953), .Z(n3955) );
  AND U4271 ( .A(n3956), .B(n3955), .Z(n4076) );
  NANDN U4272 ( .A(n3958), .B(n3957), .Z(n3961) );
  NANDN U4273 ( .A(n3959), .B(n4065), .Z(n3960) );
  NAND U4274 ( .A(n3961), .B(n3960), .Z(n4075) );
  ANDN U4275 ( .B(x[74]), .A(n5936), .Z(n4932) );
  NAND U4276 ( .A(n3962), .B(n4932), .Z(n3966) );
  NANDN U4277 ( .A(n3964), .B(n3963), .Z(n3965) );
  AND U4278 ( .A(n3966), .B(n3965), .Z(n4040) );
  NANDN U4279 ( .A(n45), .B(y[242]), .Z(n4050) );
  NANDN U4280 ( .A(n5905), .B(x[82]), .Z(n4049) );
  XOR U4281 ( .A(n4050), .B(n4049), .Z(n4051) );
  NANDN U4282 ( .A(n8626), .B(y[225]), .Z(n4071) );
  XOR U4283 ( .A(o[50]), .B(n4071), .Z(n4052) );
  XOR U4284 ( .A(n4051), .B(n4052), .Z(n4039) );
  AND U4285 ( .A(y[230]), .B(x[76]), .Z(n4143) );
  ANDN U4286 ( .B(x[67]), .A(n5936), .Z(n3968) );
  NANDN U4287 ( .A(n58), .B(y[229]), .Z(n3967) );
  XOR U4288 ( .A(n3968), .B(n3967), .Z(n4058) );
  XOR U4289 ( .A(n4143), .B(n4058), .Z(n4038) );
  XNOR U4290 ( .A(n4039), .B(n4038), .Z(n4041) );
  XOR U4291 ( .A(n4040), .B(n4041), .Z(n4092) );
  OR U4292 ( .A(n3970), .B(n3969), .Z(n3974) );
  OR U4293 ( .A(n3972), .B(n3971), .Z(n3973) );
  AND U4294 ( .A(n3974), .B(n3973), .Z(n4093) );
  XNOR U4295 ( .A(n4092), .B(n4093), .Z(n4095) );
  NANDN U4296 ( .A(n54), .B(y[240]), .Z(n4931) );
  NANDN U4297 ( .A(n4931), .B(n4044), .Z(n3978) );
  OR U4298 ( .A(n3976), .B(n3975), .Z(n3977) );
  NAND U4299 ( .A(n3978), .B(n3977), .Z(n4094) );
  XNOR U4300 ( .A(n4095), .B(n4094), .Z(n4074) );
  XNOR U4301 ( .A(n4075), .B(n4074), .Z(n4077) );
  XOR U4302 ( .A(n4076), .B(n4077), .Z(n4110) );
  XOR U4303 ( .A(n4111), .B(n4110), .Z(n4113) );
  XNOR U4304 ( .A(n4112), .B(n4113), .Z(n4107) );
  NANDN U4305 ( .A(n3980), .B(n3979), .Z(n3984) );
  OR U4306 ( .A(n3982), .B(n3981), .Z(n3983) );
  AND U4307 ( .A(n3984), .B(n3983), .Z(n4104) );
  OR U4308 ( .A(n3986), .B(n3985), .Z(n3990) );
  NAND U4309 ( .A(n3988), .B(n3987), .Z(n3989) );
  NAND U4310 ( .A(n3990), .B(n3989), .Z(n4105) );
  XOR U4311 ( .A(n4107), .B(n4106), .Z(n4012) );
  OR U4312 ( .A(n3992), .B(n3991), .Z(n3996) );
  OR U4313 ( .A(n3994), .B(n3993), .Z(n3995) );
  NAND U4314 ( .A(n3996), .B(n3995), .Z(n4010) );
  OR U4315 ( .A(n3998), .B(n3997), .Z(n4002) );
  OR U4316 ( .A(n4000), .B(n3999), .Z(n4001) );
  NAND U4317 ( .A(n4002), .B(n4001), .Z(n4009) );
  XNOR U4318 ( .A(n4010), .B(n4009), .Z(n4011) );
  XNOR U4319 ( .A(n4012), .B(n4011), .Z(n4006) );
  XOR U4320 ( .A(n4005), .B(n4006), .Z(N115) );
  NANDN U4321 ( .A(n4004), .B(n4003), .Z(n4008) );
  NANDN U4322 ( .A(n4006), .B(n4005), .Z(n4007) );
  NAND U4323 ( .A(n4008), .B(n4007), .Z(n4225) );
  OR U4324 ( .A(n4010), .B(n4009), .Z(n4014) );
  OR U4325 ( .A(n4012), .B(n4011), .Z(n4013) );
  AND U4326 ( .A(n4014), .B(n4013), .Z(n4226) );
  XNOR U4327 ( .A(n4225), .B(n4226), .Z(n4227) );
  NANDN U4328 ( .A(n4189), .B(n4524), .Z(n4018) );
  NANDN U4329 ( .A(n4016), .B(n4015), .Z(n4017) );
  AND U4330 ( .A(n4018), .B(n4017), .Z(n4221) );
  XOR U4331 ( .A(n4019), .B(n4066), .Z(n4199) );
  NANDN U4332 ( .A(n46), .B(y[242]), .Z(n4198) );
  XOR U4333 ( .A(n4199), .B(n4198), .Z(n4165) );
  AND U4334 ( .A(y[228]), .B(x[79]), .Z(n4135) );
  NANDN U4335 ( .A(n4020), .B(n4135), .Z(n4024) );
  NAND U4336 ( .A(n4022), .B(n4021), .Z(n4023) );
  NAND U4337 ( .A(n4024), .B(n4023), .Z(n4163) );
  NANDN U4338 ( .A(n47), .B(y[241]), .Z(n4146) );
  ANDN U4339 ( .B(x[76]), .A(n44), .Z(n4026) );
  NANDN U4340 ( .A(n58), .B(y[230]), .Z(n4025) );
  XOR U4341 ( .A(n4026), .B(n4025), .Z(n4145) );
  XOR U4342 ( .A(n4163), .B(n4164), .Z(n4166) );
  XNOR U4343 ( .A(n4165), .B(n4166), .Z(n4219) );
  ANDN U4344 ( .B(y[231]), .A(n8890), .Z(n4536) );
  NANDN U4345 ( .A(n4027), .B(n4536), .Z(n4031) );
  OR U4346 ( .A(n4029), .B(n4028), .Z(n4030) );
  NAND U4347 ( .A(n4031), .B(n4030), .Z(n4220) );
  XNOR U4348 ( .A(n4219), .B(n4220), .Z(n4222) );
  XOR U4349 ( .A(n4221), .B(n4222), .Z(n4128) );
  OR U4350 ( .A(n4033), .B(n4032), .Z(n4037) );
  NANDN U4351 ( .A(n4035), .B(n4034), .Z(n4036) );
  NAND U4352 ( .A(n4037), .B(n4036), .Z(n4214) );
  OR U4353 ( .A(n4039), .B(n4038), .Z(n4043) );
  OR U4354 ( .A(n4041), .B(n4040), .Z(n4042) );
  NAND U4355 ( .A(n4043), .B(n4042), .Z(n4213) );
  XOR U4356 ( .A(n4214), .B(n4213), .Z(n4215) );
  ANDN U4357 ( .B(x[74]), .A(n5874), .Z(n5333) );
  NAND U4358 ( .A(n4044), .B(n5333), .Z(n4048) );
  OR U4359 ( .A(n4046), .B(n4045), .Z(n4047) );
  NAND U4360 ( .A(n4048), .B(n4047), .Z(n4178) );
  OR U4361 ( .A(n4050), .B(n4049), .Z(n4054) );
  NANDN U4362 ( .A(n4052), .B(n4051), .Z(n4053) );
  AND U4363 ( .A(n4054), .B(n4053), .Z(n4175) );
  ANDN U4364 ( .B(x[80]), .A(n5714), .Z(n4056) );
  NANDN U4365 ( .A(n54), .B(y[234]), .Z(n4055) );
  XNOR U4366 ( .A(n4056), .B(n4055), .Z(n4136) );
  XNOR U4367 ( .A(n4135), .B(n4136), .Z(n4176) );
  XOR U4368 ( .A(n4178), .B(n4177), .Z(n4209) );
  ANDN U4369 ( .B(x[77]), .A(n5936), .Z(n5433) );
  IV U4370 ( .A(n5433), .Z(n5277) );
  NANDN U4371 ( .A(n5277), .B(n4057), .Z(n4060) );
  NANDN U4372 ( .A(n4058), .B(n4143), .Z(n4059) );
  NAND U4373 ( .A(n4060), .B(n4059), .Z(n4172) );
  ANDN U4374 ( .B(x[75]), .A(n5947), .Z(n4062) );
  NANDN U4375 ( .A(n52), .B(y[236]), .Z(n4061) );
  XOR U4376 ( .A(n4062), .B(n4061), .Z(n4151) );
  NANDN U4377 ( .A(n48), .B(y[240]), .Z(n4150) );
  XNOR U4378 ( .A(n4151), .B(n4150), .Z(n4170) );
  ANDN U4379 ( .B(y[225]), .A(n61), .Z(n4156) );
  XNOR U4380 ( .A(o[51]), .B(n4156), .Z(n4204) );
  ANDN U4381 ( .B(x[74]), .A(n5637), .Z(n4064) );
  NANDN U4382 ( .A(n8626), .B(y[226]), .Z(n4063) );
  XOR U4383 ( .A(n4064), .B(n4063), .Z(n4203) );
  XOR U4384 ( .A(n4204), .B(n4203), .Z(n4169) );
  XOR U4385 ( .A(n4172), .B(n4171), .Z(n4207) );
  NANDN U4386 ( .A(n4066), .B(n4065), .Z(n4070) );
  OR U4387 ( .A(n4068), .B(n4067), .Z(n4069) );
  NAND U4388 ( .A(n4070), .B(n4069), .Z(n4160) );
  NANDN U4389 ( .A(n4071), .B(o[50]), .Z(n4184) );
  NANDN U4390 ( .A(n45), .B(y[243]), .Z(n4182) );
  NANDN U4391 ( .A(n5905), .B(x[83]), .Z(n4181) );
  XOR U4392 ( .A(n4182), .B(n4181), .Z(n4183) );
  XOR U4393 ( .A(n4184), .B(n4183), .Z(n4158) );
  NANDN U4394 ( .A(n49), .B(y[239]), .Z(n4313) );
  ANDN U4395 ( .B(x[70]), .A(n5332), .Z(n4073) );
  NANDN U4396 ( .A(n50), .B(y[238]), .Z(n4072) );
  XOR U4397 ( .A(n4073), .B(n4072), .Z(n4190) );
  XNOR U4398 ( .A(n4158), .B(n4157), .Z(n4159) );
  XOR U4399 ( .A(n4160), .B(n4159), .Z(n4208) );
  XNOR U4400 ( .A(n4207), .B(n4208), .Z(n4210) );
  XNOR U4401 ( .A(n4209), .B(n4210), .Z(n4216) );
  XNOR U4402 ( .A(n4215), .B(n4216), .Z(n4129) );
  XNOR U4403 ( .A(n4128), .B(n4129), .Z(n4131) );
  OR U4404 ( .A(n4075), .B(n4074), .Z(n4079) );
  OR U4405 ( .A(n4077), .B(n4076), .Z(n4078) );
  NAND U4406 ( .A(n4079), .B(n4078), .Z(n4130) );
  XOR U4407 ( .A(n4131), .B(n4130), .Z(n4125) );
  OR U4408 ( .A(n4081), .B(n4080), .Z(n4085) );
  NANDN U4409 ( .A(n4083), .B(n4082), .Z(n4084) );
  NAND U4410 ( .A(n4085), .B(n4084), .Z(n4123) );
  NANDN U4411 ( .A(n4087), .B(n4086), .Z(n4091) );
  OR U4412 ( .A(n4089), .B(n4088), .Z(n4090) );
  AND U4413 ( .A(n4091), .B(n4090), .Z(n4119) );
  OR U4414 ( .A(n4093), .B(n4092), .Z(n4097) );
  OR U4415 ( .A(n4095), .B(n4094), .Z(n4096) );
  AND U4416 ( .A(n4097), .B(n4096), .Z(n4116) );
  NANDN U4417 ( .A(n4099), .B(n4098), .Z(n4103) );
  OR U4418 ( .A(n4101), .B(n4100), .Z(n4102) );
  NAND U4419 ( .A(n4103), .B(n4102), .Z(n4117) );
  XNOR U4420 ( .A(n4116), .B(n4117), .Z(n4118) );
  XOR U4421 ( .A(n4123), .B(n4122), .Z(n4124) );
  XNOR U4422 ( .A(n4125), .B(n4124), .Z(n4234) );
  OR U4423 ( .A(n4105), .B(n4104), .Z(n4109) );
  NANDN U4424 ( .A(n4107), .B(n4106), .Z(n4108) );
  NAND U4425 ( .A(n4109), .B(n4108), .Z(n4232) );
  NANDN U4426 ( .A(n4111), .B(n4110), .Z(n4115) );
  OR U4427 ( .A(n4113), .B(n4112), .Z(n4114) );
  NAND U4428 ( .A(n4115), .B(n4114), .Z(n4231) );
  XNOR U4429 ( .A(n4234), .B(n4233), .Z(n4228) );
  XOR U4430 ( .A(n4227), .B(n4228), .Z(N116) );
  OR U4431 ( .A(n4117), .B(n4116), .Z(n4121) );
  OR U4432 ( .A(n4119), .B(n4118), .Z(n4120) );
  AND U4433 ( .A(n4121), .B(n4120), .Z(n4351) );
  OR U4434 ( .A(n4123), .B(n4122), .Z(n4127) );
  NANDN U4435 ( .A(n4125), .B(n4124), .Z(n4126) );
  AND U4436 ( .A(n4127), .B(n4126), .Z(n4350) );
  OR U4437 ( .A(n4129), .B(n4128), .Z(n4133) );
  OR U4438 ( .A(n4131), .B(n4130), .Z(n4132) );
  AND U4439 ( .A(n4133), .B(n4132), .Z(n4334) );
  ANDN U4440 ( .B(x[80]), .A(n5196), .Z(n5015) );
  IV U4441 ( .A(n5015), .Z(n5089) );
  ANDN U4442 ( .B(y[227]), .A(n54), .Z(n4134) );
  NANDN U4443 ( .A(n5089), .B(n4134), .Z(n4138) );
  NAND U4444 ( .A(n4136), .B(n4135), .Z(n4137) );
  AND U4445 ( .A(n4138), .B(n4137), .Z(n4283) );
  ANDN U4446 ( .B(y[229]), .A(n60), .Z(n4140) );
  NANDN U4447 ( .A(n54), .B(y[235]), .Z(n4139) );
  XOR U4448 ( .A(n4140), .B(n4139), .Z(n4262) );
  ANDN U4449 ( .B(x[78]), .A(n5663), .Z(n4261) );
  XOR U4450 ( .A(n4262), .B(n4261), .Z(n4296) );
  NANDN U4451 ( .A(n47), .B(y[242]), .Z(n4328) );
  ANDN U4452 ( .B(y[228]), .A(n8890), .Z(n4142) );
  ANDN U4453 ( .B(x[74]), .A(n5196), .Z(n4141) );
  XNOR U4454 ( .A(n4142), .B(n4141), .Z(n4327) );
  XOR U4455 ( .A(n4328), .B(n4327), .Z(n4295) );
  ANDN U4456 ( .B(y[231]), .A(n58), .Z(n4144) );
  NAND U4457 ( .A(n4144), .B(n4143), .Z(n4148) );
  OR U4458 ( .A(n4146), .B(n4145), .Z(n4147) );
  NAND U4459 ( .A(n4148), .B(n4147), .Z(n4298) );
  XNOR U4460 ( .A(n4297), .B(n4298), .Z(n4284) );
  AND U4461 ( .A(y[236]), .B(x[75]), .Z(n4738) );
  NAND U4462 ( .A(n4738), .B(n4149), .Z(n4153) );
  OR U4463 ( .A(n4151), .B(n4150), .Z(n4152) );
  AND U4464 ( .A(n4153), .B(n4152), .Z(n4304) );
  ANDN U4465 ( .B(x[75]), .A(n5637), .Z(n4155) );
  NANDN U4466 ( .A(n46), .B(y[243]), .Z(n4154) );
  XOR U4467 ( .A(n4155), .B(n4154), .Z(n4268) );
  NANDN U4468 ( .A(n8824), .B(y[225]), .Z(n4265) );
  XNOR U4469 ( .A(n4265), .B(o[52]), .Z(n4267) );
  XOR U4470 ( .A(n4268), .B(n4267), .Z(n4302) );
  NAND U4471 ( .A(o[51]), .B(n4156), .Z(n4310) );
  NANDN U4472 ( .A(n8885), .B(y[224]), .Z(n4308) );
  NANDN U4473 ( .A(n45), .B(y[244]), .Z(n4307) );
  XNOR U4474 ( .A(n4308), .B(n4307), .Z(n4309) );
  XNOR U4475 ( .A(n4310), .B(n4309), .Z(n4301) );
  XNOR U4476 ( .A(n4302), .B(n4301), .Z(n4303) );
  XOR U4477 ( .A(n4304), .B(n4303), .Z(n4285) );
  NANDN U4478 ( .A(n4158), .B(n4157), .Z(n4162) );
  NAND U4479 ( .A(n4160), .B(n4159), .Z(n4161) );
  AND U4480 ( .A(n4162), .B(n4161), .Z(n4237) );
  NANDN U4481 ( .A(n4164), .B(n4163), .Z(n4168) );
  NANDN U4482 ( .A(n4166), .B(n4165), .Z(n4167) );
  AND U4483 ( .A(n4168), .B(n4167), .Z(n4238) );
  XOR U4484 ( .A(n4239), .B(n4240), .Z(n4280) );
  NANDN U4485 ( .A(n4170), .B(n4169), .Z(n4174) );
  NAND U4486 ( .A(n4172), .B(n4171), .Z(n4173) );
  NAND U4487 ( .A(n4174), .B(n4173), .Z(n4278) );
  OR U4488 ( .A(n4176), .B(n4175), .Z(n4180) );
  NAND U4489 ( .A(n4178), .B(n4177), .Z(n4179) );
  NAND U4490 ( .A(n4180), .B(n4179), .Z(n4246) );
  OR U4491 ( .A(n4182), .B(n4181), .Z(n4186) );
  NANDN U4492 ( .A(n4184), .B(n4183), .Z(n4185) );
  AND U4493 ( .A(n4186), .B(n4185), .Z(n4251) );
  NANDN U4494 ( .A(n8626), .B(y[227]), .Z(n4257) );
  ANDN U4495 ( .B(x[76]), .A(n5947), .Z(n4188) );
  NANDN U4496 ( .A(n61), .B(y[226]), .Z(n4187) );
  XNOR U4497 ( .A(n4188), .B(n4187), .Z(n4256) );
  XNOR U4498 ( .A(n4257), .B(n4256), .Z(n4249) );
  AND U4499 ( .A(y[238]), .B(x[70]), .Z(n4271) );
  NAND U4500 ( .A(n4271), .B(n4189), .Z(n4192) );
  OR U4501 ( .A(n4313), .B(n4190), .Z(n4191) );
  AND U4502 ( .A(n4192), .B(n4191), .Z(n4250) );
  XOR U4503 ( .A(n4249), .B(n4250), .Z(n4252) );
  NANDN U4504 ( .A(n52), .B(y[237]), .Z(n4315) );
  ANDN U4505 ( .B(x[69]), .A(n5936), .Z(n4194) );
  NANDN U4506 ( .A(n49), .B(y[240]), .Z(n4193) );
  XOR U4507 ( .A(n4194), .B(n4193), .Z(n4314) );
  XNOR U4508 ( .A(n4315), .B(n4314), .Z(n4272) );
  XOR U4509 ( .A(n4271), .B(n4272), .Z(n4274) );
  NANDN U4510 ( .A(n53), .B(y[236]), .Z(n4323) );
  ANDN U4511 ( .B(y[241]), .A(n48), .Z(n4196) );
  ANDN U4512 ( .B(x[77]), .A(n44), .Z(n4195) );
  XNOR U4513 ( .A(n4196), .B(n4195), .Z(n4322) );
  XOR U4514 ( .A(n4323), .B(n4322), .Z(n4273) );
  XNOR U4515 ( .A(n4274), .B(n4273), .Z(n4292) );
  AND U4516 ( .A(y[235]), .B(x[78]), .Z(n4820) );
  IV U4517 ( .A(n4820), .Z(n4985) );
  NANDN U4518 ( .A(n4985), .B(n4197), .Z(n4201) );
  OR U4519 ( .A(n4199), .B(n4198), .Z(n4200) );
  NAND U4520 ( .A(n4201), .B(n4200), .Z(n4290) );
  ANDN U4521 ( .B(x[81]), .A(n5637), .Z(n5104) );
  NANDN U4522 ( .A(n4202), .B(n5104), .Z(n4206) );
  OR U4523 ( .A(n4204), .B(n4203), .Z(n4205) );
  NAND U4524 ( .A(n4206), .B(n4205), .Z(n4289) );
  XOR U4525 ( .A(n4292), .B(n4291), .Z(n4244) );
  XNOR U4526 ( .A(n4243), .B(n4244), .Z(n4245) );
  XNOR U4527 ( .A(n4246), .B(n4245), .Z(n4277) );
  XOR U4528 ( .A(n4278), .B(n4277), .Z(n4279) );
  XNOR U4529 ( .A(n4280), .B(n4279), .Z(n4332) );
  OR U4530 ( .A(n4208), .B(n4207), .Z(n4212) );
  OR U4531 ( .A(n4210), .B(n4209), .Z(n4211) );
  NAND U4532 ( .A(n4212), .B(n4211), .Z(n4338) );
  OR U4533 ( .A(n4214), .B(n4213), .Z(n4218) );
  NANDN U4534 ( .A(n4216), .B(n4215), .Z(n4217) );
  NAND U4535 ( .A(n4218), .B(n4217), .Z(n4337) );
  XNOR U4536 ( .A(n4338), .B(n4337), .Z(n4339) );
  OR U4537 ( .A(n4220), .B(n4219), .Z(n4224) );
  OR U4538 ( .A(n4222), .B(n4221), .Z(n4223) );
  NAND U4539 ( .A(n4224), .B(n4223), .Z(n4340) );
  XOR U4540 ( .A(n4332), .B(n4331), .Z(n4333) );
  XNOR U4541 ( .A(n4334), .B(n4333), .Z(n4349) );
  XOR U4542 ( .A(n4351), .B(n4352), .Z(n4345) );
  NANDN U4543 ( .A(n4226), .B(n4225), .Z(n4230) );
  NANDN U4544 ( .A(n4228), .B(n4227), .Z(n4229) );
  NAND U4545 ( .A(n4230), .B(n4229), .Z(n4343) );
  OR U4546 ( .A(n4232), .B(n4231), .Z(n4236) );
  NANDN U4547 ( .A(n4234), .B(n4233), .Z(n4235) );
  NAND U4548 ( .A(n4236), .B(n4235), .Z(n4344) );
  XNOR U4549 ( .A(n4343), .B(n4344), .Z(n4346) );
  XNOR U4550 ( .A(n4345), .B(n4346), .Z(N117) );
  OR U4551 ( .A(n4238), .B(n4237), .Z(n4242) );
  NAND U4552 ( .A(n4240), .B(n4239), .Z(n4241) );
  NAND U4553 ( .A(n4242), .B(n4241), .Z(n4484) );
  NANDN U4554 ( .A(n4244), .B(n4243), .Z(n4248) );
  NANDN U4555 ( .A(n4246), .B(n4245), .Z(n4247) );
  AND U4556 ( .A(n4248), .B(n4247), .Z(n4481) );
  NANDN U4557 ( .A(n4250), .B(n4249), .Z(n4254) );
  OR U4558 ( .A(n4252), .B(n4251), .Z(n4253) );
  NAND U4559 ( .A(n4254), .B(n4253), .Z(n4406) );
  ANDN U4560 ( .B(x[82]), .A(n5947), .Z(n5003) );
  IV U4561 ( .A(n5003), .Z(n5101) );
  NANDN U4562 ( .A(n5101), .B(n4255), .Z(n4259) );
  NANDN U4563 ( .A(n4257), .B(n4256), .Z(n4258) );
  AND U4564 ( .A(n4259), .B(n4258), .Z(n4385) );
  AND U4565 ( .A(y[240]), .B(x[69]), .Z(n4444) );
  ANDN U4566 ( .B(y[229]), .A(n8890), .Z(n4443) );
  XOR U4567 ( .A(n4444), .B(n4443), .Z(n4446) );
  AND U4568 ( .A(y[230]), .B(x[79]), .Z(n4445) );
  XOR U4569 ( .A(n4446), .B(n4445), .Z(n4475) );
  ANDN U4570 ( .B(y[229]), .A(n54), .Z(n4260) );
  ANDN U4571 ( .B(y[235]), .A(n60), .Z(n5095) );
  NAND U4572 ( .A(n4260), .B(n5095), .Z(n4264) );
  NANDN U4573 ( .A(n4262), .B(n4261), .Z(n4263) );
  NAND U4574 ( .A(n4264), .B(n4263), .Z(n4476) );
  XNOR U4575 ( .A(n4475), .B(n4476), .Z(n4478) );
  AND U4576 ( .A(y[245]), .B(x[64]), .Z(n4459) );
  ANDN U4577 ( .B(o[52]), .A(n4265), .Z(n4457) );
  AND U4578 ( .A(y[224]), .B(x[85]), .Z(n4458) );
  XNOR U4579 ( .A(n4457), .B(n4458), .Z(n4460) );
  XNOR U4580 ( .A(n4459), .B(n4460), .Z(n4477) );
  XOR U4581 ( .A(n4478), .B(n4477), .Z(n4386) );
  ANDN U4582 ( .B(y[243]), .A(n56), .Z(n5848) );
  NAND U4583 ( .A(n5848), .B(n4266), .Z(n4270) );
  NANDN U4584 ( .A(n4268), .B(n4267), .Z(n4269) );
  NAND U4585 ( .A(n4270), .B(n4269), .Z(n4388) );
  XNOR U4586 ( .A(n4387), .B(n4388), .Z(n4404) );
  NANDN U4587 ( .A(n4272), .B(n4271), .Z(n4276) );
  NANDN U4588 ( .A(n4274), .B(n4273), .Z(n4275) );
  AND U4589 ( .A(n4276), .B(n4275), .Z(n4403) );
  XOR U4590 ( .A(n4406), .B(n4405), .Z(n4482) );
  XOR U4591 ( .A(n4484), .B(n4483), .Z(n4370) );
  NANDN U4592 ( .A(n4278), .B(n4277), .Z(n4282) );
  OR U4593 ( .A(n4280), .B(n4279), .Z(n4281) );
  AND U4594 ( .A(n4282), .B(n4281), .Z(n4367) );
  OR U4595 ( .A(n4284), .B(n4283), .Z(n4288) );
  NANDN U4596 ( .A(n4286), .B(n4285), .Z(n4287) );
  NAND U4597 ( .A(n4288), .B(n4287), .Z(n4376) );
  OR U4598 ( .A(n4290), .B(n4289), .Z(n4294) );
  NANDN U4599 ( .A(n4292), .B(n4291), .Z(n4293) );
  AND U4600 ( .A(n4294), .B(n4293), .Z(n4379) );
  NANDN U4601 ( .A(n4296), .B(n4295), .Z(n4300) );
  NAND U4602 ( .A(n4298), .B(n4297), .Z(n4299) );
  NAND U4603 ( .A(n4300), .B(n4299), .Z(n4380) );
  XNOR U4604 ( .A(n4379), .B(n4380), .Z(n4381) );
  OR U4605 ( .A(n4302), .B(n4301), .Z(n4306) );
  OR U4606 ( .A(n4304), .B(n4303), .Z(n4305) );
  NAND U4607 ( .A(n4306), .B(n4305), .Z(n4382) );
  OR U4608 ( .A(n4308), .B(n4307), .Z(n4312) );
  OR U4609 ( .A(n4310), .B(n4309), .Z(n4311) );
  AND U4610 ( .A(n4312), .B(n4311), .Z(n4391) );
  NANDN U4611 ( .A(n4313), .B(n4444), .Z(n4317) );
  OR U4612 ( .A(n4315), .B(n4314), .Z(n4316) );
  AND U4613 ( .A(n4317), .B(n4316), .Z(n4392) );
  XNOR U4614 ( .A(n4391), .B(n4392), .Z(n4393) );
  NANDN U4615 ( .A(n49), .B(y[241]), .Z(n4438) );
  ANDN U4616 ( .B(y[242]), .A(n48), .Z(n4319) );
  ANDN U4617 ( .B(x[77]), .A(n5947), .Z(n4318) );
  XNOR U4618 ( .A(n4319), .B(n4318), .Z(n4437) );
  XOR U4619 ( .A(n4438), .B(n4437), .Z(n4469) );
  AND U4620 ( .A(y[233]), .B(x[76]), .Z(n4423) );
  AND U4621 ( .A(y[243]), .B(x[66]), .Z(n4421) );
  AND U4622 ( .A(y[228]), .B(x[81]), .Z(n4422) );
  XNOR U4623 ( .A(n4421), .B(n4422), .Z(n4424) );
  XOR U4624 ( .A(n4423), .B(n4424), .Z(n4470) );
  XOR U4625 ( .A(n4469), .B(n4470), .Z(n4472) );
  AND U4626 ( .A(y[239]), .B(x[70]), .Z(n4451) );
  ANDN U4627 ( .B(x[71]), .A(n5473), .Z(n4449) );
  IV U4628 ( .A(n4449), .Z(n4537) );
  AND U4629 ( .A(y[231]), .B(x[78]), .Z(n4450) );
  XOR U4630 ( .A(n4537), .B(n4450), .Z(n4452) );
  XNOR U4631 ( .A(n4451), .B(n4452), .Z(n4418) );
  AND U4632 ( .A(y[237]), .B(x[72]), .Z(n4416) );
  XNOR U4633 ( .A(n4415), .B(n4416), .Z(n4417) );
  XOR U4634 ( .A(n4418), .B(n4417), .Z(n4471) );
  XNOR U4635 ( .A(n4472), .B(n4471), .Z(n4394) );
  ANDN U4636 ( .B(y[241]), .A(n58), .Z(n4321) );
  NAND U4637 ( .A(n4321), .B(n4320), .Z(n4325) );
  OR U4638 ( .A(n4323), .B(n4322), .Z(n4324) );
  AND U4639 ( .A(n4325), .B(n4324), .Z(n4399) );
  AND U4640 ( .A(y[244]), .B(x[65]), .Z(n4463) );
  AND U4641 ( .A(y[227]), .B(x[82]), .Z(n4464) );
  XNOR U4642 ( .A(n4463), .B(n4464), .Z(n4466) );
  XNOR U4643 ( .A(n4465), .B(n4466), .Z(n4397) );
  NANDN U4644 ( .A(n56), .B(y[234]), .Z(n4432) );
  ANDN U4645 ( .B(y[225]), .A(n8885), .Z(n4435) );
  XNOR U4646 ( .A(o[53]), .B(n4435), .Z(n4430) );
  NANDN U4647 ( .A(n8824), .B(y[226]), .Z(n4429) );
  XOR U4648 ( .A(n4430), .B(n4429), .Z(n4431) );
  XOR U4649 ( .A(n4432), .B(n4431), .Z(n4398) );
  XOR U4650 ( .A(n4397), .B(n4398), .Z(n4400) );
  XOR U4651 ( .A(n4399), .B(n4400), .Z(n4409) );
  NANDN U4652 ( .A(n5089), .B(n4326), .Z(n4330) );
  OR U4653 ( .A(n4328), .B(n4327), .Z(n4329) );
  NAND U4654 ( .A(n4330), .B(n4329), .Z(n4410) );
  XNOR U4655 ( .A(n4409), .B(n4410), .Z(n4412) );
  XOR U4656 ( .A(n4411), .B(n4412), .Z(n4373) );
  XNOR U4657 ( .A(n4374), .B(n4373), .Z(n4375) );
  XOR U4658 ( .A(n4376), .B(n4375), .Z(n4368) );
  XOR U4659 ( .A(n4367), .B(n4368), .Z(n4369) );
  XNOR U4660 ( .A(n4370), .B(n4369), .Z(n4363) );
  NAND U4661 ( .A(n4332), .B(n4331), .Z(n4336) );
  NANDN U4662 ( .A(n4334), .B(n4333), .Z(n4335) );
  NAND U4663 ( .A(n4336), .B(n4335), .Z(n4362) );
  OR U4664 ( .A(n4338), .B(n4337), .Z(n4342) );
  OR U4665 ( .A(n4340), .B(n4339), .Z(n4341) );
  NAND U4666 ( .A(n4342), .B(n4341), .Z(n4361) );
  XNOR U4667 ( .A(n4362), .B(n4361), .Z(n4364) );
  XOR U4668 ( .A(n4363), .B(n4364), .Z(n4358) );
  NANDN U4669 ( .A(n4344), .B(n4343), .Z(n4348) );
  NAND U4670 ( .A(n4346), .B(n4345), .Z(n4347) );
  NAND U4671 ( .A(n4348), .B(n4347), .Z(n4355) );
  OR U4672 ( .A(n4350), .B(n4349), .Z(n4354) );
  OR U4673 ( .A(n4352), .B(n4351), .Z(n4353) );
  AND U4674 ( .A(n4354), .B(n4353), .Z(n4356) );
  XNOR U4675 ( .A(n4355), .B(n4356), .Z(n4357) );
  XOR U4676 ( .A(n4358), .B(n4357), .Z(N118) );
  NANDN U4677 ( .A(n4356), .B(n4355), .Z(n4360) );
  NANDN U4678 ( .A(n4358), .B(n4357), .Z(n4359) );
  NAND U4679 ( .A(n4360), .B(n4359), .Z(n4487) );
  OR U4680 ( .A(n4362), .B(n4361), .Z(n4366) );
  NANDN U4681 ( .A(n4364), .B(n4363), .Z(n4365) );
  AND U4682 ( .A(n4366), .B(n4365), .Z(n4488) );
  XNOR U4683 ( .A(n4487), .B(n4488), .Z(n4489) );
  OR U4684 ( .A(n4368), .B(n4367), .Z(n4372) );
  NANDN U4685 ( .A(n4370), .B(n4369), .Z(n4371) );
  NAND U4686 ( .A(n4372), .B(n4371), .Z(n4496) );
  NANDN U4687 ( .A(n4374), .B(n4373), .Z(n4378) );
  NANDN U4688 ( .A(n4376), .B(n4375), .Z(n4377) );
  NAND U4689 ( .A(n4378), .B(n4377), .Z(n4506) );
  OR U4690 ( .A(n4380), .B(n4379), .Z(n4384) );
  OR U4691 ( .A(n4382), .B(n4381), .Z(n4383) );
  NAND U4692 ( .A(n4384), .B(n4383), .Z(n4505) );
  XOR U4693 ( .A(n4506), .B(n4505), .Z(n4508) );
  OR U4694 ( .A(n4386), .B(n4385), .Z(n4390) );
  NAND U4695 ( .A(n4388), .B(n4387), .Z(n4389) );
  AND U4696 ( .A(n4390), .B(n4389), .Z(n4514) );
  OR U4697 ( .A(n4392), .B(n4391), .Z(n4396) );
  OR U4698 ( .A(n4394), .B(n4393), .Z(n4395) );
  AND U4699 ( .A(n4396), .B(n4395), .Z(n4511) );
  NANDN U4700 ( .A(n4398), .B(n4397), .Z(n4402) );
  OR U4701 ( .A(n4400), .B(n4399), .Z(n4401) );
  AND U4702 ( .A(n4402), .B(n4401), .Z(n4512) );
  XOR U4703 ( .A(n4511), .B(n4512), .Z(n4513) );
  XNOR U4704 ( .A(n4514), .B(n4513), .Z(n4499) );
  OR U4705 ( .A(n4404), .B(n4403), .Z(n4408) );
  NAND U4706 ( .A(n4406), .B(n4405), .Z(n4407) );
  NAND U4707 ( .A(n4408), .B(n4407), .Z(n4500) );
  XNOR U4708 ( .A(n4499), .B(n4500), .Z(n4502) );
  OR U4709 ( .A(n4410), .B(n4409), .Z(n4414) );
  OR U4710 ( .A(n4412), .B(n4411), .Z(n4413) );
  NAND U4711 ( .A(n4414), .B(n4413), .Z(n4601) );
  OR U4712 ( .A(n4416), .B(n4415), .Z(n4420) );
  OR U4713 ( .A(n4418), .B(n4417), .Z(n4419) );
  AND U4714 ( .A(n4420), .B(n4419), .Z(n4618) );
  OR U4715 ( .A(n4422), .B(n4421), .Z(n4426) );
  OR U4716 ( .A(n4424), .B(n4423), .Z(n4425) );
  NAND U4717 ( .A(n4426), .B(n4425), .Z(n4581) );
  NANDN U4718 ( .A(n49), .B(y[242]), .Z(n4545) );
  ANDN U4719 ( .B(x[76]), .A(n5196), .Z(n4428) );
  ANDN U4720 ( .B(y[228]), .A(n61), .Z(n4427) );
  XNOR U4721 ( .A(n4428), .B(n4427), .Z(n4544) );
  XNOR U4722 ( .A(n4545), .B(n4544), .Z(n4578) );
  NANDN U4723 ( .A(n8890), .B(y[230]), .Z(n4521) );
  NANDN U4724 ( .A(n8626), .B(y[229]), .Z(n4519) );
  NANDN U4725 ( .A(n50), .B(y[241]), .Z(n4518) );
  XNOR U4726 ( .A(n4519), .B(n4518), .Z(n4520) );
  XNOR U4727 ( .A(n4521), .B(n4520), .Z(n4579) );
  XNOR U4728 ( .A(n4581), .B(n4580), .Z(n4616) );
  OR U4729 ( .A(n4430), .B(n4429), .Z(n4434) );
  NANDN U4730 ( .A(n4432), .B(n4431), .Z(n4433) );
  NAND U4731 ( .A(n4434), .B(n4433), .Z(n4617) );
  XNOR U4732 ( .A(n4616), .B(n4617), .Z(n4619) );
  XOR U4733 ( .A(n4618), .B(n4619), .Z(n4599) );
  NANDN U4734 ( .A(n8824), .B(y[227]), .Z(n4595) );
  NANDN U4735 ( .A(n48), .B(y[243]), .Z(n4593) );
  NANDN U4736 ( .A(n59), .B(y[232]), .Z(n4592) );
  XNOR U4737 ( .A(n4593), .B(n4592), .Z(n4594) );
  XNOR U4738 ( .A(n4595), .B(n4594), .Z(n4567) );
  NAND U4739 ( .A(o[53]), .B(n4435), .Z(n4589) );
  ANDN U4740 ( .B(y[245]), .A(n46), .Z(n4586) );
  XNOR U4741 ( .A(n4587), .B(n4586), .Z(n4588) );
  XOR U4742 ( .A(n4589), .B(n4588), .Z(n4566) );
  XOR U4743 ( .A(n4567), .B(n4566), .Z(n4569) );
  AND U4744 ( .A(y[242]), .B(x[77]), .Z(n5913) );
  IV U4745 ( .A(n5913), .Z(n5851) );
  NANDN U4746 ( .A(n5851), .B(n4436), .Z(n4440) );
  OR U4747 ( .A(n4438), .B(n4437), .Z(n4439) );
  AND U4748 ( .A(n4440), .B(n4439), .Z(n4568) );
  XOR U4749 ( .A(n4569), .B(n4568), .Z(n4610) );
  NANDN U4750 ( .A(n60), .B(y[231]), .Z(n4526) );
  ANDN U4751 ( .B(y[240]), .A(n51), .Z(n4442) );
  ANDN U4752 ( .B(y[236]), .A(n55), .Z(n4441) );
  XNOR U4753 ( .A(n4442), .B(n4441), .Z(n4525) );
  XNOR U4754 ( .A(n4526), .B(n4525), .Z(n4554) );
  NAND U4755 ( .A(n4444), .B(n4443), .Z(n4448) );
  NAND U4756 ( .A(n4446), .B(n4445), .Z(n4447) );
  AND U4757 ( .A(n4448), .B(n4447), .Z(n4555) );
  NANDN U4758 ( .A(n47), .B(y[244]), .Z(n4530) );
  ANDN U4759 ( .B(y[226]), .A(n8885), .Z(n4529) );
  XOR U4760 ( .A(n4530), .B(n4529), .Z(n4532) );
  ANDN U4761 ( .B(x[77]), .A(n5637), .Z(n4531) );
  XOR U4762 ( .A(n4532), .B(n4531), .Z(n4556) );
  XOR U4763 ( .A(n4557), .B(n4556), .Z(n4611) );
  XNOR U4764 ( .A(n4610), .B(n4611), .Z(n4613) );
  OR U4765 ( .A(n4450), .B(n4449), .Z(n4454) );
  OR U4766 ( .A(n4452), .B(n4451), .Z(n4453) );
  NAND U4767 ( .A(n4454), .B(n4453), .Z(n4563) );
  ANDN U4768 ( .B(y[239]), .A(n52), .Z(n4456) );
  ANDN U4769 ( .B(x[72]), .A(n5473), .Z(n4455) );
  XNOR U4770 ( .A(n4456), .B(n4455), .Z(n4540) );
  XOR U4771 ( .A(n4539), .B(n4540), .Z(n4561) );
  NANDN U4772 ( .A(n45), .B(y[246]), .Z(n4549) );
  ANDN U4773 ( .B(x[86]), .A(n5905), .Z(n4548) );
  XNOR U4774 ( .A(n4549), .B(n4548), .Z(n4551) );
  NANDN U4775 ( .A(n8827), .B(y[225]), .Z(n4517) );
  XNOR U4776 ( .A(n4517), .B(o[54]), .Z(n4550) );
  XNOR U4777 ( .A(n4551), .B(n4550), .Z(n4560) );
  XNOR U4778 ( .A(n4561), .B(n4560), .Z(n4562) );
  OR U4779 ( .A(n4458), .B(n4457), .Z(n4462) );
  OR U4780 ( .A(n4460), .B(n4459), .Z(n4461) );
  AND U4781 ( .A(n4462), .B(n4461), .Z(n4573) );
  OR U4782 ( .A(n4464), .B(n4463), .Z(n4468) );
  OR U4783 ( .A(n4466), .B(n4465), .Z(n4467) );
  AND U4784 ( .A(n4468), .B(n4467), .Z(n4572) );
  XNOR U4785 ( .A(n4573), .B(n4572), .Z(n4574) );
  XNOR U4786 ( .A(n4575), .B(n4574), .Z(n4612) );
  XNOR U4787 ( .A(n4613), .B(n4612), .Z(n4605) );
  NANDN U4788 ( .A(n4470), .B(n4469), .Z(n4474) );
  OR U4789 ( .A(n4472), .B(n4471), .Z(n4473) );
  NAND U4790 ( .A(n4474), .B(n4473), .Z(n4604) );
  XNOR U4791 ( .A(n4605), .B(n4604), .Z(n4606) );
  OR U4792 ( .A(n4476), .B(n4475), .Z(n4480) );
  OR U4793 ( .A(n4478), .B(n4477), .Z(n4479) );
  AND U4794 ( .A(n4480), .B(n4479), .Z(n4607) );
  XOR U4795 ( .A(n4599), .B(n4598), .Z(n4600) );
  XOR U4796 ( .A(n4601), .B(n4600), .Z(n4501) );
  XNOR U4797 ( .A(n4502), .B(n4501), .Z(n4507) );
  XNOR U4798 ( .A(n4508), .B(n4507), .Z(n4494) );
  OR U4799 ( .A(n4482), .B(n4481), .Z(n4486) );
  NANDN U4800 ( .A(n4484), .B(n4483), .Z(n4485) );
  NAND U4801 ( .A(n4486), .B(n4485), .Z(n4493) );
  XNOR U4802 ( .A(n4496), .B(n4495), .Z(n4490) );
  XOR U4803 ( .A(n4489), .B(n4490), .Z(N119) );
  NANDN U4804 ( .A(n4488), .B(n4487), .Z(n4492) );
  NANDN U4805 ( .A(n4490), .B(n4489), .Z(n4491) );
  NAND U4806 ( .A(n4492), .B(n4491), .Z(n4622) );
  OR U4807 ( .A(n4494), .B(n4493), .Z(n4498) );
  NANDN U4808 ( .A(n4496), .B(n4495), .Z(n4497) );
  NAND U4809 ( .A(n4498), .B(n4497), .Z(n4623) );
  XNOR U4810 ( .A(n4622), .B(n4623), .Z(n4624) );
  OR U4811 ( .A(n4500), .B(n4499), .Z(n4504) );
  OR U4812 ( .A(n4502), .B(n4501), .Z(n4503) );
  AND U4813 ( .A(n4504), .B(n4503), .Z(n4628) );
  OR U4814 ( .A(n4506), .B(n4505), .Z(n4510) );
  NAND U4815 ( .A(n4508), .B(n4507), .Z(n4509) );
  NAND U4816 ( .A(n4510), .B(n4509), .Z(n4629) );
  XOR U4817 ( .A(n4628), .B(n4629), .Z(n4631) );
  OR U4818 ( .A(n4512), .B(n4511), .Z(n4516) );
  NANDN U4819 ( .A(n4514), .B(n4513), .Z(n4515) );
  AND U4820 ( .A(n4516), .B(n4515), .Z(n4648) );
  NANDN U4821 ( .A(n8827), .B(y[226]), .Z(n4709) );
  NANDN U4822 ( .A(n47), .B(y[245]), .Z(n4707) );
  NANDN U4823 ( .A(n58), .B(y[234]), .Z(n4706) );
  XNOR U4824 ( .A(n4707), .B(n4706), .Z(n4708) );
  XNOR U4825 ( .A(n4709), .B(n4708), .Z(n4667) );
  NANDN U4826 ( .A(n4517), .B(o[54]), .Z(n4750) );
  NANDN U4827 ( .A(n46), .B(y[246]), .Z(n4748) );
  NANDN U4828 ( .A(n57), .B(y[235]), .Z(n4747) );
  XNOR U4829 ( .A(n4748), .B(n4747), .Z(n4749) );
  XNOR U4830 ( .A(n4750), .B(n4749), .Z(n4665) );
  OR U4831 ( .A(n4519), .B(n4518), .Z(n4523) );
  OR U4832 ( .A(n4521), .B(n4520), .Z(n4522) );
  AND U4833 ( .A(n4523), .B(n4522), .Z(n4664) );
  XNOR U4834 ( .A(n4665), .B(n4664), .Z(n4666) );
  XNOR U4835 ( .A(n4667), .B(n4666), .Z(n4720) );
  ANDN U4836 ( .B(y[240]), .A(n55), .Z(n5131) );
  NANDN U4837 ( .A(n4524), .B(n5131), .Z(n4528) );
  OR U4838 ( .A(n4526), .B(n4525), .Z(n4527) );
  AND U4839 ( .A(n4528), .B(n4527), .Z(n4670) );
  NANDN U4840 ( .A(n8626), .B(y[230]), .Z(n4715) );
  NANDN U4841 ( .A(n61), .B(y[229]), .Z(n4713) );
  NANDN U4842 ( .A(n50), .B(y[242]), .Z(n4712) );
  XNOR U4843 ( .A(n4713), .B(n4712), .Z(n4714) );
  XNOR U4844 ( .A(n4715), .B(n4714), .Z(n4671) );
  XOR U4845 ( .A(n4670), .B(n4671), .Z(n4672) );
  NANDN U4846 ( .A(n49), .B(y[243]), .Z(n4703) );
  NANDN U4847 ( .A(n48), .B(y[244]), .Z(n4701) );
  ANDN U4848 ( .B(x[78]), .A(n5637), .Z(n4700) );
  XOR U4849 ( .A(n4701), .B(n4700), .Z(n4702) );
  XOR U4850 ( .A(n4672), .B(n4673), .Z(n4718) );
  NANDN U4851 ( .A(n4530), .B(n4529), .Z(n4534) );
  NANDN U4852 ( .A(n4532), .B(n4531), .Z(n4533) );
  NAND U4853 ( .A(n4534), .B(n4533), .Z(n4719) );
  XOR U4854 ( .A(n4718), .B(n4719), .Z(n4721) );
  XNOR U4855 ( .A(n4720), .B(n4721), .Z(n4756) );
  ANDN U4856 ( .B(y[225]), .A(n8864), .Z(n4734) );
  XNOR U4857 ( .A(o[55]), .B(n4734), .Z(n4727) );
  NANDN U4858 ( .A(n8656), .B(y[224]), .Z(n4725) );
  NANDN U4859 ( .A(n45), .B(y[247]), .Z(n4724) );
  XNOR U4860 ( .A(n4725), .B(n4724), .Z(n4726) );
  XOR U4861 ( .A(n4727), .B(n4726), .Z(n4678) );
  AND U4862 ( .A(y[228]), .B(x[83]), .Z(n5010) );
  ANDN U4863 ( .B(x[84]), .A(n5714), .Z(n4535) );
  XNOR U4864 ( .A(n4536), .B(n4535), .Z(n4731) );
  XNOR U4865 ( .A(n5010), .B(n4731), .Z(n4676) );
  OR U4866 ( .A(n4538), .B(n4537), .Z(n4542) );
  NANDN U4867 ( .A(n4540), .B(n4539), .Z(n4541) );
  NAND U4868 ( .A(n4542), .B(n4541), .Z(n4677) );
  XNOR U4869 ( .A(n4676), .B(n4677), .Z(n4679) );
  XOR U4870 ( .A(n4678), .B(n4679), .Z(n4685) );
  AND U4871 ( .A(x[82]), .B(y[234]), .Z(n5419) );
  NANDN U4872 ( .A(n4543), .B(n5419), .Z(n4547) );
  OR U4873 ( .A(n4545), .B(n4544), .Z(n4546) );
  AND U4874 ( .A(n4547), .B(n4546), .Z(n4682) );
  NANDN U4875 ( .A(n4549), .B(n4548), .Z(n4553) );
  NAND U4876 ( .A(n4551), .B(n4550), .Z(n4552) );
  AND U4877 ( .A(n4553), .B(n4552), .Z(n4683) );
  XOR U4878 ( .A(n4682), .B(n4683), .Z(n4684) );
  XOR U4879 ( .A(n4685), .B(n4684), .Z(n4754) );
  OR U4880 ( .A(n4555), .B(n4554), .Z(n4559) );
  OR U4881 ( .A(n4557), .B(n4556), .Z(n4558) );
  AND U4882 ( .A(n4559), .B(n4558), .Z(n4753) );
  XOR U4883 ( .A(n4754), .B(n4753), .Z(n4755) );
  XOR U4884 ( .A(n4756), .B(n4755), .Z(n4647) );
  OR U4885 ( .A(n4561), .B(n4560), .Z(n4565) );
  OR U4886 ( .A(n4563), .B(n4562), .Z(n4564) );
  AND U4887 ( .A(n4565), .B(n4564), .Z(n4658) );
  NANDN U4888 ( .A(n4567), .B(n4566), .Z(n4571) );
  OR U4889 ( .A(n4569), .B(n4568), .Z(n4570) );
  AND U4890 ( .A(n4571), .B(n4570), .Z(n4659) );
  XNOR U4891 ( .A(n4658), .B(n4659), .Z(n4660) );
  OR U4892 ( .A(n4573), .B(n4572), .Z(n4577) );
  OR U4893 ( .A(n4575), .B(n4574), .Z(n4576) );
  NAND U4894 ( .A(n4577), .B(n4576), .Z(n4661) );
  OR U4895 ( .A(n4579), .B(n4578), .Z(n4583) );
  NANDN U4896 ( .A(n4581), .B(n4580), .Z(n4582) );
  AND U4897 ( .A(n4583), .B(n4582), .Z(n4634) );
  NANDN U4898 ( .A(n52), .B(y[240]), .Z(n4744) );
  ANDN U4899 ( .B(y[239]), .A(n53), .Z(n4585) );
  ANDN U4900 ( .B(x[73]), .A(n5473), .Z(n4584) );
  XNOR U4901 ( .A(n4585), .B(n4584), .Z(n4743) );
  XNOR U4902 ( .A(n4744), .B(n4743), .Z(n4695) );
  ANDN U4903 ( .B(x[74]), .A(n5332), .Z(n4694) );
  XOR U4904 ( .A(n4695), .B(n4694), .Z(n4697) );
  NANDN U4905 ( .A(n60), .B(y[232]), .Z(n4737) );
  ANDN U4906 ( .B(x[70]), .A(n5874), .Z(n4736) );
  XOR U4907 ( .A(n4737), .B(n4736), .Z(n4739) );
  XOR U4908 ( .A(n4697), .B(n4696), .Z(n4690) );
  NAND U4909 ( .A(n4587), .B(n4586), .Z(n4591) );
  OR U4910 ( .A(n4589), .B(n4588), .Z(n4590) );
  NAND U4911 ( .A(n4591), .B(n4590), .Z(n4689) );
  OR U4912 ( .A(n4593), .B(n4592), .Z(n4597) );
  OR U4913 ( .A(n4595), .B(n4594), .Z(n4596) );
  NAND U4914 ( .A(n4597), .B(n4596), .Z(n4688) );
  XNOR U4915 ( .A(n4689), .B(n4688), .Z(n4691) );
  XNOR U4916 ( .A(n4690), .B(n4691), .Z(n4635) );
  XNOR U4917 ( .A(n4634), .B(n4635), .Z(n4636) );
  XNOR U4918 ( .A(n4647), .B(n4646), .Z(n4649) );
  XNOR U4919 ( .A(n4648), .B(n4649), .Z(n4654) );
  NANDN U4920 ( .A(n4599), .B(n4598), .Z(n4603) );
  OR U4921 ( .A(n4601), .B(n4600), .Z(n4602) );
  NAND U4922 ( .A(n4603), .B(n4602), .Z(n4653) );
  OR U4923 ( .A(n4605), .B(n4604), .Z(n4609) );
  OR U4924 ( .A(n4607), .B(n4606), .Z(n4608) );
  AND U4925 ( .A(n4609), .B(n4608), .Z(n4643) );
  OR U4926 ( .A(n4611), .B(n4610), .Z(n4615) );
  OR U4927 ( .A(n4613), .B(n4612), .Z(n4614) );
  AND U4928 ( .A(n4615), .B(n4614), .Z(n4640) );
  OR U4929 ( .A(n4617), .B(n4616), .Z(n4621) );
  OR U4930 ( .A(n4619), .B(n4618), .Z(n4620) );
  AND U4931 ( .A(n4621), .B(n4620), .Z(n4641) );
  XNOR U4932 ( .A(n4640), .B(n4641), .Z(n4642) );
  XNOR U4933 ( .A(n4653), .B(n4652), .Z(n4655) );
  XNOR U4934 ( .A(n4631), .B(n4630), .Z(n4625) );
  XOR U4935 ( .A(n4624), .B(n4625), .Z(N120) );
  NANDN U4936 ( .A(n4623), .B(n4622), .Z(n4627) );
  NANDN U4937 ( .A(n4625), .B(n4624), .Z(n4626) );
  NAND U4938 ( .A(n4627), .B(n4626), .Z(n4759) );
  OR U4939 ( .A(n4629), .B(n4628), .Z(n4633) );
  NAND U4940 ( .A(n4631), .B(n4630), .Z(n4632) );
  AND U4941 ( .A(n4633), .B(n4632), .Z(n4760) );
  XNOR U4942 ( .A(n4759), .B(n4760), .Z(n4761) );
  OR U4943 ( .A(n4635), .B(n4634), .Z(n4639) );
  OR U4944 ( .A(n4637), .B(n4636), .Z(n4638) );
  NAND U4945 ( .A(n4639), .B(n4638), .Z(n4902) );
  OR U4946 ( .A(n4641), .B(n4640), .Z(n4645) );
  OR U4947 ( .A(n4643), .B(n4642), .Z(n4644) );
  AND U4948 ( .A(n4645), .B(n4644), .Z(n4901) );
  XNOR U4949 ( .A(n4902), .B(n4901), .Z(n4903) );
  OR U4950 ( .A(n4647), .B(n4646), .Z(n4651) );
  OR U4951 ( .A(n4649), .B(n4648), .Z(n4650) );
  NAND U4952 ( .A(n4651), .B(n4650), .Z(n4904) );
  OR U4953 ( .A(n4653), .B(n4652), .Z(n4657) );
  NANDN U4954 ( .A(n4655), .B(n4654), .Z(n4656) );
  AND U4955 ( .A(n4657), .B(n4656), .Z(n4765) );
  OR U4956 ( .A(n4659), .B(n4658), .Z(n4663) );
  OR U4957 ( .A(n4661), .B(n4660), .Z(n4662) );
  NAND U4958 ( .A(n4663), .B(n4662), .Z(n4772) );
  OR U4959 ( .A(n4665), .B(n4664), .Z(n4669) );
  OR U4960 ( .A(n4667), .B(n4666), .Z(n4668) );
  AND U4961 ( .A(n4669), .B(n4668), .Z(n4895) );
  OR U4962 ( .A(n4671), .B(n4670), .Z(n4675) );
  NANDN U4963 ( .A(n4673), .B(n4672), .Z(n4674) );
  NAND U4964 ( .A(n4675), .B(n4674), .Z(n4848) );
  OR U4965 ( .A(n4677), .B(n4676), .Z(n4681) );
  OR U4966 ( .A(n4679), .B(n4678), .Z(n4680) );
  AND U4967 ( .A(n4681), .B(n4680), .Z(n4845) );
  OR U4968 ( .A(n4683), .B(n4682), .Z(n4687) );
  NANDN U4969 ( .A(n4685), .B(n4684), .Z(n4686) );
  NAND U4970 ( .A(n4687), .B(n4686), .Z(n4846) );
  XOR U4971 ( .A(n4845), .B(n4846), .Z(n4847) );
  XNOR U4972 ( .A(n4848), .B(n4847), .Z(n4896) );
  XOR U4973 ( .A(n4895), .B(n4896), .Z(n4897) );
  OR U4974 ( .A(n4689), .B(n4688), .Z(n4693) );
  NANDN U4975 ( .A(n4691), .B(n4690), .Z(n4692) );
  NAND U4976 ( .A(n4693), .B(n4692), .Z(n4842) );
  NANDN U4977 ( .A(n4695), .B(n4694), .Z(n4699) );
  NANDN U4978 ( .A(n4697), .B(n4696), .Z(n4698) );
  AND U4979 ( .A(n4699), .B(n4698), .Z(n4839) );
  NANDN U4980 ( .A(n4701), .B(n4700), .Z(n4705) );
  OR U4981 ( .A(n4703), .B(n4702), .Z(n4704) );
  AND U4982 ( .A(n4705), .B(n4704), .Z(n4851) );
  OR U4983 ( .A(n4707), .B(n4706), .Z(n4711) );
  OR U4984 ( .A(n4709), .B(n4708), .Z(n4710) );
  AND U4985 ( .A(n4711), .B(n4710), .Z(n4852) );
  XOR U4986 ( .A(n4851), .B(n4852), .Z(n4853) );
  OR U4987 ( .A(n4713), .B(n4712), .Z(n4717) );
  OR U4988 ( .A(n4715), .B(n4714), .Z(n4716) );
  AND U4989 ( .A(n4717), .B(n4716), .Z(n4879) );
  NANDN U4990 ( .A(n61), .B(y[230]), .Z(n4805) );
  NANDN U4991 ( .A(n8626), .B(y[231]), .Z(n4803) );
  NANDN U4992 ( .A(n52), .B(y[241]), .Z(n4802) );
  XNOR U4993 ( .A(n4803), .B(n4802), .Z(n4804) );
  XNOR U4994 ( .A(n4805), .B(n4804), .Z(n4878) );
  NANDN U4995 ( .A(n8656), .B(y[225]), .Z(n4801) );
  XOR U4996 ( .A(o[56]), .B(n4801), .Z(n4824) );
  NANDN U4997 ( .A(n45), .B(y[248]), .Z(n4822) );
  NANDN U4998 ( .A(n8865), .B(y[224]), .Z(n4821) );
  XNOR U4999 ( .A(n4822), .B(n4821), .Z(n4823) );
  XNOR U5000 ( .A(n4824), .B(n4823), .Z(n4877) );
  XNOR U5001 ( .A(n4878), .B(n4877), .Z(n4880) );
  XNOR U5002 ( .A(n4879), .B(n4880), .Z(n4854) );
  XOR U5003 ( .A(n4853), .B(n4854), .Z(n4840) );
  XNOR U5004 ( .A(n4839), .B(n4840), .Z(n4841) );
  XOR U5005 ( .A(n4897), .B(n4898), .Z(n4771) );
  XOR U5006 ( .A(n4772), .B(n4771), .Z(n4774) );
  NANDN U5007 ( .A(n4719), .B(n4718), .Z(n4723) );
  NANDN U5008 ( .A(n4721), .B(n4720), .Z(n4722) );
  NAND U5009 ( .A(n4723), .B(n4722), .Z(n4778) );
  NANDN U5010 ( .A(n49), .B(y[244]), .Z(n4830) );
  NANDN U5011 ( .A(n48), .B(y[245]), .Z(n4828) );
  NANDN U5012 ( .A(n60), .B(y[233]), .Z(n4827) );
  XNOR U5013 ( .A(n4828), .B(n4827), .Z(n4829) );
  XNOR U5014 ( .A(n4830), .B(n4829), .Z(n4836) );
  OR U5015 ( .A(n4725), .B(n4724), .Z(n4729) );
  OR U5016 ( .A(n4727), .B(n4726), .Z(n4728) );
  AND U5017 ( .A(n4729), .B(n4728), .Z(n4833) );
  NANDN U5018 ( .A(n59), .B(y[234]), .Z(n4817) );
  NANDN U5019 ( .A(n56), .B(y[237]), .Z(n4815) );
  NANDN U5020 ( .A(n53), .B(y[240]), .Z(n4814) );
  XNOR U5021 ( .A(n4815), .B(n4814), .Z(n4816) );
  XOR U5022 ( .A(n4817), .B(n4816), .Z(n4810) );
  AND U5023 ( .A(y[239]), .B(x[73]), .Z(n4808) );
  AND U5024 ( .A(y[238]), .B(x[74]), .Z(n4809) );
  XNOR U5025 ( .A(n4808), .B(n4809), .Z(n4811) );
  XNOR U5026 ( .A(n4833), .B(n4834), .Z(n4835) );
  XNOR U5027 ( .A(n4836), .B(n4835), .Z(n4785) );
  ANDN U5028 ( .B(x[84]), .A(n44), .Z(n5177) );
  IV U5029 ( .A(n5177), .Z(n5284) );
  ANDN U5030 ( .B(y[227]), .A(n8890), .Z(n4730) );
  NANDN U5031 ( .A(n5284), .B(n4730), .Z(n4733) );
  NANDN U5032 ( .A(n4731), .B(n5010), .Z(n4732) );
  AND U5033 ( .A(n4733), .B(n4732), .Z(n4889) );
  NAND U5034 ( .A(n4734), .B(o[55]), .Z(n4792) );
  NANDN U5035 ( .A(n46), .B(y[247]), .Z(n4790) );
  XOR U5036 ( .A(n4735), .B(n4790), .Z(n4791) );
  XNOR U5037 ( .A(n4792), .B(n4791), .Z(n4890) );
  XNOR U5038 ( .A(n4889), .B(n4890), .Z(n4892) );
  NANDN U5039 ( .A(n47), .B(y[246]), .Z(n4796) );
  ANDN U5040 ( .B(y[226]), .A(n8864), .Z(n4795) );
  XOR U5041 ( .A(n4796), .B(n4795), .Z(n4798) );
  XOR U5042 ( .A(n4892), .B(n4891), .Z(n4783) );
  NANDN U5043 ( .A(n8885), .B(y[228]), .Z(n4874) );
  NANDN U5044 ( .A(n8824), .B(y[229]), .Z(n4872) );
  NANDN U5045 ( .A(n51), .B(y[242]), .Z(n4871) );
  XNOR U5046 ( .A(n4872), .B(n4871), .Z(n4873) );
  XNOR U5047 ( .A(n4874), .B(n4873), .Z(n4884) );
  NANDN U5048 ( .A(n8890), .B(y[232]), .Z(n4866) );
  NANDN U5049 ( .A(n50), .B(y[243]), .Z(n4864) );
  ANDN U5050 ( .B(x[85]), .A(n5714), .Z(n4863) );
  XOR U5051 ( .A(n4864), .B(n4863), .Z(n4865) );
  XOR U5052 ( .A(n4884), .B(n4883), .Z(n4886) );
  NANDN U5053 ( .A(n4737), .B(n4736), .Z(n4741) );
  NANDN U5054 ( .A(n4739), .B(n4738), .Z(n4740) );
  AND U5055 ( .A(n4741), .B(n4740), .Z(n4885) );
  XNOR U5056 ( .A(n4886), .B(n4885), .Z(n4857) );
  NANDN U5057 ( .A(n4742), .B(n4808), .Z(n4746) );
  OR U5058 ( .A(n4744), .B(n4743), .Z(n4745) );
  AND U5059 ( .A(n4746), .B(n4745), .Z(n4858) );
  OR U5060 ( .A(n4748), .B(n4747), .Z(n4752) );
  OR U5061 ( .A(n4750), .B(n4749), .Z(n4751) );
  AND U5062 ( .A(n4752), .B(n4751), .Z(n4859) );
  XOR U5063 ( .A(n4860), .B(n4859), .Z(n4784) );
  XOR U5064 ( .A(n4783), .B(n4784), .Z(n4786) );
  XNOR U5065 ( .A(n4785), .B(n4786), .Z(n4777) );
  XNOR U5066 ( .A(n4778), .B(n4777), .Z(n4780) );
  OR U5067 ( .A(n4754), .B(n4753), .Z(n4758) );
  NANDN U5068 ( .A(n4756), .B(n4755), .Z(n4757) );
  AND U5069 ( .A(n4758), .B(n4757), .Z(n4779) );
  XOR U5070 ( .A(n4780), .B(n4779), .Z(n4773) );
  XNOR U5071 ( .A(n4774), .B(n4773), .Z(n4766) );
  XNOR U5072 ( .A(n4765), .B(n4766), .Z(n4767) );
  XNOR U5073 ( .A(n4768), .B(n4767), .Z(n4762) );
  XOR U5074 ( .A(n4761), .B(n4762), .Z(N121) );
  NANDN U5075 ( .A(n4760), .B(n4759), .Z(n4764) );
  NANDN U5076 ( .A(n4762), .B(n4761), .Z(n4763) );
  NAND U5077 ( .A(n4764), .B(n4763), .Z(n5047) );
  OR U5078 ( .A(n4766), .B(n4765), .Z(n4770) );
  OR U5079 ( .A(n4768), .B(n4767), .Z(n4769) );
  AND U5080 ( .A(n4770), .B(n4769), .Z(n5048) );
  XNOR U5081 ( .A(n5047), .B(n5048), .Z(n5049) );
  NANDN U5082 ( .A(n4772), .B(n4771), .Z(n4776) );
  OR U5083 ( .A(n4774), .B(n4773), .Z(n4775) );
  AND U5084 ( .A(n4776), .B(n4775), .Z(n5053) );
  OR U5085 ( .A(n4778), .B(n4777), .Z(n4782) );
  OR U5086 ( .A(n4780), .B(n4779), .Z(n4781) );
  NAND U5087 ( .A(n4782), .B(n4781), .Z(n4914) );
  NANDN U5088 ( .A(n4784), .B(n4783), .Z(n4788) );
  NANDN U5089 ( .A(n4786), .B(n4785), .Z(n4787) );
  AND U5090 ( .A(n4788), .B(n4787), .Z(n5041) );
  OR U5091 ( .A(n4790), .B(n4789), .Z(n4794) );
  OR U5092 ( .A(n4792), .B(n4791), .Z(n4793) );
  AND U5093 ( .A(n4794), .B(n4793), .Z(n4939) );
  NANDN U5094 ( .A(n4796), .B(n4795), .Z(n4800) );
  NANDN U5095 ( .A(n4798), .B(n4797), .Z(n4799) );
  AND U5096 ( .A(n4800), .B(n4799), .Z(n4938) );
  NAND U5097 ( .A(y[241]), .B(x[72]), .Z(n4934) );
  XNOR U5098 ( .A(n4932), .B(n4931), .Z(n4933) );
  XOR U5099 ( .A(n4934), .B(n4933), .Z(n4919) );
  NANDN U5100 ( .A(n4801), .B(o[56]), .Z(n4928) );
  ANDN U5101 ( .B(x[89]), .A(n5905), .Z(n4926) );
  ANDN U5102 ( .B(y[249]), .A(n45), .Z(n4925) );
  XOR U5103 ( .A(n4926), .B(n4925), .Z(n4927) );
  XOR U5104 ( .A(n4928), .B(n4927), .Z(n4920) );
  XNOR U5105 ( .A(n4919), .B(n4920), .Z(n4922) );
  OR U5106 ( .A(n4803), .B(n4802), .Z(n4807) );
  OR U5107 ( .A(n4805), .B(n4804), .Z(n4806) );
  AND U5108 ( .A(n4807), .B(n4806), .Z(n4921) );
  XNOR U5109 ( .A(n4922), .B(n4921), .Z(n4937) );
  XOR U5110 ( .A(n4939), .B(n4940), .Z(n4946) );
  OR U5111 ( .A(n4809), .B(n4808), .Z(n4813) );
  OR U5112 ( .A(n4811), .B(n4810), .Z(n4812) );
  AND U5113 ( .A(n4813), .B(n4812), .Z(n4943) );
  NANDN U5114 ( .A(n46), .B(y[248]), .Z(n4992) );
  ANDN U5115 ( .B(y[236]), .A(n58), .Z(n4991) );
  XNOR U5116 ( .A(n4992), .B(n4991), .Z(n4993) );
  NANDN U5117 ( .A(n8865), .B(y[225]), .Z(n5016) );
  XOR U5118 ( .A(n5016), .B(o[57]), .Z(n4994) );
  XOR U5119 ( .A(n4993), .B(n4994), .Z(n5000) );
  NAND U5120 ( .A(y[238]), .B(x[75]), .Z(n5019) );
  NAND U5121 ( .A(y[237]), .B(x[76]), .Z(n5018) );
  NAND U5122 ( .A(x[71]), .B(y[242]), .Z(n5017) );
  XNOR U5123 ( .A(n5018), .B(n5017), .Z(n5020) );
  XNOR U5124 ( .A(n5019), .B(n5020), .Z(n4997) );
  OR U5125 ( .A(n4815), .B(n4814), .Z(n4819) );
  OR U5126 ( .A(n4817), .B(n4816), .Z(n4818) );
  AND U5127 ( .A(n4819), .B(n4818), .Z(n4998) );
  XNOR U5128 ( .A(n4997), .B(n4998), .Z(n4999) );
  XOR U5129 ( .A(n5000), .B(n4999), .Z(n4944) );
  XOR U5130 ( .A(n4943), .B(n4944), .Z(n4945) );
  XOR U5131 ( .A(n4946), .B(n4945), .Z(n5038) );
  NANDN U5132 ( .A(n48), .B(y[246]), .Z(n4988) );
  NANDN U5133 ( .A(n47), .B(y[247]), .Z(n4986) );
  XOR U5134 ( .A(n4820), .B(n4986), .Z(n4987) );
  XNOR U5135 ( .A(n4988), .B(n4987), .Z(n4980) );
  OR U5136 ( .A(n4822), .B(n4821), .Z(n4826) );
  OR U5137 ( .A(n4824), .B(n4823), .Z(n4825) );
  AND U5138 ( .A(n4826), .B(n4825), .Z(n4979) );
  XNOR U5139 ( .A(n4980), .B(n4979), .Z(n4981) );
  OR U5140 ( .A(n4828), .B(n4827), .Z(n4832) );
  OR U5141 ( .A(n4830), .B(n4829), .Z(n4831) );
  AND U5142 ( .A(n4832), .B(n4831), .Z(n4982) );
  OR U5143 ( .A(n4834), .B(n4833), .Z(n4838) );
  OR U5144 ( .A(n4836), .B(n4835), .Z(n4837) );
  AND U5145 ( .A(n4838), .B(n4837), .Z(n5035) );
  XOR U5146 ( .A(n5036), .B(n5035), .Z(n5037) );
  XOR U5147 ( .A(n5038), .B(n5037), .Z(n5042) );
  XNOR U5148 ( .A(n5041), .B(n5042), .Z(n5043) );
  OR U5149 ( .A(n4840), .B(n4839), .Z(n4844) );
  OR U5150 ( .A(n4842), .B(n4841), .Z(n4843) );
  NAND U5151 ( .A(n4844), .B(n4843), .Z(n5044) );
  XOR U5152 ( .A(n4914), .B(n4913), .Z(n4916) );
  OR U5153 ( .A(n4846), .B(n4845), .Z(n4850) );
  NANDN U5154 ( .A(n4848), .B(n4847), .Z(n4849) );
  NAND U5155 ( .A(n4850), .B(n4849), .Z(n4908) );
  OR U5156 ( .A(n4852), .B(n4851), .Z(n4856) );
  NANDN U5157 ( .A(n4854), .B(n4853), .Z(n4855) );
  NAND U5158 ( .A(n4856), .B(n4855), .Z(n4956) );
  OR U5159 ( .A(n4858), .B(n4857), .Z(n4862) );
  OR U5160 ( .A(n4860), .B(n4859), .Z(n4861) );
  NAND U5161 ( .A(n4862), .B(n4861), .Z(n4955) );
  XNOR U5162 ( .A(n4956), .B(n4955), .Z(n4957) );
  NANDN U5163 ( .A(n4864), .B(n4863), .Z(n4868) );
  OR U5164 ( .A(n4866), .B(n4865), .Z(n4867) );
  AND U5165 ( .A(n4868), .B(n4867), .Z(n4975) );
  NAND U5166 ( .A(y[227]), .B(x[86]), .Z(n5031) );
  NAND U5167 ( .A(x[69]), .B(y[244]), .Z(n5030) );
  NAND U5168 ( .A(y[232]), .B(x[81]), .Z(n5029) );
  XNOR U5169 ( .A(n5030), .B(n5029), .Z(n5032) );
  XNOR U5170 ( .A(n5031), .B(n5032), .Z(n4974) );
  NANDN U5171 ( .A(n8885), .B(y[229]), .Z(n5012) );
  ANDN U5172 ( .B(x[83]), .A(n5663), .Z(n4870) );
  ANDN U5173 ( .B(y[228]), .A(n8827), .Z(n4869) );
  XNOR U5174 ( .A(n4870), .B(n4869), .Z(n5011) );
  XOR U5175 ( .A(n5012), .B(n5011), .Z(n4973) );
  XOR U5176 ( .A(n4974), .B(n4973), .Z(n4976) );
  XOR U5177 ( .A(n4975), .B(n4976), .Z(n4949) );
  ANDN U5178 ( .B(y[226]), .A(n8656), .Z(n5025) );
  NAND U5179 ( .A(x[68]), .B(y[245]), .Z(n5024) );
  NAND U5180 ( .A(y[233]), .B(x[80]), .Z(n5023) );
  XNOR U5181 ( .A(n5024), .B(n5023), .Z(n5026) );
  XNOR U5182 ( .A(n5025), .B(n5026), .Z(n4969) );
  ANDN U5183 ( .B(x[79]), .A(n5196), .Z(n5006) );
  NAND U5184 ( .A(y[231]), .B(x[82]), .Z(n5005) );
  NAND U5185 ( .A(x[70]), .B(y[243]), .Z(n5004) );
  XNOR U5186 ( .A(n5005), .B(n5004), .Z(n5007) );
  XOR U5187 ( .A(n5006), .B(n5007), .Z(n4968) );
  OR U5188 ( .A(n4872), .B(n4871), .Z(n4876) );
  OR U5189 ( .A(n4874), .B(n4873), .Z(n4875) );
  AND U5190 ( .A(n4876), .B(n4875), .Z(n4967) );
  XNOR U5191 ( .A(n4968), .B(n4967), .Z(n4970) );
  XOR U5192 ( .A(n4969), .B(n4970), .Z(n4950) );
  XOR U5193 ( .A(n4949), .B(n4950), .Z(n4952) );
  OR U5194 ( .A(n4878), .B(n4877), .Z(n4882) );
  OR U5195 ( .A(n4880), .B(n4879), .Z(n4881) );
  AND U5196 ( .A(n4882), .B(n4881), .Z(n4951) );
  XOR U5197 ( .A(n4952), .B(n4951), .Z(n4963) );
  NANDN U5198 ( .A(n4884), .B(n4883), .Z(n4888) );
  OR U5199 ( .A(n4886), .B(n4885), .Z(n4887) );
  AND U5200 ( .A(n4888), .B(n4887), .Z(n4962) );
  OR U5201 ( .A(n4890), .B(n4889), .Z(n4894) );
  NANDN U5202 ( .A(n4892), .B(n4891), .Z(n4893) );
  AND U5203 ( .A(n4894), .B(n4893), .Z(n4961) );
  XNOR U5204 ( .A(n4962), .B(n4961), .Z(n4964) );
  XNOR U5205 ( .A(n4963), .B(n4964), .Z(n4958) );
  XNOR U5206 ( .A(n4908), .B(n4907), .Z(n4910) );
  OR U5207 ( .A(n4896), .B(n4895), .Z(n4900) );
  NANDN U5208 ( .A(n4898), .B(n4897), .Z(n4899) );
  AND U5209 ( .A(n4900), .B(n4899), .Z(n4909) );
  XOR U5210 ( .A(n4910), .B(n4909), .Z(n4915) );
  XNOR U5211 ( .A(n4916), .B(n4915), .Z(n5054) );
  XNOR U5212 ( .A(n5053), .B(n5054), .Z(n5055) );
  OR U5213 ( .A(n4902), .B(n4901), .Z(n4906) );
  OR U5214 ( .A(n4904), .B(n4903), .Z(n4905) );
  AND U5215 ( .A(n4906), .B(n4905), .Z(n5056) );
  XOR U5216 ( .A(n5049), .B(n5050), .Z(N122) );
  OR U5217 ( .A(n4908), .B(n4907), .Z(n4912) );
  OR U5218 ( .A(n4910), .B(n4909), .Z(n4911) );
  NAND U5219 ( .A(n4912), .B(n4911), .Z(n5068) );
  NANDN U5220 ( .A(n4914), .B(n4913), .Z(n4918) );
  OR U5221 ( .A(n4916), .B(n4915), .Z(n4917) );
  AND U5222 ( .A(n4918), .B(n4917), .Z(n5066) );
  OR U5223 ( .A(n4920), .B(n4919), .Z(n4924) );
  OR U5224 ( .A(n4922), .B(n4921), .Z(n4923) );
  AND U5225 ( .A(n4924), .B(n4923), .Z(n5199) );
  NANDN U5226 ( .A(n47), .B(y[248]), .Z(n5096) );
  XOR U5227 ( .A(n5095), .B(n5096), .Z(n5098) );
  NANDN U5228 ( .A(n8865), .B(y[226]), .Z(n5097) );
  XOR U5229 ( .A(n5098), .B(n5097), .Z(n5117) );
  OR U5230 ( .A(n4926), .B(n4925), .Z(n4930) );
  NAND U5231 ( .A(n4928), .B(n4927), .Z(n4929) );
  AND U5232 ( .A(n4930), .B(n4929), .Z(n5118) );
  XNOR U5233 ( .A(n5117), .B(n5118), .Z(n5120) );
  NANDN U5234 ( .A(n4932), .B(n4931), .Z(n4936) );
  NAND U5235 ( .A(n4934), .B(n4933), .Z(n4935) );
  AND U5236 ( .A(n4936), .B(n4935), .Z(n5119) );
  XOR U5237 ( .A(n5120), .B(n5119), .Z(n5198) );
  OR U5238 ( .A(n4938), .B(n4937), .Z(n4942) );
  OR U5239 ( .A(n4940), .B(n4939), .Z(n4941) );
  AND U5240 ( .A(n4942), .B(n4941), .Z(n5200) );
  XOR U5241 ( .A(n5201), .B(n5200), .Z(n5162) );
  OR U5242 ( .A(n4944), .B(n4943), .Z(n4948) );
  NANDN U5243 ( .A(n4946), .B(n4945), .Z(n4947) );
  AND U5244 ( .A(n4948), .B(n4947), .Z(n5159) );
  NANDN U5245 ( .A(n4950), .B(n4949), .Z(n4954) );
  OR U5246 ( .A(n4952), .B(n4951), .Z(n4953) );
  NAND U5247 ( .A(n4954), .B(n4953), .Z(n5160) );
  XOR U5248 ( .A(n5159), .B(n5160), .Z(n5161) );
  XOR U5249 ( .A(n5162), .B(n5161), .Z(n5074) );
  OR U5250 ( .A(n4956), .B(n4955), .Z(n4960) );
  OR U5251 ( .A(n4958), .B(n4957), .Z(n4959) );
  AND U5252 ( .A(n4960), .B(n4959), .Z(n5071) );
  OR U5253 ( .A(n4962), .B(n4961), .Z(n4966) );
  NANDN U5254 ( .A(n4964), .B(n4963), .Z(n4965) );
  AND U5255 ( .A(n4966), .B(n4965), .Z(n5155) );
  OR U5256 ( .A(n4968), .B(n4967), .Z(n4972) );
  NANDN U5257 ( .A(n4970), .B(n4969), .Z(n4971) );
  NAND U5258 ( .A(n4972), .B(n4971), .Z(n5205) );
  NANDN U5259 ( .A(n4974), .B(n4973), .Z(n4978) );
  OR U5260 ( .A(n4976), .B(n4975), .Z(n4977) );
  NAND U5261 ( .A(n4978), .B(n4977), .Z(n5204) );
  XOR U5262 ( .A(n5205), .B(n5204), .Z(n5206) );
  OR U5263 ( .A(n4980), .B(n4979), .Z(n4984) );
  OR U5264 ( .A(n4982), .B(n4981), .Z(n4983) );
  NAND U5265 ( .A(n4984), .B(n4983), .Z(n5207) );
  XNOR U5266 ( .A(n5206), .B(n5207), .Z(n5153) );
  OR U5267 ( .A(n4986), .B(n4985), .Z(n4990) );
  OR U5268 ( .A(n4988), .B(n4987), .Z(n4989) );
  NAND U5269 ( .A(n4990), .B(n4989), .Z(n5112) );
  NANDN U5270 ( .A(n4992), .B(n4991), .Z(n4996) );
  NANDN U5271 ( .A(n4994), .B(n4993), .Z(n4995) );
  NAND U5272 ( .A(n4996), .B(n4995), .Z(n5111) );
  XOR U5273 ( .A(n5112), .B(n5111), .Z(n5113) );
  ANDN U5274 ( .B(x[73]), .A(n5874), .Z(n5192) );
  NAND U5275 ( .A(x[70]), .B(y[244]), .Z(n5191) );
  NAND U5276 ( .A(x[72]), .B(y[242]), .Z(n5190) );
  XNOR U5277 ( .A(n5191), .B(n5190), .Z(n5193) );
  XNOR U5278 ( .A(n5192), .B(n5193), .Z(n5167) );
  AND U5279 ( .A(y[243]), .B(x[71]), .Z(n5165) );
  NAND U5280 ( .A(y[238]), .B(x[76]), .Z(n5130) );
  NAND U5281 ( .A(x[69]), .B(y[245]), .Z(n5129) );
  XNOR U5282 ( .A(n5130), .B(n5129), .Z(n5132) );
  XNOR U5283 ( .A(n5131), .B(n5132), .Z(n5166) );
  XNOR U5284 ( .A(n5165), .B(n5166), .Z(n5168) );
  XOR U5285 ( .A(n5113), .B(n5114), .Z(n5147) );
  OR U5286 ( .A(n4998), .B(n4997), .Z(n5002) );
  OR U5287 ( .A(n5000), .B(n4999), .Z(n5001) );
  AND U5288 ( .A(n5002), .B(n5001), .Z(n5148) );
  XOR U5289 ( .A(n5147), .B(n5148), .Z(n5150) );
  ANDN U5290 ( .B(y[246]), .A(n49), .Z(n5102) );
  XOR U5291 ( .A(n5003), .B(n5102), .Z(n5103) );
  XNOR U5292 ( .A(n5104), .B(n5103), .Z(n5083) );
  NAND U5293 ( .A(n5005), .B(n5004), .Z(n5009) );
  OR U5294 ( .A(n5007), .B(n5006), .Z(n5008) );
  NAND U5295 ( .A(n5009), .B(n5008), .Z(n5084) );
  XOR U5296 ( .A(n5083), .B(n5084), .Z(n5085) );
  NANDN U5297 ( .A(n8824), .B(y[231]), .Z(n5172) );
  NANDN U5298 ( .A(n5936), .B(x[75]), .Z(n5171) );
  XOR U5299 ( .A(n5172), .B(n5171), .Z(n5173) );
  NANDN U5300 ( .A(n48), .B(y[247]), .Z(n5174) );
  XOR U5301 ( .A(n5173), .B(n5174), .Z(n5086) );
  XNOR U5302 ( .A(n5085), .B(n5086), .Z(n5142) );
  ANDN U5303 ( .B(x[85]), .A(n5663), .Z(n5271) );
  NAND U5304 ( .A(n5010), .B(n5271), .Z(n5014) );
  OR U5305 ( .A(n5012), .B(n5011), .Z(n5013) );
  NAND U5306 ( .A(n5014), .B(n5013), .Z(n5078) );
  NAND U5307 ( .A(x[86]), .B(y[228]), .Z(n5092) );
  ANDN U5308 ( .B(x[87]), .A(n5714), .Z(n5090) );
  XOR U5309 ( .A(n5015), .B(n5090), .Z(n5091) );
  XNOR U5310 ( .A(n5092), .B(n5091), .Z(n5077) );
  XNOR U5311 ( .A(n5078), .B(n5077), .Z(n5080) );
  NAND U5312 ( .A(y[230]), .B(x[84]), .Z(n5187) );
  ANDN U5313 ( .B(y[229]), .A(n8827), .Z(n5185) );
  XOR U5314 ( .A(n5184), .B(n5185), .Z(n5186) );
  XNOR U5315 ( .A(n5187), .B(n5186), .Z(n5079) );
  XNOR U5316 ( .A(n5080), .B(n5079), .Z(n5141) );
  XNOR U5317 ( .A(n5142), .B(n5141), .Z(n5144) );
  ANDN U5318 ( .B(o[57]), .A(n5016), .Z(n5181) );
  AND U5319 ( .A(y[236]), .B(x[78]), .Z(n5179) );
  AND U5320 ( .A(y[249]), .B(x[65]), .Z(n5178) );
  XNOR U5321 ( .A(n5179), .B(n5178), .Z(n5180) );
  XNOR U5322 ( .A(n5181), .B(n5180), .Z(n5125) );
  NANDN U5323 ( .A(n45), .B(y[250]), .Z(n5136) );
  NANDN U5324 ( .A(n5905), .B(x[90]), .Z(n5135) );
  XOR U5325 ( .A(n5136), .B(n5135), .Z(n5137) );
  NANDN U5326 ( .A(n8928), .B(y[225]), .Z(n5197) );
  XOR U5327 ( .A(o[58]), .B(n5197), .Z(n5138) );
  XNOR U5328 ( .A(n5137), .B(n5138), .Z(n5123) );
  NAND U5329 ( .A(n5018), .B(n5017), .Z(n5022) );
  NANDN U5330 ( .A(n5020), .B(n5019), .Z(n5021) );
  AND U5331 ( .A(n5022), .B(n5021), .Z(n5124) );
  XNOR U5332 ( .A(n5123), .B(n5124), .Z(n5126) );
  XNOR U5333 ( .A(n5125), .B(n5126), .Z(n5109) );
  NAND U5334 ( .A(n5024), .B(n5023), .Z(n5028) );
  OR U5335 ( .A(n5026), .B(n5025), .Z(n5027) );
  NAND U5336 ( .A(n5028), .B(n5027), .Z(n5108) );
  NAND U5337 ( .A(n5030), .B(n5029), .Z(n5034) );
  NANDN U5338 ( .A(n5032), .B(n5031), .Z(n5033) );
  AND U5339 ( .A(n5034), .B(n5033), .Z(n5107) );
  XNOR U5340 ( .A(n5108), .B(n5107), .Z(n5110) );
  XOR U5341 ( .A(n5109), .B(n5110), .Z(n5143) );
  XNOR U5342 ( .A(n5144), .B(n5143), .Z(n5149) );
  XOR U5343 ( .A(n5150), .B(n5149), .Z(n5154) );
  XNOR U5344 ( .A(n5153), .B(n5154), .Z(n5156) );
  XOR U5345 ( .A(n5155), .B(n5156), .Z(n5072) );
  XNOR U5346 ( .A(n5071), .B(n5072), .Z(n5073) );
  XNOR U5347 ( .A(n5074), .B(n5073), .Z(n5213) );
  OR U5348 ( .A(n5036), .B(n5035), .Z(n5040) );
  NAND U5349 ( .A(n5038), .B(n5037), .Z(n5039) );
  NAND U5350 ( .A(n5040), .B(n5039), .Z(n5211) );
  OR U5351 ( .A(n5042), .B(n5041), .Z(n5046) );
  OR U5352 ( .A(n5044), .B(n5043), .Z(n5045) );
  AND U5353 ( .A(n5046), .B(n5045), .Z(n5210) );
  XOR U5354 ( .A(n5211), .B(n5210), .Z(n5212) );
  XNOR U5355 ( .A(n5213), .B(n5212), .Z(n5065) );
  XOR U5356 ( .A(n5066), .B(n5065), .Z(n5067) );
  XNOR U5357 ( .A(n5068), .B(n5067), .Z(n5062) );
  NANDN U5358 ( .A(n5048), .B(n5047), .Z(n5052) );
  NANDN U5359 ( .A(n5050), .B(n5049), .Z(n5051) );
  NAND U5360 ( .A(n5052), .B(n5051), .Z(n5059) );
  OR U5361 ( .A(n5054), .B(n5053), .Z(n5058) );
  OR U5362 ( .A(n5056), .B(n5055), .Z(n5057) );
  AND U5363 ( .A(n5058), .B(n5057), .Z(n5060) );
  XNOR U5364 ( .A(n5059), .B(n5060), .Z(n5061) );
  XOR U5365 ( .A(n5062), .B(n5061), .Z(N123) );
  NANDN U5366 ( .A(n5060), .B(n5059), .Z(n5064) );
  NANDN U5367 ( .A(n5062), .B(n5061), .Z(n5063) );
  NAND U5368 ( .A(n5064), .B(n5063), .Z(n5216) );
  NANDN U5369 ( .A(n5066), .B(n5065), .Z(n5070) );
  OR U5370 ( .A(n5068), .B(n5067), .Z(n5069) );
  AND U5371 ( .A(n5070), .B(n5069), .Z(n5217) );
  XNOR U5372 ( .A(n5216), .B(n5217), .Z(n5218) );
  OR U5373 ( .A(n5072), .B(n5071), .Z(n5076) );
  OR U5374 ( .A(n5074), .B(n5073), .Z(n5075) );
  AND U5375 ( .A(n5076), .B(n5075), .Z(n5222) );
  OR U5376 ( .A(n5078), .B(n5077), .Z(n5082) );
  OR U5377 ( .A(n5080), .B(n5079), .Z(n5081) );
  NAND U5378 ( .A(n5082), .B(n5081), .Z(n5241) );
  OR U5379 ( .A(n5084), .B(n5083), .Z(n5088) );
  NANDN U5380 ( .A(n5086), .B(n5085), .Z(n5087) );
  NAND U5381 ( .A(n5088), .B(n5087), .Z(n5253) );
  NANDN U5382 ( .A(n5090), .B(n5089), .Z(n5094) );
  NAND U5383 ( .A(n5092), .B(n5091), .Z(n5093) );
  AND U5384 ( .A(n5094), .B(n5093), .Z(n5320) );
  NANDN U5385 ( .A(n5096), .B(n5095), .Z(n5100) );
  OR U5386 ( .A(n5098), .B(n5097), .Z(n5099) );
  NAND U5387 ( .A(n5100), .B(n5099), .Z(n5321) );
  NANDN U5388 ( .A(n5102), .B(n5101), .Z(n5106) );
  NANDN U5389 ( .A(n5104), .B(n5103), .Z(n5105) );
  AND U5390 ( .A(n5106), .B(n5105), .Z(n5314) );
  AND U5391 ( .A(y[242]), .B(x[73]), .Z(n5274) );
  AND U5392 ( .A(y[233]), .B(x[82]), .Z(n5272) );
  XOR U5393 ( .A(n5271), .B(n5272), .Z(n5273) );
  XOR U5394 ( .A(n5274), .B(n5273), .Z(n5315) );
  AND U5395 ( .A(y[251]), .B(x[64]), .Z(n5261) );
  NANDN U5396 ( .A(n8901), .B(y[225]), .Z(n5270) );
  XNOR U5397 ( .A(n5270), .B(o[59]), .Z(n5259) );
  NAND U5398 ( .A(y[224]), .B(x[91]), .Z(n5258) );
  XOR U5399 ( .A(n5259), .B(n5258), .Z(n5260) );
  XOR U5400 ( .A(n5261), .B(n5260), .Z(n5316) );
  XNOR U5401 ( .A(n5253), .B(n5252), .Z(n5254) );
  XOR U5402 ( .A(n5254), .B(n5255), .Z(n5240) );
  XNOR U5403 ( .A(n5241), .B(n5240), .Z(n5243) );
  OR U5404 ( .A(n5112), .B(n5111), .Z(n5116) );
  NANDN U5405 ( .A(n5114), .B(n5113), .Z(n5115) );
  NAND U5406 ( .A(n5116), .B(n5115), .Z(n5242) );
  XOR U5407 ( .A(n5243), .B(n5242), .Z(n5375) );
  NAND U5408 ( .A(n5118), .B(n5117), .Z(n5122) );
  NANDN U5409 ( .A(n5120), .B(n5119), .Z(n5121) );
  NAND U5410 ( .A(n5122), .B(n5121), .Z(n5248) );
  NAND U5411 ( .A(n5124), .B(n5123), .Z(n5128) );
  NANDN U5412 ( .A(n5126), .B(n5125), .Z(n5127) );
  NAND U5413 ( .A(n5128), .B(n5127), .Z(n5247) );
  AND U5414 ( .A(y[239]), .B(x[76]), .Z(n5352) );
  AND U5415 ( .A(y[238]), .B(x[77]), .Z(n5351) );
  XNOR U5416 ( .A(n5352), .B(n5351), .Z(n5354) );
  AND U5417 ( .A(y[240]), .B(x[75]), .Z(n5336) );
  AND U5418 ( .A(y[235]), .B(x[80]), .Z(n5334) );
  XOR U5419 ( .A(n5333), .B(n5334), .Z(n5335) );
  XOR U5420 ( .A(n5336), .B(n5335), .Z(n5353) );
  XOR U5421 ( .A(n5354), .B(n5353), .Z(n5298) );
  AND U5422 ( .A(y[248]), .B(x[67]), .Z(n5360) );
  AND U5423 ( .A(y[249]), .B(x[66]), .Z(n5358) );
  AND U5424 ( .A(y[236]), .B(x[79]), .Z(n5357) );
  XNOR U5425 ( .A(n5358), .B(n5357), .Z(n5359) );
  XNOR U5426 ( .A(n5360), .B(n5359), .Z(n5296) );
  AND U5427 ( .A(y[245]), .B(x[70]), .Z(n5281) );
  AND U5428 ( .A(y[226]), .B(x[89]), .Z(n5279) );
  AND U5429 ( .A(y[232]), .B(x[83]), .Z(n5278) );
  XNOR U5430 ( .A(n5279), .B(n5278), .Z(n5280) );
  XOR U5431 ( .A(n5281), .B(n5280), .Z(n5297) );
  XOR U5432 ( .A(n5296), .B(n5297), .Z(n5299) );
  NAND U5433 ( .A(n5130), .B(n5129), .Z(n5134) );
  OR U5434 ( .A(n5132), .B(n5131), .Z(n5133) );
  AND U5435 ( .A(n5134), .B(n5133), .Z(n5326) );
  OR U5436 ( .A(n5136), .B(n5135), .Z(n5140) );
  NANDN U5437 ( .A(n5138), .B(n5137), .Z(n5139) );
  NAND U5438 ( .A(n5140), .B(n5139), .Z(n5327) );
  XOR U5439 ( .A(n5247), .B(n5246), .Z(n5249) );
  XOR U5440 ( .A(n5248), .B(n5249), .Z(n5234) );
  NAND U5441 ( .A(n5142), .B(n5141), .Z(n5146) );
  NANDN U5442 ( .A(n5144), .B(n5143), .Z(n5145) );
  AND U5443 ( .A(n5146), .B(n5145), .Z(n5235) );
  XNOR U5444 ( .A(n5234), .B(n5235), .Z(n5237) );
  NANDN U5445 ( .A(n5148), .B(n5147), .Z(n5152) );
  NANDN U5446 ( .A(n5150), .B(n5149), .Z(n5151) );
  AND U5447 ( .A(n5152), .B(n5151), .Z(n5236) );
  XOR U5448 ( .A(n5237), .B(n5236), .Z(n5376) );
  XNOR U5449 ( .A(n5375), .B(n5376), .Z(n5378) );
  OR U5450 ( .A(n5154), .B(n5153), .Z(n5158) );
  OR U5451 ( .A(n5156), .B(n5155), .Z(n5157) );
  NAND U5452 ( .A(n5158), .B(n5157), .Z(n5377) );
  XOR U5453 ( .A(n5378), .B(n5377), .Z(n5371) );
  OR U5454 ( .A(n5160), .B(n5159), .Z(n5164) );
  NANDN U5455 ( .A(n5162), .B(n5161), .Z(n5163) );
  AND U5456 ( .A(n5164), .B(n5163), .Z(n5369) );
  OR U5457 ( .A(n5166), .B(n5165), .Z(n5170) );
  OR U5458 ( .A(n5168), .B(n5167), .Z(n5169) );
  AND U5459 ( .A(n5170), .B(n5169), .Z(n5230) );
  OR U5460 ( .A(n5172), .B(n5171), .Z(n5176) );
  NANDN U5461 ( .A(n5174), .B(n5173), .Z(n5175) );
  NAND U5462 ( .A(n5176), .B(n5175), .Z(n5305) );
  AND U5463 ( .A(y[229]), .B(x[86]), .Z(n5342) );
  AND U5464 ( .A(y[228]), .B(x[87]), .Z(n5340) );
  AND U5465 ( .A(y[243]), .B(x[72]), .Z(n5339) );
  XNOR U5466 ( .A(n5340), .B(n5339), .Z(n5341) );
  XNOR U5467 ( .A(n5342), .B(n5341), .Z(n5302) );
  NAND U5468 ( .A(x[71]), .B(y[244]), .Z(n5287) );
  ANDN U5469 ( .B(x[88]), .A(n5714), .Z(n5285) );
  XOR U5470 ( .A(n5177), .B(n5285), .Z(n5286) );
  XOR U5471 ( .A(n5287), .B(n5286), .Z(n5303) );
  XNOR U5472 ( .A(n5302), .B(n5303), .Z(n5304) );
  XOR U5473 ( .A(n5305), .B(n5304), .Z(n5228) );
  OR U5474 ( .A(n5179), .B(n5178), .Z(n5183) );
  OR U5475 ( .A(n5181), .B(n5180), .Z(n5182) );
  NAND U5476 ( .A(n5183), .B(n5182), .Z(n5291) );
  OR U5477 ( .A(n5185), .B(n5184), .Z(n5189) );
  NAND U5478 ( .A(n5187), .B(n5186), .Z(n5188) );
  AND U5479 ( .A(n5189), .B(n5188), .Z(n5290) );
  XNOR U5480 ( .A(n5291), .B(n5290), .Z(n5292) );
  NAND U5481 ( .A(n5191), .B(n5190), .Z(n5195) );
  OR U5482 ( .A(n5193), .B(n5192), .Z(n5194) );
  NAND U5483 ( .A(n5195), .B(n5194), .Z(n5311) );
  NANDN U5484 ( .A(n50), .B(y[246]), .Z(n5267) );
  NANDN U5485 ( .A(n49), .B(y[247]), .Z(n5265) );
  NANDN U5486 ( .A(n5196), .B(x[81]), .Z(n5264) );
  XOR U5487 ( .A(n5265), .B(n5264), .Z(n5266) );
  XOR U5488 ( .A(n5267), .B(n5266), .Z(n5309) );
  AND U5489 ( .A(y[237]), .B(x[78]), .Z(n5348) );
  ANDN U5490 ( .B(o[58]), .A(n5197), .Z(n5345) );
  AND U5491 ( .A(y[250]), .B(x[65]), .Z(n5346) );
  XNOR U5492 ( .A(n5348), .B(n5347), .Z(n5308) );
  XNOR U5493 ( .A(n5309), .B(n5308), .Z(n5310) );
  XOR U5494 ( .A(n5311), .B(n5310), .Z(n5293) );
  XNOR U5495 ( .A(n5292), .B(n5293), .Z(n5229) );
  XNOR U5496 ( .A(n5228), .B(n5229), .Z(n5231) );
  XOR U5497 ( .A(n5230), .B(n5231), .Z(n5363) );
  OR U5498 ( .A(n5199), .B(n5198), .Z(n5203) );
  OR U5499 ( .A(n5201), .B(n5200), .Z(n5202) );
  AND U5500 ( .A(n5203), .B(n5202), .Z(n5364) );
  XNOR U5501 ( .A(n5363), .B(n5364), .Z(n5366) );
  OR U5502 ( .A(n5205), .B(n5204), .Z(n5209) );
  NANDN U5503 ( .A(n5207), .B(n5206), .Z(n5208) );
  NAND U5504 ( .A(n5209), .B(n5208), .Z(n5365) );
  XOR U5505 ( .A(n5366), .B(n5365), .Z(n5370) );
  XNOR U5506 ( .A(n5369), .B(n5370), .Z(n5372) );
  XOR U5507 ( .A(n5371), .B(n5372), .Z(n5223) );
  XNOR U5508 ( .A(n5222), .B(n5223), .Z(n5224) );
  OR U5509 ( .A(n5211), .B(n5210), .Z(n5215) );
  NANDN U5510 ( .A(n5213), .B(n5212), .Z(n5214) );
  AND U5511 ( .A(n5215), .B(n5214), .Z(n5225) );
  XOR U5512 ( .A(n5218), .B(n5219), .Z(N124) );
  NANDN U5513 ( .A(n5217), .B(n5216), .Z(n5221) );
  NANDN U5514 ( .A(n5219), .B(n5218), .Z(n5220) );
  NAND U5515 ( .A(n5221), .B(n5220), .Z(n5381) );
  OR U5516 ( .A(n5223), .B(n5222), .Z(n5227) );
  OR U5517 ( .A(n5225), .B(n5224), .Z(n5226) );
  AND U5518 ( .A(n5227), .B(n5226), .Z(n5382) );
  XNOR U5519 ( .A(n5381), .B(n5382), .Z(n5383) );
  OR U5520 ( .A(n5229), .B(n5228), .Z(n5233) );
  OR U5521 ( .A(n5231), .B(n5230), .Z(n5232) );
  AND U5522 ( .A(n5233), .B(n5232), .Z(n5543) );
  OR U5523 ( .A(n5235), .B(n5234), .Z(n5239) );
  OR U5524 ( .A(n5237), .B(n5236), .Z(n5238) );
  NAND U5525 ( .A(n5239), .B(n5238), .Z(n5541) );
  OR U5526 ( .A(n5241), .B(n5240), .Z(n5245) );
  OR U5527 ( .A(n5243), .B(n5242), .Z(n5244) );
  NAND U5528 ( .A(n5245), .B(n5244), .Z(n5540) );
  XOR U5529 ( .A(n5541), .B(n5540), .Z(n5542) );
  XNOR U5530 ( .A(n5543), .B(n5542), .Z(n5548) );
  NANDN U5531 ( .A(n5247), .B(n5246), .Z(n5251) );
  OR U5532 ( .A(n5249), .B(n5248), .Z(n5250) );
  NAND U5533 ( .A(n5251), .B(n5250), .Z(n5528) );
  NANDN U5534 ( .A(n5253), .B(n5252), .Z(n5257) );
  NAND U5535 ( .A(n5255), .B(n5254), .Z(n5256) );
  AND U5536 ( .A(n5257), .B(n5256), .Z(n5529) );
  XNOR U5537 ( .A(n5528), .B(n5529), .Z(n5530) );
  NANDN U5538 ( .A(n5259), .B(n5258), .Z(n5263) );
  OR U5539 ( .A(n5261), .B(n5260), .Z(n5262) );
  AND U5540 ( .A(n5263), .B(n5262), .Z(n5510) );
  OR U5541 ( .A(n5265), .B(n5264), .Z(n5269) );
  NANDN U5542 ( .A(n5267), .B(n5266), .Z(n5268) );
  NAND U5543 ( .A(n5269), .B(n5268), .Z(n5511) );
  ANDN U5544 ( .B(o[59]), .A(n5270), .Z(n5474) );
  AND U5545 ( .A(y[224]), .B(x[92]), .Z(n5475) );
  XNOR U5546 ( .A(n5474), .B(n5475), .Z(n5477) );
  AND U5547 ( .A(y[252]), .B(x[64]), .Z(n5476) );
  XNOR U5548 ( .A(n5477), .B(n5476), .Z(n5458) );
  OR U5549 ( .A(n5272), .B(n5271), .Z(n5276) );
  NANDN U5550 ( .A(n5274), .B(n5273), .Z(n5275) );
  AND U5551 ( .A(n5276), .B(n5275), .Z(n5456) );
  AND U5552 ( .A(y[243]), .B(x[73]), .Z(n5467) );
  AND U5553 ( .A(y[244]), .B(x[72]), .Z(n5468) );
  XNOR U5554 ( .A(n5467), .B(n5468), .Z(n5470) );
  AND U5555 ( .A(y[242]), .B(x[74]), .Z(n5469) );
  XOR U5556 ( .A(n5470), .B(n5469), .Z(n5455) );
  XOR U5557 ( .A(n5456), .B(n5455), .Z(n5457) );
  XNOR U5558 ( .A(n5458), .B(n5457), .Z(n5513) );
  XOR U5559 ( .A(n5512), .B(n5513), .Z(n5483) );
  NANDN U5560 ( .A(n50), .B(y[247]), .Z(n5413) );
  AND U5561 ( .A(y[232]), .B(x[84]), .Z(n5412) );
  NANDN U5562 ( .A(n44), .B(x[85]), .Z(n5411) );
  XOR U5563 ( .A(n5412), .B(n5411), .Z(n5414) );
  XNOR U5564 ( .A(n5413), .B(n5414), .Z(n5505) );
  AND U5565 ( .A(y[229]), .B(x[87]), .Z(n5432) );
  NANDN U5566 ( .A(n48), .B(y[249]), .Z(n5431) );
  XOR U5567 ( .A(n5432), .B(n5431), .Z(n5434) );
  XNOR U5568 ( .A(n5277), .B(n5434), .Z(n5504) );
  XOR U5569 ( .A(n5505), .B(n5504), .Z(n5506) );
  OR U5570 ( .A(n5279), .B(n5278), .Z(n5283) );
  OR U5571 ( .A(n5281), .B(n5280), .Z(n5282) );
  NAND U5572 ( .A(n5283), .B(n5282), .Z(n5507) );
  XNOR U5573 ( .A(n5506), .B(n5507), .Z(n5480) );
  AND U5574 ( .A(y[251]), .B(x[65]), .Z(n5394) );
  NANDN U5575 ( .A(n5714), .B(x[89]), .Z(n5393) );
  XOR U5576 ( .A(n5394), .B(n5393), .Z(n5396) );
  XOR U5577 ( .A(n5395), .B(n5396), .Z(n5501) );
  NANDN U5578 ( .A(n8890), .B(y[236]), .Z(n5401) );
  AND U5579 ( .A(y[250]), .B(x[66]), .Z(n5400) );
  NANDN U5580 ( .A(n8865), .B(y[228]), .Z(n5399) );
  XOR U5581 ( .A(n5400), .B(n5399), .Z(n5402) );
  XNOR U5582 ( .A(n5401), .B(n5402), .Z(n5498) );
  NANDN U5583 ( .A(n5285), .B(n5284), .Z(n5289) );
  NAND U5584 ( .A(n5287), .B(n5286), .Z(n5288) );
  NAND U5585 ( .A(n5289), .B(n5288), .Z(n5499) );
  XOR U5586 ( .A(n5498), .B(n5499), .Z(n5500) );
  XNOR U5587 ( .A(n5501), .B(n5500), .Z(n5481) );
  XOR U5588 ( .A(n5483), .B(n5482), .Z(n5534) );
  NANDN U5589 ( .A(n5291), .B(n5290), .Z(n5295) );
  NANDN U5590 ( .A(n5293), .B(n5292), .Z(n5294) );
  NAND U5591 ( .A(n5295), .B(n5294), .Z(n5489) );
  NANDN U5592 ( .A(n5297), .B(n5296), .Z(n5301) );
  OR U5593 ( .A(n5299), .B(n5298), .Z(n5300) );
  NAND U5594 ( .A(n5301), .B(n5300), .Z(n5487) );
  NANDN U5595 ( .A(n5303), .B(n5302), .Z(n5307) );
  NAND U5596 ( .A(n5305), .B(n5304), .Z(n5306) );
  NAND U5597 ( .A(n5307), .B(n5306), .Z(n5486) );
  XOR U5598 ( .A(n5489), .B(n5488), .Z(n5535) );
  NANDN U5599 ( .A(n5309), .B(n5308), .Z(n5313) );
  NANDN U5600 ( .A(n5311), .B(n5310), .Z(n5312) );
  AND U5601 ( .A(n5313), .B(n5312), .Z(n5516) );
  OR U5602 ( .A(n5315), .B(n5314), .Z(n5319) );
  NANDN U5603 ( .A(n5317), .B(n5316), .Z(n5318) );
  NAND U5604 ( .A(n5319), .B(n5318), .Z(n5517) );
  OR U5605 ( .A(n5321), .B(n5320), .Z(n5325) );
  NANDN U5606 ( .A(n5323), .B(n5322), .Z(n5324) );
  NAND U5607 ( .A(n5325), .B(n5324), .Z(n5519) );
  XOR U5608 ( .A(n5518), .B(n5519), .Z(n5524) );
  OR U5609 ( .A(n5327), .B(n5326), .Z(n5331) );
  NANDN U5610 ( .A(n5329), .B(n5328), .Z(n5330) );
  NAND U5611 ( .A(n5331), .B(n5330), .Z(n5522) );
  NANDN U5612 ( .A(n8901), .B(y[226]), .Z(n5438) );
  ANDN U5613 ( .B(x[79]), .A(n5332), .Z(n5437) );
  XNOR U5614 ( .A(n5438), .B(n5437), .Z(n5440) );
  NAND U5615 ( .A(x[91]), .B(y[225]), .Z(n5614) );
  XNOR U5616 ( .A(n5614), .B(o[60]), .Z(n5439) );
  XNOR U5617 ( .A(n5440), .B(n5439), .Z(n5428) );
  OR U5618 ( .A(n5334), .B(n5333), .Z(n5338) );
  NANDN U5619 ( .A(n5336), .B(n5335), .Z(n5337) );
  NAND U5620 ( .A(n5338), .B(n5337), .Z(n5426) );
  AND U5621 ( .A(y[245]), .B(x[71]), .Z(n5407) );
  AND U5622 ( .A(y[241]), .B(x[75]), .Z(n5405) );
  AND U5623 ( .A(y[240]), .B(x[76]), .Z(n5406) );
  XNOR U5624 ( .A(n5405), .B(n5406), .Z(n5408) );
  XOR U5625 ( .A(n5407), .B(n5408), .Z(n5425) );
  XNOR U5626 ( .A(n5426), .B(n5425), .Z(n5427) );
  XNOR U5627 ( .A(n5428), .B(n5427), .Z(n5492) );
  OR U5628 ( .A(n5340), .B(n5339), .Z(n5344) );
  OR U5629 ( .A(n5342), .B(n5341), .Z(n5343) );
  AND U5630 ( .A(n5344), .B(n5343), .Z(n5443) );
  AND U5631 ( .A(y[246]), .B(x[70]), .Z(n5421) );
  AND U5632 ( .A(y[233]), .B(x[83]), .Z(n5420) );
  XNOR U5633 ( .A(n5419), .B(n5420), .Z(n5422) );
  XNOR U5634 ( .A(n5421), .B(n5422), .Z(n5444) );
  XOR U5635 ( .A(n5443), .B(n5444), .Z(n5446) );
  NANDN U5636 ( .A(n8626), .B(y[235]), .Z(n5463) );
  AND U5637 ( .A(y[248]), .B(x[68]), .Z(n5462) );
  NANDN U5638 ( .A(n5663), .B(x[86]), .Z(n5461) );
  XOR U5639 ( .A(n5462), .B(n5461), .Z(n5464) );
  XNOR U5640 ( .A(n5463), .B(n5464), .Z(n5445) );
  XNOR U5641 ( .A(n5446), .B(n5445), .Z(n5493) );
  XOR U5642 ( .A(n5492), .B(n5493), .Z(n5495) );
  OR U5643 ( .A(n5346), .B(n5345), .Z(n5350) );
  OR U5644 ( .A(n5348), .B(n5347), .Z(n5349) );
  AND U5645 ( .A(n5350), .B(n5349), .Z(n5452) );
  OR U5646 ( .A(n5352), .B(n5351), .Z(n5356) );
  OR U5647 ( .A(n5354), .B(n5353), .Z(n5355) );
  AND U5648 ( .A(n5356), .B(n5355), .Z(n5449) );
  OR U5649 ( .A(n5358), .B(n5357), .Z(n5362) );
  OR U5650 ( .A(n5360), .B(n5359), .Z(n5361) );
  AND U5651 ( .A(n5362), .B(n5361), .Z(n5450) );
  XNOR U5652 ( .A(n5449), .B(n5450), .Z(n5451) );
  XOR U5653 ( .A(n5452), .B(n5451), .Z(n5494) );
  XOR U5654 ( .A(n5495), .B(n5494), .Z(n5523) );
  XOR U5655 ( .A(n5522), .B(n5523), .Z(n5525) );
  XOR U5656 ( .A(n5524), .B(n5525), .Z(n5536) );
  XNOR U5657 ( .A(n5537), .B(n5536), .Z(n5531) );
  XNOR U5658 ( .A(n5530), .B(n5531), .Z(n5546) );
  OR U5659 ( .A(n5364), .B(n5363), .Z(n5368) );
  OR U5660 ( .A(n5366), .B(n5365), .Z(n5367) );
  AND U5661 ( .A(n5368), .B(n5367), .Z(n5547) );
  XNOR U5662 ( .A(n5546), .B(n5547), .Z(n5549) );
  XNOR U5663 ( .A(n5548), .B(n5549), .Z(n5387) );
  OR U5664 ( .A(n5370), .B(n5369), .Z(n5374) );
  NANDN U5665 ( .A(n5372), .B(n5371), .Z(n5373) );
  AND U5666 ( .A(n5374), .B(n5373), .Z(n5388) );
  XOR U5667 ( .A(n5387), .B(n5388), .Z(n5390) );
  OR U5668 ( .A(n5376), .B(n5375), .Z(n5380) );
  OR U5669 ( .A(n5378), .B(n5377), .Z(n5379) );
  AND U5670 ( .A(n5380), .B(n5379), .Z(n5389) );
  XOR U5671 ( .A(n5390), .B(n5389), .Z(n5384) );
  XNOR U5672 ( .A(n5383), .B(n5384), .Z(N125) );
  NANDN U5673 ( .A(n5382), .B(n5381), .Z(n5386) );
  NAND U5674 ( .A(n5384), .B(n5383), .Z(n5385) );
  NAND U5675 ( .A(n5386), .B(n5385), .Z(n5552) );
  NANDN U5676 ( .A(n5388), .B(n5387), .Z(n5392) );
  OR U5677 ( .A(n5390), .B(n5389), .Z(n5391) );
  AND U5678 ( .A(n5392), .B(n5391), .Z(n5553) );
  XNOR U5679 ( .A(n5552), .B(n5553), .Z(n5554) );
  NANDN U5680 ( .A(n5394), .B(n5393), .Z(n5398) );
  OR U5681 ( .A(n5396), .B(n5395), .Z(n5397) );
  AND U5682 ( .A(n5398), .B(n5397), .Z(n5693) );
  NANDN U5683 ( .A(n5400), .B(n5399), .Z(n5404) );
  NANDN U5684 ( .A(n5402), .B(n5401), .Z(n5403) );
  AND U5685 ( .A(n5404), .B(n5403), .Z(n5690) );
  ANDN U5686 ( .B(x[87]), .A(n5663), .Z(n5625) );
  IV U5687 ( .A(n5625), .Z(n5928) );
  AND U5688 ( .A(y[229]), .B(x[88]), .Z(n5626) );
  XOR U5689 ( .A(n5928), .B(n5626), .Z(n5628) );
  AND U5690 ( .A(y[240]), .B(x[77]), .Z(n5627) );
  XNOR U5691 ( .A(n5628), .B(n5627), .Z(n5597) );
  OR U5692 ( .A(n5406), .B(n5405), .Z(n5410) );
  OR U5693 ( .A(n5408), .B(n5407), .Z(n5409) );
  AND U5694 ( .A(n5410), .B(n5409), .Z(n5595) );
  AND U5695 ( .A(y[242]), .B(x[75]), .Z(n5619) );
  AND U5696 ( .A(y[236]), .B(x[81]), .Z(n5620) );
  XNOR U5697 ( .A(n5619), .B(n5620), .Z(n5622) );
  AND U5698 ( .A(y[250]), .B(x[67]), .Z(n5621) );
  XOR U5699 ( .A(n5622), .B(n5621), .Z(n5594) );
  XOR U5700 ( .A(n5595), .B(n5594), .Z(n5596) );
  XNOR U5701 ( .A(n5597), .B(n5596), .Z(n5691) );
  XNOR U5702 ( .A(n5690), .B(n5691), .Z(n5692) );
  AND U5703 ( .A(y[235]), .B(x[82]), .Z(n5606) );
  AND U5704 ( .A(y[234]), .B(x[83]), .Z(n5607) );
  XNOR U5705 ( .A(n5606), .B(n5607), .Z(n5609) );
  AND U5706 ( .A(y[251]), .B(x[66]), .Z(n5608) );
  XNOR U5707 ( .A(n5609), .B(n5608), .Z(n5643) );
  NANDN U5708 ( .A(n5412), .B(n5411), .Z(n5416) );
  NANDN U5709 ( .A(n5414), .B(n5413), .Z(n5415) );
  AND U5710 ( .A(n5416), .B(n5415), .Z(n5641) );
  NAND U5711 ( .A(y[225]), .B(o[60]), .Z(n5417) );
  XNOR U5712 ( .A(y[226]), .B(n5417), .Z(n5418) );
  NAND U5713 ( .A(x[91]), .B(n5418), .Z(n5613) );
  AND U5714 ( .A(y[237]), .B(x[80]), .Z(n5612) );
  XOR U5715 ( .A(n5613), .B(n5612), .Z(n5640) );
  XOR U5716 ( .A(n5641), .B(n5640), .Z(n5642) );
  XNOR U5717 ( .A(n5643), .B(n5642), .Z(n5673) );
  OR U5718 ( .A(n5420), .B(n5419), .Z(n5424) );
  OR U5719 ( .A(n5422), .B(n5421), .Z(n5423) );
  NAND U5720 ( .A(n5424), .B(n5423), .Z(n5705) );
  AND U5721 ( .A(y[225]), .B(x[92]), .Z(n5662) );
  XOR U5722 ( .A(o[61]), .B(n5662), .Z(n5719) );
  AND U5723 ( .A(y[224]), .B(x[93]), .Z(n5720) );
  XNOR U5724 ( .A(n5719), .B(n5720), .Z(n5722) );
  AND U5725 ( .A(y[253]), .B(x[64]), .Z(n5721) );
  XOR U5726 ( .A(n5722), .B(n5721), .Z(n5702) );
  AND U5727 ( .A(y[228]), .B(x[89]), .Z(n5646) );
  AND U5728 ( .A(y[227]), .B(x[90]), .Z(n5647) );
  XNOR U5729 ( .A(n5646), .B(n5647), .Z(n5649) );
  AND U5730 ( .A(y[239]), .B(x[78]), .Z(n5648) );
  XOR U5731 ( .A(n5649), .B(n5648), .Z(n5703) );
  XNOR U5732 ( .A(n5702), .B(n5703), .Z(n5704) );
  XOR U5733 ( .A(n5705), .B(n5704), .Z(n5672) );
  XNOR U5734 ( .A(n5673), .B(n5672), .Z(n5674) );
  XOR U5735 ( .A(n5675), .B(n5674), .Z(n5666) );
  OR U5736 ( .A(n5426), .B(n5425), .Z(n5430) );
  OR U5737 ( .A(n5428), .B(n5427), .Z(n5429) );
  AND U5738 ( .A(n5430), .B(n5429), .Z(n5667) );
  XNOR U5739 ( .A(n5666), .B(n5667), .Z(n5669) );
  NANDN U5740 ( .A(n5432), .B(n5431), .Z(n5436) );
  OR U5741 ( .A(n5434), .B(n5433), .Z(n5435) );
  AND U5742 ( .A(n5436), .B(n5435), .Z(n5588) );
  NANDN U5743 ( .A(n5438), .B(n5437), .Z(n5442) );
  NAND U5744 ( .A(n5440), .B(n5439), .Z(n5441) );
  NAND U5745 ( .A(n5442), .B(n5441), .Z(n5589) );
  XNOR U5746 ( .A(n5588), .B(n5589), .Z(n5590) );
  AND U5747 ( .A(y[245]), .B(x[72]), .Z(n5631) );
  AND U5748 ( .A(y[246]), .B(x[71]), .Z(n5632) );
  XNOR U5749 ( .A(n5631), .B(n5632), .Z(n5634) );
  AND U5750 ( .A(y[247]), .B(x[70]), .Z(n5633) );
  XNOR U5751 ( .A(n5634), .B(n5633), .Z(n5711) );
  ANDN U5752 ( .B(y[244]), .A(n54), .Z(n5708) );
  IV U5753 ( .A(n5708), .Z(n5823) );
  AND U5754 ( .A(y[248]), .B(x[69]), .Z(n5600) );
  AND U5755 ( .A(y[243]), .B(x[74]), .Z(n5601) );
  XNOR U5756 ( .A(n5600), .B(n5601), .Z(n5603) );
  AND U5757 ( .A(y[249]), .B(x[68]), .Z(n5602) );
  XNOR U5758 ( .A(n5603), .B(n5602), .Z(n5709) );
  XOR U5759 ( .A(n5823), .B(n5709), .Z(n5710) );
  XNOR U5760 ( .A(n5711), .B(n5710), .Z(n5591) );
  XOR U5761 ( .A(n5669), .B(n5668), .Z(n5687) );
  OR U5762 ( .A(n5444), .B(n5443), .Z(n5448) );
  NAND U5763 ( .A(n5446), .B(n5445), .Z(n5447) );
  AND U5764 ( .A(n5448), .B(n5447), .Z(n5685) );
  OR U5765 ( .A(n5450), .B(n5449), .Z(n5454) );
  OR U5766 ( .A(n5452), .B(n5451), .Z(n5453) );
  AND U5767 ( .A(n5454), .B(n5453), .Z(n5734) );
  NANDN U5768 ( .A(n5456), .B(n5455), .Z(n5460) );
  OR U5769 ( .A(n5458), .B(n5457), .Z(n5459) );
  AND U5770 ( .A(n5460), .B(n5459), .Z(n5732) );
  NANDN U5771 ( .A(n5462), .B(n5461), .Z(n5466) );
  NANDN U5772 ( .A(n5464), .B(n5463), .Z(n5465) );
  AND U5773 ( .A(n5466), .B(n5465), .Z(n5725) );
  AND U5774 ( .A(x[76]), .B(y[241]), .Z(n5850) );
  AND U5775 ( .A(y[231]), .B(x[86]), .Z(n5652) );
  AND U5776 ( .A(y[252]), .B(x[65]), .Z(n5653) );
  XNOR U5777 ( .A(n5652), .B(n5653), .Z(n5654) );
  XNOR U5778 ( .A(n5850), .B(n5654), .Z(n5699) );
  OR U5779 ( .A(n5468), .B(n5467), .Z(n5472) );
  OR U5780 ( .A(n5470), .B(n5469), .Z(n5471) );
  AND U5781 ( .A(n5472), .B(n5471), .Z(n5696) );
  NANDN U5782 ( .A(n5473), .B(x[79]), .Z(n5659) );
  AND U5783 ( .A(y[233]), .B(x[84]), .Z(n5657) );
  ANDN U5784 ( .B(x[85]), .A(n5947), .Z(n5958) );
  XOR U5785 ( .A(n5657), .B(n5958), .Z(n5658) );
  XNOR U5786 ( .A(n5659), .B(n5658), .Z(n5697) );
  XNOR U5787 ( .A(n5696), .B(n5697), .Z(n5698) );
  XNOR U5788 ( .A(n5699), .B(n5698), .Z(n5726) );
  XOR U5789 ( .A(n5725), .B(n5726), .Z(n5727) );
  OR U5790 ( .A(n5475), .B(n5474), .Z(n5479) );
  OR U5791 ( .A(n5477), .B(n5476), .Z(n5478) );
  AND U5792 ( .A(n5479), .B(n5478), .Z(n5728) );
  XNOR U5793 ( .A(n5727), .B(n5728), .Z(n5731) );
  XNOR U5794 ( .A(n5732), .B(n5731), .Z(n5733) );
  XNOR U5795 ( .A(n5734), .B(n5733), .Z(n5684) );
  XOR U5796 ( .A(n5685), .B(n5684), .Z(n5686) );
  XOR U5797 ( .A(n5687), .B(n5686), .Z(n5584) );
  OR U5798 ( .A(n5481), .B(n5480), .Z(n5485) );
  NANDN U5799 ( .A(n5483), .B(n5482), .Z(n5484) );
  AND U5800 ( .A(n5485), .B(n5484), .Z(n5572) );
  OR U5801 ( .A(n5487), .B(n5486), .Z(n5491) );
  NANDN U5802 ( .A(n5489), .B(n5488), .Z(n5490) );
  AND U5803 ( .A(n5491), .B(n5490), .Z(n5570) );
  NANDN U5804 ( .A(n5493), .B(n5492), .Z(n5497) );
  NANDN U5805 ( .A(n5495), .B(n5494), .Z(n5496) );
  AND U5806 ( .A(n5497), .B(n5496), .Z(n5576) );
  OR U5807 ( .A(n5499), .B(n5498), .Z(n5503) );
  NANDN U5808 ( .A(n5501), .B(n5500), .Z(n5502) );
  AND U5809 ( .A(n5503), .B(n5502), .Z(n5678) );
  OR U5810 ( .A(n5505), .B(n5504), .Z(n5509) );
  NANDN U5811 ( .A(n5507), .B(n5506), .Z(n5508) );
  AND U5812 ( .A(n5509), .B(n5508), .Z(n5679) );
  XOR U5813 ( .A(n5678), .B(n5679), .Z(n5680) );
  OR U5814 ( .A(n5511), .B(n5510), .Z(n5515) );
  NANDN U5815 ( .A(n5513), .B(n5512), .Z(n5514) );
  NAND U5816 ( .A(n5515), .B(n5514), .Z(n5681) );
  XNOR U5817 ( .A(n5680), .B(n5681), .Z(n5577) );
  XNOR U5818 ( .A(n5576), .B(n5577), .Z(n5578) );
  OR U5819 ( .A(n5517), .B(n5516), .Z(n5521) );
  NANDN U5820 ( .A(n5519), .B(n5518), .Z(n5520) );
  NAND U5821 ( .A(n5521), .B(n5520), .Z(n5579) );
  NANDN U5822 ( .A(n5523), .B(n5522), .Z(n5527) );
  NANDN U5823 ( .A(n5525), .B(n5524), .Z(n5526) );
  NAND U5824 ( .A(n5527), .B(n5526), .Z(n5583) );
  XOR U5825 ( .A(n5582), .B(n5583), .Z(n5585) );
  XOR U5826 ( .A(n5584), .B(n5585), .Z(n5567) );
  NANDN U5827 ( .A(n5529), .B(n5528), .Z(n5533) );
  NANDN U5828 ( .A(n5531), .B(n5530), .Z(n5532) );
  NAND U5829 ( .A(n5533), .B(n5532), .Z(n5564) );
  OR U5830 ( .A(n5535), .B(n5534), .Z(n5539) );
  OR U5831 ( .A(n5537), .B(n5536), .Z(n5538) );
  AND U5832 ( .A(n5539), .B(n5538), .Z(n5565) );
  XNOR U5833 ( .A(n5564), .B(n5565), .Z(n5566) );
  XOR U5834 ( .A(n5567), .B(n5566), .Z(n5561) );
  OR U5835 ( .A(n5541), .B(n5540), .Z(n5545) );
  NANDN U5836 ( .A(n5543), .B(n5542), .Z(n5544) );
  AND U5837 ( .A(n5545), .B(n5544), .Z(n5558) );
  OR U5838 ( .A(n5547), .B(n5546), .Z(n5551) );
  OR U5839 ( .A(n5549), .B(n5548), .Z(n5550) );
  NAND U5840 ( .A(n5551), .B(n5550), .Z(n5559) );
  XNOR U5841 ( .A(n5558), .B(n5559), .Z(n5560) );
  XNOR U5842 ( .A(n5561), .B(n5560), .Z(n5555) );
  XOR U5843 ( .A(n5554), .B(n5555), .Z(N126) );
  NANDN U5844 ( .A(n5553), .B(n5552), .Z(n5557) );
  NANDN U5845 ( .A(n5555), .B(n5554), .Z(n5556) );
  AND U5846 ( .A(n5557), .B(n5556), .Z(n6028) );
  OR U5847 ( .A(n5559), .B(n5558), .Z(n5563) );
  OR U5848 ( .A(n5561), .B(n5560), .Z(n5562) );
  AND U5849 ( .A(n5563), .B(n5562), .Z(n6029) );
  XNOR U5850 ( .A(n6028), .B(n6029), .Z(n6027) );
  NANDN U5851 ( .A(n5565), .B(n5564), .Z(n5569) );
  NANDN U5852 ( .A(n5567), .B(n5566), .Z(n5568) );
  NAND U5853 ( .A(n5569), .B(n5568), .Z(n5738) );
  OR U5854 ( .A(n5571), .B(n5570), .Z(n5575) );
  OR U5855 ( .A(n5573), .B(n5572), .Z(n5574) );
  NAND U5856 ( .A(n5575), .B(n5574), .Z(n6035) );
  OR U5857 ( .A(n5577), .B(n5576), .Z(n5581) );
  OR U5858 ( .A(n5579), .B(n5578), .Z(n5580) );
  NAND U5859 ( .A(n5581), .B(n5580), .Z(n6034) );
  XNOR U5860 ( .A(n6035), .B(n6034), .Z(n6032) );
  NANDN U5861 ( .A(n5583), .B(n5582), .Z(n5587) );
  OR U5862 ( .A(n5585), .B(n5584), .Z(n5586) );
  AND U5863 ( .A(n5587), .B(n5586), .Z(n6033) );
  OR U5864 ( .A(n5589), .B(n5588), .Z(n5593) );
  OR U5865 ( .A(n5591), .B(n5590), .Z(n5592) );
  AND U5866 ( .A(n5593), .B(n5592), .Z(n5761) );
  NANDN U5867 ( .A(n5595), .B(n5594), .Z(n5599) );
  OR U5868 ( .A(n5597), .B(n5596), .Z(n5598) );
  AND U5869 ( .A(n5599), .B(n5598), .Z(n5763) );
  OR U5870 ( .A(n5601), .B(n5600), .Z(n5605) );
  OR U5871 ( .A(n5603), .B(n5602), .Z(n5604) );
  AND U5872 ( .A(n5605), .B(n5604), .Z(n5782) );
  NANDN U5873 ( .A(n51), .B(y[248]), .Z(n5861) );
  NANDN U5874 ( .A(n50), .B(y[249]), .Z(n5863) );
  NANDN U5875 ( .A(n8824), .B(y[235]), .Z(n5862) );
  XNOR U5876 ( .A(n5863), .B(n5862), .Z(n5860) );
  XNOR U5877 ( .A(n5861), .B(n5860), .Z(n5807) );
  OR U5878 ( .A(n5607), .B(n5606), .Z(n5611) );
  OR U5879 ( .A(n5609), .B(n5608), .Z(n5610) );
  AND U5880 ( .A(n5611), .B(n5610), .Z(n5809) );
  NANDN U5881 ( .A(n49), .B(y[250]), .Z(n5963) );
  NANDN U5882 ( .A(n48), .B(y[251]), .Z(n5965) );
  ANDN U5883 ( .B(y[236]), .A(n61), .Z(n5964) );
  XNOR U5884 ( .A(n5965), .B(n5964), .Z(n5962) );
  XNOR U5885 ( .A(n5963), .B(n5962), .Z(n5810) );
  XOR U5886 ( .A(n5809), .B(n5810), .Z(n5808) );
  XNOR U5887 ( .A(n5807), .B(n5808), .Z(n5781) );
  XNOR U5888 ( .A(n5782), .B(n5781), .Z(n5784) );
  OR U5889 ( .A(n5613), .B(n5612), .Z(n5618) );
  NANDN U5890 ( .A(n5614), .B(o[60]), .Z(n5616) );
  NAND U5891 ( .A(y[226]), .B(x[91]), .Z(n5615) );
  AND U5892 ( .A(n5616), .B(n5615), .Z(n5617) );
  ANDN U5893 ( .B(n5618), .A(n5617), .Z(n5783) );
  XNOR U5894 ( .A(n5763), .B(n5764), .Z(n5762) );
  XNOR U5895 ( .A(n5761), .B(n5762), .Z(n6017) );
  OR U5896 ( .A(n5620), .B(n5619), .Z(n5624) );
  OR U5897 ( .A(n5622), .B(n5621), .Z(n5623) );
  NAND U5898 ( .A(n5624), .B(n5623), .Z(n5790) );
  NANDN U5899 ( .A(n8885), .B(y[234]), .Z(n5857) );
  ANDN U5900 ( .B(y[240]), .A(n59), .Z(n5856) );
  XOR U5901 ( .A(n5857), .B(n5856), .Z(n5855) );
  ANDN U5902 ( .B(y[246]), .A(n53), .Z(n5854) );
  XOR U5903 ( .A(n5855), .B(n5854), .Z(n5792) );
  NANDN U5904 ( .A(n5905), .B(x[94]), .Z(n5829) );
  NANDN U5905 ( .A(n8893), .B(y[225]), .Z(n5912) );
  XNOR U5906 ( .A(o[62]), .B(n5912), .Z(n5828) );
  XOR U5907 ( .A(n5829), .B(n5828), .Z(n5827) );
  ANDN U5908 ( .B(y[254]), .A(n45), .Z(n5826) );
  XOR U5909 ( .A(n5827), .B(n5826), .Z(n5791) );
  XOR U5910 ( .A(n5790), .B(n5789), .Z(n5990) );
  OR U5911 ( .A(n5626), .B(n5625), .Z(n5630) );
  OR U5912 ( .A(n5628), .B(n5627), .Z(n5629) );
  AND U5913 ( .A(n5630), .B(n5629), .Z(n5991) );
  XNOR U5914 ( .A(n5990), .B(n5991), .Z(n5989) );
  OR U5915 ( .A(n5632), .B(n5631), .Z(n5636) );
  OR U5916 ( .A(n5634), .B(n5633), .Z(n5635) );
  AND U5917 ( .A(n5636), .B(n5635), .Z(n5816) );
  NANDN U5918 ( .A(n8626), .B(y[237]), .Z(n5841) );
  NANDN U5919 ( .A(n47), .B(y[252]), .Z(n5843) );
  NANDN U5920 ( .A(n8901), .B(y[228]), .Z(n5842) );
  XNOR U5921 ( .A(n5843), .B(n5842), .Z(n5840) );
  XNOR U5922 ( .A(n5841), .B(n5840), .Z(n5817) );
  NANDN U5923 ( .A(n52), .B(y[247]), .Z(n5957) );
  ANDN U5924 ( .B(y[232]), .A(n8864), .Z(n5639) );
  ANDN U5925 ( .B(x[85]), .A(n5637), .Z(n5638) );
  XNOR U5926 ( .A(n5639), .B(n5638), .Z(n5956) );
  XOR U5927 ( .A(n5957), .B(n5956), .Z(n5818) );
  XNOR U5928 ( .A(n5817), .B(n5818), .Z(n5815) );
  XOR U5929 ( .A(n5816), .B(n5815), .Z(n5988) );
  XNOR U5930 ( .A(n5989), .B(n5988), .Z(n5769) );
  NANDN U5931 ( .A(n5641), .B(n5640), .Z(n5645) );
  OR U5932 ( .A(n5643), .B(n5642), .Z(n5644) );
  NAND U5933 ( .A(n5645), .B(n5644), .Z(n5772) );
  OR U5934 ( .A(n5647), .B(n5646), .Z(n5651) );
  OR U5935 ( .A(n5649), .B(n5648), .Z(n5650) );
  AND U5936 ( .A(n5651), .B(n5650), .Z(n5775) );
  OR U5937 ( .A(n5653), .B(n5652), .Z(n5656) );
  OR U5938 ( .A(n5654), .B(n5850), .Z(n5655) );
  AND U5939 ( .A(n5656), .B(n5655), .Z(n5778) );
  OR U5940 ( .A(n5657), .B(n5958), .Z(n5661) );
  NAND U5941 ( .A(n5659), .B(n5658), .Z(n5660) );
  AND U5942 ( .A(n5661), .B(n5660), .Z(n5801) );
  NAND U5943 ( .A(n5662), .B(o[61]), .Z(n5835) );
  NANDN U5944 ( .A(n8654), .B(y[226]), .Z(n5837) );
  NANDN U5945 ( .A(n8890), .B(y[238]), .Z(n5836) );
  XNOR U5946 ( .A(n5837), .B(n5836), .Z(n5834) );
  XNOR U5947 ( .A(n5835), .B(n5834), .Z(n5803) );
  NANDN U5948 ( .A(n8928), .B(y[229]), .Z(n5927) );
  ANDN U5949 ( .B(x[88]), .A(n5663), .Z(n5665) );
  NANDN U5950 ( .A(n8656), .B(y[231]), .Z(n5664) );
  XOR U5951 ( .A(n5665), .B(n5664), .Z(n5926) );
  XOR U5952 ( .A(n5927), .B(n5926), .Z(n5804) );
  XOR U5953 ( .A(n5803), .B(n5804), .Z(n5802) );
  XNOR U5954 ( .A(n5801), .B(n5802), .Z(n5777) );
  XOR U5955 ( .A(n5775), .B(n5776), .Z(n5771) );
  XNOR U5956 ( .A(n5772), .B(n5771), .Z(n5770) );
  XNOR U5957 ( .A(n5769), .B(n5770), .Z(n6016) );
  XNOR U5958 ( .A(n6017), .B(n6016), .Z(n6015) );
  OR U5959 ( .A(n5667), .B(n5666), .Z(n5671) );
  OR U5960 ( .A(n5669), .B(n5668), .Z(n5670) );
  NAND U5961 ( .A(n5671), .B(n5670), .Z(n6014) );
  XOR U5962 ( .A(n6015), .B(n6014), .Z(n5744) );
  OR U5963 ( .A(n5673), .B(n5672), .Z(n5677) );
  OR U5964 ( .A(n5675), .B(n5674), .Z(n5676) );
  NAND U5965 ( .A(n5677), .B(n5676), .Z(n5745) );
  OR U5966 ( .A(n5679), .B(n5678), .Z(n5683) );
  NANDN U5967 ( .A(n5681), .B(n5680), .Z(n5682) );
  AND U5968 ( .A(n5683), .B(n5682), .Z(n5746) );
  XOR U5969 ( .A(n5745), .B(n5746), .Z(n5743) );
  XOR U5970 ( .A(n5744), .B(n5743), .Z(n6009) );
  NANDN U5971 ( .A(n5685), .B(n5684), .Z(n5689) );
  OR U5972 ( .A(n5687), .B(n5686), .Z(n5688) );
  NAND U5973 ( .A(n5689), .B(n5688), .Z(n6011) );
  OR U5974 ( .A(n5691), .B(n5690), .Z(n5695) );
  OR U5975 ( .A(n5693), .B(n5692), .Z(n5694) );
  AND U5976 ( .A(n5695), .B(n5694), .Z(n5757) );
  OR U5977 ( .A(n5697), .B(n5696), .Z(n5701) );
  OR U5978 ( .A(n5699), .B(n5698), .Z(n5700) );
  AND U5979 ( .A(n5701), .B(n5700), .Z(n5758) );
  XOR U5980 ( .A(n5757), .B(n5758), .Z(n5755) );
  OR U5981 ( .A(n5703), .B(n5702), .Z(n5707) );
  OR U5982 ( .A(n5705), .B(n5704), .Z(n5706) );
  NAND U5983 ( .A(n5707), .B(n5706), .Z(n5756) );
  XNOR U5984 ( .A(n5755), .B(n5756), .Z(n5752) );
  OR U5985 ( .A(n5709), .B(n5708), .Z(n5713) );
  OR U5986 ( .A(n5711), .B(n5710), .Z(n5712) );
  NAND U5987 ( .A(n5713), .B(n5712), .Z(n5985) );
  NANDN U5988 ( .A(n5714), .B(x[91]), .Z(n5923) );
  NANDN U5989 ( .A(n46), .B(y[253]), .Z(n5922) );
  XOR U5990 ( .A(n5923), .B(n5922), .Z(n5921) );
  XOR U5991 ( .A(n5920), .B(n5921), .Z(n5795) );
  ANDN U5992 ( .B(y[242]), .A(n57), .Z(n5716) );
  ANDN U5993 ( .B(x[77]), .A(n5874), .Z(n5715) );
  XNOR U5994 ( .A(n5716), .B(n5715), .Z(n5849) );
  XOR U5995 ( .A(n5848), .B(n5849), .Z(n5822) );
  ANDN U5996 ( .B(y[244]), .A(n55), .Z(n5718) );
  ANDN U5997 ( .B(y[245]), .A(n54), .Z(n5717) );
  XNOR U5998 ( .A(n5718), .B(n5717), .Z(n5821) );
  XOR U5999 ( .A(n5822), .B(n5821), .Z(n5797) );
  OR U6000 ( .A(n5720), .B(n5719), .Z(n5724) );
  OR U6001 ( .A(n5722), .B(n5721), .Z(n5723) );
  AND U6002 ( .A(n5724), .B(n5723), .Z(n5798) );
  XNOR U6003 ( .A(n5797), .B(n5798), .Z(n5796) );
  XOR U6004 ( .A(n5795), .B(n5796), .Z(n5984) );
  XNOR U6005 ( .A(n5985), .B(n5984), .Z(n5983) );
  OR U6006 ( .A(n5726), .B(n5725), .Z(n5730) );
  NANDN U6007 ( .A(n5728), .B(n5727), .Z(n5729) );
  NAND U6008 ( .A(n5730), .B(n5729), .Z(n5982) );
  XOR U6009 ( .A(n5983), .B(n5982), .Z(n5751) );
  XOR U6010 ( .A(n5752), .B(n5751), .Z(n5750) );
  NANDN U6011 ( .A(n5732), .B(n5731), .Z(n5736) );
  NANDN U6012 ( .A(n5734), .B(n5733), .Z(n5735) );
  NAND U6013 ( .A(n5736), .B(n5735), .Z(n5749) );
  XNOR U6014 ( .A(n5750), .B(n5749), .Z(n6010) );
  XNOR U6015 ( .A(n6011), .B(n6010), .Z(n6008) );
  XOR U6016 ( .A(n6009), .B(n6008), .Z(n5740) );
  XOR U6017 ( .A(n5739), .B(n5740), .Z(n5737) );
  XNOR U6018 ( .A(n5738), .B(n5737), .Z(n6026) );
  XNOR U6019 ( .A(n6027), .B(n6026), .Z(N127) );
  NAND U6020 ( .A(n5738), .B(n5737), .Z(n5742) );
  OR U6021 ( .A(n5740), .B(n5739), .Z(n5741) );
  AND U6022 ( .A(n5742), .B(n5741), .Z(n6043) );
  NANDN U6023 ( .A(n5744), .B(n5743), .Z(n5748) );
  NOR U6024 ( .A(n5746), .B(n5745), .Z(n5747) );
  ANDN U6025 ( .B(n5748), .A(n5747), .Z(n6025) );
  OR U6026 ( .A(n5750), .B(n5749), .Z(n5754) );
  NANDN U6027 ( .A(n5752), .B(n5751), .Z(n5753) );
  AND U6028 ( .A(n5754), .B(n5753), .Z(n6007) );
  NANDN U6029 ( .A(n5756), .B(n5755), .Z(n5760) );
  OR U6030 ( .A(n5758), .B(n5757), .Z(n5759) );
  AND U6031 ( .A(n5760), .B(n5759), .Z(n5768) );
  OR U6032 ( .A(n5762), .B(n5761), .Z(n5766) );
  OR U6033 ( .A(n5764), .B(n5763), .Z(n5765) );
  NAND U6034 ( .A(n5766), .B(n5765), .Z(n5767) );
  XNOR U6035 ( .A(n5768), .B(n5767), .Z(n6005) );
  NANDN U6036 ( .A(n5770), .B(n5769), .Z(n5774) );
  OR U6037 ( .A(n5772), .B(n5771), .Z(n5773) );
  AND U6038 ( .A(n5774), .B(n5773), .Z(n6003) );
  OR U6039 ( .A(n5776), .B(n5775), .Z(n5780) );
  OR U6040 ( .A(n5778), .B(n5777), .Z(n5779) );
  AND U6041 ( .A(n5780), .B(n5779), .Z(n5788) );
  NOR U6042 ( .A(n5782), .B(n5781), .Z(n5786) );
  NOR U6043 ( .A(n5784), .B(n5783), .Z(n5785) );
  OR U6044 ( .A(n5786), .B(n5785), .Z(n5787) );
  XNOR U6045 ( .A(n5788), .B(n5787), .Z(n6001) );
  OR U6046 ( .A(n5790), .B(n5789), .Z(n5794) );
  OR U6047 ( .A(n5792), .B(n5791), .Z(n5793) );
  AND U6048 ( .A(n5794), .B(n5793), .Z(n5999) );
  OR U6049 ( .A(n5796), .B(n5795), .Z(n5800) );
  OR U6050 ( .A(n5798), .B(n5797), .Z(n5799) );
  AND U6051 ( .A(n5800), .B(n5799), .Z(n5981) );
  OR U6052 ( .A(n5802), .B(n5801), .Z(n5806) );
  NANDN U6053 ( .A(n5804), .B(n5803), .Z(n5805) );
  AND U6054 ( .A(n5806), .B(n5805), .Z(n5814) );
  NAND U6055 ( .A(n5808), .B(n5807), .Z(n5812) );
  OR U6056 ( .A(n5810), .B(n5809), .Z(n5811) );
  NAND U6057 ( .A(n5812), .B(n5811), .Z(n5813) );
  XNOR U6058 ( .A(n5814), .B(n5813), .Z(n5979) );
  NANDN U6059 ( .A(n5816), .B(n5815), .Z(n5820) );
  NANDN U6060 ( .A(n5818), .B(n5817), .Z(n5819) );
  AND U6061 ( .A(n5820), .B(n5819), .Z(n5977) );
  OR U6062 ( .A(n5822), .B(n5821), .Z(n5825) );
  NANDN U6063 ( .A(n55), .B(y[245]), .Z(n5953) );
  OR U6064 ( .A(n5953), .B(n5823), .Z(n5824) );
  AND U6065 ( .A(n5825), .B(n5824), .Z(n5833) );
  NANDN U6066 ( .A(n5827), .B(n5826), .Z(n5831) );
  NANDN U6067 ( .A(n5829), .B(n5828), .Z(n5830) );
  NAND U6068 ( .A(n5831), .B(n5830), .Z(n5832) );
  XNOR U6069 ( .A(n5833), .B(n5832), .Z(n5975) );
  OR U6070 ( .A(n5835), .B(n5834), .Z(n5839) );
  OR U6071 ( .A(n5837), .B(n5836), .Z(n5838) );
  AND U6072 ( .A(n5839), .B(n5838), .Z(n5847) );
  OR U6073 ( .A(n5841), .B(n5840), .Z(n5845) );
  OR U6074 ( .A(n5843), .B(n5842), .Z(n5844) );
  NAND U6075 ( .A(n5845), .B(n5844), .Z(n5846) );
  XNOR U6076 ( .A(n5847), .B(n5846), .Z(n5888) );
  NANDN U6077 ( .A(n5849), .B(n5848), .Z(n5853) );
  NANDN U6078 ( .A(n5851), .B(n5850), .Z(n5852) );
  AND U6079 ( .A(n5853), .B(n5852), .Z(n5886) );
  NANDN U6080 ( .A(n5855), .B(n5854), .Z(n5859) );
  NANDN U6081 ( .A(n5857), .B(n5856), .Z(n5858) );
  AND U6082 ( .A(n5859), .B(n5858), .Z(n5867) );
  OR U6083 ( .A(n5861), .B(n5860), .Z(n5865) );
  OR U6084 ( .A(n5863), .B(n5862), .Z(n5864) );
  NAND U6085 ( .A(n5865), .B(n5864), .Z(n5866) );
  XNOR U6086 ( .A(n5867), .B(n5866), .Z(n5884) );
  ANDN U6087 ( .B(y[246]), .A(n54), .Z(n5869) );
  NANDN U6088 ( .A(n45), .B(y[255]), .Z(n5868) );
  XNOR U6089 ( .A(n5869), .B(n5868), .Z(n5873) );
  ANDN U6090 ( .B(y[240]), .A(n60), .Z(n5871) );
  NANDN U6091 ( .A(n46), .B(y[254]), .Z(n5870) );
  XNOR U6092 ( .A(n5871), .B(n5870), .Z(n5872) );
  XOR U6093 ( .A(n5873), .B(n5872), .Z(n5882) );
  ANDN U6094 ( .B(x[78]), .A(n5874), .Z(n5876) );
  NANDN U6095 ( .A(n8928), .B(y[230]), .Z(n5875) );
  XNOR U6096 ( .A(n5876), .B(n5875), .Z(n5880) );
  ANDN U6097 ( .B(y[226]), .A(n8893), .Z(n5878) );
  NAND U6098 ( .A(y[225]), .B(x[94]), .Z(n5877) );
  XNOR U6099 ( .A(n5878), .B(n5877), .Z(n5879) );
  XNOR U6100 ( .A(n5880), .B(n5879), .Z(n5881) );
  XNOR U6101 ( .A(n5882), .B(n5881), .Z(n5883) );
  XNOR U6102 ( .A(n5884), .B(n5883), .Z(n5885) );
  XNOR U6103 ( .A(n5886), .B(n5885), .Z(n5887) );
  XOR U6104 ( .A(n5888), .B(n5887), .Z(n5973) );
  ANDN U6105 ( .B(y[243]), .A(n57), .Z(n5890) );
  NANDN U6106 ( .A(n8654), .B(y[227]), .Z(n5889) );
  XNOR U6107 ( .A(n5890), .B(n5889), .Z(n5894) );
  ANDN U6108 ( .B(y[244]), .A(n56), .Z(n5892) );
  NANDN U6109 ( .A(n8901), .B(y[229]), .Z(n5891) );
  XNOR U6110 ( .A(n5892), .B(n5891), .Z(n5893) );
  XOR U6111 ( .A(n5894), .B(n5893), .Z(n5902) );
  ANDN U6112 ( .B(y[253]), .A(n47), .Z(n5896) );
  NAND U6113 ( .A(x[91]), .B(y[228]), .Z(n5895) );
  XNOR U6114 ( .A(n5896), .B(n5895), .Z(n5900) );
  ANDN U6115 ( .B(y[251]), .A(n49), .Z(n5898) );
  NANDN U6116 ( .A(n8626), .B(y[238]), .Z(n5897) );
  XNOR U6117 ( .A(n5898), .B(n5897), .Z(n5899) );
  XNOR U6118 ( .A(n5900), .B(n5899), .Z(n5901) );
  XNOR U6119 ( .A(n5902), .B(n5901), .Z(n5911) );
  ANDN U6120 ( .B(y[249]), .A(n51), .Z(n5904) );
  NANDN U6121 ( .A(n50), .B(y[250]), .Z(n5903) );
  XNOR U6122 ( .A(n5904), .B(n5903), .Z(n5909) );
  ANDN U6123 ( .B(x[95]), .A(n5905), .Z(n5907) );
  NANDN U6124 ( .A(n52), .B(y[248]), .Z(n5906) );
  XNOR U6125 ( .A(n5907), .B(n5906), .Z(n5908) );
  XNOR U6126 ( .A(n5909), .B(n5908), .Z(n5910) );
  XNOR U6127 ( .A(n5911), .B(n5910), .Z(n5946) );
  ANDN U6128 ( .B(y[236]), .A(n8824), .Z(n5919) );
  ANDN U6129 ( .B(o[62]), .A(n5912), .Z(n5917) );
  XOR U6130 ( .A(n5913), .B(o[63]), .Z(n5915) );
  NANDN U6131 ( .A(n8864), .B(y[233]), .Z(n5959) );
  NANDN U6132 ( .A(n8865), .B(y[231]), .Z(n5929) );
  XNOR U6133 ( .A(n5959), .B(n5929), .Z(n5914) );
  XNOR U6134 ( .A(n5915), .B(n5914), .Z(n5916) );
  XNOR U6135 ( .A(n5917), .B(n5916), .Z(n5918) );
  XNOR U6136 ( .A(n5919), .B(n5918), .Z(n5935) );
  NAND U6137 ( .A(n5921), .B(n5920), .Z(n5925) );
  OR U6138 ( .A(n5923), .B(n5922), .Z(n5924) );
  AND U6139 ( .A(n5925), .B(n5924), .Z(n5933) );
  OR U6140 ( .A(n5927), .B(n5926), .Z(n5931) );
  OR U6141 ( .A(n5929), .B(n5928), .Z(n5930) );
  NAND U6142 ( .A(n5931), .B(n5930), .Z(n5932) );
  XNOR U6143 ( .A(n5933), .B(n5932), .Z(n5934) );
  XOR U6144 ( .A(n5935), .B(n5934), .Z(n5944) );
  ANDN U6145 ( .B(x[80]), .A(n5936), .Z(n5938) );
  NANDN U6146 ( .A(n8885), .B(y[235]), .Z(n5937) );
  XNOR U6147 ( .A(n5938), .B(n5937), .Z(n5942) );
  ANDN U6148 ( .B(y[247]), .A(n53), .Z(n5940) );
  NANDN U6149 ( .A(n8827), .B(y[234]), .Z(n5939) );
  XNOR U6150 ( .A(n5940), .B(n5939), .Z(n5941) );
  XNOR U6151 ( .A(n5942), .B(n5941), .Z(n5943) );
  XNOR U6152 ( .A(n5944), .B(n5943), .Z(n5945) );
  XOR U6153 ( .A(n5946), .B(n5945), .Z(n5955) );
  ANDN U6154 ( .B(x[87]), .A(n5947), .Z(n5949) );
  NANDN U6155 ( .A(n61), .B(y[237]), .Z(n5948) );
  XNOR U6156 ( .A(n5949), .B(n5948), .Z(n5951) );
  NANDN U6157 ( .A(n48), .B(y[252]), .Z(n5950) );
  XNOR U6158 ( .A(n5951), .B(n5950), .Z(n5952) );
  XOR U6159 ( .A(n5953), .B(n5952), .Z(n5954) );
  XNOR U6160 ( .A(n5955), .B(n5954), .Z(n5971) );
  OR U6161 ( .A(n5957), .B(n5956), .Z(n5961) );
  NANDN U6162 ( .A(n5959), .B(n5958), .Z(n5960) );
  AND U6163 ( .A(n5961), .B(n5960), .Z(n5969) );
  NANDN U6164 ( .A(n5963), .B(n5962), .Z(n5967) );
  NANDN U6165 ( .A(n5965), .B(n5964), .Z(n5966) );
  NAND U6166 ( .A(n5967), .B(n5966), .Z(n5968) );
  XNOR U6167 ( .A(n5969), .B(n5968), .Z(n5970) );
  XNOR U6168 ( .A(n5971), .B(n5970), .Z(n5972) );
  XNOR U6169 ( .A(n5973), .B(n5972), .Z(n5974) );
  XNOR U6170 ( .A(n5975), .B(n5974), .Z(n5976) );
  XNOR U6171 ( .A(n5977), .B(n5976), .Z(n5978) );
  XNOR U6172 ( .A(n5979), .B(n5978), .Z(n5980) );
  XNOR U6173 ( .A(n5981), .B(n5980), .Z(n5997) );
  OR U6174 ( .A(n5983), .B(n5982), .Z(n5987) );
  OR U6175 ( .A(n5985), .B(n5984), .Z(n5986) );
  AND U6176 ( .A(n5987), .B(n5986), .Z(n5995) );
  OR U6177 ( .A(n5989), .B(n5988), .Z(n5993) );
  OR U6178 ( .A(n5991), .B(n5990), .Z(n5992) );
  NAND U6179 ( .A(n5993), .B(n5992), .Z(n5994) );
  XNOR U6180 ( .A(n5995), .B(n5994), .Z(n5996) );
  XNOR U6181 ( .A(n5997), .B(n5996), .Z(n5998) );
  XNOR U6182 ( .A(n5999), .B(n5998), .Z(n6000) );
  XNOR U6183 ( .A(n6001), .B(n6000), .Z(n6002) );
  XNOR U6184 ( .A(n6003), .B(n6002), .Z(n6004) );
  XNOR U6185 ( .A(n6005), .B(n6004), .Z(n6006) );
  XNOR U6186 ( .A(n6007), .B(n6006), .Z(n6023) );
  OR U6187 ( .A(n6009), .B(n6008), .Z(n6013) );
  OR U6188 ( .A(n6011), .B(n6010), .Z(n6012) );
  AND U6189 ( .A(n6013), .B(n6012), .Z(n6021) );
  OR U6190 ( .A(n6015), .B(n6014), .Z(n6019) );
  OR U6191 ( .A(n6017), .B(n6016), .Z(n6018) );
  NAND U6192 ( .A(n6019), .B(n6018), .Z(n6020) );
  XNOR U6193 ( .A(n6021), .B(n6020), .Z(n6022) );
  XNOR U6194 ( .A(n6023), .B(n6022), .Z(n6024) );
  XNOR U6195 ( .A(n6025), .B(n6024), .Z(n6041) );
  OR U6196 ( .A(n6027), .B(n6026), .Z(n6031) );
  OR U6197 ( .A(n6029), .B(n6028), .Z(n6030) );
  AND U6198 ( .A(n6031), .B(n6030), .Z(n6039) );
  OR U6199 ( .A(n6033), .B(n6032), .Z(n6037) );
  OR U6200 ( .A(n6035), .B(n6034), .Z(n6036) );
  NAND U6201 ( .A(n6037), .B(n6036), .Z(n6038) );
  XNOR U6202 ( .A(n6039), .B(n6038), .Z(n6040) );
  XNOR U6203 ( .A(n6041), .B(n6040), .Z(n6042) );
  XNOR U6204 ( .A(n6043), .B(n6042), .Z(N128) );
  IV U6205 ( .A(y[256]), .Z(n8872) );
  ANDN U6206 ( .B(x[64]), .A(n8872), .Z(n6748) );
  XOR U6207 ( .A(n6748), .B(o[64]), .Z(N161) );
  ANDN U6208 ( .B(x[65]), .A(n8872), .Z(n6044) );
  NANDN U6209 ( .A(n45), .B(y[257]), .Z(n6050) );
  XNOR U6210 ( .A(n6050), .B(o[65]), .Z(n6045) );
  XOR U6211 ( .A(n6044), .B(n6045), .Z(n6046) );
  AND U6212 ( .A(o[64]), .B(n6748), .Z(n6047) );
  XOR U6213 ( .A(n6046), .B(n6047), .Z(N162) );
  OR U6214 ( .A(n6045), .B(n6044), .Z(n6049) );
  NANDN U6215 ( .A(n6047), .B(n6046), .Z(n6048) );
  NAND U6216 ( .A(n6049), .B(n6048), .Z(n6052) );
  NANDN U6217 ( .A(n45), .B(y[258]), .Z(n6063) );
  XOR U6218 ( .A(n6063), .B(o[66]), .Z(n6051) );
  XNOR U6219 ( .A(n6052), .B(n6051), .Z(n6054) );
  ANDN U6220 ( .B(o[65]), .A(n6050), .Z(n6057) );
  AND U6221 ( .A(y[256]), .B(x[66]), .Z(n6058) );
  XNOR U6222 ( .A(n6057), .B(n6058), .Z(n6060) );
  AND U6223 ( .A(y[257]), .B(x[65]), .Z(n6059) );
  XNOR U6224 ( .A(n6060), .B(n6059), .Z(n6053) );
  XNOR U6225 ( .A(n6054), .B(n6053), .Z(N163) );
  NAND U6226 ( .A(n6052), .B(n6051), .Z(n6056) );
  OR U6227 ( .A(n6054), .B(n6053), .Z(n6055) );
  NAND U6228 ( .A(n6056), .B(n6055), .Z(n6067) );
  OR U6229 ( .A(n6058), .B(n6057), .Z(n6062) );
  OR U6230 ( .A(n6060), .B(n6059), .Z(n6061) );
  AND U6231 ( .A(n6062), .B(n6061), .Z(n6068) );
  XNOR U6232 ( .A(n6067), .B(n6068), .Z(n6069) );
  NANDN U6233 ( .A(n47), .B(y[257]), .Z(n6075) );
  XNOR U6234 ( .A(n6075), .B(o[67]), .Z(n6073) );
  NANDN U6235 ( .A(n6063), .B(o[66]), .Z(n6079) );
  ANDN U6236 ( .B(x[67]), .A(n8872), .Z(n6065) );
  NANDN U6237 ( .A(n45), .B(y[259]), .Z(n6064) );
  XOR U6238 ( .A(n6065), .B(n6064), .Z(n6078) );
  XNOR U6239 ( .A(n6079), .B(n6078), .Z(n6074) );
  AND U6240 ( .A(y[258]), .B(x[65]), .Z(n6103) );
  XOR U6241 ( .A(n6074), .B(n6103), .Z(n6066) );
  XOR U6242 ( .A(n6073), .B(n6066), .Z(n6070) );
  XNOR U6243 ( .A(n6069), .B(n6070), .Z(N164) );
  NANDN U6244 ( .A(n6068), .B(n6067), .Z(n6072) );
  NAND U6245 ( .A(n6070), .B(n6069), .Z(n6071) );
  NAND U6246 ( .A(n6072), .B(n6071), .Z(n6084) );
  XNOR U6247 ( .A(n6084), .B(n6085), .Z(n6086) );
  NANDN U6248 ( .A(n6075), .B(o[67]), .Z(n6100) );
  ANDN U6249 ( .B(x[68]), .A(n8872), .Z(n6077) );
  ANDN U6250 ( .B(y[260]), .A(n45), .Z(n6076) );
  XNOR U6251 ( .A(n6077), .B(n6076), .Z(n6099) );
  XOR U6252 ( .A(n6100), .B(n6099), .Z(n6092) );
  AND U6253 ( .A(y[259]), .B(x[67]), .Z(n6156) );
  NAND U6254 ( .A(n6748), .B(n6156), .Z(n6081) );
  OR U6255 ( .A(n6079), .B(n6078), .Z(n6080) );
  AND U6256 ( .A(n6081), .B(n6080), .Z(n6090) );
  IV U6257 ( .A(y[259]), .Z(n8881) );
  ANDN U6258 ( .B(x[65]), .A(n8881), .Z(n6083) );
  NANDN U6259 ( .A(n47), .B(y[258]), .Z(n6082) );
  XOR U6260 ( .A(n6083), .B(n6082), .Z(n6105) );
  NANDN U6261 ( .A(n48), .B(y[257]), .Z(n6096) );
  XNOR U6262 ( .A(n6096), .B(o[68]), .Z(n6104) );
  XOR U6263 ( .A(n6105), .B(n6104), .Z(n6091) );
  XOR U6264 ( .A(n6092), .B(n6093), .Z(n6087) );
  XOR U6265 ( .A(n6086), .B(n6087), .Z(N165) );
  NANDN U6266 ( .A(n6085), .B(n6084), .Z(n6089) );
  NANDN U6267 ( .A(n6087), .B(n6086), .Z(n6088) );
  NAND U6268 ( .A(n6089), .B(n6088), .Z(n6108) );
  OR U6269 ( .A(n6091), .B(n6090), .Z(n6095) );
  NAND U6270 ( .A(n6093), .B(n6092), .Z(n6094) );
  NAND U6271 ( .A(n6095), .B(n6094), .Z(n6109) );
  XNOR U6272 ( .A(n6108), .B(n6109), .Z(n6110) );
  NANDN U6273 ( .A(n6096), .B(o[68]), .Z(n6127) );
  ANDN U6274 ( .B(x[69]), .A(n8872), .Z(n6098) );
  IV U6275 ( .A(y[261]), .Z(n7989) );
  ANDN U6276 ( .B(x[64]), .A(n7989), .Z(n6097) );
  XNOR U6277 ( .A(n6098), .B(n6097), .Z(n6126) );
  XOR U6278 ( .A(n6127), .B(n6126), .Z(n6122) );
  AND U6279 ( .A(y[259]), .B(x[66]), .Z(n6120) );
  AND U6280 ( .A(y[260]), .B(x[65]), .Z(n6135) );
  NANDN U6281 ( .A(n49), .B(y[257]), .Z(n6130) );
  XNOR U6282 ( .A(o[69]), .B(n6130), .Z(n6133) );
  AND U6283 ( .A(y[258]), .B(x[67]), .Z(n6134) );
  XNOR U6284 ( .A(n6133), .B(n6134), .Z(n6136) );
  XNOR U6285 ( .A(n6135), .B(n6136), .Z(n6121) );
  XNOR U6286 ( .A(n6120), .B(n6121), .Z(n6123) );
  XNOR U6287 ( .A(n6122), .B(n6123), .Z(n6117) );
  AND U6288 ( .A(y[260]), .B(x[68]), .Z(n6245) );
  NAND U6289 ( .A(n6748), .B(n6245), .Z(n6102) );
  OR U6290 ( .A(n6100), .B(n6099), .Z(n6101) );
  NAND U6291 ( .A(n6102), .B(n6101), .Z(n6115) );
  NAND U6292 ( .A(n6103), .B(n6120), .Z(n6107) );
  NANDN U6293 ( .A(n6105), .B(n6104), .Z(n6106) );
  NAND U6294 ( .A(n6107), .B(n6106), .Z(n6114) );
  XNOR U6295 ( .A(n6115), .B(n6114), .Z(n6116) );
  XNOR U6296 ( .A(n6117), .B(n6116), .Z(n6111) );
  XOR U6297 ( .A(n6110), .B(n6111), .Z(N166) );
  NANDN U6298 ( .A(n6109), .B(n6108), .Z(n6113) );
  NANDN U6299 ( .A(n6111), .B(n6110), .Z(n6112) );
  NAND U6300 ( .A(n6113), .B(n6112), .Z(n6139) );
  OR U6301 ( .A(n6115), .B(n6114), .Z(n6119) );
  OR U6302 ( .A(n6117), .B(n6116), .Z(n6118) );
  AND U6303 ( .A(n6119), .B(n6118), .Z(n6140) );
  XNOR U6304 ( .A(n6139), .B(n6140), .Z(n6141) );
  OR U6305 ( .A(n6121), .B(n6120), .Z(n6125) );
  OR U6306 ( .A(n6123), .B(n6122), .Z(n6124) );
  AND U6307 ( .A(n6125), .B(n6124), .Z(n6145) );
  NANDN U6308 ( .A(n50), .B(y[261]), .Z(n6518) );
  NANDN U6309 ( .A(n6518), .B(n6748), .Z(n6129) );
  OR U6310 ( .A(n6127), .B(n6126), .Z(n6128) );
  NAND U6311 ( .A(n6129), .B(n6128), .Z(n6168) );
  NANDN U6312 ( .A(n6130), .B(o[69]), .Z(n6153) );
  ANDN U6313 ( .B(x[70]), .A(n8872), .Z(n6132) );
  NANDN U6314 ( .A(n45), .B(y[262]), .Z(n6131) );
  XNOR U6315 ( .A(n6132), .B(n6131), .Z(n6152) );
  XNOR U6316 ( .A(n6153), .B(n6152), .Z(n6167) );
  XNOR U6317 ( .A(n6168), .B(n6167), .Z(n6170) );
  AND U6318 ( .A(y[261]), .B(x[65]), .Z(n6444) );
  NANDN U6319 ( .A(n50), .B(y[257]), .Z(n6166) );
  XOR U6320 ( .A(o[70]), .B(n6166), .Z(n6161) );
  XNOR U6321 ( .A(n6444), .B(n6161), .Z(n6162) );
  NANDN U6322 ( .A(n49), .B(y[258]), .Z(n6163) );
  XNOR U6323 ( .A(n6162), .B(n6163), .Z(n6157) );
  ANDN U6324 ( .B(y[260]), .A(n47), .Z(n6500) );
  XNOR U6325 ( .A(n6156), .B(n6500), .Z(n6158) );
  XOR U6326 ( .A(n6170), .B(n6169), .Z(n6146) );
  XNOR U6327 ( .A(n6145), .B(n6146), .Z(n6147) );
  OR U6328 ( .A(n6134), .B(n6133), .Z(n6138) );
  OR U6329 ( .A(n6136), .B(n6135), .Z(n6137) );
  AND U6330 ( .A(n6138), .B(n6137), .Z(n6148) );
  XOR U6331 ( .A(n6141), .B(n6142), .Z(N167) );
  NANDN U6332 ( .A(n6140), .B(n6139), .Z(n6144) );
  NANDN U6333 ( .A(n6142), .B(n6141), .Z(n6143) );
  NAND U6334 ( .A(n6144), .B(n6143), .Z(n6173) );
  OR U6335 ( .A(n6146), .B(n6145), .Z(n6150) );
  OR U6336 ( .A(n6148), .B(n6147), .Z(n6149) );
  AND U6337 ( .A(n6150), .B(n6149), .Z(n6174) );
  XNOR U6338 ( .A(n6173), .B(n6174), .Z(n6175) );
  ANDN U6339 ( .B(y[262]), .A(n51), .Z(n6151) );
  NAND U6340 ( .A(n6748), .B(n6151), .Z(n6155) );
  NANDN U6341 ( .A(n6153), .B(n6152), .Z(n6154) );
  NAND U6342 ( .A(n6155), .B(n6154), .Z(n6185) );
  AND U6343 ( .A(y[258]), .B(x[69]), .Z(n6363) );
  AND U6344 ( .A(y[262]), .B(x[65]), .Z(n6565) );
  NANDN U6345 ( .A(n51), .B(y[257]), .Z(n6191) );
  XOR U6346 ( .A(o[71]), .B(n6191), .Z(n6193) );
  XNOR U6347 ( .A(n6565), .B(n6193), .Z(n6194) );
  XNOR U6348 ( .A(n6363), .B(n6194), .Z(n6186) );
  XOR U6349 ( .A(n6185), .B(n6186), .Z(n6188) );
  OR U6350 ( .A(n6156), .B(n6500), .Z(n6160) );
  OR U6351 ( .A(n6158), .B(n6157), .Z(n6159) );
  AND U6352 ( .A(n6160), .B(n6159), .Z(n6187) );
  XNOR U6353 ( .A(n6188), .B(n6187), .Z(n6179) );
  NANDN U6354 ( .A(n6161), .B(n6444), .Z(n6165) );
  NANDN U6355 ( .A(n6163), .B(n6162), .Z(n6164) );
  NAND U6356 ( .A(n6165), .B(n6164), .Z(n6200) );
  ANDN U6357 ( .B(x[66]), .A(n7989), .Z(n6212) );
  IV U6358 ( .A(n6212), .Z(n6637) );
  AND U6359 ( .A(y[259]), .B(x[68]), .Z(n6349) );
  NANDN U6360 ( .A(n48), .B(y[260]), .Z(n6211) );
  XOR U6361 ( .A(n6349), .B(n6211), .Z(n6213) );
  XNOR U6362 ( .A(n6637), .B(n6213), .Z(n6198) );
  NANDN U6363 ( .A(n45), .B(y[263]), .Z(n6207) );
  NANDN U6364 ( .A(n6166), .B(o[70]), .Z(n6205) );
  NANDN U6365 ( .A(n8872), .B(x[71]), .Z(n6206) );
  XNOR U6366 ( .A(n6205), .B(n6206), .Z(n6208) );
  XNOR U6367 ( .A(n6207), .B(n6208), .Z(n6197) );
  XOR U6368 ( .A(n6198), .B(n6197), .Z(n6199) );
  XOR U6369 ( .A(n6200), .B(n6199), .Z(n6180) );
  XNOR U6370 ( .A(n6179), .B(n6180), .Z(n6182) );
  OR U6371 ( .A(n6168), .B(n6167), .Z(n6172) );
  NANDN U6372 ( .A(n6170), .B(n6169), .Z(n6171) );
  AND U6373 ( .A(n6172), .B(n6171), .Z(n6181) );
  XOR U6374 ( .A(n6182), .B(n6181), .Z(n6176) );
  XNOR U6375 ( .A(n6175), .B(n6176), .Z(N168) );
  NANDN U6376 ( .A(n6174), .B(n6173), .Z(n6178) );
  NAND U6377 ( .A(n6176), .B(n6175), .Z(n6177) );
  NAND U6378 ( .A(n6178), .B(n6177), .Z(n6257) );
  OR U6379 ( .A(n6180), .B(n6179), .Z(n6184) );
  OR U6380 ( .A(n6182), .B(n6181), .Z(n6183) );
  AND U6381 ( .A(n6184), .B(n6183), .Z(n6258) );
  XNOR U6382 ( .A(n6257), .B(n6258), .Z(n6259) );
  NANDN U6383 ( .A(n6186), .B(n6185), .Z(n6190) );
  NANDN U6384 ( .A(n6188), .B(n6187), .Z(n6189) );
  NAND U6385 ( .A(n6190), .B(n6189), .Z(n6264) );
  AND U6386 ( .A(y[258]), .B(x[70]), .Z(n6246) );
  XNOR U6387 ( .A(n6245), .B(n6246), .Z(n6248) );
  IV U6388 ( .A(y[262]), .Z(n8655) );
  ANDN U6389 ( .B(x[66]), .A(n8655), .Z(n6247) );
  IV U6390 ( .A(n6247), .Z(n6758) );
  XOR U6391 ( .A(n6248), .B(n6758), .Z(n6252) );
  ANDN U6392 ( .B(x[67]), .A(n7989), .Z(n6251) );
  IV U6393 ( .A(n6251), .Z(n7061) );
  XOR U6394 ( .A(n6252), .B(n7061), .Z(n6254) );
  NANDN U6395 ( .A(n6191), .B(o[71]), .Z(n6242) );
  ANDN U6396 ( .B(y[263]), .A(n46), .Z(n6743) );
  ANDN U6397 ( .B(x[69]), .A(n8881), .Z(n6192) );
  XNOR U6398 ( .A(n6743), .B(n6192), .Z(n6241) );
  XOR U6399 ( .A(n6242), .B(n6241), .Z(n6253) );
  XNOR U6400 ( .A(n6254), .B(n6253), .Z(n6216) );
  NANDN U6401 ( .A(n6193), .B(n6565), .Z(n6196) );
  NAND U6402 ( .A(n6194), .B(n6363), .Z(n6195) );
  AND U6403 ( .A(n6196), .B(n6195), .Z(n6217) );
  XOR U6404 ( .A(n6216), .B(n6217), .Z(n6219) );
  OR U6405 ( .A(n6198), .B(n6197), .Z(n6202) );
  NAND U6406 ( .A(n6200), .B(n6199), .Z(n6201) );
  AND U6407 ( .A(n6202), .B(n6201), .Z(n6218) );
  XOR U6408 ( .A(n6219), .B(n6218), .Z(n6263) );
  XNOR U6409 ( .A(n6264), .B(n6263), .Z(n6265) );
  ANDN U6410 ( .B(x[72]), .A(n8872), .Z(n6204) );
  NANDN U6411 ( .A(n45), .B(y[264]), .Z(n6203) );
  XOR U6412 ( .A(n6204), .B(n6203), .Z(n6230) );
  NANDN U6413 ( .A(n52), .B(y[257]), .Z(n6233) );
  XOR U6414 ( .A(n6233), .B(o[72]), .Z(n6229) );
  XNOR U6415 ( .A(n6230), .B(n6229), .Z(n6223) );
  NAND U6416 ( .A(n6206), .B(n6205), .Z(n6210) );
  NANDN U6417 ( .A(n6208), .B(n6207), .Z(n6209) );
  NAND U6418 ( .A(n6210), .B(n6209), .Z(n6222) );
  XNOR U6419 ( .A(n6223), .B(n6222), .Z(n6224) );
  NANDN U6420 ( .A(n6349), .B(n6211), .Z(n6215) );
  OR U6421 ( .A(n6213), .B(n6212), .Z(n6214) );
  NAND U6422 ( .A(n6215), .B(n6214), .Z(n6225) );
  XOR U6423 ( .A(n6265), .B(n6266), .Z(n6260) );
  XOR U6424 ( .A(n6259), .B(n6260), .Z(N169) );
  NANDN U6425 ( .A(n6217), .B(n6216), .Z(n6221) );
  OR U6426 ( .A(n6219), .B(n6218), .Z(n6220) );
  NAND U6427 ( .A(n6221), .B(n6220), .Z(n6276) );
  OR U6428 ( .A(n6223), .B(n6222), .Z(n6227) );
  OR U6429 ( .A(n6225), .B(n6224), .Z(n6226) );
  NAND U6430 ( .A(n6227), .B(n6226), .Z(n6275) );
  XOR U6431 ( .A(n6276), .B(n6275), .Z(n6277) );
  ANDN U6432 ( .B(y[264]), .A(n53), .Z(n6228) );
  NAND U6433 ( .A(n6748), .B(n6228), .Z(n6232) );
  OR U6434 ( .A(n6230), .B(n6229), .Z(n6231) );
  NAND U6435 ( .A(n6232), .B(n6231), .Z(n6290) );
  NANDN U6436 ( .A(n6233), .B(o[72]), .Z(n6314) );
  ANDN U6437 ( .B(y[258]), .A(n52), .Z(n6235) );
  NANDN U6438 ( .A(n50), .B(y[260]), .Z(n6234) );
  XNOR U6439 ( .A(n6235), .B(n6234), .Z(n6313) );
  XNOR U6440 ( .A(n6314), .B(n6313), .Z(n6288) );
  ANDN U6441 ( .B(x[73]), .A(n8872), .Z(n6237) );
  NANDN U6442 ( .A(n45), .B(y[265]), .Z(n6236) );
  XOR U6443 ( .A(n6237), .B(n6236), .Z(n6310) );
  NANDN U6444 ( .A(n53), .B(y[257]), .Z(n6303) );
  XOR U6445 ( .A(n6303), .B(o[73]), .Z(n6309) );
  XNOR U6446 ( .A(n6310), .B(n6309), .Z(n6287) );
  XNOR U6447 ( .A(n6288), .B(n6287), .Z(n6289) );
  XNOR U6448 ( .A(n6290), .B(n6289), .Z(n6283) );
  NANDN U6449 ( .A(n49), .B(y[261]), .Z(n6739) );
  IV U6450 ( .A(y[264]), .Z(n8927) );
  ANDN U6451 ( .B(x[65]), .A(n8927), .Z(n6239) );
  NANDN U6452 ( .A(n51), .B(y[259]), .Z(n6238) );
  XNOR U6453 ( .A(n6239), .B(n6238), .Z(n6305) );
  XNOR U6454 ( .A(n6739), .B(n6305), .Z(n6293) );
  AND U6455 ( .A(y[262]), .B(x[67]), .Z(n6663) );
  AND U6456 ( .A(y[263]), .B(x[66]), .Z(n6969) );
  XNOR U6457 ( .A(n6663), .B(n6969), .Z(n6294) );
  XNOR U6458 ( .A(n6293), .B(n6294), .Z(n6281) );
  NANDN U6459 ( .A(n46), .B(y[259]), .Z(n6304) );
  ANDN U6460 ( .B(y[263]), .A(n50), .Z(n6240) );
  NANDN U6461 ( .A(n6304), .B(n6240), .Z(n6244) );
  OR U6462 ( .A(n6242), .B(n6241), .Z(n6243) );
  AND U6463 ( .A(n6244), .B(n6243), .Z(n6282) );
  XOR U6464 ( .A(n6281), .B(n6282), .Z(n6284) );
  XNOR U6465 ( .A(n6283), .B(n6284), .Z(n6299) );
  OR U6466 ( .A(n6246), .B(n6245), .Z(n6250) );
  OR U6467 ( .A(n6248), .B(n6247), .Z(n6249) );
  AND U6468 ( .A(n6250), .B(n6249), .Z(n6298) );
  OR U6469 ( .A(n6252), .B(n6251), .Z(n6256) );
  OR U6470 ( .A(n6254), .B(n6253), .Z(n6255) );
  AND U6471 ( .A(n6256), .B(n6255), .Z(n6297) );
  XNOR U6472 ( .A(n6298), .B(n6297), .Z(n6300) );
  XOR U6473 ( .A(n6299), .B(n6300), .Z(n6278) );
  XOR U6474 ( .A(n6277), .B(n6278), .Z(n6272) );
  NANDN U6475 ( .A(n6258), .B(n6257), .Z(n6262) );
  NANDN U6476 ( .A(n6260), .B(n6259), .Z(n6261) );
  NAND U6477 ( .A(n6262), .B(n6261), .Z(n6269) );
  NAND U6478 ( .A(n6264), .B(n6263), .Z(n6268) );
  OR U6479 ( .A(n6266), .B(n6265), .Z(n6267) );
  NAND U6480 ( .A(n6268), .B(n6267), .Z(n6270) );
  XNOR U6481 ( .A(n6269), .B(n6270), .Z(n6271) );
  XOR U6482 ( .A(n6272), .B(n6271), .Z(N170) );
  NANDN U6483 ( .A(n6270), .B(n6269), .Z(n6274) );
  NANDN U6484 ( .A(n6272), .B(n6271), .Z(n6273) );
  NAND U6485 ( .A(n6274), .B(n6273), .Z(n6320) );
  OR U6486 ( .A(n6276), .B(n6275), .Z(n6280) );
  NANDN U6487 ( .A(n6278), .B(n6277), .Z(n6279) );
  AND U6488 ( .A(n6280), .B(n6279), .Z(n6321) );
  XNOR U6489 ( .A(n6320), .B(n6321), .Z(n6322) );
  NANDN U6490 ( .A(n6282), .B(n6281), .Z(n6286) );
  OR U6491 ( .A(n6284), .B(n6283), .Z(n6285) );
  AND U6492 ( .A(n6286), .B(n6285), .Z(n6383) );
  NANDN U6493 ( .A(n6288), .B(n6287), .Z(n6292) );
  NANDN U6494 ( .A(n6290), .B(n6289), .Z(n6291) );
  NAND U6495 ( .A(n6292), .B(n6291), .Z(n6381) );
  OR U6496 ( .A(n6969), .B(n6663), .Z(n6296) );
  OR U6497 ( .A(n6294), .B(n6293), .Z(n6295) );
  NAND U6498 ( .A(n6296), .B(n6295), .Z(n6380) );
  XOR U6499 ( .A(n6381), .B(n6380), .Z(n6382) );
  XNOR U6500 ( .A(n6383), .B(n6382), .Z(n6328) );
  OR U6501 ( .A(n6298), .B(n6297), .Z(n6302) );
  NANDN U6502 ( .A(n6300), .B(n6299), .Z(n6301) );
  AND U6503 ( .A(n6302), .B(n6301), .Z(n6327) );
  AND U6504 ( .A(y[266]), .B(x[64]), .Z(n6346) );
  ANDN U6505 ( .B(o[73]), .A(n6303), .Z(n6343) );
  AND U6506 ( .A(y[256]), .B(x[74]), .Z(n6344) );
  XNOR U6507 ( .A(n6346), .B(n6345), .Z(n6335) );
  IV U6508 ( .A(y[265]), .Z(n8627) );
  ANDN U6509 ( .B(x[65]), .A(n8627), .Z(n6360) );
  IV U6510 ( .A(n6360), .Z(n7257) );
  AND U6511 ( .A(y[264]), .B(x[66]), .Z(n6358) );
  ANDN U6512 ( .B(y[263]), .A(n48), .Z(n7287) );
  XOR U6513 ( .A(n6358), .B(n7287), .Z(n6359) );
  XOR U6514 ( .A(n7257), .B(n6359), .Z(n6333) );
  AND U6515 ( .A(y[264]), .B(x[70]), .Z(n6634) );
  NANDN U6516 ( .A(n6304), .B(n6634), .Z(n6307) );
  NANDN U6517 ( .A(n6739), .B(n6305), .Z(n6306) );
  AND U6518 ( .A(n6307), .B(n6306), .Z(n6332) );
  XOR U6519 ( .A(n6333), .B(n6332), .Z(n6334) );
  XOR U6520 ( .A(n6335), .B(n6334), .Z(n6374) );
  ANDN U6521 ( .B(y[265]), .A(n54), .Z(n6308) );
  NAND U6522 ( .A(n6748), .B(n6308), .Z(n6312) );
  OR U6523 ( .A(n6310), .B(n6309), .Z(n6311) );
  NAND U6524 ( .A(n6312), .B(n6311), .Z(n6375) );
  XNOR U6525 ( .A(n6374), .B(n6375), .Z(n6377) );
  ANDN U6526 ( .B(y[260]), .A(n52), .Z(n6357) );
  NAND U6527 ( .A(n6357), .B(n6363), .Z(n6316) );
  NANDN U6528 ( .A(n6314), .B(n6313), .Z(n6315) );
  NAND U6529 ( .A(n6316), .B(n6315), .Z(n6371) );
  AND U6530 ( .A(y[260]), .B(x[70]), .Z(n6578) );
  ANDN U6531 ( .B(x[71]), .A(n8881), .Z(n6318) );
  NANDN U6532 ( .A(n49), .B(y[262]), .Z(n6317) );
  XOR U6533 ( .A(n6318), .B(n6317), .Z(n6351) );
  XNOR U6534 ( .A(n6578), .B(n6351), .Z(n6368) );
  ANDN U6535 ( .B(y[258]), .A(n53), .Z(n6319) );
  XOR U6536 ( .A(n6319), .B(n6518), .Z(n6365) );
  NANDN U6537 ( .A(n54), .B(y[257]), .Z(n6338) );
  XOR U6538 ( .A(o[74]), .B(n6338), .Z(n6364) );
  XOR U6539 ( .A(n6365), .B(n6364), .Z(n6369) );
  XOR U6540 ( .A(n6371), .B(n6370), .Z(n6376) );
  XNOR U6541 ( .A(n6377), .B(n6376), .Z(n6326) );
  XNOR U6542 ( .A(n6328), .B(n6329), .Z(n6323) );
  XOR U6543 ( .A(n6322), .B(n6323), .Z(N171) );
  NANDN U6544 ( .A(n6321), .B(n6320), .Z(n6325) );
  NANDN U6545 ( .A(n6323), .B(n6322), .Z(n6324) );
  NAND U6546 ( .A(n6325), .B(n6324), .Z(n6386) );
  OR U6547 ( .A(n6327), .B(n6326), .Z(n6331) );
  OR U6548 ( .A(n6329), .B(n6328), .Z(n6330) );
  AND U6549 ( .A(n6331), .B(n6330), .Z(n6387) );
  XNOR U6550 ( .A(n6386), .B(n6387), .Z(n6388) );
  OR U6551 ( .A(n6333), .B(n6332), .Z(n6337) );
  NAND U6552 ( .A(n6335), .B(n6334), .Z(n6336) );
  NAND U6553 ( .A(n6337), .B(n6336), .Z(n6401) );
  NANDN U6554 ( .A(n6338), .B(o[74]), .Z(n6422) );
  ANDN U6555 ( .B(x[75]), .A(n8872), .Z(n6340) );
  NANDN U6556 ( .A(n45), .B(y[267]), .Z(n6339) );
  XOR U6557 ( .A(n6340), .B(n6339), .Z(n6421) );
  IV U6558 ( .A(y[266]), .Z(n7862) );
  ANDN U6559 ( .B(x[65]), .A(n7862), .Z(n6342) );
  NANDN U6560 ( .A(n51), .B(y[261]), .Z(n6341) );
  XOR U6561 ( .A(n6342), .B(n6341), .Z(n6447) );
  NANDN U6562 ( .A(n55), .B(y[257]), .Z(n6429) );
  XOR U6563 ( .A(o[75]), .B(n6429), .Z(n6446) );
  XOR U6564 ( .A(n6447), .B(n6446), .Z(n6404) );
  OR U6565 ( .A(n6344), .B(n6343), .Z(n6348) );
  OR U6566 ( .A(n6346), .B(n6345), .Z(n6347) );
  NAND U6567 ( .A(n6348), .B(n6347), .Z(n6407) );
  XNOR U6568 ( .A(n6406), .B(n6407), .Z(n6398) );
  ANDN U6569 ( .B(y[262]), .A(n52), .Z(n6350) );
  NAND U6570 ( .A(n6350), .B(n6349), .Z(n6353) );
  NANDN U6571 ( .A(n6351), .B(n6578), .Z(n6352) );
  NAND U6572 ( .A(n6353), .B(n6352), .Z(n6399) );
  XOR U6573 ( .A(n6401), .B(n6400), .Z(n6453) );
  ANDN U6574 ( .B(y[264]), .A(n48), .Z(n7420) );
  ANDN U6575 ( .B(x[66]), .A(n8627), .Z(n6355) );
  NANDN U6576 ( .A(n50), .B(y[262]), .Z(n6354) );
  XOR U6577 ( .A(n6355), .B(n6354), .Z(n6441) );
  NANDN U6578 ( .A(n49), .B(y[263]), .Z(n6440) );
  XNOR U6579 ( .A(n6441), .B(n6440), .Z(n6410) );
  XOR U6580 ( .A(n7420), .B(n6410), .Z(n6412) );
  NANDN U6581 ( .A(n54), .B(y[258]), .Z(n6356) );
  XOR U6582 ( .A(n6357), .B(n6356), .Z(n6426) );
  NANDN U6583 ( .A(n8881), .B(x[72]), .Z(n6425) );
  XOR U6584 ( .A(n6426), .B(n6425), .Z(n6411) );
  XNOR U6585 ( .A(n6412), .B(n6411), .Z(n6418) );
  OR U6586 ( .A(n6358), .B(n7287), .Z(n6362) );
  NANDN U6587 ( .A(n6360), .B(n6359), .Z(n6361) );
  AND U6588 ( .A(n6362), .B(n6361), .Z(n6415) );
  AND U6589 ( .A(y[261]), .B(x[72]), .Z(n7153) );
  NAND U6590 ( .A(n7153), .B(n6363), .Z(n6367) );
  OR U6591 ( .A(n6365), .B(n6364), .Z(n6366) );
  NAND U6592 ( .A(n6367), .B(n6366), .Z(n6416) );
  XNOR U6593 ( .A(n6418), .B(n6417), .Z(n6450) );
  OR U6594 ( .A(n6369), .B(n6368), .Z(n6373) );
  NANDN U6595 ( .A(n6371), .B(n6370), .Z(n6372) );
  NAND U6596 ( .A(n6373), .B(n6372), .Z(n6451) );
  XOR U6597 ( .A(n6450), .B(n6451), .Z(n6452) );
  XOR U6598 ( .A(n6453), .B(n6452), .Z(n6392) );
  OR U6599 ( .A(n6375), .B(n6374), .Z(n6379) );
  OR U6600 ( .A(n6377), .B(n6376), .Z(n6378) );
  AND U6601 ( .A(n6379), .B(n6378), .Z(n6393) );
  XNOR U6602 ( .A(n6392), .B(n6393), .Z(n6395) );
  OR U6603 ( .A(n6381), .B(n6380), .Z(n6385) );
  NANDN U6604 ( .A(n6383), .B(n6382), .Z(n6384) );
  NAND U6605 ( .A(n6385), .B(n6384), .Z(n6394) );
  XOR U6606 ( .A(n6395), .B(n6394), .Z(n6389) );
  XNOR U6607 ( .A(n6388), .B(n6389), .Z(N172) );
  NANDN U6608 ( .A(n6387), .B(n6386), .Z(n6391) );
  NAND U6609 ( .A(n6389), .B(n6388), .Z(n6390) );
  NAND U6610 ( .A(n6391), .B(n6390), .Z(n6456) );
  OR U6611 ( .A(n6393), .B(n6392), .Z(n6397) );
  OR U6612 ( .A(n6395), .B(n6394), .Z(n6396) );
  AND U6613 ( .A(n6397), .B(n6396), .Z(n6457) );
  XNOR U6614 ( .A(n6456), .B(n6457), .Z(n6458) );
  OR U6615 ( .A(n6399), .B(n6398), .Z(n6403) );
  NANDN U6616 ( .A(n6401), .B(n6400), .Z(n6402) );
  NAND U6617 ( .A(n6403), .B(n6402), .Z(n6526) );
  NANDN U6618 ( .A(n6405), .B(n6404), .Z(n6409) );
  NANDN U6619 ( .A(n6407), .B(n6406), .Z(n6408) );
  AND U6620 ( .A(n6409), .B(n6408), .Z(n6523) );
  NANDN U6621 ( .A(n6410), .B(n7420), .Z(n6414) );
  NANDN U6622 ( .A(n6412), .B(n6411), .Z(n6413) );
  AND U6623 ( .A(n6414), .B(n6413), .Z(n6524) );
  XOR U6624 ( .A(n6526), .B(n6525), .Z(n6464) );
  OR U6625 ( .A(n6416), .B(n6415), .Z(n6420) );
  NANDN U6626 ( .A(n6418), .B(n6417), .Z(n6419) );
  NAND U6627 ( .A(n6420), .B(n6419), .Z(n6531) );
  AND U6628 ( .A(y[267]), .B(x[75]), .Z(n7574) );
  NAND U6629 ( .A(n6748), .B(n7574), .Z(n6424) );
  OR U6630 ( .A(n6422), .B(n6421), .Z(n6423) );
  AND U6631 ( .A(n6424), .B(n6423), .Z(n6470) );
  NANDN U6632 ( .A(n52), .B(y[258]), .Z(n6641) );
  NANDN U6633 ( .A(n54), .B(y[260]), .Z(n7021) );
  OR U6634 ( .A(n6641), .B(n7021), .Z(n6428) );
  OR U6635 ( .A(n6426), .B(n6425), .Z(n6427) );
  AND U6636 ( .A(n6428), .B(n6427), .Z(n6468) );
  NANDN U6637 ( .A(n6429), .B(o[75]), .Z(n6475) );
  ANDN U6638 ( .B(y[267]), .A(n46), .Z(n6431) );
  NANDN U6639 ( .A(n51), .B(y[262]), .Z(n6430) );
  XOR U6640 ( .A(n6431), .B(n6430), .Z(n6474) );
  XNOR U6641 ( .A(n6475), .B(n6474), .Z(n6469) );
  XNOR U6642 ( .A(n6468), .B(n6469), .Z(n6471) );
  XOR U6643 ( .A(n6470), .B(n6471), .Z(n6529) );
  ANDN U6644 ( .B(x[71]), .A(n7989), .Z(n6433) );
  NANDN U6645 ( .A(n50), .B(y[263]), .Z(n6432) );
  XOR U6646 ( .A(n6433), .B(n6432), .Z(n6520) );
  NANDN U6647 ( .A(n49), .B(y[264]), .Z(n6491) );
  ANDN U6648 ( .B(y[258]), .A(n55), .Z(n6435) );
  NANDN U6649 ( .A(n54), .B(y[259]), .Z(n6434) );
  XOR U6650 ( .A(n6435), .B(n6434), .Z(n6490) );
  XNOR U6651 ( .A(n6491), .B(n6490), .Z(n6519) );
  XNOR U6652 ( .A(n6520), .B(n6519), .Z(n6514) );
  ANDN U6653 ( .B(x[76]), .A(n8872), .Z(n6437) );
  NANDN U6654 ( .A(n45), .B(y[268]), .Z(n6436) );
  XOR U6655 ( .A(n6437), .B(n6436), .Z(n6479) );
  NANDN U6656 ( .A(n56), .B(y[257]), .Z(n6508) );
  XOR U6657 ( .A(o[76]), .B(n6508), .Z(n6478) );
  XOR U6658 ( .A(n6479), .B(n6478), .Z(n6511) );
  ANDN U6659 ( .B(x[66]), .A(n7862), .Z(n6439) );
  NANDN U6660 ( .A(n53), .B(y[260]), .Z(n6438) );
  XOR U6661 ( .A(n6439), .B(n6438), .Z(n6503) );
  NANDN U6662 ( .A(n8627), .B(x[67]), .Z(n6502) );
  XNOR U6663 ( .A(n6503), .B(n6502), .Z(n6512) );
  XOR U6664 ( .A(n6511), .B(n6512), .Z(n6513) );
  XOR U6665 ( .A(n6514), .B(n6513), .Z(n6497) );
  AND U6666 ( .A(y[265]), .B(x[69]), .Z(n6664) );
  NANDN U6667 ( .A(n6758), .B(n6664), .Z(n6443) );
  OR U6668 ( .A(n6441), .B(n6440), .Z(n6442) );
  NAND U6669 ( .A(n6443), .B(n6442), .Z(n6495) );
  ANDN U6670 ( .B(y[266]), .A(n51), .Z(n6445) );
  NAND U6671 ( .A(n6445), .B(n6444), .Z(n6449) );
  OR U6672 ( .A(n6447), .B(n6446), .Z(n6448) );
  NAND U6673 ( .A(n6449), .B(n6448), .Z(n6494) );
  XOR U6674 ( .A(n6495), .B(n6494), .Z(n6496) );
  XOR U6675 ( .A(n6497), .B(n6496), .Z(n6530) );
  XOR U6676 ( .A(n6531), .B(n6532), .Z(n6462) );
  OR U6677 ( .A(n6451), .B(n6450), .Z(n6455) );
  NAND U6678 ( .A(n6453), .B(n6452), .Z(n6454) );
  AND U6679 ( .A(n6455), .B(n6454), .Z(n6463) );
  XOR U6680 ( .A(n6462), .B(n6463), .Z(n6465) );
  XOR U6681 ( .A(n6464), .B(n6465), .Z(n6459) );
  XOR U6682 ( .A(n6458), .B(n6459), .Z(N173) );
  NANDN U6683 ( .A(n6457), .B(n6456), .Z(n6461) );
  NANDN U6684 ( .A(n6459), .B(n6458), .Z(n6460) );
  NAND U6685 ( .A(n6461), .B(n6460), .Z(n6601) );
  NANDN U6686 ( .A(n6463), .B(n6462), .Z(n6467) );
  OR U6687 ( .A(n6465), .B(n6464), .Z(n6466) );
  NAND U6688 ( .A(n6467), .B(n6466), .Z(n6602) );
  XNOR U6689 ( .A(n6601), .B(n6602), .Z(n6603) );
  OR U6690 ( .A(n6469), .B(n6468), .Z(n6473) );
  OR U6691 ( .A(n6471), .B(n6470), .Z(n6472) );
  NAND U6692 ( .A(n6473), .B(n6472), .Z(n6550) );
  AND U6693 ( .A(y[267]), .B(x[70]), .Z(n6976) );
  NAND U6694 ( .A(n6976), .B(n6565), .Z(n6477) );
  OR U6695 ( .A(n6475), .B(n6474), .Z(n6476) );
  NAND U6696 ( .A(n6477), .B(n6476), .Z(n6556) );
  AND U6697 ( .A(y[268]), .B(x[76]), .Z(n7793) );
  NAND U6698 ( .A(n6748), .B(n7793), .Z(n6481) );
  OR U6699 ( .A(n6479), .B(n6478), .Z(n6480) );
  AND U6700 ( .A(n6481), .B(n6480), .Z(n6553) );
  ANDN U6701 ( .B(y[258]), .A(n56), .Z(n6483) );
  NANDN U6702 ( .A(n55), .B(y[259]), .Z(n6482) );
  XNOR U6703 ( .A(n6483), .B(n6482), .Z(n6571) );
  XNOR U6704 ( .A(n7153), .B(n6571), .Z(n6554) );
  XOR U6705 ( .A(n6556), .B(n6555), .Z(n6548) );
  ANDN U6706 ( .B(x[67]), .A(n7862), .Z(n6485) );
  NANDN U6707 ( .A(n50), .B(y[264]), .Z(n6484) );
  XOR U6708 ( .A(n6485), .B(n6484), .Z(n6588) );
  NANDN U6709 ( .A(n8627), .B(x[68]), .Z(n6587) );
  XNOR U6710 ( .A(n6588), .B(n6587), .Z(n6595) );
  ANDN U6711 ( .B(x[77]), .A(n8872), .Z(n6487) );
  NANDN U6712 ( .A(n45), .B(y[269]), .Z(n6486) );
  XOR U6713 ( .A(n6487), .B(n6486), .Z(n6592) );
  NANDN U6714 ( .A(n57), .B(y[257]), .Z(n6584) );
  XOR U6715 ( .A(o[77]), .B(n6584), .Z(n6591) );
  XNOR U6716 ( .A(n6592), .B(n6591), .Z(n6596) );
  ANDN U6717 ( .B(y[258]), .A(n54), .Z(n6489) );
  ANDN U6718 ( .B(y[259]), .A(n55), .Z(n6488) );
  NAND U6719 ( .A(n6489), .B(n6488), .Z(n6493) );
  OR U6720 ( .A(n6491), .B(n6490), .Z(n6492) );
  AND U6721 ( .A(n6493), .B(n6492), .Z(n6597) );
  XNOR U6722 ( .A(n6598), .B(n6597), .Z(n6547) );
  XOR U6723 ( .A(n6548), .B(n6547), .Z(n6549) );
  XNOR U6724 ( .A(n6550), .B(n6549), .Z(n6544) );
  OR U6725 ( .A(n6495), .B(n6494), .Z(n6499) );
  NANDN U6726 ( .A(n6497), .B(n6496), .Z(n6498) );
  AND U6727 ( .A(n6499), .B(n6498), .Z(n6541) );
  ANDN U6728 ( .B(y[266]), .A(n53), .Z(n6501) );
  NAND U6729 ( .A(n6501), .B(n6500), .Z(n6505) );
  OR U6730 ( .A(n6503), .B(n6502), .Z(n6504) );
  NAND U6731 ( .A(n6505), .B(n6504), .Z(n6562) );
  NANDN U6732 ( .A(n47), .B(y[267]), .Z(n6580) );
  ANDN U6733 ( .B(y[263]), .A(n51), .Z(n6507) );
  ANDN U6734 ( .B(y[260]), .A(n54), .Z(n6506) );
  XNOR U6735 ( .A(n6507), .B(n6506), .Z(n6579) );
  XNOR U6736 ( .A(n6580), .B(n6579), .Z(n6560) );
  NANDN U6737 ( .A(n6508), .B(o[76]), .Z(n6568) );
  ANDN U6738 ( .B(y[268]), .A(n46), .Z(n6510) );
  NANDN U6739 ( .A(n52), .B(y[262]), .Z(n6509) );
  XOR U6740 ( .A(n6510), .B(n6509), .Z(n6567) );
  XNOR U6741 ( .A(n6562), .B(n6561), .Z(n6538) );
  NANDN U6742 ( .A(n6512), .B(n6511), .Z(n6516) );
  OR U6743 ( .A(n6514), .B(n6513), .Z(n6515) );
  AND U6744 ( .A(n6516), .B(n6515), .Z(n6535) );
  ANDN U6745 ( .B(y[263]), .A(n52), .Z(n6517) );
  NANDN U6746 ( .A(n6518), .B(n6517), .Z(n6522) );
  OR U6747 ( .A(n6520), .B(n6519), .Z(n6521) );
  AND U6748 ( .A(n6522), .B(n6521), .Z(n6536) );
  XOR U6749 ( .A(n6535), .B(n6536), .Z(n6537) );
  XNOR U6750 ( .A(n6538), .B(n6537), .Z(n6542) );
  XOR U6751 ( .A(n6541), .B(n6542), .Z(n6543) );
  XNOR U6752 ( .A(n6544), .B(n6543), .Z(n6610) );
  OR U6753 ( .A(n6524), .B(n6523), .Z(n6528) );
  NANDN U6754 ( .A(n6526), .B(n6525), .Z(n6527) );
  AND U6755 ( .A(n6528), .B(n6527), .Z(n6607) );
  OR U6756 ( .A(n6530), .B(n6529), .Z(n6534) );
  NANDN U6757 ( .A(n6532), .B(n6531), .Z(n6533) );
  NAND U6758 ( .A(n6534), .B(n6533), .Z(n6608) );
  XNOR U6759 ( .A(n6610), .B(n6609), .Z(n6604) );
  XOR U6760 ( .A(n6603), .B(n6604), .Z(N174) );
  OR U6761 ( .A(n6536), .B(n6535), .Z(n6540) );
  NANDN U6762 ( .A(n6538), .B(n6537), .Z(n6539) );
  NAND U6763 ( .A(n6540), .B(n6539), .Z(n6622) );
  OR U6764 ( .A(n6542), .B(n6541), .Z(n6546) );
  NANDN U6765 ( .A(n6544), .B(n6543), .Z(n6545) );
  AND U6766 ( .A(n6546), .B(n6545), .Z(n6619) );
  NANDN U6767 ( .A(n6548), .B(n6547), .Z(n6552) );
  OR U6768 ( .A(n6550), .B(n6549), .Z(n6551) );
  AND U6769 ( .A(n6552), .B(n6551), .Z(n6699) );
  OR U6770 ( .A(n6554), .B(n6553), .Z(n6558) );
  NAND U6771 ( .A(n6556), .B(n6555), .Z(n6557) );
  NAND U6772 ( .A(n6558), .B(n6557), .Z(n6692) );
  NANDN U6773 ( .A(n6560), .B(n6559), .Z(n6564) );
  NAND U6774 ( .A(n6562), .B(n6561), .Z(n6563) );
  AND U6775 ( .A(n6564), .B(n6563), .Z(n6690) );
  ANDN U6776 ( .B(y[268]), .A(n52), .Z(n6566) );
  NAND U6777 ( .A(n6566), .B(n6565), .Z(n6570) );
  OR U6778 ( .A(n6568), .B(n6567), .Z(n6569) );
  AND U6779 ( .A(n6570), .B(n6569), .Z(n6684) );
  NANDN U6780 ( .A(n55), .B(y[258]), .Z(n7158) );
  ANDN U6781 ( .B(x[75]), .A(n8881), .Z(n6632) );
  IV U6782 ( .A(n6632), .Z(n6779) );
  OR U6783 ( .A(n7158), .B(n6779), .Z(n6573) );
  NAND U6784 ( .A(n6571), .B(n7153), .Z(n6572) );
  AND U6785 ( .A(n6573), .B(n6572), .Z(n6685) );
  XOR U6786 ( .A(n6684), .B(n6685), .Z(n6687) );
  AND U6787 ( .A(y[266]), .B(x[68]), .Z(n6678) );
  AND U6788 ( .A(y[260]), .B(x[74]), .Z(n7293) );
  ANDN U6789 ( .B(y[268]), .A(n47), .Z(n6575) );
  NANDN U6790 ( .A(n54), .B(y[261]), .Z(n6574) );
  XOR U6791 ( .A(n6575), .B(n6574), .Z(n6638) );
  XNOR U6792 ( .A(n7293), .B(n6638), .Z(n6679) );
  XNOR U6793 ( .A(n6678), .B(n6679), .Z(n6681) );
  ANDN U6794 ( .B(y[267]), .A(n48), .Z(n6577) );
  ANDN U6795 ( .B(x[72]), .A(n8655), .Z(n6576) );
  XNOR U6796 ( .A(n6577), .B(n6576), .Z(n6665) );
  XNOR U6797 ( .A(n6664), .B(n6665), .Z(n6680) );
  XNOR U6798 ( .A(n6681), .B(n6680), .Z(n6686) );
  XNOR U6799 ( .A(n6687), .B(n6686), .Z(n6691) );
  XOR U6800 ( .A(n6692), .B(n6693), .Z(n6696) );
  ANDN U6801 ( .B(y[263]), .A(n54), .Z(n6775) );
  NAND U6802 ( .A(n6775), .B(n6578), .Z(n6582) );
  OR U6803 ( .A(n6580), .B(n6579), .Z(n6581) );
  NAND U6804 ( .A(n6582), .B(n6581), .Z(n6653) );
  ANDN U6805 ( .B(y[257]), .A(n58), .Z(n6646) );
  XNOR U6806 ( .A(o[78]), .B(n6646), .Z(n6643) );
  ANDN U6807 ( .B(y[258]), .A(n57), .Z(n7252) );
  NANDN U6808 ( .A(n52), .B(y[263]), .Z(n6583) );
  XNOR U6809 ( .A(n7252), .B(n6583), .Z(n6642) );
  XOR U6810 ( .A(n6643), .B(n6642), .Z(n6652) );
  NANDN U6811 ( .A(n6584), .B(o[77]), .Z(n6669) );
  ANDN U6812 ( .B(x[78]), .A(n8872), .Z(n6586) );
  NANDN U6813 ( .A(n45), .B(y[270]), .Z(n6585) );
  XOR U6814 ( .A(n6586), .B(n6585), .Z(n6668) );
  XOR U6815 ( .A(n6652), .B(n6651), .Z(n6654) );
  XNOR U6816 ( .A(n6653), .B(n6654), .Z(n6625) );
  AND U6817 ( .A(y[266]), .B(x[69]), .Z(n6732) );
  NAND U6818 ( .A(n7420), .B(n6732), .Z(n6590) );
  OR U6819 ( .A(n6588), .B(n6587), .Z(n6589) );
  NAND U6820 ( .A(n6590), .B(n6589), .Z(n6660) );
  NAND U6821 ( .A(y[269]), .B(x[65]), .Z(n6631) );
  XOR U6822 ( .A(n6632), .B(n6631), .Z(n6633) );
  XOR U6823 ( .A(n6634), .B(n6633), .Z(n6658) );
  IV U6824 ( .A(y[269]), .Z(n8815) );
  NANDN U6825 ( .A(n8815), .B(x[77]), .Z(n8173) );
  NANDN U6826 ( .A(n8173), .B(n6748), .Z(n6594) );
  OR U6827 ( .A(n6592), .B(n6591), .Z(n6593) );
  AND U6828 ( .A(n6594), .B(n6593), .Z(n6657) );
  XOR U6829 ( .A(n6658), .B(n6657), .Z(n6659) );
  XOR U6830 ( .A(n6660), .B(n6659), .Z(n6626) );
  XNOR U6831 ( .A(n6625), .B(n6626), .Z(n6628) );
  OR U6832 ( .A(n6596), .B(n6595), .Z(n6600) );
  OR U6833 ( .A(n6598), .B(n6597), .Z(n6599) );
  NAND U6834 ( .A(n6600), .B(n6599), .Z(n6627) );
  XNOR U6835 ( .A(n6628), .B(n6627), .Z(n6697) );
  XNOR U6836 ( .A(n6696), .B(n6697), .Z(n6698) );
  XOR U6837 ( .A(n6699), .B(n6698), .Z(n6620) );
  XNOR U6838 ( .A(n6619), .B(n6620), .Z(n6621) );
  XNOR U6839 ( .A(n6622), .B(n6621), .Z(n6616) );
  NANDN U6840 ( .A(n6602), .B(n6601), .Z(n6606) );
  NANDN U6841 ( .A(n6604), .B(n6603), .Z(n6605) );
  NAND U6842 ( .A(n6606), .B(n6605), .Z(n6613) );
  OR U6843 ( .A(n6608), .B(n6607), .Z(n6612) );
  NANDN U6844 ( .A(n6610), .B(n6609), .Z(n6611) );
  NAND U6845 ( .A(n6612), .B(n6611), .Z(n6614) );
  XNOR U6846 ( .A(n6613), .B(n6614), .Z(n6615) );
  XOR U6847 ( .A(n6616), .B(n6615), .Z(N175) );
  NANDN U6848 ( .A(n6614), .B(n6613), .Z(n6618) );
  NANDN U6849 ( .A(n6616), .B(n6615), .Z(n6617) );
  NAND U6850 ( .A(n6618), .B(n6617), .Z(n6702) );
  OR U6851 ( .A(n6620), .B(n6619), .Z(n6624) );
  OR U6852 ( .A(n6622), .B(n6621), .Z(n6623) );
  AND U6853 ( .A(n6624), .B(n6623), .Z(n6703) );
  XNOR U6854 ( .A(n6702), .B(n6703), .Z(n6704) );
  OR U6855 ( .A(n6626), .B(n6625), .Z(n6630) );
  OR U6856 ( .A(n6628), .B(n6627), .Z(n6629) );
  AND U6857 ( .A(n6630), .B(n6629), .Z(n6709) );
  NANDN U6858 ( .A(n6632), .B(n6631), .Z(n6636) );
  OR U6859 ( .A(n6634), .B(n6633), .Z(n6635) );
  AND U6860 ( .A(n6636), .B(n6635), .Z(n6728) );
  AND U6861 ( .A(y[268]), .B(x[73]), .Z(n7383) );
  NANDN U6862 ( .A(n6637), .B(n7383), .Z(n6640) );
  NANDN U6863 ( .A(n6638), .B(n7293), .Z(n6639) );
  NAND U6864 ( .A(n6640), .B(n6639), .Z(n6727) );
  ANDN U6865 ( .B(y[263]), .A(n57), .Z(n7027) );
  NANDN U6866 ( .A(n6641), .B(n7027), .Z(n6645) );
  NANDN U6867 ( .A(n6643), .B(n6642), .Z(n6644) );
  NAND U6868 ( .A(n6645), .B(n6644), .Z(n6787) );
  NAND U6869 ( .A(n6646), .B(o[78]), .Z(n6750) );
  ANDN U6870 ( .B(x[79]), .A(n8872), .Z(n6648) );
  ANDN U6871 ( .B(y[271]), .A(n45), .Z(n6647) );
  XNOR U6872 ( .A(n6648), .B(n6647), .Z(n6749) );
  XOR U6873 ( .A(n6750), .B(n6749), .Z(n6784) );
  NANDN U6874 ( .A(n58), .B(y[258]), .Z(n6781) );
  ANDN U6875 ( .B(x[76]), .A(n8881), .Z(n6650) );
  NANDN U6876 ( .A(n56), .B(y[260]), .Z(n6649) );
  XOR U6877 ( .A(n6650), .B(n6649), .Z(n6780) );
  XOR U6878 ( .A(n6781), .B(n6780), .Z(n6785) );
  XNOR U6879 ( .A(n6784), .B(n6785), .Z(n6786) );
  XNOR U6880 ( .A(n6787), .B(n6786), .Z(n6726) );
  XNOR U6881 ( .A(n6727), .B(n6726), .Z(n6729) );
  XOR U6882 ( .A(n6728), .B(n6729), .Z(n6714) );
  NANDN U6883 ( .A(n6652), .B(n6651), .Z(n6656) );
  NANDN U6884 ( .A(n6654), .B(n6653), .Z(n6655) );
  AND U6885 ( .A(n6656), .B(n6655), .Z(n6715) );
  XNOR U6886 ( .A(n6714), .B(n6715), .Z(n6717) );
  OR U6887 ( .A(n6658), .B(n6657), .Z(n6662) );
  NAND U6888 ( .A(n6660), .B(n6659), .Z(n6661) );
  AND U6889 ( .A(n6662), .B(n6661), .Z(n6716) );
  XNOR U6890 ( .A(n6717), .B(n6716), .Z(n6792) );
  NANDN U6891 ( .A(n53), .B(y[267]), .Z(n7068) );
  NANDN U6892 ( .A(n7068), .B(n6663), .Z(n6667) );
  NANDN U6893 ( .A(n6665), .B(n6664), .Z(n6666) );
  NAND U6894 ( .A(n6667), .B(n6666), .Z(n6764) );
  IV U6895 ( .A(y[270]), .Z(n8861) );
  ANDN U6896 ( .B(x[78]), .A(n8861), .Z(n8392) );
  NAND U6897 ( .A(n6748), .B(n8392), .Z(n6671) );
  OR U6898 ( .A(n6669), .B(n6668), .Z(n6670) );
  NAND U6899 ( .A(n6671), .B(n6670), .Z(n6763) );
  XNOR U6900 ( .A(n6764), .B(n6763), .Z(n6765) );
  ANDN U6901 ( .B(y[257]), .A(n59), .Z(n6753) );
  XNOR U6902 ( .A(o[79]), .B(n6753), .Z(n6745) );
  ANDN U6903 ( .B(y[270]), .A(n46), .Z(n6673) );
  ANDN U6904 ( .B(y[263]), .A(n53), .Z(n6672) );
  XNOR U6905 ( .A(n6673), .B(n6672), .Z(n6744) );
  XOR U6906 ( .A(n6745), .B(n6744), .Z(n6769) );
  NANDN U6907 ( .A(n48), .B(y[268]), .Z(n6760) );
  ANDN U6908 ( .B(x[66]), .A(n8815), .Z(n6675) );
  NANDN U6909 ( .A(n54), .B(y[262]), .Z(n6674) );
  XOR U6910 ( .A(n6675), .B(n6674), .Z(n6759) );
  XOR U6911 ( .A(n6760), .B(n6759), .Z(n6770) );
  XNOR U6912 ( .A(n6769), .B(n6770), .Z(n6772) );
  AND U6913 ( .A(y[264]), .B(x[71]), .Z(n7184) );
  ANDN U6914 ( .B(x[74]), .A(n7989), .Z(n6677) );
  ANDN U6915 ( .B(y[267]), .A(n49), .Z(n6676) );
  XNOR U6916 ( .A(n6677), .B(n6676), .Z(n6740) );
  XNOR U6917 ( .A(n7184), .B(n6740), .Z(n6733) );
  ANDN U6918 ( .B(x[70]), .A(n8627), .Z(n6864) );
  XNOR U6919 ( .A(n6732), .B(n6864), .Z(n6734) );
  XNOR U6920 ( .A(n6733), .B(n6734), .Z(n6771) );
  XNOR U6921 ( .A(n6772), .B(n6771), .Z(n6766) );
  OR U6922 ( .A(n6679), .B(n6678), .Z(n6683) );
  OR U6923 ( .A(n6681), .B(n6680), .Z(n6682) );
  NAND U6924 ( .A(n6683), .B(n6682), .Z(n6721) );
  XNOR U6925 ( .A(n6720), .B(n6721), .Z(n6723) );
  OR U6926 ( .A(n6685), .B(n6684), .Z(n6689) );
  NAND U6927 ( .A(n6687), .B(n6686), .Z(n6688) );
  AND U6928 ( .A(n6689), .B(n6688), .Z(n6722) );
  XNOR U6929 ( .A(n6723), .B(n6722), .Z(n6790) );
  OR U6930 ( .A(n6691), .B(n6690), .Z(n6695) );
  NANDN U6931 ( .A(n6693), .B(n6692), .Z(n6694) );
  NAND U6932 ( .A(n6695), .B(n6694), .Z(n6791) );
  XOR U6933 ( .A(n6790), .B(n6791), .Z(n6793) );
  XOR U6934 ( .A(n6792), .B(n6793), .Z(n6708) );
  NANDN U6935 ( .A(n6697), .B(n6696), .Z(n6701) );
  NANDN U6936 ( .A(n6699), .B(n6698), .Z(n6700) );
  AND U6937 ( .A(n6701), .B(n6700), .Z(n6710) );
  XNOR U6938 ( .A(n6711), .B(n6710), .Z(n6705) );
  XOR U6939 ( .A(n6704), .B(n6705), .Z(N176) );
  NANDN U6940 ( .A(n6703), .B(n6702), .Z(n6707) );
  NANDN U6941 ( .A(n6705), .B(n6704), .Z(n6706) );
  NAND U6942 ( .A(n6707), .B(n6706), .Z(n6796) );
  OR U6943 ( .A(n6709), .B(n6708), .Z(n6713) );
  OR U6944 ( .A(n6711), .B(n6710), .Z(n6712) );
  AND U6945 ( .A(n6713), .B(n6712), .Z(n6797) );
  XNOR U6946 ( .A(n6796), .B(n6797), .Z(n6798) );
  OR U6947 ( .A(n6715), .B(n6714), .Z(n6719) );
  OR U6948 ( .A(n6717), .B(n6716), .Z(n6718) );
  NAND U6949 ( .A(n6719), .B(n6718), .Z(n6886) );
  OR U6950 ( .A(n6721), .B(n6720), .Z(n6725) );
  OR U6951 ( .A(n6723), .B(n6722), .Z(n6724) );
  NAND U6952 ( .A(n6725), .B(n6724), .Z(n6884) );
  OR U6953 ( .A(n6727), .B(n6726), .Z(n6731) );
  OR U6954 ( .A(n6729), .B(n6728), .Z(n6730) );
  AND U6955 ( .A(n6731), .B(n6730), .Z(n6883) );
  XOR U6956 ( .A(n6884), .B(n6883), .Z(n6885) );
  XNOR U6957 ( .A(n6886), .B(n6885), .Z(n6805) );
  OR U6958 ( .A(n6732), .B(n6864), .Z(n6736) );
  OR U6959 ( .A(n6734), .B(n6733), .Z(n6735) );
  AND U6960 ( .A(n6736), .B(n6735), .Z(n6842) );
  NANDN U6961 ( .A(n8890), .B(y[256]), .Z(n6871) );
  IV U6962 ( .A(y[272]), .Z(n8884) );
  ANDN U6963 ( .B(x[64]), .A(n8884), .Z(n6870) );
  XNOR U6964 ( .A(n6871), .B(n6870), .Z(n6873) );
  NANDN U6965 ( .A(n60), .B(y[257]), .Z(n6876) );
  XNOR U6966 ( .A(n6876), .B(o[80]), .Z(n6872) );
  XNOR U6967 ( .A(n6873), .B(n6872), .Z(n6855) );
  NANDN U6968 ( .A(n55), .B(y[262]), .Z(n6866) );
  ANDN U6969 ( .B(x[71]), .A(n8627), .Z(n6738) );
  NANDN U6970 ( .A(n51), .B(y[266]), .Z(n6737) );
  XOR U6971 ( .A(n6738), .B(n6737), .Z(n6865) );
  XNOR U6972 ( .A(n6866), .B(n6865), .Z(n6854) );
  XNOR U6973 ( .A(n6855), .B(n6854), .Z(n6857) );
  AND U6974 ( .A(y[267]), .B(x[74]), .Z(n7415) );
  NANDN U6975 ( .A(n6739), .B(n7415), .Z(n6742) );
  NANDN U6976 ( .A(n6740), .B(n7184), .Z(n6741) );
  AND U6977 ( .A(n6742), .B(n6741), .Z(n6856) );
  XOR U6978 ( .A(n6857), .B(n6856), .Z(n6827) );
  NANDN U6979 ( .A(n53), .B(y[270]), .Z(n7678) );
  NANDN U6980 ( .A(n7678), .B(n6743), .Z(n6747) );
  OR U6981 ( .A(n6745), .B(n6744), .Z(n6746) );
  AND U6982 ( .A(n6747), .B(n6746), .Z(n6824) );
  ANDN U6983 ( .B(y[271]), .A(n60), .Z(n8957) );
  NAND U6984 ( .A(n6748), .B(n8957), .Z(n6752) );
  OR U6985 ( .A(n6750), .B(n6749), .Z(n6751) );
  AND U6986 ( .A(n6752), .B(n6751), .Z(n6825) );
  XOR U6987 ( .A(n6824), .B(n6825), .Z(n6826) );
  XOR U6988 ( .A(n6827), .B(n6826), .Z(n6843) );
  XOR U6989 ( .A(n6842), .B(n6843), .Z(n6844) );
  NAND U6990 ( .A(o[79]), .B(n6753), .Z(n6861) );
  ANDN U6991 ( .B(y[271]), .A(n46), .Z(n6755) );
  ANDN U6992 ( .B(x[72]), .A(n8927), .Z(n6754) );
  XNOR U6993 ( .A(n6755), .B(n6754), .Z(n6860) );
  XNOR U6994 ( .A(n6861), .B(n6860), .Z(n6850) );
  NANDN U6995 ( .A(n49), .B(y[268]), .Z(n6815) );
  ANDN U6996 ( .B(x[75]), .A(n7989), .Z(n6757) );
  ANDN U6997 ( .B(y[258]), .A(n59), .Z(n6756) );
  XNOR U6998 ( .A(n6757), .B(n6756), .Z(n6814) );
  XOR U6999 ( .A(n6815), .B(n6814), .Z(n6849) );
  AND U7000 ( .A(y[269]), .B(x[73]), .Z(n7515) );
  NANDN U7001 ( .A(n6758), .B(n7515), .Z(n6762) );
  OR U7002 ( .A(n6760), .B(n6759), .Z(n6761) );
  NAND U7003 ( .A(n6762), .B(n6761), .Z(n6848) );
  XNOR U7004 ( .A(n6849), .B(n6848), .Z(n6851) );
  XOR U7005 ( .A(n6850), .B(n6851), .Z(n6845) );
  XOR U7006 ( .A(n6844), .B(n6845), .Z(n6837) );
  OR U7007 ( .A(n6764), .B(n6763), .Z(n6768) );
  OR U7008 ( .A(n6766), .B(n6765), .Z(n6767) );
  AND U7009 ( .A(n6768), .B(n6767), .Z(n6836) );
  XOR U7010 ( .A(n6837), .B(n6836), .Z(n6838) );
  OR U7011 ( .A(n6770), .B(n6769), .Z(n6774) );
  OR U7012 ( .A(n6772), .B(n6771), .Z(n6773) );
  NAND U7013 ( .A(n6774), .B(n6773), .Z(n6831) );
  NANDN U7014 ( .A(n48), .B(y[269]), .Z(n6810) );
  ANDN U7015 ( .B(y[270]), .A(n47), .Z(n6776) );
  XNOR U7016 ( .A(n6776), .B(n6775), .Z(n6809) );
  XOR U7017 ( .A(n6810), .B(n6809), .Z(n6819) );
  ANDN U7018 ( .B(y[260]), .A(n57), .Z(n7519) );
  ANDN U7019 ( .B(x[77]), .A(n8881), .Z(n6778) );
  NANDN U7020 ( .A(n50), .B(y[267]), .Z(n6777) );
  XOR U7021 ( .A(n6778), .B(n6777), .Z(n6880) );
  XNOR U7022 ( .A(n7519), .B(n6880), .Z(n6818) );
  XNOR U7023 ( .A(n6819), .B(n6818), .Z(n6821) );
  NANDN U7024 ( .A(n6779), .B(n7519), .Z(n6783) );
  OR U7025 ( .A(n6781), .B(n6780), .Z(n6782) );
  AND U7026 ( .A(n6783), .B(n6782), .Z(n6820) );
  XNOR U7027 ( .A(n6821), .B(n6820), .Z(n6830) );
  XNOR U7028 ( .A(n6831), .B(n6830), .Z(n6833) );
  OR U7029 ( .A(n6785), .B(n6784), .Z(n6789) );
  OR U7030 ( .A(n6787), .B(n6786), .Z(n6788) );
  NAND U7031 ( .A(n6789), .B(n6788), .Z(n6832) );
  XOR U7032 ( .A(n6833), .B(n6832), .Z(n6839) );
  XNOR U7033 ( .A(n6838), .B(n6839), .Z(n6802) );
  NANDN U7034 ( .A(n6791), .B(n6790), .Z(n6795) );
  NANDN U7035 ( .A(n6793), .B(n6792), .Z(n6794) );
  NAND U7036 ( .A(n6795), .B(n6794), .Z(n6803) );
  XOR U7037 ( .A(n6802), .B(n6803), .Z(n6804) );
  XNOR U7038 ( .A(n6805), .B(n6804), .Z(n6799) );
  XOR U7039 ( .A(n6798), .B(n6799), .Z(N177) );
  NANDN U7040 ( .A(n6797), .B(n6796), .Z(n6801) );
  NANDN U7041 ( .A(n6799), .B(n6798), .Z(n6800) );
  NAND U7042 ( .A(n6801), .B(n6800), .Z(n6889) );
  OR U7043 ( .A(n6803), .B(n6802), .Z(n6807) );
  NANDN U7044 ( .A(n6805), .B(n6804), .Z(n6806) );
  NAND U7045 ( .A(n6807), .B(n6806), .Z(n6890) );
  XNOR U7046 ( .A(n6889), .B(n6890), .Z(n6891) );
  ANDN U7047 ( .B(y[266]), .A(n52), .Z(n7067) );
  AND U7048 ( .A(y[265]), .B(x[72]), .Z(n6977) );
  XNOR U7049 ( .A(n6976), .B(n6977), .Z(n6979) );
  AND U7050 ( .A(y[268]), .B(x[69]), .Z(n6978) );
  XOR U7051 ( .A(n6979), .B(n6978), .Z(n6964) );
  AND U7052 ( .A(y[269]), .B(x[68]), .Z(n6933) );
  AND U7053 ( .A(y[262]), .B(x[75]), .Z(n6931) );
  AND U7054 ( .A(y[260]), .B(x[77]), .Z(n6932) );
  XNOR U7055 ( .A(n6931), .B(n6932), .Z(n6934) );
  XOR U7056 ( .A(n6933), .B(n6934), .Z(n6965) );
  XOR U7057 ( .A(n6964), .B(n6965), .Z(n6966) );
  XNOR U7058 ( .A(n7067), .B(n6966), .Z(n6960) );
  ANDN U7059 ( .B(y[270]), .A(n54), .Z(n6808) );
  NAND U7060 ( .A(n6808), .B(n6969), .Z(n6812) );
  OR U7061 ( .A(n6810), .B(n6809), .Z(n6811) );
  NAND U7062 ( .A(n6812), .B(n6811), .Z(n6959) );
  NANDN U7063 ( .A(n56), .B(y[258]), .Z(n7029) );
  ANDN U7064 ( .B(y[261]), .A(n59), .Z(n6813) );
  NANDN U7065 ( .A(n7029), .B(n6813), .Z(n6817) );
  OR U7066 ( .A(n6815), .B(n6814), .Z(n6816) );
  NAND U7067 ( .A(n6817), .B(n6816), .Z(n6958) );
  XOR U7068 ( .A(n6959), .B(n6958), .Z(n6961) );
  XNOR U7069 ( .A(n6960), .B(n6961), .Z(n6908) );
  NAND U7070 ( .A(n6819), .B(n6818), .Z(n6823) );
  OR U7071 ( .A(n6821), .B(n6820), .Z(n6822) );
  NAND U7072 ( .A(n6823), .B(n6822), .Z(n6907) );
  XOR U7073 ( .A(n6908), .B(n6907), .Z(n6909) );
  OR U7074 ( .A(n6825), .B(n6824), .Z(n6829) );
  NAND U7075 ( .A(n6827), .B(n6826), .Z(n6828) );
  NAND U7076 ( .A(n6829), .B(n6828), .Z(n6910) );
  XNOR U7077 ( .A(n6909), .B(n6910), .Z(n6986) );
  OR U7078 ( .A(n6831), .B(n6830), .Z(n6835) );
  OR U7079 ( .A(n6833), .B(n6832), .Z(n6834) );
  AND U7080 ( .A(n6835), .B(n6834), .Z(n6987) );
  XNOR U7081 ( .A(n6986), .B(n6987), .Z(n6989) );
  OR U7082 ( .A(n6837), .B(n6836), .Z(n6841) );
  NANDN U7083 ( .A(n6839), .B(n6838), .Z(n6840) );
  NAND U7084 ( .A(n6841), .B(n6840), .Z(n6988) );
  XOR U7085 ( .A(n6989), .B(n6988), .Z(n6895) );
  OR U7086 ( .A(n6843), .B(n6842), .Z(n6847) );
  NANDN U7087 ( .A(n6845), .B(n6844), .Z(n6846) );
  NAND U7088 ( .A(n6847), .B(n6846), .Z(n6995) );
  OR U7089 ( .A(n6849), .B(n6848), .Z(n6853) );
  NANDN U7090 ( .A(n6851), .B(n6850), .Z(n6852) );
  NAND U7091 ( .A(n6853), .B(n6852), .Z(n6993) );
  OR U7092 ( .A(n6855), .B(n6854), .Z(n6859) );
  OR U7093 ( .A(n6857), .B(n6856), .Z(n6858) );
  NAND U7094 ( .A(n6859), .B(n6858), .Z(n6904) );
  NANDN U7095 ( .A(n53), .B(y[271]), .Z(n7514) );
  AND U7096 ( .A(y[264]), .B(x[65]), .Z(n7054) );
  NANDN U7097 ( .A(n7514), .B(n7054), .Z(n6863) );
  OR U7098 ( .A(n6861), .B(n6860), .Z(n6862) );
  AND U7099 ( .A(n6863), .B(n6862), .Z(n6925) );
  NAND U7100 ( .A(n7067), .B(n6864), .Z(n6868) );
  OR U7101 ( .A(n6866), .B(n6865), .Z(n6867) );
  AND U7102 ( .A(n6868), .B(n6867), .Z(n6926) );
  XNOR U7103 ( .A(n6925), .B(n6926), .Z(n6928) );
  NANDN U7104 ( .A(n45), .B(y[273]), .Z(n6945) );
  ANDN U7105 ( .B(y[257]), .A(n8890), .Z(n6937) );
  XNOR U7106 ( .A(o[81]), .B(n6937), .Z(n6943) );
  NANDN U7107 ( .A(n8626), .B(y[256]), .Z(n6942) );
  XOR U7108 ( .A(n6943), .B(n6942), .Z(n6944) );
  XOR U7109 ( .A(n6945), .B(n6944), .Z(n6922) );
  NANDN U7110 ( .A(n48), .B(y[270]), .Z(n6971) );
  ANDN U7111 ( .B(y[271]), .A(n47), .Z(n6869) );
  ANDN U7112 ( .B(y[263]), .A(n55), .Z(n7543) );
  XNOR U7113 ( .A(n6869), .B(n7543), .Z(n6970) );
  XNOR U7114 ( .A(n6971), .B(n6970), .Z(n6919) );
  NANDN U7115 ( .A(n6871), .B(n6870), .Z(n6875) );
  NAND U7116 ( .A(n6873), .B(n6872), .Z(n6874) );
  AND U7117 ( .A(n6875), .B(n6874), .Z(n6920) );
  XOR U7118 ( .A(n6922), .B(n6921), .Z(n6927) );
  NANDN U7119 ( .A(n6876), .B(o[80]), .Z(n6983) );
  ANDN U7120 ( .B(y[272]), .A(n46), .Z(n6878) );
  ANDN U7121 ( .B(x[73]), .A(n8927), .Z(n6877) );
  XNOR U7122 ( .A(n6878), .B(n6877), .Z(n6982) );
  XOR U7123 ( .A(n6983), .B(n6982), .Z(n6913) );
  AND U7124 ( .A(y[261]), .B(x[76]), .Z(n6954) );
  AND U7125 ( .A(y[259]), .B(x[78]), .Z(n6952) );
  AND U7126 ( .A(y[258]), .B(x[79]), .Z(n6953) );
  XNOR U7127 ( .A(n6952), .B(n6953), .Z(n6955) );
  XOR U7128 ( .A(n6954), .B(n6955), .Z(n6914) );
  XOR U7129 ( .A(n6913), .B(n6914), .Z(n6916) );
  AND U7130 ( .A(y[267]), .B(x[77]), .Z(n7695) );
  IV U7131 ( .A(n7695), .Z(n7797) );
  ANDN U7132 ( .B(y[259]), .A(n50), .Z(n6879) );
  NANDN U7133 ( .A(n7797), .B(n6879), .Z(n6882) );
  NANDN U7134 ( .A(n6880), .B(n7519), .Z(n6881) );
  AND U7135 ( .A(n6882), .B(n6881), .Z(n6915) );
  XNOR U7136 ( .A(n6916), .B(n6915), .Z(n6902) );
  XOR U7137 ( .A(n6901), .B(n6902), .Z(n6903) );
  XNOR U7138 ( .A(n6904), .B(n6903), .Z(n6992) );
  XNOR U7139 ( .A(n6993), .B(n6992), .Z(n6994) );
  XOR U7140 ( .A(n6995), .B(n6994), .Z(n6896) );
  XNOR U7141 ( .A(n6895), .B(n6896), .Z(n6898) );
  OR U7142 ( .A(n6884), .B(n6883), .Z(n6888) );
  NANDN U7143 ( .A(n6886), .B(n6885), .Z(n6887) );
  AND U7144 ( .A(n6888), .B(n6887), .Z(n6897) );
  XOR U7145 ( .A(n6898), .B(n6897), .Z(n6892) );
  XNOR U7146 ( .A(n6891), .B(n6892), .Z(N178) );
  NANDN U7147 ( .A(n6890), .B(n6889), .Z(n6894) );
  NAND U7148 ( .A(n6892), .B(n6891), .Z(n6893) );
  NAND U7149 ( .A(n6894), .B(n6893), .Z(n6998) );
  OR U7150 ( .A(n6896), .B(n6895), .Z(n6900) );
  OR U7151 ( .A(n6898), .B(n6897), .Z(n6899) );
  AND U7152 ( .A(n6900), .B(n6899), .Z(n6999) );
  XNOR U7153 ( .A(n6998), .B(n6999), .Z(n7000) );
  NAND U7154 ( .A(n6902), .B(n6901), .Z(n6906) );
  NANDN U7155 ( .A(n6904), .B(n6903), .Z(n6905) );
  AND U7156 ( .A(n6906), .B(n6905), .Z(n7106) );
  OR U7157 ( .A(n6908), .B(n6907), .Z(n6912) );
  NANDN U7158 ( .A(n6910), .B(n6909), .Z(n6911) );
  AND U7159 ( .A(n6912), .B(n6911), .Z(n7107) );
  XOR U7160 ( .A(n7106), .B(n7107), .Z(n7109) );
  NANDN U7161 ( .A(n6914), .B(n6913), .Z(n6918) );
  OR U7162 ( .A(n6916), .B(n6915), .Z(n6917) );
  AND U7163 ( .A(n6918), .B(n6917), .Z(n7082) );
  OR U7164 ( .A(n6920), .B(n6919), .Z(n6924) );
  OR U7165 ( .A(n6922), .B(n6921), .Z(n6923) );
  AND U7166 ( .A(n6924), .B(n6923), .Z(n7083) );
  XNOR U7167 ( .A(n7082), .B(n7083), .Z(n7084) );
  OR U7168 ( .A(n6926), .B(n6925), .Z(n6930) );
  NANDN U7169 ( .A(n6928), .B(n6927), .Z(n6929) );
  AND U7170 ( .A(n6930), .B(n6929), .Z(n7085) );
  OR U7171 ( .A(n6932), .B(n6931), .Z(n6936) );
  OR U7172 ( .A(n6934), .B(n6933), .Z(n6935) );
  NAND U7173 ( .A(n6936), .B(n6935), .Z(n7037) );
  NAND U7174 ( .A(o[81]), .B(n6937), .Z(n7056) );
  ANDN U7175 ( .B(y[273]), .A(n46), .Z(n6939) );
  ANDN U7176 ( .B(x[74]), .A(n8927), .Z(n6938) );
  XNOR U7177 ( .A(n6939), .B(n6938), .Z(n7055) );
  XOR U7178 ( .A(n7056), .B(n7055), .Z(n7034) );
  NANDN U7179 ( .A(n60), .B(y[259]), .Z(n7023) );
  ANDN U7180 ( .B(y[260]), .A(n59), .Z(n6941) );
  ANDN U7181 ( .B(x[73]), .A(n8627), .Z(n6940) );
  XNOR U7182 ( .A(n6941), .B(n6940), .Z(n7022) );
  XNOR U7183 ( .A(n7023), .B(n7022), .Z(n7035) );
  XOR U7184 ( .A(n7034), .B(n7035), .Z(n7036) );
  XNOR U7185 ( .A(n7037), .B(n7036), .Z(n7101) );
  OR U7186 ( .A(n6943), .B(n6942), .Z(n6947) );
  NANDN U7187 ( .A(n6945), .B(n6944), .Z(n6946) );
  NAND U7188 ( .A(n6947), .B(n6946), .Z(n7089) );
  NANDN U7189 ( .A(n49), .B(y[270]), .Z(n7070) );
  ANDN U7190 ( .B(y[267]), .A(n52), .Z(n6949) );
  ANDN U7191 ( .B(x[72]), .A(n7862), .Z(n6948) );
  XNOR U7192 ( .A(n6949), .B(n6948), .Z(n7069) );
  XNOR U7193 ( .A(n7070), .B(n7069), .Z(n7018) );
  AND U7194 ( .A(y[268]), .B(x[70]), .Z(n7016) );
  ANDN U7195 ( .B(x[69]), .A(n8815), .Z(n7138) );
  XOR U7196 ( .A(n7016), .B(n7138), .Z(n7017) );
  XOR U7197 ( .A(n7018), .B(n7017), .Z(n7088) );
  XOR U7198 ( .A(n7089), .B(n7088), .Z(n7091) );
  NANDN U7199 ( .A(n47), .B(y[272]), .Z(n7031) );
  ANDN U7200 ( .B(y[263]), .A(n56), .Z(n6951) );
  ANDN U7201 ( .B(y[258]), .A(n8890), .Z(n6950) );
  XNOR U7202 ( .A(n6951), .B(n6950), .Z(n7030) );
  XOR U7203 ( .A(n7031), .B(n7030), .Z(n7090) );
  XNOR U7204 ( .A(n7091), .B(n7090), .Z(n7100) );
  XOR U7205 ( .A(n7101), .B(n7100), .Z(n7103) );
  OR U7206 ( .A(n6953), .B(n6952), .Z(n6957) );
  OR U7207 ( .A(n6955), .B(n6954), .Z(n6956) );
  NAND U7208 ( .A(n6957), .B(n6956), .Z(n7102) );
  XOR U7209 ( .A(n7103), .B(n7102), .Z(n7011) );
  OR U7210 ( .A(n6959), .B(n6958), .Z(n6963) );
  NAND U7211 ( .A(n6961), .B(n6960), .Z(n6962) );
  NAND U7212 ( .A(n6963), .B(n6962), .Z(n7079) );
  OR U7213 ( .A(n6965), .B(n6964), .Z(n6968) );
  NAND U7214 ( .A(n6966), .B(n7067), .Z(n6967) );
  AND U7215 ( .A(n6968), .B(n6967), .Z(n7076) );
  ANDN U7216 ( .B(y[271]), .A(n55), .Z(n7935) );
  NAND U7217 ( .A(n6969), .B(n7935), .Z(n6973) );
  OR U7218 ( .A(n6971), .B(n6970), .Z(n6972) );
  AND U7219 ( .A(n6973), .B(n6972), .Z(n7042) );
  ANDN U7220 ( .B(y[257]), .A(n8626), .Z(n7073) );
  XNOR U7221 ( .A(o[82]), .B(n7073), .Z(n7051) );
  NANDN U7222 ( .A(n45), .B(y[274]), .Z(n7049) );
  NANDN U7223 ( .A(n61), .B(y[256]), .Z(n7048) );
  XNOR U7224 ( .A(n7049), .B(n7048), .Z(n7050) );
  XNOR U7225 ( .A(n7051), .B(n7050), .Z(n7041) );
  ANDN U7226 ( .B(y[262]), .A(n57), .Z(n7178) );
  ANDN U7227 ( .B(y[271]), .A(n48), .Z(n6975) );
  NANDN U7228 ( .A(n58), .B(y[261]), .Z(n6974) );
  XOR U7229 ( .A(n6975), .B(n6974), .Z(n7062) );
  XNOR U7230 ( .A(n7178), .B(n7062), .Z(n7040) );
  XOR U7231 ( .A(n7041), .B(n7040), .Z(n7043) );
  XOR U7232 ( .A(n7042), .B(n7043), .Z(n7094) );
  OR U7233 ( .A(n6977), .B(n6976), .Z(n6981) );
  OR U7234 ( .A(n6979), .B(n6978), .Z(n6980) );
  AND U7235 ( .A(n6981), .B(n6980), .Z(n7095) );
  XNOR U7236 ( .A(n7094), .B(n7095), .Z(n7097) );
  ANDN U7237 ( .B(x[73]), .A(n8884), .Z(n7803) );
  IV U7238 ( .A(n7803), .Z(n7934) );
  NANDN U7239 ( .A(n7934), .B(n7054), .Z(n6985) );
  OR U7240 ( .A(n6983), .B(n6982), .Z(n6984) );
  NAND U7241 ( .A(n6985), .B(n6984), .Z(n7096) );
  XOR U7242 ( .A(n7097), .B(n7096), .Z(n7077) );
  XNOR U7243 ( .A(n7076), .B(n7077), .Z(n7078) );
  XNOR U7244 ( .A(n7079), .B(n7078), .Z(n7010) );
  XOR U7245 ( .A(n7011), .B(n7010), .Z(n7013) );
  XNOR U7246 ( .A(n7109), .B(n7108), .Z(n7007) );
  OR U7247 ( .A(n6987), .B(n6986), .Z(n6991) );
  OR U7248 ( .A(n6989), .B(n6988), .Z(n6990) );
  NAND U7249 ( .A(n6991), .B(n6990), .Z(n7005) );
  OR U7250 ( .A(n6993), .B(n6992), .Z(n6997) );
  OR U7251 ( .A(n6995), .B(n6994), .Z(n6996) );
  NAND U7252 ( .A(n6997), .B(n6996), .Z(n7004) );
  XNOR U7253 ( .A(n7005), .B(n7004), .Z(n7006) );
  XNOR U7254 ( .A(n7007), .B(n7006), .Z(n7001) );
  XOR U7255 ( .A(n7000), .B(n7001), .Z(N179) );
  NANDN U7256 ( .A(n6999), .B(n6998), .Z(n7003) );
  NANDN U7257 ( .A(n7001), .B(n7000), .Z(n7002) );
  NAND U7258 ( .A(n7003), .B(n7002), .Z(n7222) );
  OR U7259 ( .A(n7005), .B(n7004), .Z(n7009) );
  OR U7260 ( .A(n7007), .B(n7006), .Z(n7008) );
  AND U7261 ( .A(n7009), .B(n7008), .Z(n7223) );
  XNOR U7262 ( .A(n7222), .B(n7223), .Z(n7224) );
  NANDN U7263 ( .A(n7011), .B(n7010), .Z(n7015) );
  NANDN U7264 ( .A(n7013), .B(n7012), .Z(n7014) );
  AND U7265 ( .A(n7015), .B(n7014), .Z(n7228) );
  OR U7266 ( .A(n7016), .B(n7138), .Z(n7020) );
  NAND U7267 ( .A(n7018), .B(n7017), .Z(n7019) );
  AND U7268 ( .A(n7020), .B(n7019), .Z(n7218) );
  NANDN U7269 ( .A(n8627), .B(x[78]), .Z(n7721) );
  OR U7270 ( .A(n7021), .B(n7721), .Z(n7025) );
  OR U7271 ( .A(n7023), .B(n7022), .Z(n7024) );
  AND U7272 ( .A(n7025), .B(n7024), .Z(n7199) );
  NANDN U7273 ( .A(n47), .B(y[273]), .Z(n7181) );
  ANDN U7274 ( .B(x[77]), .A(n8655), .Z(n7026) );
  XNOR U7275 ( .A(n7027), .B(n7026), .Z(n7180) );
  XNOR U7276 ( .A(n7181), .B(n7180), .Z(n7198) );
  NANDN U7277 ( .A(n46), .B(y[274]), .Z(n7155) );
  ANDN U7278 ( .B(x[78]), .A(n7989), .Z(n7028) );
  XOR U7279 ( .A(n7028), .B(n7068), .Z(n7154) );
  XNOR U7280 ( .A(n7155), .B(n7154), .Z(n7200) );
  XOR U7281 ( .A(n7201), .B(n7200), .Z(n7216) );
  ANDN U7282 ( .B(y[263]), .A(n8890), .Z(n7512) );
  NANDN U7283 ( .A(n7029), .B(n7512), .Z(n7033) );
  OR U7284 ( .A(n7031), .B(n7030), .Z(n7032) );
  NAND U7285 ( .A(n7033), .B(n7032), .Z(n7217) );
  XNOR U7286 ( .A(n7216), .B(n7217), .Z(n7219) );
  XOR U7287 ( .A(n7218), .B(n7219), .Z(n7124) );
  NANDN U7288 ( .A(n7035), .B(n7034), .Z(n7039) );
  OR U7289 ( .A(n7037), .B(n7036), .Z(n7038) );
  NAND U7290 ( .A(n7039), .B(n7038), .Z(n7211) );
  NANDN U7291 ( .A(n7041), .B(n7040), .Z(n7045) );
  OR U7292 ( .A(n7043), .B(n7042), .Z(n7044) );
  NAND U7293 ( .A(n7045), .B(n7044), .Z(n7210) );
  XOR U7294 ( .A(n7211), .B(n7210), .Z(n7212) );
  ANDN U7295 ( .B(x[80]), .A(n8881), .Z(n7047) );
  NANDN U7296 ( .A(n54), .B(y[266]), .Z(n7046) );
  XOR U7297 ( .A(n7047), .B(n7046), .Z(n7171) );
  ANDN U7298 ( .B(y[260]), .A(n60), .Z(n7170) );
  XOR U7299 ( .A(n7171), .B(n7170), .Z(n7130) );
  OR U7300 ( .A(n7049), .B(n7048), .Z(n7053) );
  OR U7301 ( .A(n7051), .B(n7050), .Z(n7052) );
  AND U7302 ( .A(n7053), .B(n7052), .Z(n7131) );
  IV U7303 ( .A(y[273]), .Z(n8904) );
  ANDN U7304 ( .B(x[74]), .A(n8904), .Z(n8306) );
  NAND U7305 ( .A(n7054), .B(n8306), .Z(n7058) );
  OR U7306 ( .A(n7056), .B(n7055), .Z(n7057) );
  AND U7307 ( .A(n7058), .B(n7057), .Z(n7132) );
  XOR U7308 ( .A(n7133), .B(n7132), .Z(n7206) );
  ANDN U7309 ( .B(y[257]), .A(n61), .Z(n7191) );
  XNOR U7310 ( .A(o[83]), .B(n7191), .Z(n7160) );
  ANDN U7311 ( .B(x[74]), .A(n8627), .Z(n7060) );
  ANDN U7312 ( .B(y[258]), .A(n8626), .Z(n7059) );
  XNOR U7313 ( .A(n7060), .B(n7059), .Z(n7159) );
  XNOR U7314 ( .A(n7160), .B(n7159), .Z(n7166) );
  AND U7315 ( .A(y[271]), .B(x[77]), .Z(n8430) );
  NANDN U7316 ( .A(n7061), .B(n8430), .Z(n7064) );
  NANDN U7317 ( .A(n7062), .B(n7178), .Z(n7063) );
  AND U7318 ( .A(n7064), .B(n7063), .Z(n7163) );
  NANDN U7319 ( .A(n48), .B(y[272]), .Z(n7186) );
  ANDN U7320 ( .B(x[75]), .A(n8927), .Z(n7066) );
  NANDN U7321 ( .A(n52), .B(y[268]), .Z(n7065) );
  XOR U7322 ( .A(n7066), .B(n7065), .Z(n7185) );
  XNOR U7323 ( .A(n7186), .B(n7185), .Z(n7164) );
  XNOR U7324 ( .A(n7163), .B(n7164), .Z(n7165) );
  XOR U7325 ( .A(n7166), .B(n7165), .Z(n7205) );
  NANDN U7326 ( .A(n7068), .B(n7067), .Z(n7072) );
  OR U7327 ( .A(n7070), .B(n7069), .Z(n7071) );
  AND U7328 ( .A(n7072), .B(n7071), .Z(n7195) );
  NAND U7329 ( .A(n7073), .B(o[82]), .Z(n7145) );
  NANDN U7330 ( .A(n8824), .B(y[256]), .Z(n7143) );
  NANDN U7331 ( .A(n45), .B(y[275]), .Z(n7142) );
  XNOR U7332 ( .A(n7143), .B(n7142), .Z(n7144) );
  XNOR U7333 ( .A(n7145), .B(n7144), .Z(n7193) );
  ANDN U7334 ( .B(y[271]), .A(n49), .Z(n7280) );
  ANDN U7335 ( .B(y[269]), .A(n51), .Z(n7075) );
  ANDN U7336 ( .B(x[69]), .A(n8861), .Z(n7074) );
  XNOR U7337 ( .A(n7075), .B(n7074), .Z(n7139) );
  XOR U7338 ( .A(n7280), .B(n7139), .Z(n7192) );
  XOR U7339 ( .A(n7193), .B(n7192), .Z(n7194) );
  XOR U7340 ( .A(n7195), .B(n7194), .Z(n7204) );
  XOR U7341 ( .A(n7205), .B(n7204), .Z(n7207) );
  XNOR U7342 ( .A(n7206), .B(n7207), .Z(n7213) );
  XNOR U7343 ( .A(n7212), .B(n7213), .Z(n7125) );
  XNOR U7344 ( .A(n7124), .B(n7125), .Z(n7127) );
  OR U7345 ( .A(n7077), .B(n7076), .Z(n7081) );
  OR U7346 ( .A(n7079), .B(n7078), .Z(n7080) );
  AND U7347 ( .A(n7081), .B(n7080), .Z(n7126) );
  XOR U7348 ( .A(n7127), .B(n7126), .Z(n7121) );
  OR U7349 ( .A(n7083), .B(n7082), .Z(n7087) );
  OR U7350 ( .A(n7085), .B(n7084), .Z(n7086) );
  NAND U7351 ( .A(n7087), .B(n7086), .Z(n7119) );
  NANDN U7352 ( .A(n7089), .B(n7088), .Z(n7093) );
  OR U7353 ( .A(n7091), .B(n7090), .Z(n7092) );
  AND U7354 ( .A(n7093), .B(n7092), .Z(n7114) );
  OR U7355 ( .A(n7095), .B(n7094), .Z(n7099) );
  OR U7356 ( .A(n7097), .B(n7096), .Z(n7098) );
  AND U7357 ( .A(n7099), .B(n7098), .Z(n7112) );
  NANDN U7358 ( .A(n7101), .B(n7100), .Z(n7105) );
  OR U7359 ( .A(n7103), .B(n7102), .Z(n7104) );
  NAND U7360 ( .A(n7105), .B(n7104), .Z(n7113) );
  XNOR U7361 ( .A(n7112), .B(n7113), .Z(n7115) );
  XNOR U7362 ( .A(n7114), .B(n7115), .Z(n7118) );
  XOR U7363 ( .A(n7119), .B(n7118), .Z(n7120) );
  XOR U7364 ( .A(n7121), .B(n7120), .Z(n7229) );
  XNOR U7365 ( .A(n7228), .B(n7229), .Z(n7230) );
  OR U7366 ( .A(n7107), .B(n7106), .Z(n7111) );
  NAND U7367 ( .A(n7109), .B(n7108), .Z(n7110) );
  AND U7368 ( .A(n7111), .B(n7110), .Z(n7231) );
  XOR U7369 ( .A(n7224), .B(n7225), .Z(N180) );
  OR U7370 ( .A(n7113), .B(n7112), .Z(n7117) );
  OR U7371 ( .A(n7115), .B(n7114), .Z(n7116) );
  AND U7372 ( .A(n7117), .B(n7116), .Z(n7348) );
  OR U7373 ( .A(n7119), .B(n7118), .Z(n7123) );
  NANDN U7374 ( .A(n7121), .B(n7120), .Z(n7122) );
  AND U7375 ( .A(n7123), .B(n7122), .Z(n7346) );
  OR U7376 ( .A(n7125), .B(n7124), .Z(n7129) );
  OR U7377 ( .A(n7127), .B(n7126), .Z(n7128) );
  AND U7378 ( .A(n7129), .B(n7128), .Z(n7337) );
  OR U7379 ( .A(n7131), .B(n7130), .Z(n7135) );
  OR U7380 ( .A(n7133), .B(n7132), .Z(n7134) );
  NAND U7381 ( .A(n7135), .B(n7134), .Z(n7237) );
  NANDN U7382 ( .A(n8626), .B(y[259]), .Z(n7254) );
  ANDN U7383 ( .B(x[76]), .A(n8927), .Z(n7137) );
  ANDN U7384 ( .B(y[258]), .A(n61), .Z(n7136) );
  XNOR U7385 ( .A(n7137), .B(n7136), .Z(n7253) );
  XNOR U7386 ( .A(n7254), .B(n7253), .Z(n7262) );
  NOR U7387 ( .A(n8861), .B(n51), .Z(n7150) );
  IV U7388 ( .A(n7150), .Z(n7240) );
  NANDN U7389 ( .A(n7240), .B(n7138), .Z(n7141) );
  NANDN U7390 ( .A(n7139), .B(n7280), .Z(n7140) );
  AND U7391 ( .A(n7141), .B(n7140), .Z(n7263) );
  OR U7392 ( .A(n7143), .B(n7142), .Z(n7147) );
  OR U7393 ( .A(n7145), .B(n7144), .Z(n7146) );
  AND U7394 ( .A(n7147), .B(n7146), .Z(n7264) );
  XNOR U7395 ( .A(n7265), .B(n7264), .Z(n7234) );
  NANDN U7396 ( .A(n52), .B(y[269]), .Z(n7282) );
  ANDN U7397 ( .B(y[271]), .A(n50), .Z(n7149) );
  NANDN U7398 ( .A(n49), .B(y[272]), .Z(n7148) );
  XOR U7399 ( .A(n7149), .B(n7148), .Z(n7281) );
  XNOR U7400 ( .A(n7282), .B(n7281), .Z(n7241) );
  XOR U7401 ( .A(n7150), .B(n7241), .Z(n7243) );
  NANDN U7402 ( .A(n53), .B(y[268]), .Z(n7290) );
  ANDN U7403 ( .B(x[67]), .A(n8904), .Z(n7152) );
  NANDN U7404 ( .A(n58), .B(y[263]), .Z(n7151) );
  XOR U7405 ( .A(n7152), .B(n7151), .Z(n7289) );
  XNOR U7406 ( .A(n7290), .B(n7289), .Z(n7242) );
  XNOR U7407 ( .A(n7243), .B(n7242), .Z(n7300) );
  AND U7408 ( .A(y[267]), .B(x[78]), .Z(n7811) );
  IV U7409 ( .A(n7811), .Z(n7995) );
  NANDN U7410 ( .A(n7995), .B(n7153), .Z(n7157) );
  OR U7411 ( .A(n7155), .B(n7154), .Z(n7156) );
  NAND U7412 ( .A(n7157), .B(n7156), .Z(n7299) );
  ANDN U7413 ( .B(x[81]), .A(n8627), .Z(n8103) );
  NANDN U7414 ( .A(n7158), .B(n8103), .Z(n7162) );
  OR U7415 ( .A(n7160), .B(n7159), .Z(n7161) );
  NAND U7416 ( .A(n7162), .B(n7161), .Z(n7298) );
  XNOR U7417 ( .A(n7299), .B(n7298), .Z(n7301) );
  XOR U7418 ( .A(n7300), .B(n7301), .Z(n7235) );
  XOR U7419 ( .A(n7237), .B(n7236), .Z(n7323) );
  OR U7420 ( .A(n7164), .B(n7163), .Z(n7168) );
  OR U7421 ( .A(n7166), .B(n7165), .Z(n7167) );
  NAND U7422 ( .A(n7168), .B(n7167), .Z(n7322) );
  XOR U7423 ( .A(n7323), .B(n7322), .Z(n7325) );
  ANDN U7424 ( .B(y[259]), .A(n54), .Z(n7169) );
  ANDN U7425 ( .B(x[80]), .A(n7862), .Z(n8090) );
  NAND U7426 ( .A(n7169), .B(n8090), .Z(n7173) );
  NANDN U7427 ( .A(n7171), .B(n7170), .Z(n7172) );
  AND U7428 ( .A(n7173), .B(n7172), .Z(n7317) );
  ANDN U7429 ( .B(x[79]), .A(n7989), .Z(n7175) );
  NANDN U7430 ( .A(n54), .B(y[267]), .Z(n7174) );
  XOR U7431 ( .A(n7175), .B(n7174), .Z(n7248) );
  ANDN U7432 ( .B(x[78]), .A(n8655), .Z(n7247) );
  XNOR U7433 ( .A(n7248), .B(n7247), .Z(n7304) );
  NANDN U7434 ( .A(n47), .B(y[274]), .Z(n7295) );
  ANDN U7435 ( .B(y[260]), .A(n8890), .Z(n7177) );
  NANDN U7436 ( .A(n55), .B(y[266]), .Z(n7176) );
  XOR U7437 ( .A(n7177), .B(n7176), .Z(n7294) );
  XNOR U7438 ( .A(n7295), .B(n7294), .Z(n7305) );
  XOR U7439 ( .A(n7304), .B(n7305), .Z(n7307) );
  ANDN U7440 ( .B(y[263]), .A(n58), .Z(n7179) );
  NAND U7441 ( .A(n7179), .B(n7178), .Z(n7183) );
  OR U7442 ( .A(n7181), .B(n7180), .Z(n7182) );
  AND U7443 ( .A(n7183), .B(n7182), .Z(n7306) );
  XNOR U7444 ( .A(n7307), .B(n7306), .Z(n7316) );
  AND U7445 ( .A(y[268]), .B(x[75]), .Z(n7685) );
  NAND U7446 ( .A(n7184), .B(n7685), .Z(n7188) );
  OR U7447 ( .A(n7186), .B(n7185), .Z(n7187) );
  AND U7448 ( .A(n7188), .B(n7187), .Z(n7313) );
  ANDN U7449 ( .B(y[257]), .A(n8824), .Z(n7251) );
  XNOR U7450 ( .A(o[84]), .B(n7251), .Z(n7259) );
  ANDN U7451 ( .B(x[75]), .A(n8627), .Z(n7190) );
  ANDN U7452 ( .B(y[275]), .A(n46), .Z(n7189) );
  XNOR U7453 ( .A(n7190), .B(n7189), .Z(n7258) );
  XNOR U7454 ( .A(n7259), .B(n7258), .Z(n7311) );
  NAND U7455 ( .A(o[83]), .B(n7191), .Z(n7277) );
  NANDN U7456 ( .A(n8885), .B(y[256]), .Z(n7275) );
  NANDN U7457 ( .A(n45), .B(y[276]), .Z(n7274) );
  XNOR U7458 ( .A(n7275), .B(n7274), .Z(n7276) );
  XNOR U7459 ( .A(n7277), .B(n7276), .Z(n7310) );
  XOR U7460 ( .A(n7311), .B(n7310), .Z(n7312) );
  XOR U7461 ( .A(n7313), .B(n7312), .Z(n7318) );
  XNOR U7462 ( .A(n7319), .B(n7318), .Z(n7270) );
  OR U7463 ( .A(n7193), .B(n7192), .Z(n7197) );
  NANDN U7464 ( .A(n7195), .B(n7194), .Z(n7196) );
  NAND U7465 ( .A(n7197), .B(n7196), .Z(n7269) );
  OR U7466 ( .A(n7199), .B(n7198), .Z(n7203) );
  OR U7467 ( .A(n7201), .B(n7200), .Z(n7202) );
  NAND U7468 ( .A(n7203), .B(n7202), .Z(n7268) );
  XNOR U7469 ( .A(n7269), .B(n7268), .Z(n7271) );
  XNOR U7470 ( .A(n7270), .B(n7271), .Z(n7324) );
  XNOR U7471 ( .A(n7325), .B(n7324), .Z(n7334) );
  NANDN U7472 ( .A(n7205), .B(n7204), .Z(n7209) );
  OR U7473 ( .A(n7207), .B(n7206), .Z(n7208) );
  NAND U7474 ( .A(n7209), .B(n7208), .Z(n7329) );
  OR U7475 ( .A(n7211), .B(n7210), .Z(n7215) );
  NANDN U7476 ( .A(n7213), .B(n7212), .Z(n7214) );
  NAND U7477 ( .A(n7215), .B(n7214), .Z(n7328) );
  XNOR U7478 ( .A(n7329), .B(n7328), .Z(n7330) );
  OR U7479 ( .A(n7217), .B(n7216), .Z(n7221) );
  OR U7480 ( .A(n7219), .B(n7218), .Z(n7220) );
  NAND U7481 ( .A(n7221), .B(n7220), .Z(n7331) );
  XNOR U7482 ( .A(n7334), .B(n7335), .Z(n7336) );
  XNOR U7483 ( .A(n7337), .B(n7336), .Z(n7347) );
  XNOR U7484 ( .A(n7346), .B(n7347), .Z(n7349) );
  XOR U7485 ( .A(n7348), .B(n7349), .Z(n7342) );
  NANDN U7486 ( .A(n7223), .B(n7222), .Z(n7227) );
  NANDN U7487 ( .A(n7225), .B(n7224), .Z(n7226) );
  NAND U7488 ( .A(n7227), .B(n7226), .Z(n7340) );
  OR U7489 ( .A(n7229), .B(n7228), .Z(n7233) );
  OR U7490 ( .A(n7231), .B(n7230), .Z(n7232) );
  AND U7491 ( .A(n7233), .B(n7232), .Z(n7341) );
  XNOR U7492 ( .A(n7340), .B(n7341), .Z(n7343) );
  XNOR U7493 ( .A(n7342), .B(n7343), .Z(N181) );
  NANDN U7494 ( .A(n7235), .B(n7234), .Z(n7239) );
  NANDN U7495 ( .A(n7237), .B(n7236), .Z(n7238) );
  NAND U7496 ( .A(n7239), .B(n7238), .Z(n7476) );
  OR U7497 ( .A(n7241), .B(n7240), .Z(n7245) );
  OR U7498 ( .A(n7243), .B(n7242), .Z(n7244) );
  AND U7499 ( .A(n7245), .B(n7244), .Z(n7464) );
  ANDN U7500 ( .B(y[272]), .A(n50), .Z(n7427) );
  NANDN U7501 ( .A(n7989), .B(x[80]), .Z(n7428) );
  XOR U7502 ( .A(n7427), .B(n7428), .Z(n7430) );
  NANDN U7503 ( .A(n8655), .B(x[79]), .Z(n7429) );
  XOR U7504 ( .A(n7430), .B(n7429), .Z(n7433) );
  ANDN U7505 ( .B(y[261]), .A(n54), .Z(n7246) );
  AND U7506 ( .A(y[267]), .B(x[79]), .Z(n8095) );
  NAND U7507 ( .A(n7246), .B(n8095), .Z(n7250) );
  NANDN U7508 ( .A(n7248), .B(n7247), .Z(n7249) );
  NAND U7509 ( .A(n7250), .B(n7249), .Z(n7434) );
  XNOR U7510 ( .A(n7433), .B(n7434), .Z(n7436) );
  IV U7511 ( .A(y[277]), .Z(n8703) );
  NANDN U7512 ( .A(n8703), .B(x[64]), .Z(n7410) );
  AND U7513 ( .A(n7251), .B(o[84]), .Z(n7408) );
  NANDN U7514 ( .A(n8872), .B(x[85]), .Z(n7407) );
  XNOR U7515 ( .A(n7408), .B(n7407), .Z(n7409) );
  XNOR U7516 ( .A(n7410), .B(n7409), .Z(n7435) );
  XNOR U7517 ( .A(n7436), .B(n7435), .Z(n7457) );
  ANDN U7518 ( .B(x[82]), .A(n8927), .Z(n8102) );
  NAND U7519 ( .A(n7252), .B(n8102), .Z(n7256) );
  OR U7520 ( .A(n7254), .B(n7253), .Z(n7255) );
  AND U7521 ( .A(n7256), .B(n7255), .Z(n7458) );
  XOR U7522 ( .A(n7457), .B(n7458), .Z(n7460) );
  AND U7523 ( .A(y[275]), .B(x[75]), .Z(n8836) );
  NANDN U7524 ( .A(n7257), .B(n8836), .Z(n7261) );
  OR U7525 ( .A(n7259), .B(n7258), .Z(n7260) );
  AND U7526 ( .A(n7261), .B(n7260), .Z(n7459) );
  XNOR U7527 ( .A(n7460), .B(n7459), .Z(n7463) );
  OR U7528 ( .A(n7263), .B(n7262), .Z(n7267) );
  OR U7529 ( .A(n7265), .B(n7264), .Z(n7266) );
  AND U7530 ( .A(n7267), .B(n7266), .Z(n7465) );
  XOR U7531 ( .A(n7466), .B(n7465), .Z(n7475) );
  XOR U7532 ( .A(n7476), .B(n7475), .Z(n7478) );
  OR U7533 ( .A(n7269), .B(n7268), .Z(n7273) );
  NANDN U7534 ( .A(n7271), .B(n7270), .Z(n7272) );
  NAND U7535 ( .A(n7273), .B(n7272), .Z(n7477) );
  XOR U7536 ( .A(n7478), .B(n7477), .Z(n7471) );
  OR U7537 ( .A(n7275), .B(n7274), .Z(n7279) );
  OR U7538 ( .A(n7277), .B(n7276), .Z(n7278) );
  AND U7539 ( .A(n7279), .B(n7278), .Z(n7445) );
  NAND U7540 ( .A(n7280), .B(n7427), .Z(n7284) );
  OR U7541 ( .A(n7282), .B(n7281), .Z(n7283) );
  AND U7542 ( .A(n7284), .B(n7283), .Z(n7446) );
  XNOR U7543 ( .A(n7445), .B(n7446), .Z(n7447) );
  AND U7544 ( .A(y[271]), .B(x[70]), .Z(n7402) );
  AND U7545 ( .A(y[270]), .B(x[71]), .Z(n7513) );
  AND U7546 ( .A(y[263]), .B(x[78]), .Z(n7401) );
  XNOR U7547 ( .A(n7513), .B(n7401), .Z(n7403) );
  XNOR U7548 ( .A(n7402), .B(n7403), .Z(n7385) );
  NANDN U7549 ( .A(n8815), .B(x[72]), .Z(n7382) );
  XOR U7550 ( .A(n7383), .B(n7382), .Z(n7384) );
  XNOR U7551 ( .A(n7385), .B(n7384), .Z(n7442) );
  NANDN U7552 ( .A(n49), .B(y[273]), .Z(n7422) );
  ANDN U7553 ( .B(y[274]), .A(n48), .Z(n7286) );
  ANDN U7554 ( .B(x[77]), .A(n8927), .Z(n7285) );
  XNOR U7555 ( .A(n7286), .B(n7285), .Z(n7421) );
  XNOR U7556 ( .A(n7422), .B(n7421), .Z(n7439) );
  NANDN U7557 ( .A(n8627), .B(x[76]), .Z(n7390) );
  AND U7558 ( .A(y[275]), .B(x[66]), .Z(n7389) );
  NANDN U7559 ( .A(n8626), .B(y[260]), .Z(n7388) );
  XOR U7560 ( .A(n7389), .B(n7388), .Z(n7391) );
  XNOR U7561 ( .A(n7390), .B(n7391), .Z(n7440) );
  XNOR U7562 ( .A(n7442), .B(n7441), .Z(n7448) );
  ANDN U7563 ( .B(y[273]), .A(n58), .Z(n7288) );
  NAND U7564 ( .A(n7288), .B(n7287), .Z(n7292) );
  OR U7565 ( .A(n7290), .B(n7289), .Z(n7291) );
  AND U7566 ( .A(n7292), .B(n7291), .Z(n7453) );
  AND U7567 ( .A(y[276]), .B(x[65]), .Z(n7413) );
  AND U7568 ( .A(y[259]), .B(x[82]), .Z(n7414) );
  XNOR U7569 ( .A(n7413), .B(n7414), .Z(n7416) );
  XOR U7570 ( .A(n7415), .B(n7416), .Z(n7451) );
  ANDN U7571 ( .B(y[266]), .A(n56), .Z(n7786) );
  NANDN U7572 ( .A(n8885), .B(y[257]), .Z(n7419) );
  XOR U7573 ( .A(o[85]), .B(n7419), .Z(n7397) );
  NANDN U7574 ( .A(n8824), .B(y[258]), .Z(n7396) );
  XNOR U7575 ( .A(n7397), .B(n7396), .Z(n7398) );
  XOR U7576 ( .A(n7786), .B(n7398), .Z(n7452) );
  XNOR U7577 ( .A(n7451), .B(n7452), .Z(n7454) );
  XOR U7578 ( .A(n7453), .B(n7454), .Z(n7376) );
  NAND U7579 ( .A(n7293), .B(n8090), .Z(n7297) );
  OR U7580 ( .A(n7295), .B(n7294), .Z(n7296) );
  NAND U7581 ( .A(n7297), .B(n7296), .Z(n7377) );
  XNOR U7582 ( .A(n7376), .B(n7377), .Z(n7379) );
  XNOR U7583 ( .A(n7378), .B(n7379), .Z(n7365) );
  OR U7584 ( .A(n7299), .B(n7298), .Z(n7303) );
  NANDN U7585 ( .A(n7301), .B(n7300), .Z(n7302) );
  AND U7586 ( .A(n7303), .B(n7302), .Z(n7370) );
  NANDN U7587 ( .A(n7305), .B(n7304), .Z(n7309) );
  OR U7588 ( .A(n7307), .B(n7306), .Z(n7308) );
  NAND U7589 ( .A(n7309), .B(n7308), .Z(n7371) );
  XNOR U7590 ( .A(n7370), .B(n7371), .Z(n7372) );
  OR U7591 ( .A(n7311), .B(n7310), .Z(n7315) );
  NANDN U7592 ( .A(n7313), .B(n7312), .Z(n7314) );
  NAND U7593 ( .A(n7315), .B(n7314), .Z(n7373) );
  XOR U7594 ( .A(n7365), .B(n7364), .Z(n7367) );
  OR U7595 ( .A(n7317), .B(n7316), .Z(n7321) );
  OR U7596 ( .A(n7319), .B(n7318), .Z(n7320) );
  NAND U7597 ( .A(n7321), .B(n7320), .Z(n7366) );
  XNOR U7598 ( .A(n7367), .B(n7366), .Z(n7469) );
  OR U7599 ( .A(n7323), .B(n7322), .Z(n7327) );
  NAND U7600 ( .A(n7325), .B(n7324), .Z(n7326) );
  AND U7601 ( .A(n7327), .B(n7326), .Z(n7470) );
  XNOR U7602 ( .A(n7471), .B(n7472), .Z(n7361) );
  OR U7603 ( .A(n7329), .B(n7328), .Z(n7333) );
  OR U7604 ( .A(n7331), .B(n7330), .Z(n7332) );
  NAND U7605 ( .A(n7333), .B(n7332), .Z(n7359) );
  NANDN U7606 ( .A(n7335), .B(n7334), .Z(n7339) );
  NANDN U7607 ( .A(n7337), .B(n7336), .Z(n7338) );
  NAND U7608 ( .A(n7339), .B(n7338), .Z(n7358) );
  XNOR U7609 ( .A(n7359), .B(n7358), .Z(n7360) );
  XNOR U7610 ( .A(n7361), .B(n7360), .Z(n7355) );
  NANDN U7611 ( .A(n7341), .B(n7340), .Z(n7345) );
  NAND U7612 ( .A(n7343), .B(n7342), .Z(n7344) );
  NAND U7613 ( .A(n7345), .B(n7344), .Z(n7352) );
  OR U7614 ( .A(n7347), .B(n7346), .Z(n7351) );
  OR U7615 ( .A(n7349), .B(n7348), .Z(n7350) );
  AND U7616 ( .A(n7351), .B(n7350), .Z(n7353) );
  XNOR U7617 ( .A(n7352), .B(n7353), .Z(n7354) );
  XOR U7618 ( .A(n7355), .B(n7354), .Z(N182) );
  NANDN U7619 ( .A(n7353), .B(n7352), .Z(n7357) );
  NANDN U7620 ( .A(n7355), .B(n7354), .Z(n7356) );
  NAND U7621 ( .A(n7357), .B(n7356), .Z(n7481) );
  OR U7622 ( .A(n7359), .B(n7358), .Z(n7363) );
  OR U7623 ( .A(n7361), .B(n7360), .Z(n7362) );
  AND U7624 ( .A(n7363), .B(n7362), .Z(n7482) );
  XNOR U7625 ( .A(n7481), .B(n7482), .Z(n7483) );
  NANDN U7626 ( .A(n7365), .B(n7364), .Z(n7369) );
  OR U7627 ( .A(n7367), .B(n7366), .Z(n7368) );
  AND U7628 ( .A(n7369), .B(n7368), .Z(n7493) );
  OR U7629 ( .A(n7371), .B(n7370), .Z(n7375) );
  OR U7630 ( .A(n7373), .B(n7372), .Z(n7374) );
  AND U7631 ( .A(n7375), .B(n7374), .Z(n7494) );
  XOR U7632 ( .A(n7493), .B(n7494), .Z(n7495) );
  OR U7633 ( .A(n7377), .B(n7376), .Z(n7381) );
  OR U7634 ( .A(n7379), .B(n7378), .Z(n7380) );
  NAND U7635 ( .A(n7381), .B(n7380), .Z(n7595) );
  NANDN U7636 ( .A(n7383), .B(n7382), .Z(n7387) );
  OR U7637 ( .A(n7385), .B(n7384), .Z(n7386) );
  AND U7638 ( .A(n7387), .B(n7386), .Z(n7612) );
  NANDN U7639 ( .A(n7389), .B(n7388), .Z(n7393) );
  NANDN U7640 ( .A(n7391), .B(n7390), .Z(n7392) );
  NAND U7641 ( .A(n7393), .B(n7392), .Z(n7569) );
  ANDN U7642 ( .B(x[76]), .A(n7862), .Z(n7395) );
  NANDN U7643 ( .A(n61), .B(y[260]), .Z(n7394) );
  XOR U7644 ( .A(n7395), .B(n7394), .Z(n7521) );
  NANDN U7645 ( .A(n49), .B(y[274]), .Z(n7520) );
  XNOR U7646 ( .A(n7521), .B(n7520), .Z(n7566) );
  NANDN U7647 ( .A(n50), .B(y[273]), .Z(n7537) );
  NANDN U7648 ( .A(n7989), .B(x[81]), .Z(n7536) );
  XOR U7649 ( .A(n7537), .B(n7536), .Z(n7538) );
  NANDN U7650 ( .A(n8655), .B(x[80]), .Z(n7539) );
  XOR U7651 ( .A(n7538), .B(n7539), .Z(n7567) );
  XOR U7652 ( .A(n7569), .B(n7568), .Z(n7610) );
  OR U7653 ( .A(n7397), .B(n7396), .Z(n7400) );
  NANDN U7654 ( .A(n7398), .B(n7786), .Z(n7399) );
  NAND U7655 ( .A(n7400), .B(n7399), .Z(n7611) );
  XNOR U7656 ( .A(n7610), .B(n7611), .Z(n7613) );
  XOR U7657 ( .A(n7612), .B(n7613), .Z(n7593) );
  OR U7658 ( .A(n7401), .B(n7513), .Z(n7405) );
  OR U7659 ( .A(n7403), .B(n7402), .Z(n7404) );
  NAND U7660 ( .A(n7405), .B(n7404), .Z(n7551) );
  ANDN U7661 ( .B(y[271]), .A(n52), .Z(n7406) );
  XOR U7662 ( .A(n7406), .B(n7678), .Z(n7516) );
  NANDN U7663 ( .A(n45), .B(y[278]), .Z(n7525) );
  NANDN U7664 ( .A(n8872), .B(x[86]), .Z(n7524) );
  XNOR U7665 ( .A(n7525), .B(n7524), .Z(n7527) );
  ANDN U7666 ( .B(y[257]), .A(n8827), .Z(n7542) );
  XOR U7667 ( .A(o[86]), .B(n7542), .Z(n7526) );
  XNOR U7668 ( .A(n7549), .B(n7548), .Z(n7550) );
  XOR U7669 ( .A(n7551), .B(n7550), .Z(n7563) );
  NANDN U7670 ( .A(n7408), .B(n7407), .Z(n7412) );
  NAND U7671 ( .A(n7410), .B(n7409), .Z(n7411) );
  AND U7672 ( .A(n7412), .B(n7411), .Z(n7560) );
  OR U7673 ( .A(n7414), .B(n7413), .Z(n7418) );
  OR U7674 ( .A(n7416), .B(n7415), .Z(n7417) );
  AND U7675 ( .A(n7418), .B(n7417), .Z(n7561) );
  XNOR U7676 ( .A(n7560), .B(n7561), .Z(n7562) );
  NANDN U7677 ( .A(n59), .B(y[264]), .Z(n7581) );
  NANDN U7678 ( .A(n48), .B(y[275]), .Z(n7580) );
  XOR U7679 ( .A(n7581), .B(n7580), .Z(n7582) );
  NANDN U7680 ( .A(n8881), .B(x[83]), .Z(n7583) );
  XOR U7681 ( .A(n7582), .B(n7583), .Z(n7555) );
  NANDN U7682 ( .A(n7419), .B(o[85]), .Z(n7577) );
  NANDN U7683 ( .A(n8703), .B(x[65]), .Z(n7575) );
  XOR U7684 ( .A(n7574), .B(n7575), .Z(n7576) );
  XNOR U7685 ( .A(n7577), .B(n7576), .Z(n7554) );
  XNOR U7686 ( .A(n7555), .B(n7554), .Z(n7557) );
  AND U7687 ( .A(y[274]), .B(x[77]), .Z(n8863) );
  NAND U7688 ( .A(n7420), .B(n8863), .Z(n7424) );
  OR U7689 ( .A(n7422), .B(n7421), .Z(n7423) );
  AND U7690 ( .A(n7424), .B(n7423), .Z(n7556) );
  XNOR U7691 ( .A(n7557), .B(n7556), .Z(n7605) );
  NANDN U7692 ( .A(n8885), .B(y[258]), .Z(n7531) );
  IV U7693 ( .A(y[276]), .Z(n8900) );
  NANDN U7694 ( .A(n8900), .B(x[66]), .Z(n7530) );
  XOR U7695 ( .A(n7531), .B(n7530), .Z(n7532) );
  NANDN U7696 ( .A(n58), .B(y[265]), .Z(n7533) );
  XOR U7697 ( .A(n7532), .B(n7533), .Z(n7508) );
  ANDN U7698 ( .B(y[263]), .A(n60), .Z(n7426) );
  NANDN U7699 ( .A(n55), .B(y[268]), .Z(n7425) );
  XOR U7700 ( .A(n7426), .B(n7425), .Z(n7545) );
  NANDN U7701 ( .A(n51), .B(y[272]), .Z(n7544) );
  XOR U7702 ( .A(n7545), .B(n7544), .Z(n7505) );
  NANDN U7703 ( .A(n7428), .B(n7427), .Z(n7432) );
  OR U7704 ( .A(n7430), .B(n7429), .Z(n7431) );
  NAND U7705 ( .A(n7432), .B(n7431), .Z(n7506) );
  XOR U7706 ( .A(n7508), .B(n7507), .Z(n7604) );
  XNOR U7707 ( .A(n7605), .B(n7604), .Z(n7607) );
  XOR U7708 ( .A(n7606), .B(n7607), .Z(n7601) );
  OR U7709 ( .A(n7434), .B(n7433), .Z(n7438) );
  OR U7710 ( .A(n7436), .B(n7435), .Z(n7437) );
  AND U7711 ( .A(n7438), .B(n7437), .Z(n7598) );
  OR U7712 ( .A(n7440), .B(n7439), .Z(n7444) );
  NAND U7713 ( .A(n7442), .B(n7441), .Z(n7443) );
  NAND U7714 ( .A(n7444), .B(n7443), .Z(n7599) );
  XOR U7715 ( .A(n7598), .B(n7599), .Z(n7600) );
  XOR U7716 ( .A(n7601), .B(n7600), .Z(n7592) );
  XOR U7717 ( .A(n7593), .B(n7592), .Z(n7594) );
  XNOR U7718 ( .A(n7595), .B(n7594), .Z(n7501) );
  OR U7719 ( .A(n7446), .B(n7445), .Z(n7450) );
  OR U7720 ( .A(n7448), .B(n7447), .Z(n7449) );
  AND U7721 ( .A(n7450), .B(n7449), .Z(n7586) );
  OR U7722 ( .A(n7452), .B(n7451), .Z(n7456) );
  OR U7723 ( .A(n7454), .B(n7453), .Z(n7455) );
  AND U7724 ( .A(n7456), .B(n7455), .Z(n7587) );
  XNOR U7725 ( .A(n7586), .B(n7587), .Z(n7588) );
  NANDN U7726 ( .A(n7458), .B(n7457), .Z(n7462) );
  OR U7727 ( .A(n7460), .B(n7459), .Z(n7461) );
  AND U7728 ( .A(n7462), .B(n7461), .Z(n7589) );
  OR U7729 ( .A(n7464), .B(n7463), .Z(n7468) );
  OR U7730 ( .A(n7466), .B(n7465), .Z(n7467) );
  NAND U7731 ( .A(n7468), .B(n7467), .Z(n7500) );
  XOR U7732 ( .A(n7499), .B(n7500), .Z(n7502) );
  XOR U7733 ( .A(n7501), .B(n7502), .Z(n7496) );
  XOR U7734 ( .A(n7495), .B(n7496), .Z(n7490) );
  OR U7735 ( .A(n7470), .B(n7469), .Z(n7474) );
  OR U7736 ( .A(n7472), .B(n7471), .Z(n7473) );
  AND U7737 ( .A(n7474), .B(n7473), .Z(n7487) );
  NANDN U7738 ( .A(n7476), .B(n7475), .Z(n7480) );
  OR U7739 ( .A(n7478), .B(n7477), .Z(n7479) );
  NAND U7740 ( .A(n7480), .B(n7479), .Z(n7488) );
  XNOR U7741 ( .A(n7487), .B(n7488), .Z(n7489) );
  XOR U7742 ( .A(n7490), .B(n7489), .Z(n7484) );
  XNOR U7743 ( .A(n7483), .B(n7484), .Z(N183) );
  NANDN U7744 ( .A(n7482), .B(n7481), .Z(n7486) );
  NAND U7745 ( .A(n7484), .B(n7483), .Z(n7485) );
  NAND U7746 ( .A(n7486), .B(n7485), .Z(n7616) );
  OR U7747 ( .A(n7488), .B(n7487), .Z(n7492) );
  OR U7748 ( .A(n7490), .B(n7489), .Z(n7491) );
  AND U7749 ( .A(n7492), .B(n7491), .Z(n7617) );
  XNOR U7750 ( .A(n7616), .B(n7617), .Z(n7618) );
  OR U7751 ( .A(n7494), .B(n7493), .Z(n7498) );
  NANDN U7752 ( .A(n7496), .B(n7495), .Z(n7497) );
  AND U7753 ( .A(n7498), .B(n7497), .Z(n7622) );
  NANDN U7754 ( .A(n7500), .B(n7499), .Z(n7504) );
  NANDN U7755 ( .A(n7502), .B(n7501), .Z(n7503) );
  AND U7756 ( .A(n7504), .B(n7503), .Z(n7623) );
  XOR U7757 ( .A(n7622), .B(n7623), .Z(n7625) );
  OR U7758 ( .A(n7506), .B(n7505), .Z(n7510) );
  NAND U7759 ( .A(n7508), .B(n7507), .Z(n7509) );
  NAND U7760 ( .A(n7510), .B(n7509), .Z(n7653) );
  ANDN U7761 ( .B(y[257]), .A(n8864), .Z(n7694) );
  XNOR U7762 ( .A(o[87]), .B(n7694), .Z(n7669) );
  NANDN U7763 ( .A(n45), .B(y[279]), .Z(n7667) );
  ANDN U7764 ( .B(x[87]), .A(n8872), .Z(n7666) );
  XNOR U7765 ( .A(n7667), .B(n7666), .Z(n7668) );
  XNOR U7766 ( .A(n7669), .B(n7668), .Z(n7752) );
  NANDN U7767 ( .A(n8885), .B(y[259]), .Z(n7511) );
  XOR U7768 ( .A(n7512), .B(n7511), .Z(n7691) );
  NANDN U7769 ( .A(n8824), .B(y[260]), .Z(n7690) );
  XNOR U7770 ( .A(n7691), .B(n7690), .Z(n7750) );
  NANDN U7771 ( .A(n7514), .B(n7513), .Z(n7518) );
  NANDN U7772 ( .A(n7516), .B(n7515), .Z(n7517) );
  NAND U7773 ( .A(n7518), .B(n7517), .Z(n7751) );
  XOR U7774 ( .A(n7750), .B(n7751), .Z(n7753) );
  XOR U7775 ( .A(n7752), .B(n7753), .Z(n7747) );
  ANDN U7776 ( .B(x[82]), .A(n7862), .Z(n8416) );
  IV U7777 ( .A(n8416), .Z(n8317) );
  NANDN U7778 ( .A(n8317), .B(n7519), .Z(n7523) );
  OR U7779 ( .A(n7521), .B(n7520), .Z(n7522) );
  AND U7780 ( .A(n7523), .B(n7522), .Z(n7744) );
  OR U7781 ( .A(n7525), .B(n7524), .Z(n7529) );
  NANDN U7782 ( .A(n7527), .B(n7526), .Z(n7528) );
  AND U7783 ( .A(n7529), .B(n7528), .Z(n7745) );
  XNOR U7784 ( .A(n7747), .B(n7746), .Z(n7652) );
  XOR U7785 ( .A(n7653), .B(n7652), .Z(n7655) );
  OR U7786 ( .A(n7531), .B(n7530), .Z(n7535) );
  NANDN U7787 ( .A(n7533), .B(n7532), .Z(n7534) );
  NAND U7788 ( .A(n7535), .B(n7534), .Z(n7659) );
  NANDN U7789 ( .A(n58), .B(y[266]), .Z(n7727) );
  NANDN U7790 ( .A(n8703), .B(x[66]), .Z(n7726) );
  XOR U7791 ( .A(n7727), .B(n7726), .Z(n7728) );
  NANDN U7792 ( .A(n8827), .B(y[258]), .Z(n7729) );
  XOR U7793 ( .A(n7728), .B(n7729), .Z(n7735) );
  OR U7794 ( .A(n7537), .B(n7536), .Z(n7541) );
  NANDN U7795 ( .A(n7539), .B(n7538), .Z(n7540) );
  AND U7796 ( .A(n7541), .B(n7540), .Z(n7732) );
  NAND U7797 ( .A(n7542), .B(o[86]), .Z(n7675) );
  NANDN U7798 ( .A(n57), .B(y[267]), .Z(n7673) );
  IV U7799 ( .A(y[278]), .Z(n8613) );
  NANDN U7800 ( .A(n8613), .B(x[65]), .Z(n7672) );
  XOR U7801 ( .A(n7673), .B(n7672), .Z(n7674) );
  XOR U7802 ( .A(n7675), .B(n7674), .Z(n7733) );
  XOR U7803 ( .A(n7732), .B(n7733), .Z(n7734) );
  XNOR U7804 ( .A(n7735), .B(n7734), .Z(n7658) );
  XNOR U7805 ( .A(n7659), .B(n7658), .Z(n7661) );
  AND U7806 ( .A(y[268]), .B(x[79]), .Z(n8299) );
  NAND U7807 ( .A(n7543), .B(n8299), .Z(n7547) );
  OR U7808 ( .A(n7545), .B(n7544), .Z(n7546) );
  AND U7809 ( .A(n7547), .B(n7546), .Z(n7741) );
  NANDN U7810 ( .A(n50), .B(y[274]), .Z(n7715) );
  ANDN U7811 ( .B(x[82]), .A(n7989), .Z(n7714) );
  XOR U7812 ( .A(n7715), .B(n7714), .Z(n7717) );
  ANDN U7813 ( .B(x[81]), .A(n8655), .Z(n7716) );
  XOR U7814 ( .A(n7717), .B(n7716), .Z(n7739) );
  ANDN U7815 ( .B(x[67]), .A(n8900), .Z(n7720) );
  XOR U7816 ( .A(n7721), .B(n7720), .Z(n7723) );
  ANDN U7817 ( .B(y[275]), .A(n49), .Z(n7722) );
  XNOR U7818 ( .A(n7723), .B(n7722), .Z(n7738) );
  XOR U7819 ( .A(n7739), .B(n7738), .Z(n7740) );
  XOR U7820 ( .A(n7741), .B(n7740), .Z(n7660) );
  XNOR U7821 ( .A(n7661), .B(n7660), .Z(n7654) );
  XNOR U7822 ( .A(n7655), .B(n7654), .Z(n7640) );
  NAND U7823 ( .A(n7549), .B(n7548), .Z(n7553) );
  OR U7824 ( .A(n7551), .B(n7550), .Z(n7552) );
  AND U7825 ( .A(n7553), .B(n7552), .Z(n7696) );
  OR U7826 ( .A(n7555), .B(n7554), .Z(n7559) );
  OR U7827 ( .A(n7557), .B(n7556), .Z(n7558) );
  AND U7828 ( .A(n7559), .B(n7558), .Z(n7697) );
  XNOR U7829 ( .A(n7696), .B(n7697), .Z(n7698) );
  OR U7830 ( .A(n7561), .B(n7560), .Z(n7565) );
  OR U7831 ( .A(n7563), .B(n7562), .Z(n7564) );
  NAND U7832 ( .A(n7565), .B(n7564), .Z(n7699) );
  OR U7833 ( .A(n7567), .B(n7566), .Z(n7571) );
  OR U7834 ( .A(n7569), .B(n7568), .Z(n7570) );
  AND U7835 ( .A(n7571), .B(n7570), .Z(n7628) );
  ANDN U7836 ( .B(y[271]), .A(n53), .Z(n7573) );
  NANDN U7837 ( .A(n54), .B(y[270]), .Z(n7572) );
  XOR U7838 ( .A(n7573), .B(n7572), .Z(n7680) );
  NANDN U7839 ( .A(n8884), .B(x[71]), .Z(n7679) );
  XNOR U7840 ( .A(n7680), .B(n7679), .Z(n7709) );
  ANDN U7841 ( .B(x[74]), .A(n8815), .Z(n7708) );
  XOR U7842 ( .A(n7709), .B(n7708), .Z(n7711) );
  NANDN U7843 ( .A(n51), .B(y[273]), .Z(n7684) );
  NANDN U7844 ( .A(n8927), .B(x[79]), .Z(n7683) );
  XOR U7845 ( .A(n7684), .B(n7683), .Z(n7686) );
  XNOR U7846 ( .A(n7685), .B(n7686), .Z(n7710) );
  XOR U7847 ( .A(n7711), .B(n7710), .Z(n7705) );
  NANDN U7848 ( .A(n7575), .B(n7574), .Z(n7579) );
  OR U7849 ( .A(n7577), .B(n7576), .Z(n7578) );
  NAND U7850 ( .A(n7579), .B(n7578), .Z(n7703) );
  OR U7851 ( .A(n7581), .B(n7580), .Z(n7585) );
  NANDN U7852 ( .A(n7583), .B(n7582), .Z(n7584) );
  NAND U7853 ( .A(n7585), .B(n7584), .Z(n7702) );
  XNOR U7854 ( .A(n7705), .B(n7704), .Z(n7629) );
  XNOR U7855 ( .A(n7628), .B(n7629), .Z(n7630) );
  XOR U7856 ( .A(n7640), .B(n7641), .Z(n7643) );
  OR U7857 ( .A(n7587), .B(n7586), .Z(n7591) );
  OR U7858 ( .A(n7589), .B(n7588), .Z(n7590) );
  AND U7859 ( .A(n7591), .B(n7590), .Z(n7642) );
  XNOR U7860 ( .A(n7643), .B(n7642), .Z(n7648) );
  NANDN U7861 ( .A(n7593), .B(n7592), .Z(n7597) );
  OR U7862 ( .A(n7595), .B(n7594), .Z(n7596) );
  NAND U7863 ( .A(n7597), .B(n7596), .Z(n7647) );
  OR U7864 ( .A(n7599), .B(n7598), .Z(n7603) );
  NANDN U7865 ( .A(n7601), .B(n7600), .Z(n7602) );
  AND U7866 ( .A(n7603), .B(n7602), .Z(n7637) );
  OR U7867 ( .A(n7605), .B(n7604), .Z(n7609) );
  OR U7868 ( .A(n7607), .B(n7606), .Z(n7608) );
  NAND U7869 ( .A(n7609), .B(n7608), .Z(n7635) );
  OR U7870 ( .A(n7611), .B(n7610), .Z(n7615) );
  OR U7871 ( .A(n7613), .B(n7612), .Z(n7614) );
  AND U7872 ( .A(n7615), .B(n7614), .Z(n7634) );
  XNOR U7873 ( .A(n7635), .B(n7634), .Z(n7636) );
  XNOR U7874 ( .A(n7647), .B(n7646), .Z(n7649) );
  XNOR U7875 ( .A(n7625), .B(n7624), .Z(n7619) );
  XOR U7876 ( .A(n7618), .B(n7619), .Z(N184) );
  NANDN U7877 ( .A(n7617), .B(n7616), .Z(n7621) );
  NANDN U7878 ( .A(n7619), .B(n7618), .Z(n7620) );
  NAND U7879 ( .A(n7621), .B(n7620), .Z(n7756) );
  OR U7880 ( .A(n7623), .B(n7622), .Z(n7627) );
  NAND U7881 ( .A(n7625), .B(n7624), .Z(n7626) );
  AND U7882 ( .A(n7627), .B(n7626), .Z(n7757) );
  XNOR U7883 ( .A(n7756), .B(n7757), .Z(n7758) );
  OR U7884 ( .A(n7629), .B(n7628), .Z(n7633) );
  OR U7885 ( .A(n7631), .B(n7630), .Z(n7632) );
  NAND U7886 ( .A(n7633), .B(n7632), .Z(n7893) );
  OR U7887 ( .A(n7635), .B(n7634), .Z(n7639) );
  OR U7888 ( .A(n7637), .B(n7636), .Z(n7638) );
  AND U7889 ( .A(n7639), .B(n7638), .Z(n7892) );
  XNOR U7890 ( .A(n7893), .B(n7892), .Z(n7894) );
  NANDN U7891 ( .A(n7641), .B(n7640), .Z(n7645) );
  OR U7892 ( .A(n7643), .B(n7642), .Z(n7644) );
  NAND U7893 ( .A(n7645), .B(n7644), .Z(n7895) );
  OR U7894 ( .A(n7647), .B(n7646), .Z(n7651) );
  NANDN U7895 ( .A(n7649), .B(n7648), .Z(n7650) );
  AND U7896 ( .A(n7651), .B(n7650), .Z(n7763) );
  NANDN U7897 ( .A(n7653), .B(n7652), .Z(n7657) );
  NANDN U7898 ( .A(n7655), .B(n7654), .Z(n7656) );
  NAND U7899 ( .A(n7657), .B(n7656), .Z(n7770) );
  NAND U7900 ( .A(n7659), .B(n7658), .Z(n7663) );
  NANDN U7901 ( .A(n7661), .B(n7660), .Z(n7662) );
  AND U7902 ( .A(n7663), .B(n7662), .Z(n7768) );
  NANDN U7903 ( .A(n53), .B(y[272]), .Z(n7788) );
  ANDN U7904 ( .B(x[75]), .A(n8815), .Z(n7665) );
  NANDN U7905 ( .A(n59), .B(y[266]), .Z(n7664) );
  XOR U7906 ( .A(n7665), .B(n7664), .Z(n7787) );
  XNOR U7907 ( .A(n7788), .B(n7787), .Z(n7783) );
  AND U7908 ( .A(y[271]), .B(x[73]), .Z(n7781) );
  NAND U7909 ( .A(y[270]), .B(x[74]), .Z(n7780) );
  XNOR U7910 ( .A(n7781), .B(n7780), .Z(n7782) );
  XOR U7911 ( .A(n7783), .B(n7782), .Z(n7826) );
  NANDN U7912 ( .A(n7667), .B(n7666), .Z(n7671) );
  NANDN U7913 ( .A(n7669), .B(n7668), .Z(n7670) );
  AND U7914 ( .A(n7671), .B(n7670), .Z(n7824) );
  NANDN U7915 ( .A(n49), .B(y[276]), .Z(n7821) );
  NANDN U7916 ( .A(n48), .B(y[277]), .Z(n7819) );
  NANDN U7917 ( .A(n8627), .B(x[79]), .Z(n7818) );
  XOR U7918 ( .A(n7819), .B(n7818), .Z(n7820) );
  XOR U7919 ( .A(n7821), .B(n7820), .Z(n7825) );
  XOR U7920 ( .A(n7826), .B(n7827), .Z(n7832) );
  OR U7921 ( .A(n7673), .B(n7672), .Z(n7677) );
  NANDN U7922 ( .A(n7675), .B(n7674), .Z(n7676) );
  NAND U7923 ( .A(n7677), .B(n7676), .Z(n7850) );
  NANDN U7924 ( .A(n7678), .B(n7781), .Z(n7682) );
  OR U7925 ( .A(n7680), .B(n7679), .Z(n7681) );
  AND U7926 ( .A(n7682), .B(n7681), .Z(n7848) );
  NANDN U7927 ( .A(n8890), .B(y[264]), .Z(n7857) );
  NANDN U7928 ( .A(n50), .B(y[275]), .Z(n7855) );
  NANDN U7929 ( .A(n8827), .B(y[259]), .Z(n7854) );
  XNOR U7930 ( .A(n7855), .B(n7854), .Z(n7856) );
  XNOR U7931 ( .A(n7857), .B(n7856), .Z(n7877) );
  OR U7932 ( .A(n7684), .B(n7683), .Z(n7688) );
  NAND U7933 ( .A(n7686), .B(n7685), .Z(n7687) );
  AND U7934 ( .A(n7688), .B(n7687), .Z(n7875) );
  AND U7935 ( .A(y[260]), .B(x[84]), .Z(n7990) );
  NANDN U7936 ( .A(n8824), .B(y[261]), .Z(n7864) );
  ANDN U7937 ( .B(y[274]), .A(n51), .Z(n7863) );
  XNOR U7938 ( .A(n7864), .B(n7863), .Z(n7865) );
  XOR U7939 ( .A(n7990), .B(n7865), .Z(n7874) );
  XOR U7940 ( .A(n7875), .B(n7874), .Z(n7876) );
  XNOR U7941 ( .A(n7877), .B(n7876), .Z(n7849) );
  XOR U7942 ( .A(n7850), .B(n7851), .Z(n7830) );
  NANDN U7943 ( .A(n47), .B(y[278]), .Z(n7792) );
  NANDN U7944 ( .A(n8864), .B(y[258]), .Z(n7791) );
  XNOR U7945 ( .A(n7792), .B(n7791), .Z(n7794) );
  XOR U7946 ( .A(n7793), .B(n7794), .Z(n7883) );
  ANDN U7947 ( .B(y[259]), .A(n8890), .Z(n7689) );
  AND U7948 ( .A(y[263]), .B(x[84]), .Z(n8242) );
  NAND U7949 ( .A(n7689), .B(n8242), .Z(n7693) );
  OR U7950 ( .A(n7691), .B(n7690), .Z(n7692) );
  AND U7951 ( .A(n7693), .B(n7692), .Z(n7880) );
  NAND U7952 ( .A(n7694), .B(o[87]), .Z(n7800) );
  NANDN U7953 ( .A(n46), .B(y[279]), .Z(n7798) );
  XNOR U7954 ( .A(n7695), .B(n7798), .Z(n7799) );
  XOR U7955 ( .A(n7800), .B(n7799), .Z(n7881) );
  XNOR U7956 ( .A(n7883), .B(n7882), .Z(n7831) );
  XOR U7957 ( .A(n7830), .B(n7831), .Z(n7833) );
  XOR U7958 ( .A(n7832), .B(n7833), .Z(n7769) );
  XOR U7959 ( .A(n7770), .B(n7771), .Z(n7900) );
  OR U7960 ( .A(n7697), .B(n7696), .Z(n7701) );
  OR U7961 ( .A(n7699), .B(n7698), .Z(n7700) );
  NAND U7962 ( .A(n7701), .B(n7700), .Z(n7899) );
  OR U7963 ( .A(n7703), .B(n7702), .Z(n7707) );
  NANDN U7964 ( .A(n7705), .B(n7704), .Z(n7706) );
  NAND U7965 ( .A(n7707), .B(n7706), .Z(n7777) );
  NANDN U7966 ( .A(n7709), .B(n7708), .Z(n7713) );
  OR U7967 ( .A(n7711), .B(n7710), .Z(n7712) );
  AND U7968 ( .A(n7713), .B(n7712), .Z(n7775) );
  NANDN U7969 ( .A(n7715), .B(n7714), .Z(n7719) );
  NANDN U7970 ( .A(n7717), .B(n7716), .Z(n7718) );
  AND U7971 ( .A(n7719), .B(n7718), .Z(n7870) );
  AND U7972 ( .A(y[257]), .B(x[87]), .Z(n7804) );
  XOR U7973 ( .A(o[88]), .B(n7804), .Z(n7814) );
  NANDN U7974 ( .A(n45), .B(y[280]), .Z(n7813) );
  NANDN U7975 ( .A(n8865), .B(y[256]), .Z(n7812) );
  XNOR U7976 ( .A(n7813), .B(n7812), .Z(n7815) );
  XOR U7977 ( .A(n7814), .B(n7815), .Z(n7869) );
  NANDN U7978 ( .A(n61), .B(y[262]), .Z(n7808) );
  NANDN U7979 ( .A(n8626), .B(y[263]), .Z(n7806) );
  ANDN U7980 ( .B(x[71]), .A(n8904), .Z(n7805) );
  XOR U7981 ( .A(n7806), .B(n7805), .Z(n7807) );
  XOR U7982 ( .A(n7869), .B(n7868), .Z(n7871) );
  XNOR U7983 ( .A(n7870), .B(n7871), .Z(n7845) );
  NANDN U7984 ( .A(n7721), .B(n7720), .Z(n7725) );
  NANDN U7985 ( .A(n7723), .B(n7722), .Z(n7724) );
  AND U7986 ( .A(n7725), .B(n7724), .Z(n7842) );
  OR U7987 ( .A(n7727), .B(n7726), .Z(n7731) );
  NANDN U7988 ( .A(n7729), .B(n7728), .Z(n7730) );
  AND U7989 ( .A(n7731), .B(n7730), .Z(n7843) );
  XOR U7990 ( .A(n7775), .B(n7774), .Z(n7776) );
  XOR U7991 ( .A(n7777), .B(n7776), .Z(n7888) );
  OR U7992 ( .A(n7733), .B(n7732), .Z(n7737) );
  NANDN U7993 ( .A(n7735), .B(n7734), .Z(n7736) );
  AND U7994 ( .A(n7737), .B(n7736), .Z(n7886) );
  NANDN U7995 ( .A(n7739), .B(n7738), .Z(n7743) );
  OR U7996 ( .A(n7741), .B(n7740), .Z(n7742) );
  NAND U7997 ( .A(n7743), .B(n7742), .Z(n7839) );
  OR U7998 ( .A(n7745), .B(n7744), .Z(n7749) );
  NANDN U7999 ( .A(n7747), .B(n7746), .Z(n7748) );
  AND U8000 ( .A(n7749), .B(n7748), .Z(n7836) );
  NANDN U8001 ( .A(n7751), .B(n7750), .Z(n7755) );
  OR U8002 ( .A(n7753), .B(n7752), .Z(n7754) );
  NAND U8003 ( .A(n7755), .B(n7754), .Z(n7837) );
  XNOR U8004 ( .A(n7839), .B(n7838), .Z(n7887) );
  XOR U8005 ( .A(n7888), .B(n7889), .Z(n7898) );
  XNOR U8006 ( .A(n7899), .B(n7898), .Z(n7901) );
  XNOR U8007 ( .A(n7900), .B(n7901), .Z(n7762) );
  XOR U8008 ( .A(n7763), .B(n7762), .Z(n7764) );
  XNOR U8009 ( .A(n7765), .B(n7764), .Z(n7759) );
  XOR U8010 ( .A(n7758), .B(n7759), .Z(N185) );
  NANDN U8011 ( .A(n7757), .B(n7756), .Z(n7761) );
  NANDN U8012 ( .A(n7759), .B(n7758), .Z(n7760) );
  NAND U8013 ( .A(n7761), .B(n7760), .Z(n7904) );
  NANDN U8014 ( .A(n7763), .B(n7762), .Z(n7767) );
  OR U8015 ( .A(n7765), .B(n7764), .Z(n7766) );
  AND U8016 ( .A(n7767), .B(n7766), .Z(n7905) );
  XNOR U8017 ( .A(n7904), .B(n7905), .Z(n7906) );
  OR U8018 ( .A(n7769), .B(n7768), .Z(n7773) );
  NANDN U8019 ( .A(n7771), .B(n7770), .Z(n7772) );
  NAND U8020 ( .A(n7773), .B(n7772), .Z(n8052) );
  NANDN U8021 ( .A(n7775), .B(n7774), .Z(n7779) );
  OR U8022 ( .A(n7777), .B(n7776), .Z(n7778) );
  AND U8023 ( .A(n7779), .B(n7778), .Z(n8040) );
  NANDN U8024 ( .A(n7781), .B(n7780), .Z(n7785) );
  NAND U8025 ( .A(n7783), .B(n7782), .Z(n7784) );
  NAND U8026 ( .A(n7785), .B(n7784), .Z(n7947) );
  NANDN U8027 ( .A(n46), .B(y[280]), .Z(n8002) );
  ANDN U8028 ( .B(y[268]), .A(n58), .Z(n8001) );
  XNOR U8029 ( .A(n8002), .B(n8001), .Z(n8004) );
  NANDN U8030 ( .A(n8865), .B(y[257]), .Z(n7964) );
  XNOR U8031 ( .A(n7964), .B(o[89]), .Z(n8003) );
  XNOR U8032 ( .A(n8004), .B(n8003), .Z(n8010) );
  NAND U8033 ( .A(y[270]), .B(x[75]), .Z(n7967) );
  NAND U8034 ( .A(y[269]), .B(x[76]), .Z(n7965) );
  NAND U8035 ( .A(x[71]), .B(y[274]), .Z(n7966) );
  XNOR U8036 ( .A(n7965), .B(n7966), .Z(n7968) );
  XNOR U8037 ( .A(n7967), .B(n7968), .Z(n8007) );
  ANDN U8038 ( .B(x[78]), .A(n8815), .Z(n8289) );
  NAND U8039 ( .A(n7786), .B(n8289), .Z(n7790) );
  OR U8040 ( .A(n7788), .B(n7787), .Z(n7789) );
  AND U8041 ( .A(n7790), .B(n7789), .Z(n8008) );
  XNOR U8042 ( .A(n8007), .B(n8008), .Z(n8009) );
  XNOR U8043 ( .A(n8010), .B(n8009), .Z(n7946) );
  XNOR U8044 ( .A(n7947), .B(n7946), .Z(n7949) );
  OR U8045 ( .A(n7792), .B(n7791), .Z(n7796) );
  NANDN U8046 ( .A(n7794), .B(n7793), .Z(n7795) );
  AND U8047 ( .A(n7796), .B(n7795), .Z(n7940) );
  OR U8048 ( .A(n7798), .B(n7797), .Z(n7802) );
  NANDN U8049 ( .A(n7800), .B(n7799), .Z(n7801) );
  AND U8050 ( .A(n7802), .B(n7801), .Z(n7941) );
  XOR U8051 ( .A(n7940), .B(n7941), .Z(n7942) );
  NAND U8052 ( .A(y[273]), .B(x[72]), .Z(n7936) );
  XNOR U8053 ( .A(n7935), .B(n7803), .Z(n7937) );
  XNOR U8054 ( .A(n7936), .B(n7937), .Z(n7922) );
  AND U8055 ( .A(n7804), .B(o[88]), .Z(n7931) );
  NAND U8056 ( .A(y[256]), .B(x[89]), .Z(n7928) );
  NANDN U8057 ( .A(n45), .B(y[281]), .Z(n7929) );
  XNOR U8058 ( .A(n7928), .B(n7929), .Z(n7930) );
  XOR U8059 ( .A(n7931), .B(n7930), .Z(n7923) );
  XNOR U8060 ( .A(n7922), .B(n7923), .Z(n7925) );
  NANDN U8061 ( .A(n7806), .B(n7805), .Z(n7810) );
  OR U8062 ( .A(n7808), .B(n7807), .Z(n7809) );
  AND U8063 ( .A(n7810), .B(n7809), .Z(n7924) );
  XNOR U8064 ( .A(n7925), .B(n7924), .Z(n7943) );
  XOR U8065 ( .A(n7942), .B(n7943), .Z(n7948) );
  XOR U8066 ( .A(n7949), .B(n7948), .Z(n8045) );
  NANDN U8067 ( .A(n47), .B(y[279]), .Z(n7998) );
  NANDN U8068 ( .A(n48), .B(y[278]), .Z(n7996) );
  XNOR U8069 ( .A(n7811), .B(n7996), .Z(n7997) );
  XOR U8070 ( .A(n7998), .B(n7997), .Z(n8026) );
  OR U8071 ( .A(n7813), .B(n7812), .Z(n7817) );
  NANDN U8072 ( .A(n7815), .B(n7814), .Z(n7816) );
  AND U8073 ( .A(n7817), .B(n7816), .Z(n8025) );
  XOR U8074 ( .A(n8026), .B(n8025), .Z(n8027) );
  OR U8075 ( .A(n7819), .B(n7818), .Z(n7823) );
  NANDN U8076 ( .A(n7821), .B(n7820), .Z(n7822) );
  AND U8077 ( .A(n7823), .B(n7822), .Z(n8028) );
  XNOR U8078 ( .A(n8027), .B(n8028), .Z(n8043) );
  OR U8079 ( .A(n7825), .B(n7824), .Z(n7829) );
  OR U8080 ( .A(n7827), .B(n7826), .Z(n7828) );
  NAND U8081 ( .A(n7829), .B(n7828), .Z(n8044) );
  XNOR U8082 ( .A(n8043), .B(n8044), .Z(n8046) );
  XNOR U8083 ( .A(n8045), .B(n8046), .Z(n8037) );
  NANDN U8084 ( .A(n7831), .B(n7830), .Z(n7835) );
  OR U8085 ( .A(n7833), .B(n7832), .Z(n7834) );
  NAND U8086 ( .A(n7835), .B(n7834), .Z(n8038) );
  XNOR U8087 ( .A(n8037), .B(n8038), .Z(n8039) );
  XOR U8088 ( .A(n8040), .B(n8039), .Z(n8049) );
  OR U8089 ( .A(n7837), .B(n7836), .Z(n7841) );
  NAND U8090 ( .A(n7839), .B(n7838), .Z(n7840) );
  NAND U8091 ( .A(n7841), .B(n7840), .Z(n7917) );
  OR U8092 ( .A(n7843), .B(n7842), .Z(n7847) );
  NANDN U8093 ( .A(n7845), .B(n7844), .Z(n7846) );
  NAND U8094 ( .A(n7847), .B(n7846), .Z(n7959) );
  OR U8095 ( .A(n7849), .B(n7848), .Z(n7853) );
  NANDN U8096 ( .A(n7851), .B(n7850), .Z(n7852) );
  NAND U8097 ( .A(n7853), .B(n7852), .Z(n7958) );
  XNOR U8098 ( .A(n7959), .B(n7958), .Z(n7960) );
  OR U8099 ( .A(n7855), .B(n7854), .Z(n7859) );
  OR U8100 ( .A(n7857), .B(n7856), .Z(n7858) );
  AND U8101 ( .A(n7859), .B(n7858), .Z(n8021) );
  NAND U8102 ( .A(y[259]), .B(x[86]), .Z(n7973) );
  NAND U8103 ( .A(y[276]), .B(x[69]), .Z(n7971) );
  NAND U8104 ( .A(y[264]), .B(x[81]), .Z(n7972) );
  XNOR U8105 ( .A(n7971), .B(n7972), .Z(n7974) );
  XNOR U8106 ( .A(n7973), .B(n7974), .Z(n8020) );
  NANDN U8107 ( .A(n8824), .B(y[262]), .Z(n7992) );
  ANDN U8108 ( .B(x[84]), .A(n7989), .Z(n7861) );
  ANDN U8109 ( .B(y[260]), .A(n8827), .Z(n7860) );
  XNOR U8110 ( .A(n7861), .B(n7860), .Z(n7991) );
  XOR U8111 ( .A(n7992), .B(n7991), .Z(n8019) );
  XOR U8112 ( .A(n8020), .B(n8019), .Z(n8022) );
  XOR U8113 ( .A(n8021), .B(n8022), .Z(n7952) );
  ANDN U8114 ( .B(y[258]), .A(n8656), .Z(n7979) );
  NAND U8115 ( .A(y[277]), .B(x[68]), .Z(n7977) );
  NAND U8116 ( .A(y[265]), .B(x[80]), .Z(n7978) );
  XNOR U8117 ( .A(n7977), .B(n7978), .Z(n7980) );
  XNOR U8118 ( .A(n7979), .B(n7980), .Z(n8015) );
  ANDN U8119 ( .B(x[79]), .A(n7862), .Z(n7985) );
  NAND U8120 ( .A(x[82]), .B(y[263]), .Z(n7983) );
  NAND U8121 ( .A(x[70]), .B(y[275]), .Z(n7984) );
  XNOR U8122 ( .A(n7983), .B(n7984), .Z(n7986) );
  XOR U8123 ( .A(n7985), .B(n7986), .Z(n8014) );
  NANDN U8124 ( .A(n7864), .B(n7863), .Z(n7867) );
  NAND U8125 ( .A(n7865), .B(n7990), .Z(n7866) );
  AND U8126 ( .A(n7867), .B(n7866), .Z(n8013) );
  XNOR U8127 ( .A(n8014), .B(n8013), .Z(n8016) );
  XOR U8128 ( .A(n8015), .B(n8016), .Z(n7953) );
  XOR U8129 ( .A(n7952), .B(n7953), .Z(n7955) );
  NANDN U8130 ( .A(n7869), .B(n7868), .Z(n7873) );
  OR U8131 ( .A(n7871), .B(n7870), .Z(n7872) );
  AND U8132 ( .A(n7873), .B(n7872), .Z(n7954) );
  XNOR U8133 ( .A(n7955), .B(n7954), .Z(n8031) );
  NANDN U8134 ( .A(n7875), .B(n7874), .Z(n7879) );
  OR U8135 ( .A(n7877), .B(n7876), .Z(n7878) );
  AND U8136 ( .A(n7879), .B(n7878), .Z(n8032) );
  OR U8137 ( .A(n7881), .B(n7880), .Z(n7885) );
  NANDN U8138 ( .A(n7883), .B(n7882), .Z(n7884) );
  AND U8139 ( .A(n7885), .B(n7884), .Z(n8033) );
  XOR U8140 ( .A(n8034), .B(n8033), .Z(n7961) );
  XOR U8141 ( .A(n7917), .B(n7916), .Z(n7919) );
  OR U8142 ( .A(n7887), .B(n7886), .Z(n7891) );
  NAND U8143 ( .A(n7889), .B(n7888), .Z(n7890) );
  NAND U8144 ( .A(n7891), .B(n7890), .Z(n7918) );
  XNOR U8145 ( .A(n7919), .B(n7918), .Z(n8050) );
  XOR U8146 ( .A(n8052), .B(n8051), .Z(n7913) );
  OR U8147 ( .A(n7893), .B(n7892), .Z(n7897) );
  OR U8148 ( .A(n7895), .B(n7894), .Z(n7896) );
  AND U8149 ( .A(n7897), .B(n7896), .Z(n7911) );
  OR U8150 ( .A(n7899), .B(n7898), .Z(n7903) );
  NANDN U8151 ( .A(n7901), .B(n7900), .Z(n7902) );
  AND U8152 ( .A(n7903), .B(n7902), .Z(n7910) );
  XNOR U8153 ( .A(n7911), .B(n7910), .Z(n7912) );
  XNOR U8154 ( .A(n7913), .B(n7912), .Z(n7907) );
  XOR U8155 ( .A(n7906), .B(n7907), .Z(N186) );
  NANDN U8156 ( .A(n7905), .B(n7904), .Z(n7909) );
  NANDN U8157 ( .A(n7907), .B(n7906), .Z(n7908) );
  NAND U8158 ( .A(n7909), .B(n7908), .Z(n8055) );
  OR U8159 ( .A(n7911), .B(n7910), .Z(n7915) );
  OR U8160 ( .A(n7913), .B(n7912), .Z(n7914) );
  AND U8161 ( .A(n7915), .B(n7914), .Z(n8056) );
  XNOR U8162 ( .A(n8055), .B(n8056), .Z(n8057) );
  NANDN U8163 ( .A(n7917), .B(n7916), .Z(n7921) );
  OR U8164 ( .A(n7919), .B(n7918), .Z(n7920) );
  NAND U8165 ( .A(n7921), .B(n7920), .Z(n8064) );
  OR U8166 ( .A(n7923), .B(n7922), .Z(n7927) );
  OR U8167 ( .A(n7925), .B(n7924), .Z(n7926) );
  AND U8168 ( .A(n7927), .B(n7926), .Z(n8192) );
  NANDN U8169 ( .A(n47), .B(y[280]), .Z(n8096) );
  XNOR U8170 ( .A(n8096), .B(n8095), .Z(n8098) );
  AND U8171 ( .A(y[258]), .B(x[88]), .Z(n8097) );
  XOR U8172 ( .A(n8098), .B(n8097), .Z(n8119) );
  NAND U8173 ( .A(n7929), .B(n7928), .Z(n7933) );
  OR U8174 ( .A(n7931), .B(n7930), .Z(n7932) );
  AND U8175 ( .A(n7933), .B(n7932), .Z(n8120) );
  XNOR U8176 ( .A(n8119), .B(n8120), .Z(n8122) );
  NANDN U8177 ( .A(n7935), .B(n7934), .Z(n7939) );
  NANDN U8178 ( .A(n7937), .B(n7936), .Z(n7938) );
  AND U8179 ( .A(n7939), .B(n7938), .Z(n8121) );
  XOR U8180 ( .A(n8122), .B(n8121), .Z(n8193) );
  XNOR U8181 ( .A(n8192), .B(n8193), .Z(n8195) );
  OR U8182 ( .A(n7941), .B(n7940), .Z(n7945) );
  NANDN U8183 ( .A(n7943), .B(n7942), .Z(n7944) );
  AND U8184 ( .A(n7945), .B(n7944), .Z(n8194) );
  XOR U8185 ( .A(n8195), .B(n8194), .Z(n8158) );
  OR U8186 ( .A(n7947), .B(n7946), .Z(n7951) );
  OR U8187 ( .A(n7949), .B(n7948), .Z(n7950) );
  NAND U8188 ( .A(n7951), .B(n7950), .Z(n8156) );
  NANDN U8189 ( .A(n7953), .B(n7952), .Z(n7957) );
  OR U8190 ( .A(n7955), .B(n7954), .Z(n7956) );
  NAND U8191 ( .A(n7957), .B(n7956), .Z(n8155) );
  XOR U8192 ( .A(n8156), .B(n8155), .Z(n8157) );
  XOR U8193 ( .A(n8158), .B(n8157), .Z(n8070) );
  OR U8194 ( .A(n7959), .B(n7958), .Z(n7963) );
  OR U8195 ( .A(n7961), .B(n7960), .Z(n7962) );
  AND U8196 ( .A(n7963), .B(n7962), .Z(n8067) );
  NANDN U8197 ( .A(n7964), .B(o[89]), .Z(n8169) );
  NAND U8198 ( .A(x[78]), .B(y[268]), .Z(n8167) );
  NAND U8199 ( .A(x[65]), .B(y[281]), .Z(n8168) );
  XNOR U8200 ( .A(n8167), .B(n8168), .Z(n8170) );
  XNOR U8201 ( .A(n8169), .B(n8170), .Z(n8125) );
  NANDN U8202 ( .A(n45), .B(y[282]), .Z(n8138) );
  AND U8203 ( .A(y[256]), .B(x[90]), .Z(n8137) );
  XNOR U8204 ( .A(n8138), .B(n8137), .Z(n8140) );
  NANDN U8205 ( .A(n8928), .B(y[257]), .Z(n8179) );
  XNOR U8206 ( .A(n8179), .B(o[90]), .Z(n8139) );
  XNOR U8207 ( .A(n8140), .B(n8139), .Z(n8126) );
  XNOR U8208 ( .A(n8125), .B(n8126), .Z(n8128) );
  NAND U8209 ( .A(n7966), .B(n7965), .Z(n7970) );
  NANDN U8210 ( .A(n7968), .B(n7967), .Z(n7969) );
  NAND U8211 ( .A(n7970), .B(n7969), .Z(n8127) );
  XOR U8212 ( .A(n8128), .B(n8127), .Z(n8082) );
  NAND U8213 ( .A(n7972), .B(n7971), .Z(n7976) );
  NANDN U8214 ( .A(n7974), .B(n7973), .Z(n7975) );
  NAND U8215 ( .A(n7976), .B(n7975), .Z(n8079) );
  NAND U8216 ( .A(n7978), .B(n7977), .Z(n7982) );
  OR U8217 ( .A(n7980), .B(n7979), .Z(n7981) );
  AND U8218 ( .A(n7982), .B(n7981), .Z(n8080) );
  XNOR U8219 ( .A(n8079), .B(n8080), .Z(n8081) );
  XOR U8220 ( .A(n8082), .B(n8081), .Z(n8146) );
  NAND U8221 ( .A(y[278]), .B(x[68]), .Z(n8101) );
  XOR U8222 ( .A(n8102), .B(n8101), .Z(n8104) );
  XNOR U8223 ( .A(n8103), .B(n8104), .Z(n8083) );
  NAND U8224 ( .A(n7984), .B(n7983), .Z(n7988) );
  OR U8225 ( .A(n7986), .B(n7985), .Z(n7987) );
  NAND U8226 ( .A(n7988), .B(n7987), .Z(n8084) );
  XOR U8227 ( .A(n8083), .B(n8084), .Z(n8086) );
  NANDN U8228 ( .A(n8824), .B(y[263]), .Z(n8162) );
  AND U8229 ( .A(y[271]), .B(x[75]), .Z(n8161) );
  XNOR U8230 ( .A(n8162), .B(n8161), .Z(n8163) );
  NANDN U8231 ( .A(n48), .B(y[279]), .Z(n8164) );
  XNOR U8232 ( .A(n8163), .B(n8164), .Z(n8085) );
  XOR U8233 ( .A(n8086), .B(n8085), .Z(n8143) );
  ANDN U8234 ( .B(x[85]), .A(n7989), .Z(n8174) );
  NAND U8235 ( .A(n7990), .B(n8174), .Z(n7994) );
  OR U8236 ( .A(n7992), .B(n7991), .Z(n7993) );
  NAND U8237 ( .A(n7994), .B(n7993), .Z(n8074) );
  NANDN U8238 ( .A(n8864), .B(y[260]), .Z(n8092) );
  NANDN U8239 ( .A(n8881), .B(x[87]), .Z(n8089) );
  XNOR U8240 ( .A(n8090), .B(n8089), .Z(n8091) );
  XNOR U8241 ( .A(n8092), .B(n8091), .Z(n8073) );
  XNOR U8242 ( .A(n8074), .B(n8073), .Z(n8076) );
  NAND U8243 ( .A(y[262]), .B(x[84]), .Z(n8175) );
  XOR U8244 ( .A(n8174), .B(n8173), .Z(n8176) );
  XOR U8245 ( .A(n8175), .B(n8176), .Z(n8075) );
  XNOR U8246 ( .A(n8076), .B(n8075), .Z(n8144) );
  XOR U8247 ( .A(n8143), .B(n8144), .Z(n8145) );
  XOR U8248 ( .A(n8146), .B(n8145), .Z(n8151) );
  OR U8249 ( .A(n7996), .B(n7995), .Z(n8000) );
  NANDN U8250 ( .A(n7998), .B(n7997), .Z(n7999) );
  NAND U8251 ( .A(n8000), .B(n7999), .Z(n8108) );
  NANDN U8252 ( .A(n8002), .B(n8001), .Z(n8006) );
  NAND U8253 ( .A(n8004), .B(n8003), .Z(n8005) );
  NAND U8254 ( .A(n8006), .B(n8005), .Z(n8107) );
  XNOR U8255 ( .A(n8108), .B(n8107), .Z(n8109) );
  NAND U8256 ( .A(y[273]), .B(x[73]), .Z(n8182) );
  NAND U8257 ( .A(y[276]), .B(x[70]), .Z(n8180) );
  NAND U8258 ( .A(x[72]), .B(y[274]), .Z(n8181) );
  XNOR U8259 ( .A(n8180), .B(n8181), .Z(n8183) );
  XOR U8260 ( .A(n8182), .B(n8183), .Z(n8189) );
  AND U8261 ( .A(y[275]), .B(x[71]), .Z(n8186) );
  NAND U8262 ( .A(y[272]), .B(x[74]), .Z(n8133) );
  NAND U8263 ( .A(y[270]), .B(x[76]), .Z(n8131) );
  NAND U8264 ( .A(y[277]), .B(x[69]), .Z(n8132) );
  XNOR U8265 ( .A(n8131), .B(n8132), .Z(n8134) );
  XOR U8266 ( .A(n8133), .B(n8134), .Z(n8187) );
  XNOR U8267 ( .A(n8186), .B(n8187), .Z(n8188) );
  XNOR U8268 ( .A(n8189), .B(n8188), .Z(n8110) );
  OR U8269 ( .A(n8008), .B(n8007), .Z(n8012) );
  OR U8270 ( .A(n8010), .B(n8009), .Z(n8011) );
  AND U8271 ( .A(n8012), .B(n8011), .Z(n8150) );
  XNOR U8272 ( .A(n8149), .B(n8150), .Z(n8152) );
  XNOR U8273 ( .A(n8151), .B(n8152), .Z(n8113) );
  OR U8274 ( .A(n8014), .B(n8013), .Z(n8018) );
  NANDN U8275 ( .A(n8016), .B(n8015), .Z(n8017) );
  NAND U8276 ( .A(n8018), .B(n8017), .Z(n8199) );
  NANDN U8277 ( .A(n8020), .B(n8019), .Z(n8024) );
  OR U8278 ( .A(n8022), .B(n8021), .Z(n8023) );
  NAND U8279 ( .A(n8024), .B(n8023), .Z(n8198) );
  XNOR U8280 ( .A(n8199), .B(n8198), .Z(n8200) );
  OR U8281 ( .A(n8026), .B(n8025), .Z(n8030) );
  NANDN U8282 ( .A(n8028), .B(n8027), .Z(n8029) );
  NAND U8283 ( .A(n8030), .B(n8029), .Z(n8201) );
  XOR U8284 ( .A(n8113), .B(n8114), .Z(n8116) );
  OR U8285 ( .A(n8032), .B(n8031), .Z(n8036) );
  OR U8286 ( .A(n8034), .B(n8033), .Z(n8035) );
  NAND U8287 ( .A(n8036), .B(n8035), .Z(n8115) );
  XNOR U8288 ( .A(n8116), .B(n8115), .Z(n8068) );
  XNOR U8289 ( .A(n8067), .B(n8068), .Z(n8069) );
  XNOR U8290 ( .A(n8070), .B(n8069), .Z(n8207) );
  NANDN U8291 ( .A(n8038), .B(n8037), .Z(n8042) );
  NANDN U8292 ( .A(n8040), .B(n8039), .Z(n8041) );
  NAND U8293 ( .A(n8042), .B(n8041), .Z(n8205) );
  OR U8294 ( .A(n8044), .B(n8043), .Z(n8048) );
  OR U8295 ( .A(n8046), .B(n8045), .Z(n8047) );
  AND U8296 ( .A(n8048), .B(n8047), .Z(n8204) );
  XOR U8297 ( .A(n8205), .B(n8204), .Z(n8206) );
  XNOR U8298 ( .A(n8207), .B(n8206), .Z(n8061) );
  NANDN U8299 ( .A(n8050), .B(n8049), .Z(n8054) );
  NANDN U8300 ( .A(n8052), .B(n8051), .Z(n8053) );
  NAND U8301 ( .A(n8054), .B(n8053), .Z(n8062) );
  XOR U8302 ( .A(n8061), .B(n8062), .Z(n8063) );
  XNOR U8303 ( .A(n8064), .B(n8063), .Z(n8058) );
  XOR U8304 ( .A(n8057), .B(n8058), .Z(N187) );
  NANDN U8305 ( .A(n8056), .B(n8055), .Z(n8060) );
  NANDN U8306 ( .A(n8058), .B(n8057), .Z(n8059) );
  NAND U8307 ( .A(n8060), .B(n8059), .Z(n8210) );
  OR U8308 ( .A(n8062), .B(n8061), .Z(n8066) );
  NANDN U8309 ( .A(n8064), .B(n8063), .Z(n8065) );
  NAND U8310 ( .A(n8066), .B(n8065), .Z(n8211) );
  XNOR U8311 ( .A(n8210), .B(n8211), .Z(n8212) );
  OR U8312 ( .A(n8068), .B(n8067), .Z(n8072) );
  OR U8313 ( .A(n8070), .B(n8069), .Z(n8071) );
  AND U8314 ( .A(n8072), .B(n8071), .Z(n8216) );
  OR U8315 ( .A(n8074), .B(n8073), .Z(n8078) );
  OR U8316 ( .A(n8076), .B(n8075), .Z(n8077) );
  NAND U8317 ( .A(n8078), .B(n8077), .Z(n8349) );
  NANDN U8318 ( .A(n8084), .B(n8083), .Z(n8088) );
  NANDN U8319 ( .A(n8086), .B(n8085), .Z(n8087) );
  NAND U8320 ( .A(n8088), .B(n8087), .Z(n8325) );
  NANDN U8321 ( .A(n8090), .B(n8089), .Z(n8094) );
  NAND U8322 ( .A(n8092), .B(n8091), .Z(n8093) );
  NAND U8323 ( .A(n8094), .B(n8093), .Z(n8279) );
  NANDN U8324 ( .A(n8096), .B(n8095), .Z(n8100) );
  NAND U8325 ( .A(n8098), .B(n8097), .Z(n8099) );
  NAND U8326 ( .A(n8100), .B(n8099), .Z(n8280) );
  XNOR U8327 ( .A(n8279), .B(n8280), .Z(n8281) );
  NANDN U8328 ( .A(n8102), .B(n8101), .Z(n8106) );
  OR U8329 ( .A(n8104), .B(n8103), .Z(n8105) );
  NAND U8330 ( .A(n8106), .B(n8105), .Z(n8275) );
  NAND U8331 ( .A(x[73]), .B(y[274]), .Z(n8237) );
  NAND U8332 ( .A(y[265]), .B(x[82]), .Z(n8235) );
  NAND U8333 ( .A(y[262]), .B(x[85]), .Z(n8236) );
  XNOR U8334 ( .A(n8235), .B(n8236), .Z(n8238) );
  XOR U8335 ( .A(n8237), .B(n8238), .Z(n8276) );
  XNOR U8336 ( .A(n8275), .B(n8276), .Z(n8277) );
  NANDN U8337 ( .A(n45), .B(y[283]), .Z(n8225) );
  AND U8338 ( .A(y[257]), .B(x[90]), .Z(n8234) );
  XOR U8339 ( .A(o[91]), .B(n8234), .Z(n8223) );
  NANDN U8340 ( .A(n8872), .B(x[91]), .Z(n8222) );
  XNOR U8341 ( .A(n8223), .B(n8222), .Z(n8224) );
  XNOR U8342 ( .A(n8225), .B(n8224), .Z(n8278) );
  XOR U8343 ( .A(n8277), .B(n8278), .Z(n8282) );
  XNOR U8344 ( .A(n8281), .B(n8282), .Z(n8324) );
  XOR U8345 ( .A(n8325), .B(n8324), .Z(n8327) );
  XNOR U8346 ( .A(n8326), .B(n8327), .Z(n8348) );
  XNOR U8347 ( .A(n8349), .B(n8348), .Z(n8351) );
  OR U8348 ( .A(n8108), .B(n8107), .Z(n8112) );
  OR U8349 ( .A(n8110), .B(n8109), .Z(n8111) );
  NAND U8350 ( .A(n8112), .B(n8111), .Z(n8350) );
  XNOR U8351 ( .A(n8351), .B(n8350), .Z(n8360) );
  NANDN U8352 ( .A(n8114), .B(n8113), .Z(n8118) );
  OR U8353 ( .A(n8116), .B(n8115), .Z(n8117) );
  NAND U8354 ( .A(n8118), .B(n8117), .Z(n8361) );
  NAND U8355 ( .A(n8120), .B(n8119), .Z(n8124) );
  NANDN U8356 ( .A(n8122), .B(n8121), .Z(n8123) );
  NAND U8357 ( .A(n8124), .B(n8123), .Z(n8321) );
  OR U8358 ( .A(n8126), .B(n8125), .Z(n8130) );
  OR U8359 ( .A(n8128), .B(n8127), .Z(n8129) );
  NAND U8360 ( .A(n8130), .B(n8129), .Z(n8319) );
  AND U8361 ( .A(y[271]), .B(x[76]), .Z(n8293) );
  AND U8362 ( .A(y[270]), .B(x[77]), .Z(n8294) );
  XNOR U8363 ( .A(n8293), .B(n8294), .Z(n8296) );
  NANDN U8364 ( .A(n8884), .B(x[75]), .Z(n8308) );
  NANDN U8365 ( .A(n8890), .B(y[267]), .Z(n8305) );
  XNOR U8366 ( .A(n8306), .B(n8305), .Z(n8307) );
  XNOR U8367 ( .A(n8308), .B(n8307), .Z(n8295) );
  XNOR U8368 ( .A(n8296), .B(n8295), .Z(n8259) );
  AND U8369 ( .A(y[280]), .B(x[67]), .Z(n8301) );
  AND U8370 ( .A(y[281]), .B(x[66]), .Z(n8300) );
  XNOR U8371 ( .A(n8299), .B(n8300), .Z(n8302) );
  XOR U8372 ( .A(n8301), .B(n8302), .Z(n8257) );
  NANDN U8373 ( .A(n8703), .B(x[70]), .Z(n8249) );
  AND U8374 ( .A(y[258]), .B(x[89]), .Z(n8248) );
  NANDN U8375 ( .A(n8927), .B(x[83]), .Z(n8247) );
  XOR U8376 ( .A(n8248), .B(n8247), .Z(n8250) );
  XNOR U8377 ( .A(n8249), .B(n8250), .Z(n8258) );
  XNOR U8378 ( .A(n8257), .B(n8258), .Z(n8260) );
  XNOR U8379 ( .A(n8259), .B(n8260), .Z(n8286) );
  NAND U8380 ( .A(n8132), .B(n8131), .Z(n8136) );
  NANDN U8381 ( .A(n8134), .B(n8133), .Z(n8135) );
  NAND U8382 ( .A(n8136), .B(n8135), .Z(n8283) );
  NANDN U8383 ( .A(n8138), .B(n8137), .Z(n8142) );
  NAND U8384 ( .A(n8140), .B(n8139), .Z(n8141) );
  NAND U8385 ( .A(n8142), .B(n8141), .Z(n8284) );
  XNOR U8386 ( .A(n8283), .B(n8284), .Z(n8285) );
  XOR U8387 ( .A(n8286), .B(n8285), .Z(n8318) );
  XNOR U8388 ( .A(n8319), .B(n8318), .Z(n8320) );
  XNOR U8389 ( .A(n8321), .B(n8320), .Z(n8342) );
  NANDN U8390 ( .A(n8144), .B(n8143), .Z(n8148) );
  OR U8391 ( .A(n8146), .B(n8145), .Z(n8147) );
  NAND U8392 ( .A(n8148), .B(n8147), .Z(n8343) );
  XOR U8393 ( .A(n8342), .B(n8343), .Z(n8345) );
  OR U8394 ( .A(n8150), .B(n8149), .Z(n8154) );
  OR U8395 ( .A(n8152), .B(n8151), .Z(n8153) );
  AND U8396 ( .A(n8154), .B(n8153), .Z(n8344) );
  XNOR U8397 ( .A(n8345), .B(n8344), .Z(n8362) );
  XOR U8398 ( .A(n8363), .B(n8362), .Z(n8357) );
  OR U8399 ( .A(n8156), .B(n8155), .Z(n8160) );
  NANDN U8400 ( .A(n8158), .B(n8157), .Z(n8159) );
  AND U8401 ( .A(n8160), .B(n8159), .Z(n8354) );
  NANDN U8402 ( .A(n8162), .B(n8161), .Z(n8166) );
  NANDN U8403 ( .A(n8164), .B(n8163), .Z(n8165) );
  NAND U8404 ( .A(n8166), .B(n8165), .Z(n8265) );
  AND U8405 ( .A(y[261]), .B(x[86]), .Z(n8313) );
  AND U8406 ( .A(y[260]), .B(x[87]), .Z(n8311) );
  AND U8407 ( .A(y[275]), .B(x[72]), .Z(n8312) );
  XNOR U8408 ( .A(n8311), .B(n8312), .Z(n8314) );
  XOR U8409 ( .A(n8313), .B(n8314), .Z(n8263) );
  NANDN U8410 ( .A(n8900), .B(x[71]), .Z(n8243) );
  NANDN U8411 ( .A(n8881), .B(x[88]), .Z(n8241) );
  XOR U8412 ( .A(n8242), .B(n8241), .Z(n8244) );
  XNOR U8413 ( .A(n8243), .B(n8244), .Z(n8264) );
  XNOR U8414 ( .A(n8263), .B(n8264), .Z(n8266) );
  XNOR U8415 ( .A(n8265), .B(n8266), .Z(n8336) );
  NAND U8416 ( .A(n8168), .B(n8167), .Z(n8172) );
  NANDN U8417 ( .A(n8170), .B(n8169), .Z(n8171) );
  NAND U8418 ( .A(n8172), .B(n8171), .Z(n8254) );
  NANDN U8419 ( .A(n8174), .B(n8173), .Z(n8178) );
  NANDN U8420 ( .A(n8176), .B(n8175), .Z(n8177) );
  AND U8421 ( .A(n8178), .B(n8177), .Z(n8253) );
  XNOR U8422 ( .A(n8254), .B(n8253), .Z(n8256) );
  ANDN U8423 ( .B(o[90]), .A(n8179), .Z(n8287) );
  AND U8424 ( .A(y[282]), .B(x[65]), .Z(n8288) );
  XNOR U8425 ( .A(n8287), .B(n8288), .Z(n8290) );
  XNOR U8426 ( .A(n8289), .B(n8290), .Z(n8269) );
  NANDN U8427 ( .A(n8626), .B(y[266]), .Z(n8229) );
  ANDN U8428 ( .B(y[279]), .A(n49), .Z(n8228) );
  XOR U8429 ( .A(n8229), .B(n8228), .Z(n8231) );
  ANDN U8430 ( .B(x[69]), .A(n8613), .Z(n8230) );
  XOR U8431 ( .A(n8231), .B(n8230), .Z(n8270) );
  XOR U8432 ( .A(n8269), .B(n8270), .Z(n8272) );
  NAND U8433 ( .A(n8181), .B(n8180), .Z(n8185) );
  NANDN U8434 ( .A(n8183), .B(n8182), .Z(n8184) );
  NAND U8435 ( .A(n8185), .B(n8184), .Z(n8271) );
  XOR U8436 ( .A(n8272), .B(n8271), .Z(n8255) );
  XOR U8437 ( .A(n8256), .B(n8255), .Z(n8337) );
  XNOR U8438 ( .A(n8336), .B(n8337), .Z(n8339) );
  OR U8439 ( .A(n8187), .B(n8186), .Z(n8191) );
  OR U8440 ( .A(n8189), .B(n8188), .Z(n8190) );
  AND U8441 ( .A(n8191), .B(n8190), .Z(n8338) );
  XOR U8442 ( .A(n8339), .B(n8338), .Z(n8330) );
  OR U8443 ( .A(n8193), .B(n8192), .Z(n8197) );
  OR U8444 ( .A(n8195), .B(n8194), .Z(n8196) );
  AND U8445 ( .A(n8197), .B(n8196), .Z(n8331) );
  XNOR U8446 ( .A(n8330), .B(n8331), .Z(n8333) );
  OR U8447 ( .A(n8199), .B(n8198), .Z(n8203) );
  OR U8448 ( .A(n8201), .B(n8200), .Z(n8202) );
  NAND U8449 ( .A(n8203), .B(n8202), .Z(n8332) );
  XOR U8450 ( .A(n8333), .B(n8332), .Z(n8355) );
  XOR U8451 ( .A(n8354), .B(n8355), .Z(n8356) );
  XOR U8452 ( .A(n8357), .B(n8356), .Z(n8217) );
  XNOR U8453 ( .A(n8216), .B(n8217), .Z(n8218) );
  OR U8454 ( .A(n8205), .B(n8204), .Z(n8209) );
  NANDN U8455 ( .A(n8207), .B(n8206), .Z(n8208) );
  AND U8456 ( .A(n8209), .B(n8208), .Z(n8219) );
  XOR U8457 ( .A(n8212), .B(n8213), .Z(N188) );
  NANDN U8458 ( .A(n8211), .B(n8210), .Z(n8215) );
  NANDN U8459 ( .A(n8213), .B(n8212), .Z(n8214) );
  NAND U8460 ( .A(n8215), .B(n8214), .Z(n8366) );
  OR U8461 ( .A(n8217), .B(n8216), .Z(n8221) );
  OR U8462 ( .A(n8219), .B(n8218), .Z(n8220) );
  AND U8463 ( .A(n8221), .B(n8220), .Z(n8367) );
  XNOR U8464 ( .A(n8366), .B(n8367), .Z(n8368) );
  NANDN U8465 ( .A(n8223), .B(n8222), .Z(n8227) );
  NAND U8466 ( .A(n8225), .B(n8224), .Z(n8226) );
  AND U8467 ( .A(n8227), .B(n8226), .Z(n8494) );
  NANDN U8468 ( .A(n8229), .B(n8228), .Z(n8233) );
  NANDN U8469 ( .A(n8231), .B(n8230), .Z(n8232) );
  NAND U8470 ( .A(n8233), .B(n8232), .Z(n8495) );
  XOR U8471 ( .A(n8494), .B(n8495), .Z(n8497) );
  AND U8472 ( .A(n8234), .B(o[91]), .Z(n8464) );
  AND U8473 ( .A(y[256]), .B(x[92]), .Z(n8465) );
  XNOR U8474 ( .A(n8464), .B(n8465), .Z(n8467) );
  AND U8475 ( .A(y[284]), .B(x[64]), .Z(n8466) );
  XNOR U8476 ( .A(n8467), .B(n8466), .Z(n8449) );
  NAND U8477 ( .A(n8236), .B(n8235), .Z(n8240) );
  NANDN U8478 ( .A(n8238), .B(n8237), .Z(n8239) );
  AND U8479 ( .A(n8240), .B(n8239), .Z(n8446) );
  AND U8480 ( .A(y[275]), .B(x[73]), .Z(n8458) );
  AND U8481 ( .A(y[276]), .B(x[72]), .Z(n8459) );
  XNOR U8482 ( .A(n8458), .B(n8459), .Z(n8461) );
  AND U8483 ( .A(y[274]), .B(x[74]), .Z(n8460) );
  XNOR U8484 ( .A(n8461), .B(n8460), .Z(n8447) );
  XNOR U8485 ( .A(n8446), .B(n8447), .Z(n8448) );
  XNOR U8486 ( .A(n8497), .B(n8496), .Z(n8479) );
  AND U8487 ( .A(y[283]), .B(x[65]), .Z(n8390) );
  AND U8488 ( .A(y[259]), .B(x[89]), .Z(n8391) );
  XNOR U8489 ( .A(n8390), .B(n8391), .Z(n8393) );
  XNOR U8490 ( .A(n8392), .B(n8393), .Z(n8490) );
  AND U8491 ( .A(y[268]), .B(x[80]), .Z(n8398) );
  AND U8492 ( .A(y[282]), .B(x[66]), .Z(n8396) );
  AND U8493 ( .A(y[260]), .B(x[88]), .Z(n8397) );
  XNOR U8494 ( .A(n8396), .B(n8397), .Z(n8399) );
  XOR U8495 ( .A(n8398), .B(n8399), .Z(n8488) );
  NANDN U8496 ( .A(n8242), .B(n8241), .Z(n8246) );
  NANDN U8497 ( .A(n8244), .B(n8243), .Z(n8245) );
  NAND U8498 ( .A(n8246), .B(n8245), .Z(n8489) );
  XNOR U8499 ( .A(n8488), .B(n8489), .Z(n8491) );
  XNOR U8500 ( .A(n8490), .B(n8491), .Z(n8477) );
  AND U8501 ( .A(y[261]), .B(x[87]), .Z(n8428) );
  AND U8502 ( .A(y[281]), .B(x[67]), .Z(n8429) );
  XNOR U8503 ( .A(n8428), .B(n8429), .Z(n8431) );
  XOR U8504 ( .A(n8430), .B(n8431), .Z(n8502) );
  AND U8505 ( .A(y[279]), .B(x[69]), .Z(n8410) );
  AND U8506 ( .A(y[264]), .B(x[84]), .Z(n8408) );
  AND U8507 ( .A(y[263]), .B(x[85]), .Z(n8409) );
  XNOR U8508 ( .A(n8408), .B(n8409), .Z(n8411) );
  XOR U8509 ( .A(n8410), .B(n8411), .Z(n8500) );
  NANDN U8510 ( .A(n8248), .B(n8247), .Z(n8252) );
  NANDN U8511 ( .A(n8250), .B(n8249), .Z(n8251) );
  NAND U8512 ( .A(n8252), .B(n8251), .Z(n8501) );
  XNOR U8513 ( .A(n8500), .B(n8501), .Z(n8503) );
  XNOR U8514 ( .A(n8502), .B(n8503), .Z(n8476) );
  XNOR U8515 ( .A(n8477), .B(n8476), .Z(n8478) );
  XNOR U8516 ( .A(n8479), .B(n8478), .Z(n8528) );
  OR U8517 ( .A(n8258), .B(n8257), .Z(n8262) );
  NANDN U8518 ( .A(n8260), .B(n8259), .Z(n8261) );
  NAND U8519 ( .A(n8262), .B(n8261), .Z(n8513) );
  OR U8520 ( .A(n8264), .B(n8263), .Z(n8268) );
  NANDN U8521 ( .A(n8266), .B(n8265), .Z(n8267) );
  NAND U8522 ( .A(n8268), .B(n8267), .Z(n8512) );
  XOR U8523 ( .A(n8513), .B(n8512), .Z(n8514) );
  XNOR U8524 ( .A(n8515), .B(n8514), .Z(n8529) );
  XNOR U8525 ( .A(n8528), .B(n8529), .Z(n8531) );
  NANDN U8526 ( .A(n8270), .B(n8269), .Z(n8274) );
  OR U8527 ( .A(n8272), .B(n8271), .Z(n8273) );
  AND U8528 ( .A(n8274), .B(n8273), .Z(n8506) );
  XOR U8529 ( .A(n8506), .B(n8507), .Z(n8508) );
  XNOR U8530 ( .A(n8508), .B(n8509), .Z(n8521) );
  OR U8531 ( .A(n8288), .B(n8287), .Z(n8292) );
  OR U8532 ( .A(n8290), .B(n8289), .Z(n8291) );
  AND U8533 ( .A(n8292), .B(n8291), .Z(n8473) );
  OR U8534 ( .A(n8294), .B(n8293), .Z(n8298) );
  OR U8535 ( .A(n8296), .B(n8295), .Z(n8297) );
  AND U8536 ( .A(n8298), .B(n8297), .Z(n8470) );
  OR U8537 ( .A(n8300), .B(n8299), .Z(n8304) );
  OR U8538 ( .A(n8302), .B(n8301), .Z(n8303) );
  AND U8539 ( .A(n8304), .B(n8303), .Z(n8471) );
  XNOR U8540 ( .A(n8470), .B(n8471), .Z(n8472) );
  NANDN U8541 ( .A(n8901), .B(y[258]), .Z(n8435) );
  ANDN U8542 ( .B(x[79]), .A(n8815), .Z(n8434) );
  XNOR U8543 ( .A(n8435), .B(n8434), .Z(n8437) );
  NAND U8544 ( .A(x[91]), .B(y[257]), .Z(n8602) );
  XNOR U8545 ( .A(n8602), .B(o[92]), .Z(n8436) );
  XNOR U8546 ( .A(n8437), .B(n8436), .Z(n8425) );
  NANDN U8547 ( .A(n8306), .B(n8305), .Z(n8310) );
  NAND U8548 ( .A(n8308), .B(n8307), .Z(n8309) );
  NAND U8549 ( .A(n8310), .B(n8309), .Z(n8423) );
  NANDN U8550 ( .A(n8703), .B(x[71]), .Z(n8404) );
  AND U8551 ( .A(y[273]), .B(x[75]), .Z(n8403) );
  NANDN U8552 ( .A(n8884), .B(x[76]), .Z(n8402) );
  XOR U8553 ( .A(n8403), .B(n8402), .Z(n8405) );
  XNOR U8554 ( .A(n8404), .B(n8405), .Z(n8422) );
  XNOR U8555 ( .A(n8423), .B(n8422), .Z(n8424) );
  XNOR U8556 ( .A(n8425), .B(n8424), .Z(n8483) );
  OR U8557 ( .A(n8312), .B(n8311), .Z(n8316) );
  OR U8558 ( .A(n8314), .B(n8313), .Z(n8315) );
  AND U8559 ( .A(n8316), .B(n8315), .Z(n8440) );
  AND U8560 ( .A(y[278]), .B(x[70]), .Z(n8418) );
  AND U8561 ( .A(y[265]), .B(x[83]), .Z(n8417) );
  XOR U8562 ( .A(n8317), .B(n8417), .Z(n8419) );
  XNOR U8563 ( .A(n8418), .B(n8419), .Z(n8441) );
  XNOR U8564 ( .A(n8440), .B(n8441), .Z(n8442) );
  AND U8565 ( .A(y[267]), .B(x[81]), .Z(n8454) );
  AND U8566 ( .A(y[280]), .B(x[68]), .Z(n8452) );
  AND U8567 ( .A(y[262]), .B(x[86]), .Z(n8453) );
  XNOR U8568 ( .A(n8452), .B(n8453), .Z(n8455) );
  XNOR U8569 ( .A(n8454), .B(n8455), .Z(n8443) );
  XNOR U8570 ( .A(n8483), .B(n8482), .Z(n8484) );
  XNOR U8571 ( .A(n8485), .B(n8484), .Z(n8519) );
  XNOR U8572 ( .A(n8518), .B(n8519), .Z(n8520) );
  XNOR U8573 ( .A(n8521), .B(n8520), .Z(n8530) );
  XNOR U8574 ( .A(n8531), .B(n8530), .Z(n8527) );
  OR U8575 ( .A(n8319), .B(n8318), .Z(n8323) );
  OR U8576 ( .A(n8321), .B(n8320), .Z(n8322) );
  NAND U8577 ( .A(n8323), .B(n8322), .Z(n8524) );
  NANDN U8578 ( .A(n8325), .B(n8324), .Z(n8329) );
  NANDN U8579 ( .A(n8327), .B(n8326), .Z(n8328) );
  AND U8580 ( .A(n8329), .B(n8328), .Z(n8525) );
  XNOR U8581 ( .A(n8524), .B(n8525), .Z(n8526) );
  XOR U8582 ( .A(n8527), .B(n8526), .Z(n8384) );
  OR U8583 ( .A(n8331), .B(n8330), .Z(n8335) );
  OR U8584 ( .A(n8333), .B(n8332), .Z(n8334) );
  AND U8585 ( .A(n8335), .B(n8334), .Z(n8385) );
  XOR U8586 ( .A(n8384), .B(n8385), .Z(n8387) );
  OR U8587 ( .A(n8337), .B(n8336), .Z(n8341) );
  OR U8588 ( .A(n8339), .B(n8338), .Z(n8340) );
  AND U8589 ( .A(n8341), .B(n8340), .Z(n8381) );
  NANDN U8590 ( .A(n8343), .B(n8342), .Z(n8347) );
  OR U8591 ( .A(n8345), .B(n8344), .Z(n8346) );
  NAND U8592 ( .A(n8347), .B(n8346), .Z(n8379) );
  OR U8593 ( .A(n8349), .B(n8348), .Z(n8353) );
  OR U8594 ( .A(n8351), .B(n8350), .Z(n8352) );
  NAND U8595 ( .A(n8353), .B(n8352), .Z(n8378) );
  XOR U8596 ( .A(n8379), .B(n8378), .Z(n8380) );
  XNOR U8597 ( .A(n8381), .B(n8380), .Z(n8386) );
  XNOR U8598 ( .A(n8387), .B(n8386), .Z(n8372) );
  OR U8599 ( .A(n8355), .B(n8354), .Z(n8359) );
  NANDN U8600 ( .A(n8357), .B(n8356), .Z(n8358) );
  AND U8601 ( .A(n8359), .B(n8358), .Z(n8373) );
  XOR U8602 ( .A(n8372), .B(n8373), .Z(n8375) );
  OR U8603 ( .A(n8361), .B(n8360), .Z(n8365) );
  OR U8604 ( .A(n8363), .B(n8362), .Z(n8364) );
  NAND U8605 ( .A(n8365), .B(n8364), .Z(n8374) );
  XOR U8606 ( .A(n8375), .B(n8374), .Z(n8369) );
  XNOR U8607 ( .A(n8368), .B(n8369), .Z(N189) );
  NANDN U8608 ( .A(n8367), .B(n8366), .Z(n8371) );
  NAND U8609 ( .A(n8369), .B(n8368), .Z(n8370) );
  NAND U8610 ( .A(n8371), .B(n8370), .Z(n8534) );
  NANDN U8611 ( .A(n8373), .B(n8372), .Z(n8377) );
  OR U8612 ( .A(n8375), .B(n8374), .Z(n8376) );
  AND U8613 ( .A(n8377), .B(n8376), .Z(n8535) );
  XNOR U8614 ( .A(n8534), .B(n8535), .Z(n8536) );
  OR U8615 ( .A(n8379), .B(n8378), .Z(n8383) );
  NANDN U8616 ( .A(n8381), .B(n8380), .Z(n8382) );
  AND U8617 ( .A(n8383), .B(n8382), .Z(n8540) );
  NANDN U8618 ( .A(n8385), .B(n8384), .Z(n8389) );
  OR U8619 ( .A(n8387), .B(n8386), .Z(n8388) );
  NAND U8620 ( .A(n8389), .B(n8388), .Z(n8541) );
  XOR U8621 ( .A(n8540), .B(n8541), .Z(n8542) );
  OR U8622 ( .A(n8391), .B(n8390), .Z(n8395) );
  OR U8623 ( .A(n8393), .B(n8392), .Z(n8394) );
  AND U8624 ( .A(n8395), .B(n8394), .Z(n8686) );
  OR U8625 ( .A(n8397), .B(n8396), .Z(n8401) );
  OR U8626 ( .A(n8399), .B(n8398), .Z(n8400) );
  AND U8627 ( .A(n8401), .B(n8400), .Z(n8683) );
  ANDN U8628 ( .B(x[87]), .A(n8655), .Z(n8614) );
  IV U8629 ( .A(n8614), .Z(n8945) );
  AND U8630 ( .A(y[261]), .B(x[88]), .Z(n8615) );
  XOR U8631 ( .A(n8945), .B(n8615), .Z(n8617) );
  AND U8632 ( .A(y[272]), .B(x[77]), .Z(n8616) );
  XNOR U8633 ( .A(n8617), .B(n8616), .Z(n8585) );
  NANDN U8634 ( .A(n8403), .B(n8402), .Z(n8407) );
  NANDN U8635 ( .A(n8405), .B(n8404), .Z(n8406) );
  AND U8636 ( .A(n8407), .B(n8406), .Z(n8583) );
  AND U8637 ( .A(y[274]), .B(x[75]), .Z(n8607) );
  AND U8638 ( .A(y[268]), .B(x[81]), .Z(n8608) );
  XNOR U8639 ( .A(n8607), .B(n8608), .Z(n8610) );
  AND U8640 ( .A(y[282]), .B(x[67]), .Z(n8609) );
  XOR U8641 ( .A(n8610), .B(n8609), .Z(n8582) );
  XOR U8642 ( .A(n8583), .B(n8582), .Z(n8584) );
  XNOR U8643 ( .A(n8585), .B(n8584), .Z(n8684) );
  XNOR U8644 ( .A(n8683), .B(n8684), .Z(n8685) );
  AND U8645 ( .A(y[267]), .B(x[82]), .Z(n8594) );
  AND U8646 ( .A(y[266]), .B(x[83]), .Z(n8595) );
  XNOR U8647 ( .A(n8594), .B(n8595), .Z(n8597) );
  AND U8648 ( .A(y[283]), .B(x[66]), .Z(n8596) );
  XNOR U8649 ( .A(n8597), .B(n8596), .Z(n8633) );
  OR U8650 ( .A(n8409), .B(n8408), .Z(n8413) );
  OR U8651 ( .A(n8411), .B(n8410), .Z(n8412) );
  AND U8652 ( .A(n8413), .B(n8412), .Z(n8631) );
  NAND U8653 ( .A(y[257]), .B(o[92]), .Z(n8414) );
  XNOR U8654 ( .A(y[258]), .B(n8414), .Z(n8415) );
  NAND U8655 ( .A(x[91]), .B(n8415), .Z(n8601) );
  AND U8656 ( .A(y[269]), .B(x[80]), .Z(n8600) );
  XOR U8657 ( .A(n8601), .B(n8600), .Z(n8630) );
  XOR U8658 ( .A(n8631), .B(n8630), .Z(n8632) );
  XNOR U8659 ( .A(n8633), .B(n8632), .Z(n8666) );
  OR U8660 ( .A(n8417), .B(n8416), .Z(n8421) );
  OR U8661 ( .A(n8419), .B(n8418), .Z(n8420) );
  NAND U8662 ( .A(n8421), .B(n8420), .Z(n8692) );
  AND U8663 ( .A(y[257]), .B(x[92]), .Z(n8653) );
  XOR U8664 ( .A(o[93]), .B(n8653), .Z(n8706) );
  AND U8665 ( .A(y[256]), .B(x[93]), .Z(n8707) );
  XNOR U8666 ( .A(n8706), .B(n8707), .Z(n8709) );
  AND U8667 ( .A(y[285]), .B(x[64]), .Z(n8708) );
  XOR U8668 ( .A(n8709), .B(n8708), .Z(n8689) );
  AND U8669 ( .A(y[260]), .B(x[89]), .Z(n8636) );
  AND U8670 ( .A(y[259]), .B(x[90]), .Z(n8637) );
  XNOR U8671 ( .A(n8636), .B(n8637), .Z(n8639) );
  AND U8672 ( .A(y[271]), .B(x[78]), .Z(n8638) );
  XOR U8673 ( .A(n8639), .B(n8638), .Z(n8690) );
  XNOR U8674 ( .A(n8689), .B(n8690), .Z(n8691) );
  XOR U8675 ( .A(n8692), .B(n8691), .Z(n8665) );
  XNOR U8676 ( .A(n8666), .B(n8665), .Z(n8667) );
  XOR U8677 ( .A(n8668), .B(n8667), .Z(n8659) );
  OR U8678 ( .A(n8423), .B(n8422), .Z(n8427) );
  OR U8679 ( .A(n8425), .B(n8424), .Z(n8426) );
  AND U8680 ( .A(n8427), .B(n8426), .Z(n8660) );
  XNOR U8681 ( .A(n8659), .B(n8660), .Z(n8662) );
  OR U8682 ( .A(n8429), .B(n8428), .Z(n8433) );
  OR U8683 ( .A(n8431), .B(n8430), .Z(n8432) );
  AND U8684 ( .A(n8433), .B(n8432), .Z(n8576) );
  NANDN U8685 ( .A(n8435), .B(n8434), .Z(n8439) );
  NAND U8686 ( .A(n8437), .B(n8436), .Z(n8438) );
  NAND U8687 ( .A(n8439), .B(n8438), .Z(n8577) );
  XNOR U8688 ( .A(n8576), .B(n8577), .Z(n8578) );
  AND U8689 ( .A(y[277]), .B(x[72]), .Z(n8620) );
  AND U8690 ( .A(y[278]), .B(x[71]), .Z(n8621) );
  XNOR U8691 ( .A(n8620), .B(n8621), .Z(n8623) );
  AND U8692 ( .A(y[279]), .B(x[70]), .Z(n8622) );
  XNOR U8693 ( .A(n8623), .B(n8622), .Z(n8698) );
  ANDN U8694 ( .B(x[73]), .A(n8900), .Z(n8695) );
  IV U8695 ( .A(n8695), .Z(n8804) );
  AND U8696 ( .A(y[280]), .B(x[69]), .Z(n8588) );
  AND U8697 ( .A(y[275]), .B(x[74]), .Z(n8589) );
  XNOR U8698 ( .A(n8588), .B(n8589), .Z(n8591) );
  AND U8699 ( .A(y[281]), .B(x[68]), .Z(n8590) );
  XNOR U8700 ( .A(n8591), .B(n8590), .Z(n8696) );
  XOR U8701 ( .A(n8804), .B(n8696), .Z(n8697) );
  XNOR U8702 ( .A(n8698), .B(n8697), .Z(n8579) );
  XOR U8703 ( .A(n8662), .B(n8661), .Z(n8673) );
  OR U8704 ( .A(n8441), .B(n8440), .Z(n8445) );
  OR U8705 ( .A(n8443), .B(n8442), .Z(n8444) );
  AND U8706 ( .A(n8445), .B(n8444), .Z(n8671) );
  OR U8707 ( .A(n8447), .B(n8446), .Z(n8451) );
  OR U8708 ( .A(n8449), .B(n8448), .Z(n8450) );
  AND U8709 ( .A(n8451), .B(n8450), .Z(n8718) );
  OR U8710 ( .A(n8453), .B(n8452), .Z(n8457) );
  OR U8711 ( .A(n8455), .B(n8454), .Z(n8456) );
  AND U8712 ( .A(n8457), .B(n8456), .Z(n8712) );
  ANDN U8713 ( .B(x[76]), .A(n8904), .Z(n8644) );
  IV U8714 ( .A(n8644), .Z(n8838) );
  AND U8715 ( .A(y[263]), .B(x[86]), .Z(n8642) );
  AND U8716 ( .A(y[284]), .B(x[65]), .Z(n8643) );
  XNOR U8717 ( .A(n8642), .B(n8643), .Z(n8645) );
  XOR U8718 ( .A(n8838), .B(n8645), .Z(n8680) );
  OR U8719 ( .A(n8459), .B(n8458), .Z(n8463) );
  OR U8720 ( .A(n8461), .B(n8460), .Z(n8462) );
  AND U8721 ( .A(n8463), .B(n8462), .Z(n8677) );
  NANDN U8722 ( .A(n8861), .B(x[79]), .Z(n8650) );
  AND U8723 ( .A(y[265]), .B(x[84]), .Z(n8648) );
  ANDN U8724 ( .B(x[85]), .A(n8927), .Z(n8965) );
  XOR U8725 ( .A(n8648), .B(n8965), .Z(n8649) );
  XNOR U8726 ( .A(n8650), .B(n8649), .Z(n8678) );
  XNOR U8727 ( .A(n8677), .B(n8678), .Z(n8679) );
  XNOR U8728 ( .A(n8680), .B(n8679), .Z(n8713) );
  XNOR U8729 ( .A(n8712), .B(n8713), .Z(n8714) );
  OR U8730 ( .A(n8465), .B(n8464), .Z(n8469) );
  OR U8731 ( .A(n8467), .B(n8466), .Z(n8468) );
  AND U8732 ( .A(n8469), .B(n8468), .Z(n8715) );
  XNOR U8733 ( .A(n8718), .B(n8719), .Z(n8721) );
  OR U8734 ( .A(n8471), .B(n8470), .Z(n8475) );
  OR U8735 ( .A(n8473), .B(n8472), .Z(n8474) );
  AND U8736 ( .A(n8475), .B(n8474), .Z(n8720) );
  XNOR U8737 ( .A(n8721), .B(n8720), .Z(n8672) );
  XNOR U8738 ( .A(n8671), .B(n8672), .Z(n8674) );
  XOR U8739 ( .A(n8673), .B(n8674), .Z(n8566) );
  NANDN U8740 ( .A(n8477), .B(n8476), .Z(n8481) );
  NANDN U8741 ( .A(n8479), .B(n8478), .Z(n8480) );
  AND U8742 ( .A(n8481), .B(n8480), .Z(n8554) );
  NAND U8743 ( .A(n8483), .B(n8482), .Z(n8487) );
  OR U8744 ( .A(n8485), .B(n8484), .Z(n8486) );
  NAND U8745 ( .A(n8487), .B(n8486), .Z(n8559) );
  OR U8746 ( .A(n8489), .B(n8488), .Z(n8493) );
  NANDN U8747 ( .A(n8491), .B(n8490), .Z(n8492) );
  NAND U8748 ( .A(n8493), .B(n8492), .Z(n8573) );
  OR U8749 ( .A(n8495), .B(n8494), .Z(n8499) );
  NAND U8750 ( .A(n8497), .B(n8496), .Z(n8498) );
  AND U8751 ( .A(n8499), .B(n8498), .Z(n8570) );
  OR U8752 ( .A(n8501), .B(n8500), .Z(n8505) );
  OR U8753 ( .A(n8503), .B(n8502), .Z(n8504) );
  NAND U8754 ( .A(n8505), .B(n8504), .Z(n8571) );
  XNOR U8755 ( .A(n8570), .B(n8571), .Z(n8572) );
  XOR U8756 ( .A(n8573), .B(n8572), .Z(n8558) );
  XNOR U8757 ( .A(n8559), .B(n8558), .Z(n8561) );
  OR U8758 ( .A(n8507), .B(n8506), .Z(n8511) );
  NANDN U8759 ( .A(n8509), .B(n8508), .Z(n8510) );
  AND U8760 ( .A(n8511), .B(n8510), .Z(n8560) );
  XOR U8761 ( .A(n8561), .B(n8560), .Z(n8552) );
  OR U8762 ( .A(n8513), .B(n8512), .Z(n8517) );
  NANDN U8763 ( .A(n8515), .B(n8514), .Z(n8516) );
  AND U8764 ( .A(n8517), .B(n8516), .Z(n8553) );
  XNOR U8765 ( .A(n8552), .B(n8553), .Z(n8555) );
  XOR U8766 ( .A(n8554), .B(n8555), .Z(n8564) );
  OR U8767 ( .A(n8519), .B(n8518), .Z(n8523) );
  OR U8768 ( .A(n8521), .B(n8520), .Z(n8522) );
  NAND U8769 ( .A(n8523), .B(n8522), .Z(n8565) );
  XNOR U8770 ( .A(n8564), .B(n8565), .Z(n8567) );
  XOR U8771 ( .A(n8566), .B(n8567), .Z(n8549) );
  OR U8772 ( .A(n8529), .B(n8528), .Z(n8533) );
  NANDN U8773 ( .A(n8531), .B(n8530), .Z(n8532) );
  NAND U8774 ( .A(n8533), .B(n8532), .Z(n8547) );
  XNOR U8775 ( .A(n8546), .B(n8547), .Z(n8548) );
  XOR U8776 ( .A(n8549), .B(n8548), .Z(n8543) );
  XOR U8777 ( .A(n8542), .B(n8543), .Z(n8537) );
  XOR U8778 ( .A(n8536), .B(n8537), .Z(N190) );
  NANDN U8779 ( .A(n8535), .B(n8534), .Z(n8539) );
  NANDN U8780 ( .A(n8537), .B(n8536), .Z(n8538) );
  AND U8781 ( .A(n8539), .B(n8538), .Z(n8726) );
  OR U8782 ( .A(n8541), .B(n8540), .Z(n8545) );
  NANDN U8783 ( .A(n8543), .B(n8542), .Z(n8544) );
  AND U8784 ( .A(n8545), .B(n8544), .Z(n8727) );
  XNOR U8785 ( .A(n8726), .B(n8727), .Z(n8725) );
  NANDN U8786 ( .A(n8547), .B(n8546), .Z(n8551) );
  NANDN U8787 ( .A(n8549), .B(n8548), .Z(n8550) );
  AND U8788 ( .A(n8551), .B(n8550), .Z(n9027) );
  OR U8789 ( .A(n8553), .B(n8552), .Z(n8557) );
  OR U8790 ( .A(n8555), .B(n8554), .Z(n8556) );
  NAND U8791 ( .A(n8557), .B(n8556), .Z(n9036) );
  OR U8792 ( .A(n8559), .B(n8558), .Z(n8563) );
  OR U8793 ( .A(n8561), .B(n8560), .Z(n8562) );
  AND U8794 ( .A(n8563), .B(n8562), .Z(n9035) );
  XOR U8795 ( .A(n9036), .B(n9035), .Z(n9033) );
  OR U8796 ( .A(n8565), .B(n8564), .Z(n8569) );
  OR U8797 ( .A(n8567), .B(n8566), .Z(n8568) );
  AND U8798 ( .A(n8569), .B(n8568), .Z(n9034) );
  XNOR U8799 ( .A(n9033), .B(n9034), .Z(n9029) );
  OR U8800 ( .A(n8571), .B(n8570), .Z(n8575) );
  OR U8801 ( .A(n8573), .B(n8572), .Z(n8574) );
  NAND U8802 ( .A(n8575), .B(n8574), .Z(n8733) );
  OR U8803 ( .A(n8577), .B(n8576), .Z(n8581) );
  OR U8804 ( .A(n8579), .B(n8578), .Z(n8580) );
  AND U8805 ( .A(n8581), .B(n8580), .Z(n8742) );
  NANDN U8806 ( .A(n8583), .B(n8582), .Z(n8587) );
  OR U8807 ( .A(n8585), .B(n8584), .Z(n8586) );
  AND U8808 ( .A(n8587), .B(n8586), .Z(n8744) );
  OR U8809 ( .A(n8589), .B(n8588), .Z(n8593) );
  OR U8810 ( .A(n8591), .B(n8590), .Z(n8592) );
  AND U8811 ( .A(n8593), .B(n8592), .Z(n8769) );
  NANDN U8812 ( .A(n51), .B(y[280]), .Z(n8842) );
  NANDN U8813 ( .A(n50), .B(y[281]), .Z(n8844) );
  NANDN U8814 ( .A(n8824), .B(y[267]), .Z(n8843) );
  XNOR U8815 ( .A(n8844), .B(n8843), .Z(n8841) );
  XNOR U8816 ( .A(n8842), .B(n8841), .Z(n8788) );
  OR U8817 ( .A(n8595), .B(n8594), .Z(n8599) );
  OR U8818 ( .A(n8597), .B(n8596), .Z(n8598) );
  AND U8819 ( .A(n8599), .B(n8598), .Z(n8790) );
  NANDN U8820 ( .A(n49), .B(y[282]), .Z(n8950) );
  NANDN U8821 ( .A(n48), .B(y[283]), .Z(n8952) );
  ANDN U8822 ( .B(y[268]), .A(n61), .Z(n8951) );
  XNOR U8823 ( .A(n8952), .B(n8951), .Z(n8949) );
  XNOR U8824 ( .A(n8950), .B(n8949), .Z(n8791) );
  XOR U8825 ( .A(n8790), .B(n8791), .Z(n8789) );
  XNOR U8826 ( .A(n8788), .B(n8789), .Z(n8768) );
  XNOR U8827 ( .A(n8769), .B(n8768), .Z(n8771) );
  OR U8828 ( .A(n8601), .B(n8600), .Z(n8606) );
  NANDN U8829 ( .A(n8602), .B(o[92]), .Z(n8604) );
  NAND U8830 ( .A(y[258]), .B(x[91]), .Z(n8603) );
  AND U8831 ( .A(n8604), .B(n8603), .Z(n8605) );
  ANDN U8832 ( .B(n8606), .A(n8605), .Z(n8770) );
  XNOR U8833 ( .A(n8744), .B(n8745), .Z(n8743) );
  XNOR U8834 ( .A(n8742), .B(n8743), .Z(n9018) );
  OR U8835 ( .A(n8608), .B(n8607), .Z(n8612) );
  OR U8836 ( .A(n8610), .B(n8609), .Z(n8611) );
  NAND U8837 ( .A(n8612), .B(n8611), .Z(n8797) );
  NANDN U8838 ( .A(n8885), .B(y[266]), .Z(n8920) );
  ANDN U8839 ( .B(x[78]), .A(n8884), .Z(n8919) );
  XOR U8840 ( .A(n8920), .B(n8919), .Z(n8918) );
  ANDN U8841 ( .B(x[72]), .A(n8613), .Z(n8917) );
  XOR U8842 ( .A(n8918), .B(n8917), .Z(n8799) );
  NANDN U8843 ( .A(n8872), .B(x[94]), .Z(n8810) );
  NANDN U8844 ( .A(n8893), .B(y[257]), .Z(n8862) );
  XNOR U8845 ( .A(o[94]), .B(n8862), .Z(n8809) );
  XOR U8846 ( .A(n8810), .B(n8809), .Z(n8808) );
  ANDN U8847 ( .B(y[286]), .A(n45), .Z(n8807) );
  XOR U8848 ( .A(n8808), .B(n8807), .Z(n8798) );
  XOR U8849 ( .A(n8797), .B(n8796), .Z(n8752) );
  OR U8850 ( .A(n8615), .B(n8614), .Z(n8619) );
  OR U8851 ( .A(n8617), .B(n8616), .Z(n8618) );
  AND U8852 ( .A(n8619), .B(n8618), .Z(n8753) );
  XNOR U8853 ( .A(n8752), .B(n8753), .Z(n8751) );
  OR U8854 ( .A(n8621), .B(n8620), .Z(n8625) );
  OR U8855 ( .A(n8623), .B(n8622), .Z(n8624) );
  AND U8856 ( .A(n8625), .B(n8624), .Z(n8783) );
  NANDN U8857 ( .A(n8626), .B(y[269]), .Z(n8820) );
  NANDN U8858 ( .A(n47), .B(y[284]), .Z(n8819) );
  NANDN U8859 ( .A(n8901), .B(y[260]), .Z(n8818) );
  XNOR U8860 ( .A(n8819), .B(n8818), .Z(n8821) );
  XNOR U8861 ( .A(n8820), .B(n8821), .Z(n8784) );
  NANDN U8862 ( .A(n52), .B(y[279]), .Z(n8964) );
  ANDN U8863 ( .B(x[86]), .A(n8927), .Z(n8629) );
  ANDN U8864 ( .B(x[85]), .A(n8627), .Z(n8628) );
  XNOR U8865 ( .A(n8629), .B(n8628), .Z(n8963) );
  XOR U8866 ( .A(n8964), .B(n8963), .Z(n8785) );
  XNOR U8867 ( .A(n8784), .B(n8785), .Z(n8782) );
  XOR U8868 ( .A(n8783), .B(n8782), .Z(n8750) );
  XNOR U8869 ( .A(n8751), .B(n8750), .Z(n8736) );
  NANDN U8870 ( .A(n8631), .B(n8630), .Z(n8635) );
  OR U8871 ( .A(n8633), .B(n8632), .Z(n8634) );
  NAND U8872 ( .A(n8635), .B(n8634), .Z(n8739) );
  OR U8873 ( .A(n8637), .B(n8636), .Z(n8641) );
  OR U8874 ( .A(n8639), .B(n8638), .Z(n8640) );
  AND U8875 ( .A(n8641), .B(n8640), .Z(n8762) );
  OR U8876 ( .A(n8643), .B(n8642), .Z(n8647) );
  OR U8877 ( .A(n8645), .B(n8644), .Z(n8646) );
  AND U8878 ( .A(n8647), .B(n8646), .Z(n8765) );
  OR U8879 ( .A(n8648), .B(n8965), .Z(n8652) );
  NAND U8880 ( .A(n8650), .B(n8649), .Z(n8651) );
  AND U8881 ( .A(n8652), .B(n8651), .Z(n8855) );
  NAND U8882 ( .A(n8653), .B(o[93]), .Z(n8912) );
  NANDN U8883 ( .A(n8654), .B(y[258]), .Z(n8914) );
  NANDN U8884 ( .A(n8890), .B(y[270]), .Z(n8913) );
  XNOR U8885 ( .A(n8914), .B(n8913), .Z(n8911) );
  XNOR U8886 ( .A(n8912), .B(n8911), .Z(n8857) );
  NANDN U8887 ( .A(n8928), .B(y[261]), .Z(n8944) );
  ANDN U8888 ( .B(x[88]), .A(n8655), .Z(n8658) );
  NANDN U8889 ( .A(n8656), .B(y[263]), .Z(n8657) );
  XOR U8890 ( .A(n8658), .B(n8657), .Z(n8943) );
  XOR U8891 ( .A(n8944), .B(n8943), .Z(n8858) );
  XOR U8892 ( .A(n8857), .B(n8858), .Z(n8856) );
  XNOR U8893 ( .A(n8855), .B(n8856), .Z(n8764) );
  XOR U8894 ( .A(n8762), .B(n8763), .Z(n8738) );
  XNOR U8895 ( .A(n8739), .B(n8738), .Z(n8737) );
  XNOR U8896 ( .A(n8736), .B(n8737), .Z(n9017) );
  XNOR U8897 ( .A(n9018), .B(n9017), .Z(n9016) );
  OR U8898 ( .A(n8660), .B(n8659), .Z(n8664) );
  OR U8899 ( .A(n8662), .B(n8661), .Z(n8663) );
  NAND U8900 ( .A(n8664), .B(n8663), .Z(n9015) );
  XOR U8901 ( .A(n9016), .B(n9015), .Z(n8732) );
  XNOR U8902 ( .A(n8733), .B(n8732), .Z(n8731) );
  OR U8903 ( .A(n8666), .B(n8665), .Z(n8670) );
  OR U8904 ( .A(n8668), .B(n8667), .Z(n8669) );
  NAND U8905 ( .A(n8670), .B(n8669), .Z(n8730) );
  XOR U8906 ( .A(n8731), .B(n8730), .Z(n9010) );
  OR U8907 ( .A(n8672), .B(n8671), .Z(n8676) );
  OR U8908 ( .A(n8674), .B(n8673), .Z(n8675) );
  AND U8909 ( .A(n8676), .B(n8675), .Z(n9011) );
  OR U8910 ( .A(n8678), .B(n8677), .Z(n8682) );
  OR U8911 ( .A(n8680), .B(n8679), .Z(n8681) );
  AND U8912 ( .A(n8682), .B(n8681), .Z(n8995) );
  OR U8913 ( .A(n8684), .B(n8683), .Z(n8688) );
  OR U8914 ( .A(n8686), .B(n8685), .Z(n8687) );
  AND U8915 ( .A(n8688), .B(n8687), .Z(n8996) );
  XOR U8916 ( .A(n8995), .B(n8996), .Z(n8993) );
  OR U8917 ( .A(n8690), .B(n8689), .Z(n8694) );
  OR U8918 ( .A(n8692), .B(n8691), .Z(n8693) );
  NAND U8919 ( .A(n8694), .B(n8693), .Z(n8994) );
  XNOR U8920 ( .A(n8993), .B(n8994), .Z(n8990) );
  OR U8921 ( .A(n8696), .B(n8695), .Z(n8700) );
  OR U8922 ( .A(n8698), .B(n8697), .Z(n8699) );
  NAND U8923 ( .A(n8700), .B(n8699), .Z(n8759) );
  NANDN U8924 ( .A(n8881), .B(x[91]), .Z(n8960) );
  NANDN U8925 ( .A(n46), .B(y[285]), .Z(n8959) );
  XNOR U8926 ( .A(n8960), .B(n8959), .Z(n8958) );
  XNOR U8927 ( .A(n8957), .B(n8958), .Z(n8776) );
  ANDN U8928 ( .B(y[274]), .A(n57), .Z(n8702) );
  ANDN U8929 ( .B(x[77]), .A(n8904), .Z(n8701) );
  XNOR U8930 ( .A(n8702), .B(n8701), .Z(n8837) );
  XNOR U8931 ( .A(n8836), .B(n8837), .Z(n8802) );
  ANDN U8932 ( .B(x[74]), .A(n8900), .Z(n8705) );
  ANDN U8933 ( .B(x[73]), .A(n8703), .Z(n8704) );
  XNOR U8934 ( .A(n8705), .B(n8704), .Z(n8803) );
  XNOR U8935 ( .A(n8802), .B(n8803), .Z(n8778) );
  OR U8936 ( .A(n8707), .B(n8706), .Z(n8711) );
  OR U8937 ( .A(n8709), .B(n8708), .Z(n8710) );
  AND U8938 ( .A(n8711), .B(n8710), .Z(n8779) );
  XNOR U8939 ( .A(n8778), .B(n8779), .Z(n8777) );
  XOR U8940 ( .A(n8776), .B(n8777), .Z(n8758) );
  XNOR U8941 ( .A(n8759), .B(n8758), .Z(n8757) );
  OR U8942 ( .A(n8713), .B(n8712), .Z(n8717) );
  OR U8943 ( .A(n8715), .B(n8714), .Z(n8716) );
  NAND U8944 ( .A(n8717), .B(n8716), .Z(n8756) );
  XOR U8945 ( .A(n8757), .B(n8756), .Z(n8989) );
  XOR U8946 ( .A(n8990), .B(n8989), .Z(n8988) );
  OR U8947 ( .A(n8719), .B(n8718), .Z(n8723) );
  OR U8948 ( .A(n8721), .B(n8720), .Z(n8722) );
  NAND U8949 ( .A(n8723), .B(n8722), .Z(n8987) );
  XOR U8950 ( .A(n8988), .B(n8987), .Z(n9012) );
  XOR U8951 ( .A(n9011), .B(n9012), .Z(n9009) );
  XOR U8952 ( .A(n9010), .B(n9009), .Z(n9030) );
  XNOR U8953 ( .A(n9029), .B(n9030), .Z(n9028) );
  XOR U8954 ( .A(n9027), .B(n9028), .Z(n8724) );
  XOR U8955 ( .A(n8725), .B(n8724), .Z(N191) );
  NANDN U8956 ( .A(n8725), .B(n8724), .Z(n8729) );
  OR U8957 ( .A(n8727), .B(n8726), .Z(n8728) );
  AND U8958 ( .A(n8729), .B(n8728), .Z(n9026) );
  OR U8959 ( .A(n8731), .B(n8730), .Z(n8735) );
  OR U8960 ( .A(n8733), .B(n8732), .Z(n8734) );
  AND U8961 ( .A(n8735), .B(n8734), .Z(n9008) );
  NANDN U8962 ( .A(n8737), .B(n8736), .Z(n8741) );
  OR U8963 ( .A(n8739), .B(n8738), .Z(n8740) );
  AND U8964 ( .A(n8741), .B(n8740), .Z(n8749) );
  OR U8965 ( .A(n8743), .B(n8742), .Z(n8747) );
  OR U8966 ( .A(n8745), .B(n8744), .Z(n8746) );
  NAND U8967 ( .A(n8747), .B(n8746), .Z(n8748) );
  XNOR U8968 ( .A(n8749), .B(n8748), .Z(n9006) );
  OR U8969 ( .A(n8751), .B(n8750), .Z(n8755) );
  OR U8970 ( .A(n8753), .B(n8752), .Z(n8754) );
  AND U8971 ( .A(n8755), .B(n8754), .Z(n9004) );
  OR U8972 ( .A(n8757), .B(n8756), .Z(n8761) );
  OR U8973 ( .A(n8759), .B(n8758), .Z(n8760) );
  AND U8974 ( .A(n8761), .B(n8760), .Z(n8986) );
  OR U8975 ( .A(n8763), .B(n8762), .Z(n8767) );
  OR U8976 ( .A(n8765), .B(n8764), .Z(n8766) );
  AND U8977 ( .A(n8767), .B(n8766), .Z(n8775) );
  NOR U8978 ( .A(n8769), .B(n8768), .Z(n8773) );
  NOR U8979 ( .A(n8771), .B(n8770), .Z(n8772) );
  OR U8980 ( .A(n8773), .B(n8772), .Z(n8774) );
  XNOR U8981 ( .A(n8775), .B(n8774), .Z(n8984) );
  OR U8982 ( .A(n8777), .B(n8776), .Z(n8781) );
  OR U8983 ( .A(n8779), .B(n8778), .Z(n8780) );
  AND U8984 ( .A(n8781), .B(n8780), .Z(n8982) );
  NANDN U8985 ( .A(n8783), .B(n8782), .Z(n8787) );
  NANDN U8986 ( .A(n8785), .B(n8784), .Z(n8786) );
  AND U8987 ( .A(n8787), .B(n8786), .Z(n8795) );
  NAND U8988 ( .A(n8789), .B(n8788), .Z(n8793) );
  OR U8989 ( .A(n8791), .B(n8790), .Z(n8792) );
  NAND U8990 ( .A(n8793), .B(n8792), .Z(n8794) );
  XNOR U8991 ( .A(n8795), .B(n8794), .Z(n8980) );
  OR U8992 ( .A(n8797), .B(n8796), .Z(n8801) );
  OR U8993 ( .A(n8799), .B(n8798), .Z(n8800) );
  AND U8994 ( .A(n8801), .B(n8800), .Z(n8978) );
  NANDN U8995 ( .A(n8803), .B(n8802), .Z(n8806) );
  NANDN U8996 ( .A(n55), .B(y[277]), .Z(n8934) );
  OR U8997 ( .A(n8934), .B(n8804), .Z(n8805) );
  AND U8998 ( .A(n8806), .B(n8805), .Z(n8814) );
  NANDN U8999 ( .A(n8808), .B(n8807), .Z(n8812) );
  NANDN U9000 ( .A(n8810), .B(n8809), .Z(n8811) );
  NAND U9001 ( .A(n8812), .B(n8811), .Z(n8813) );
  XNOR U9002 ( .A(n8814), .B(n8813), .Z(n8976) );
  ANDN U9003 ( .B(x[82]), .A(n8815), .Z(n8817) );
  NANDN U9004 ( .A(n49), .B(y[283]), .Z(n8816) );
  XNOR U9005 ( .A(n8817), .B(n8816), .Z(n8835) );
  NOR U9006 ( .A(n8819), .B(n8818), .Z(n8823) );
  NOR U9007 ( .A(n8821), .B(n8820), .Z(n8822) );
  NOR U9008 ( .A(n8823), .B(n8822), .Z(n8833) );
  ANDN U9009 ( .B(y[268]), .A(n8824), .Z(n8826) );
  ANDN U9010 ( .B(y[279]), .A(n53), .Z(n8825) );
  XNOR U9011 ( .A(n8826), .B(n8825), .Z(n8831) );
  ANDN U9012 ( .B(y[286]), .A(n46), .Z(n8829) );
  NANDN U9013 ( .A(n8827), .B(y[266]), .Z(n8828) );
  XNOR U9014 ( .A(n8829), .B(n8828), .Z(n8830) );
  XOR U9015 ( .A(n8831), .B(n8830), .Z(n8832) );
  XNOR U9016 ( .A(n8833), .B(n8832), .Z(n8834) );
  XOR U9017 ( .A(n8835), .B(n8834), .Z(n8854) );
  NANDN U9018 ( .A(n8837), .B(n8836), .Z(n8840) );
  NANDN U9019 ( .A(n8838), .B(n8863), .Z(n8839) );
  AND U9020 ( .A(n8840), .B(n8839), .Z(n8848) );
  OR U9021 ( .A(n8842), .B(n8841), .Z(n8846) );
  OR U9022 ( .A(n8844), .B(n8843), .Z(n8845) );
  NAND U9023 ( .A(n8846), .B(n8845), .Z(n8847) );
  XNOR U9024 ( .A(n8848), .B(n8847), .Z(n8852) );
  ANDN U9025 ( .B(y[285]), .A(n47), .Z(n8850) );
  NANDN U9026 ( .A(n48), .B(y[284]), .Z(n8849) );
  XNOR U9027 ( .A(n8850), .B(n8849), .Z(n8851) );
  XNOR U9028 ( .A(n8852), .B(n8851), .Z(n8853) );
  XNOR U9029 ( .A(n8854), .B(n8853), .Z(n8942) );
  OR U9030 ( .A(n8856), .B(n8855), .Z(n8860) );
  NANDN U9031 ( .A(n8858), .B(n8857), .Z(n8859) );
  AND U9032 ( .A(n8860), .B(n8859), .Z(n8940) );
  ANDN U9033 ( .B(x[81]), .A(n8861), .Z(n8871) );
  ANDN U9034 ( .B(o[94]), .A(n8862), .Z(n8869) );
  XOR U9035 ( .A(n8863), .B(o[95]), .Z(n8867) );
  NANDN U9036 ( .A(n8864), .B(y[265]), .Z(n8966) );
  NANDN U9037 ( .A(n8865), .B(y[263]), .Z(n8946) );
  XNOR U9038 ( .A(n8966), .B(n8946), .Z(n8866) );
  XNOR U9039 ( .A(n8867), .B(n8866), .Z(n8868) );
  XNOR U9040 ( .A(n8869), .B(n8868), .Z(n8870) );
  XNOR U9041 ( .A(n8871), .B(n8870), .Z(n8880) );
  ANDN U9042 ( .B(x[95]), .A(n8872), .Z(n8874) );
  NANDN U9043 ( .A(n51), .B(y[281]), .Z(n8873) );
  XNOR U9044 ( .A(n8874), .B(n8873), .Z(n8878) );
  ANDN U9045 ( .B(y[280]), .A(n52), .Z(n8876) );
  NANDN U9046 ( .A(n50), .B(y[282]), .Z(n8875) );
  XNOR U9047 ( .A(n8876), .B(n8875), .Z(n8877) );
  XNOR U9048 ( .A(n8878), .B(n8877), .Z(n8879) );
  XNOR U9049 ( .A(n8880), .B(n8879), .Z(n8938) );
  ANDN U9050 ( .B(x[92]), .A(n8881), .Z(n8883) );
  NANDN U9051 ( .A(n45), .B(y[287]), .Z(n8882) );
  XNOR U9052 ( .A(n8883), .B(n8882), .Z(n8889) );
  ANDN U9053 ( .B(x[79]), .A(n8884), .Z(n8887) );
  NANDN U9054 ( .A(n8885), .B(y[267]), .Z(n8886) );
  XNOR U9055 ( .A(n8887), .B(n8886), .Z(n8888) );
  XOR U9056 ( .A(n8889), .B(n8888), .Z(n8899) );
  AND U9057 ( .A(x[94]), .B(y[257]), .Z(n8892) );
  NANDN U9058 ( .A(n8890), .B(y[271]), .Z(n8891) );
  XNOR U9059 ( .A(n8892), .B(n8891), .Z(n8897) );
  ANDN U9060 ( .B(y[258]), .A(n8893), .Z(n8895) );
  NANDN U9061 ( .A(n57), .B(y[275]), .Z(n8894) );
  XNOR U9062 ( .A(n8895), .B(n8894), .Z(n8896) );
  XNOR U9063 ( .A(n8897), .B(n8896), .Z(n8898) );
  XNOR U9064 ( .A(n8899), .B(n8898), .Z(n8910) );
  ANDN U9065 ( .B(x[75]), .A(n8900), .Z(n8903) );
  NANDN U9066 ( .A(n8901), .B(y[261]), .Z(n8902) );
  XNOR U9067 ( .A(n8903), .B(n8902), .Z(n8908) );
  ANDN U9068 ( .B(x[78]), .A(n8904), .Z(n8906) );
  NANDN U9069 ( .A(n54), .B(y[278]), .Z(n8905) );
  XNOR U9070 ( .A(n8906), .B(n8905), .Z(n8907) );
  XNOR U9071 ( .A(n8908), .B(n8907), .Z(n8909) );
  XNOR U9072 ( .A(n8910), .B(n8909), .Z(n8926) );
  OR U9073 ( .A(n8912), .B(n8911), .Z(n8916) );
  OR U9074 ( .A(n8914), .B(n8913), .Z(n8915) );
  AND U9075 ( .A(n8916), .B(n8915), .Z(n8924) );
  NANDN U9076 ( .A(n8918), .B(n8917), .Z(n8922) );
  NANDN U9077 ( .A(n8920), .B(n8919), .Z(n8921) );
  NAND U9078 ( .A(n8922), .B(n8921), .Z(n8923) );
  XNOR U9079 ( .A(n8924), .B(n8923), .Z(n8925) );
  XOR U9080 ( .A(n8926), .B(n8925), .Z(n8936) );
  ANDN U9081 ( .B(x[87]), .A(n8927), .Z(n8930) );
  NANDN U9082 ( .A(n8928), .B(y[262]), .Z(n8929) );
  XNOR U9083 ( .A(n8930), .B(n8929), .Z(n8932) );
  NAND U9084 ( .A(x[91]), .B(y[260]), .Z(n8931) );
  XNOR U9085 ( .A(n8932), .B(n8931), .Z(n8933) );
  XOR U9086 ( .A(n8934), .B(n8933), .Z(n8935) );
  XNOR U9087 ( .A(n8936), .B(n8935), .Z(n8937) );
  XNOR U9088 ( .A(n8938), .B(n8937), .Z(n8939) );
  XNOR U9089 ( .A(n8940), .B(n8939), .Z(n8941) );
  XOR U9090 ( .A(n8942), .B(n8941), .Z(n8974) );
  OR U9091 ( .A(n8944), .B(n8943), .Z(n8948) );
  OR U9092 ( .A(n8946), .B(n8945), .Z(n8947) );
  AND U9093 ( .A(n8948), .B(n8947), .Z(n8956) );
  NANDN U9094 ( .A(n8950), .B(n8949), .Z(n8954) );
  NANDN U9095 ( .A(n8952), .B(n8951), .Z(n8953) );
  NAND U9096 ( .A(n8954), .B(n8953), .Z(n8955) );
  XNOR U9097 ( .A(n8956), .B(n8955), .Z(n8972) );
  NANDN U9098 ( .A(n8958), .B(n8957), .Z(n8962) );
  OR U9099 ( .A(n8960), .B(n8959), .Z(n8961) );
  AND U9100 ( .A(n8962), .B(n8961), .Z(n8970) );
  OR U9101 ( .A(n8964), .B(n8963), .Z(n8968) );
  NANDN U9102 ( .A(n8966), .B(n8965), .Z(n8967) );
  NAND U9103 ( .A(n8968), .B(n8967), .Z(n8969) );
  XNOR U9104 ( .A(n8970), .B(n8969), .Z(n8971) );
  XNOR U9105 ( .A(n8972), .B(n8971), .Z(n8973) );
  XNOR U9106 ( .A(n8974), .B(n8973), .Z(n8975) );
  XNOR U9107 ( .A(n8976), .B(n8975), .Z(n8977) );
  XNOR U9108 ( .A(n8978), .B(n8977), .Z(n8979) );
  XNOR U9109 ( .A(n8980), .B(n8979), .Z(n8981) );
  XNOR U9110 ( .A(n8982), .B(n8981), .Z(n8983) );
  XNOR U9111 ( .A(n8984), .B(n8983), .Z(n8985) );
  XNOR U9112 ( .A(n8986), .B(n8985), .Z(n9002) );
  OR U9113 ( .A(n8988), .B(n8987), .Z(n8992) );
  NANDN U9114 ( .A(n8990), .B(n8989), .Z(n8991) );
  AND U9115 ( .A(n8992), .B(n8991), .Z(n9000) );
  NANDN U9116 ( .A(n8994), .B(n8993), .Z(n8998) );
  OR U9117 ( .A(n8996), .B(n8995), .Z(n8997) );
  NAND U9118 ( .A(n8998), .B(n8997), .Z(n8999) );
  XNOR U9119 ( .A(n9000), .B(n8999), .Z(n9001) );
  XNOR U9120 ( .A(n9002), .B(n9001), .Z(n9003) );
  XNOR U9121 ( .A(n9004), .B(n9003), .Z(n9005) );
  XNOR U9122 ( .A(n9006), .B(n9005), .Z(n9007) );
  XNOR U9123 ( .A(n9008), .B(n9007), .Z(n9024) );
  NANDN U9124 ( .A(n9010), .B(n9009), .Z(n9014) );
  OR U9125 ( .A(n9012), .B(n9011), .Z(n9013) );
  AND U9126 ( .A(n9014), .B(n9013), .Z(n9022) );
  OR U9127 ( .A(n9016), .B(n9015), .Z(n9020) );
  OR U9128 ( .A(n9018), .B(n9017), .Z(n9019) );
  NAND U9129 ( .A(n9020), .B(n9019), .Z(n9021) );
  XNOR U9130 ( .A(n9022), .B(n9021), .Z(n9023) );
  XNOR U9131 ( .A(n9024), .B(n9023), .Z(n9025) );
  XNOR U9132 ( .A(n9026), .B(n9025), .Z(n9042) );
  OR U9133 ( .A(n9028), .B(n9027), .Z(n9032) );
  OR U9134 ( .A(n9030), .B(n9029), .Z(n9031) );
  AND U9135 ( .A(n9032), .B(n9031), .Z(n9040) );
  NANDN U9136 ( .A(n9034), .B(n9033), .Z(n9038) );
  OR U9137 ( .A(n9036), .B(n9035), .Z(n9037) );
  NAND U9138 ( .A(n9038), .B(n9037), .Z(n9039) );
  XNOR U9139 ( .A(n9040), .B(n9039), .Z(n9041) );
  XNOR U9140 ( .A(n9042), .B(n9041), .Z(N192) );
endmodule

