
module hamming_N16000_CC8 ( clk, rst, x, y, o );
  input [1999:0] x;
  input [1999:0] y;
  output [13:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011;
  wire   [13:0] oglobal;

  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NAND U2003 ( .A(n11046), .B(n11047), .Z(n1) );
  NANDN U2004 ( .A(n11045), .B(n11044), .Z(n2) );
  NAND U2005 ( .A(n1), .B(n2), .Z(n11611) );
  XNOR U2006 ( .A(n10829), .B(n10828), .Z(n10830) );
  NAND U2007 ( .A(n11125), .B(n11126), .Z(n3) );
  XOR U2008 ( .A(n11125), .B(n11126), .Z(n4) );
  NANDN U2009 ( .A(n11124), .B(n4), .Z(n5) );
  NAND U2010 ( .A(n3), .B(n5), .Z(n11612) );
  NAND U2011 ( .A(n11052), .B(n11053), .Z(n6) );
  XOR U2012 ( .A(n11052), .B(n11053), .Z(n7) );
  NANDN U2013 ( .A(n11051), .B(n7), .Z(n8) );
  NAND U2014 ( .A(n6), .B(n8), .Z(n11609) );
  XNOR U2015 ( .A(n6553), .B(n6552), .Z(n6555) );
  XNOR U2016 ( .A(n6547), .B(n6546), .Z(n6548) );
  XNOR U2017 ( .A(n11313), .B(n11312), .Z(n11354) );
  XNOR U2018 ( .A(n11347), .B(n11346), .Z(n11348) );
  XOR U2019 ( .A(n11662), .B(n11661), .Z(n11664) );
  XNOR U2020 ( .A(n11836), .B(n11835), .Z(n11837) );
  XNOR U2021 ( .A(n11974), .B(n11973), .Z(n11990) );
  NAND U2022 ( .A(n10332), .B(n10333), .Z(n9) );
  XOR U2023 ( .A(n10332), .B(n10333), .Z(n10) );
  NANDN U2024 ( .A(n10331), .B(n10), .Z(n11) );
  NAND U2025 ( .A(n9), .B(n11), .Z(n10634) );
  NAND U2026 ( .A(n11705), .B(n11706), .Z(n12) );
  XOR U2027 ( .A(n11705), .B(n11706), .Z(n13) );
  NANDN U2028 ( .A(n11704), .B(n13), .Z(n14) );
  NAND U2029 ( .A(n12), .B(n14), .Z(n11919) );
  NAND U2030 ( .A(n261), .B(n260), .Z(n15) );
  NAND U2031 ( .A(n258), .B(n259), .Z(n16) );
  AND U2032 ( .A(n15), .B(n16), .Z(n8470) );
  NAND U2033 ( .A(n1772), .B(n1771), .Z(n17) );
  NANDN U2034 ( .A(n1774), .B(n1773), .Z(n18) );
  AND U2035 ( .A(n17), .B(n18), .Z(n7721) );
  NAND U2036 ( .A(n11049), .B(n11050), .Z(n19) );
  XOR U2037 ( .A(n11049), .B(n11050), .Z(n20) );
  NANDN U2038 ( .A(n11048), .B(n20), .Z(n21) );
  NAND U2039 ( .A(n19), .B(n21), .Z(n11610) );
  XOR U2040 ( .A(n11222), .B(n11221), .Z(n22) );
  NANDN U2041 ( .A(n11223), .B(n22), .Z(n23) );
  NAND U2042 ( .A(n11222), .B(n11221), .Z(n24) );
  AND U2043 ( .A(n23), .B(n24), .Z(n11583) );
  NAND U2044 ( .A(n11613), .B(n11614), .Z(n25) );
  XOR U2045 ( .A(n11613), .B(n11614), .Z(n26) );
  NANDN U2046 ( .A(n11612), .B(n26), .Z(n27) );
  NAND U2047 ( .A(n25), .B(n27), .Z(n11749) );
  XNOR U2048 ( .A(n10835), .B(n10834), .Z(n10837) );
  XNOR U2049 ( .A(n10568), .B(n10567), .Z(n10569) );
  XOR U2050 ( .A(n9372), .B(n9371), .Z(n10442) );
  XOR U2051 ( .A(n10831), .B(n10830), .Z(n11263) );
  XNOR U2052 ( .A(n11640), .B(n11639), .Z(n11641) );
  XNOR U2053 ( .A(n11353), .B(n11352), .Z(n11355) );
  XNOR U2054 ( .A(n11656), .B(n11655), .Z(n11657) );
  XNOR U2055 ( .A(n11909), .B(n11908), .Z(n11900) );
  XNOR U2056 ( .A(n11710), .B(n11709), .Z(n11649) );
  XOR U2057 ( .A(n11699), .B(n11698), .Z(n11701) );
  NAND U2058 ( .A(n11645), .B(n11647), .Z(n28) );
  XOR U2059 ( .A(n11645), .B(n11647), .Z(n29) );
  NAND U2060 ( .A(n29), .B(n11646), .Z(n30) );
  NAND U2061 ( .A(n28), .B(n30), .Z(n11704) );
  NAND U2062 ( .A(n11934), .B(n11936), .Z(n31) );
  XOR U2063 ( .A(n11934), .B(n11936), .Z(n32) );
  NAND U2064 ( .A(n32), .B(n11935), .Z(n33) );
  NAND U2065 ( .A(n31), .B(n33), .Z(n11989) );
  NAND U2066 ( .A(n257), .B(n256), .Z(n34) );
  NAND U2067 ( .A(n254), .B(n255), .Z(n35) );
  AND U2068 ( .A(n34), .B(n35), .Z(n8472) );
  NAND U2069 ( .A(n7675), .B(n7674), .Z(n36) );
  NAND U2070 ( .A(n7672), .B(n7673), .Z(n37) );
  AND U2071 ( .A(n36), .B(n37), .Z(n9281) );
  NAND U2072 ( .A(n7721), .B(n7720), .Z(n38) );
  NAND U2073 ( .A(n7718), .B(n7719), .Z(n39) );
  AND U2074 ( .A(n38), .B(n39), .Z(n9264) );
  NAND U2075 ( .A(n6903), .B(n6902), .Z(n40) );
  NAND U2076 ( .A(n6900), .B(n6901), .Z(n41) );
  AND U2077 ( .A(n40), .B(n41), .Z(n9321) );
  XOR U2078 ( .A(n7915), .B(n7914), .Z(n42) );
  NANDN U2079 ( .A(n7916), .B(n42), .Z(n43) );
  NAND U2080 ( .A(n7915), .B(n7914), .Z(n44) );
  AND U2081 ( .A(n43), .B(n44), .Z(n10150) );
  NAND U2082 ( .A(n9582), .B(n9581), .Z(n45) );
  NAND U2083 ( .A(n9579), .B(n9580), .Z(n46) );
  AND U2084 ( .A(n45), .B(n46), .Z(n11134) );
  NAND U2085 ( .A(n9333), .B(n9332), .Z(n47) );
  XOR U2086 ( .A(n9333), .B(n9332), .Z(n48) );
  NANDN U2087 ( .A(n9334), .B(n48), .Z(n49) );
  NAND U2088 ( .A(n47), .B(n49), .Z(n10648) );
  NAND U2089 ( .A(n10541), .B(n10540), .Z(n50) );
  NAND U2090 ( .A(n10538), .B(n10539), .Z(n51) );
  NAND U2091 ( .A(n50), .B(n51), .Z(n10714) );
  NAND U2092 ( .A(n9299), .B(n9298), .Z(n52) );
  NANDN U2093 ( .A(n9301), .B(n9300), .Z(n53) );
  NAND U2094 ( .A(n52), .B(n53), .Z(n10822) );
  NAND U2095 ( .A(n9349), .B(n9350), .Z(n54) );
  NANDN U2096 ( .A(n9348), .B(n9347), .Z(n55) );
  NAND U2097 ( .A(n54), .B(n55), .Z(n10678) );
  XOR U2098 ( .A(n11122), .B(n11121), .Z(n56) );
  NANDN U2099 ( .A(n11123), .B(n56), .Z(n57) );
  NAND U2100 ( .A(n11122), .B(n11121), .Z(n58) );
  AND U2101 ( .A(n57), .B(n58), .Z(n11613) );
  NAND U2102 ( .A(n11143), .B(n11142), .Z(n59) );
  NANDN U2103 ( .A(n11141), .B(n11140), .Z(n60) );
  AND U2104 ( .A(n59), .B(n60), .Z(n11604) );
  NAND U2105 ( .A(n660), .B(n659), .Z(n61) );
  NAND U2106 ( .A(n657), .B(n658), .Z(n62) );
  AND U2107 ( .A(n61), .B(n62), .Z(n8637) );
  XNOR U2108 ( .A(n9382), .B(n9381), .Z(n9384) );
  XOR U2109 ( .A(n11611), .B(n11609), .Z(n63) );
  NAND U2110 ( .A(n63), .B(n11610), .Z(n64) );
  NAND U2111 ( .A(n11611), .B(n11609), .Z(n65) );
  AND U2112 ( .A(n64), .B(n65), .Z(n11750) );
  NAND U2113 ( .A(n11583), .B(n11584), .Z(n66) );
  XOR U2114 ( .A(n11583), .B(n11584), .Z(n67) );
  NANDN U2115 ( .A(n11582), .B(n67), .Z(n68) );
  NAND U2116 ( .A(n66), .B(n68), .Z(n11756) );
  XNOR U2117 ( .A(n9370), .B(n9369), .Z(n9371) );
  XNOR U2118 ( .A(n9107), .B(n9106), .Z(n9109) );
  XNOR U2119 ( .A(n6549), .B(n6548), .Z(n6660) );
  XNOR U2120 ( .A(n11311), .B(n11310), .Z(n11312) );
  XNOR U2121 ( .A(n11287), .B(n11286), .Z(n11288) );
  XOR U2122 ( .A(n11642), .B(n11641), .Z(n11365) );
  XNOR U2123 ( .A(n9378), .B(n9377), .Z(n10444) );
  XOR U2124 ( .A(n9067), .B(n9066), .Z(n10549) );
  XNOR U2125 ( .A(n11829), .B(n11828), .Z(n11831) );
  NAND U2126 ( .A(n11963), .B(n11962), .Z(n69) );
  NAND U2127 ( .A(n11960), .B(n11961), .Z(n70) );
  AND U2128 ( .A(n69), .B(n70), .Z(n11983) );
  XOR U2129 ( .A(n11361), .B(n11360), .Z(n11371) );
  XOR U2130 ( .A(n11349), .B(n11348), .Z(n11377) );
  XNOR U2131 ( .A(n11842), .B(n11841), .Z(n11843) );
  XNOR U2132 ( .A(n11650), .B(n11649), .Z(n11652) );
  NAND U2133 ( .A(n10634), .B(n10635), .Z(n71) );
  XOR U2134 ( .A(n10634), .B(n10635), .Z(n72) );
  NANDN U2135 ( .A(n10633), .B(n72), .Z(n73) );
  NAND U2136 ( .A(n71), .B(n73), .Z(n11646) );
  NAND U2137 ( .A(n11918), .B(n11920), .Z(n74) );
  XOR U2138 ( .A(n11918), .B(n11920), .Z(n75) );
  NAND U2139 ( .A(n75), .B(n11919), .Z(n76) );
  NAND U2140 ( .A(n74), .B(n76), .Z(n11935) );
  NAND U2141 ( .A(n11997), .B(n11998), .Z(n77) );
  XOR U2142 ( .A(n11997), .B(n11998), .Z(n78) );
  NANDN U2143 ( .A(n11996), .B(n78), .Z(n79) );
  NAND U2144 ( .A(n77), .B(n79), .Z(n12006) );
  XOR U2145 ( .A(x[816]), .B(y[816]), .Z(n3296) );
  XOR U2146 ( .A(x[818]), .B(y[818]), .Z(n3294) );
  XOR U2147 ( .A(x[1935]), .B(y[1935]), .Z(n3293) );
  XOR U2148 ( .A(n3294), .B(n3293), .Z(n3295) );
  XOR U2149 ( .A(n3296), .B(n3295), .Z(n2402) );
  XOR U2150 ( .A(x[1382]), .B(y[1382]), .Z(n5169) );
  XOR U2151 ( .A(x[1384]), .B(y[1384]), .Z(n5167) );
  XOR U2152 ( .A(x[1386]), .B(y[1386]), .Z(n5166) );
  XOR U2153 ( .A(n5167), .B(n5166), .Z(n5168) );
  XOR U2154 ( .A(n5169), .B(n5168), .Z(n2400) );
  XOR U2155 ( .A(x[812]), .B(y[812]), .Z(n3284) );
  XOR U2156 ( .A(x[387]), .B(y[387]), .Z(n3282) );
  XOR U2157 ( .A(x[814]), .B(y[814]), .Z(n3281) );
  XOR U2158 ( .A(n3282), .B(n3281), .Z(n3283) );
  XNOR U2159 ( .A(n3284), .B(n3283), .Z(n2399) );
  XNOR U2160 ( .A(n2400), .B(n2399), .Z(n2401) );
  XNOR U2161 ( .A(n2402), .B(n2401), .Z(n4092) );
  XOR U2162 ( .A(x[808]), .B(y[808]), .Z(n3272) );
  XOR U2163 ( .A(x[810]), .B(y[810]), .Z(n3269) );
  XNOR U2164 ( .A(x[1933]), .B(y[1933]), .Z(n3270) );
  XNOR U2165 ( .A(n3269), .B(n3270), .Z(n3271) );
  XOR U2166 ( .A(n3272), .B(n3271), .Z(n2174) );
  XOR U2167 ( .A(x[1870]), .B(y[1870]), .Z(n2546) );
  XOR U2168 ( .A(x[628]), .B(y[628]), .Z(n2543) );
  XNOR U2169 ( .A(x[1872]), .B(y[1872]), .Z(n2544) );
  XNOR U2170 ( .A(n2543), .B(n2544), .Z(n2545) );
  XOR U2171 ( .A(n2546), .B(n2545), .Z(n2172) );
  XOR U2172 ( .A(x[804]), .B(y[804]), .Z(n3278) );
  XOR U2173 ( .A(x[393]), .B(y[393]), .Z(n3275) );
  XNOR U2174 ( .A(x[806]), .B(y[806]), .Z(n3276) );
  XNOR U2175 ( .A(n3275), .B(n3276), .Z(n3277) );
  XNOR U2176 ( .A(n3278), .B(n3277), .Z(n2171) );
  XNOR U2177 ( .A(n2172), .B(n2171), .Z(n2173) );
  XOR U2178 ( .A(n2174), .B(n2173), .Z(n4093) );
  XNOR U2179 ( .A(n4092), .B(n4093), .Z(n4095) );
  XOR U2180 ( .A(x[800]), .B(y[800]), .Z(n4791) );
  XOR U2181 ( .A(x[397]), .B(y[397]), .Z(n4788) );
  XNOR U2182 ( .A(x[802]), .B(y[802]), .Z(n4789) );
  XNOR U2183 ( .A(n4788), .B(n4789), .Z(n4790) );
  XOR U2184 ( .A(n4791), .B(n4790), .Z(n2150) );
  XOR U2185 ( .A(x[1374]), .B(y[1374]), .Z(n5331) );
  XOR U2186 ( .A(x[19]), .B(y[19]), .Z(n5328) );
  XNOR U2187 ( .A(x[1376]), .B(y[1376]), .Z(n5329) );
  XNOR U2188 ( .A(n5328), .B(n5329), .Z(n5330) );
  XOR U2189 ( .A(n5331), .B(n5330), .Z(n2148) );
  XOR U2190 ( .A(x[794]), .B(y[794]), .Z(n4779) );
  XOR U2191 ( .A(x[761]), .B(y[761]), .Z(n4776) );
  XNOR U2192 ( .A(x[796]), .B(y[796]), .Z(n4777) );
  XNOR U2193 ( .A(n4776), .B(n4777), .Z(n4778) );
  XNOR U2194 ( .A(n4779), .B(n4778), .Z(n2147) );
  XNOR U2195 ( .A(n2148), .B(n2147), .Z(n2149) );
  XNOR U2196 ( .A(n2150), .B(n2149), .Z(n4094) );
  XNOR U2197 ( .A(n4095), .B(n4094), .Z(n4443) );
  XOR U2198 ( .A(x[790]), .B(y[790]), .Z(n4785) );
  XOR U2199 ( .A(x[403]), .B(y[403]), .Z(n4782) );
  XNOR U2200 ( .A(x[792]), .B(y[792]), .Z(n4783) );
  XNOR U2201 ( .A(n4782), .B(n4783), .Z(n4784) );
  XOR U2202 ( .A(n4785), .B(n4784), .Z(n2438) );
  XOR U2203 ( .A(x[1874]), .B(y[1874]), .Z(n3206) );
  XOR U2204 ( .A(x[632]), .B(y[632]), .Z(n3204) );
  XOR U2205 ( .A(x[1876]), .B(y[1876]), .Z(n3203) );
  XOR U2206 ( .A(n3204), .B(n3203), .Z(n3205) );
  XOR U2207 ( .A(n3206), .B(n3205), .Z(n2436) );
  XOR U2208 ( .A(x[784]), .B(y[784]), .Z(n3404) );
  XOR U2209 ( .A(x[767]), .B(y[767]), .Z(n3402) );
  XOR U2210 ( .A(x[788]), .B(y[788]), .Z(n3401) );
  XOR U2211 ( .A(n3402), .B(n3401), .Z(n3403) );
  XNOR U2212 ( .A(n3404), .B(n3403), .Z(n2435) );
  XNOR U2213 ( .A(n2436), .B(n2435), .Z(n2437) );
  XNOR U2214 ( .A(n2438), .B(n2437), .Z(n1811) );
  XOR U2215 ( .A(x[778]), .B(y[778]), .Z(n3392) );
  XOR U2216 ( .A(x[780]), .B(y[780]), .Z(n3389) );
  XNOR U2217 ( .A(x[1931]), .B(y[1931]), .Z(n3390) );
  XNOR U2218 ( .A(n3389), .B(n3390), .Z(n3391) );
  XOR U2219 ( .A(n3392), .B(n3391), .Z(n2204) );
  XOR U2220 ( .A(x[1366]), .B(y[1366]), .Z(n5361) );
  XOR U2221 ( .A(x[421]), .B(y[421]), .Z(n5358) );
  XNOR U2222 ( .A(x[1368]), .B(y[1368]), .Z(n5359) );
  XNOR U2223 ( .A(n5358), .B(n5359), .Z(n5360) );
  XOR U2224 ( .A(n5361), .B(n5360), .Z(n2202) );
  XOR U2225 ( .A(x[774]), .B(y[774]), .Z(n3398) );
  XOR U2226 ( .A(x[409]), .B(y[409]), .Z(n3395) );
  XNOR U2227 ( .A(x[776]), .B(y[776]), .Z(n3396) );
  XNOR U2228 ( .A(n3395), .B(n3396), .Z(n3397) );
  XNOR U2229 ( .A(n3398), .B(n3397), .Z(n2201) );
  XNOR U2230 ( .A(n2202), .B(n2201), .Z(n2203) );
  XOR U2231 ( .A(n2204), .B(n2203), .Z(n1812) );
  XNOR U2232 ( .A(n1811), .B(n1812), .Z(n1814) );
  XOR U2233 ( .A(x[770]), .B(y[770]), .Z(n3176) );
  XOR U2234 ( .A(x[772]), .B(y[772]), .Z(n3173) );
  XNOR U2235 ( .A(x[1929]), .B(y[1929]), .Z(n3174) );
  XNOR U2236 ( .A(n3173), .B(n3174), .Z(n3175) );
  XOR U2237 ( .A(n3176), .B(n3175), .Z(n2234) );
  XOR U2238 ( .A(x[1878]), .B(y[1878]), .Z(n3674) );
  XOR U2239 ( .A(x[636]), .B(y[636]), .Z(n3671) );
  XNOR U2240 ( .A(x[1880]), .B(y[1880]), .Z(n3672) );
  XNOR U2241 ( .A(n3671), .B(n3672), .Z(n3673) );
  XOR U2242 ( .A(n3674), .B(n3673), .Z(n2232) );
  XOR U2243 ( .A(x[764]), .B(y[764]), .Z(n3164) );
  XOR U2244 ( .A(x[415]), .B(y[415]), .Z(n3161) );
  XNOR U2245 ( .A(x[766]), .B(y[766]), .Z(n3162) );
  XNOR U2246 ( .A(n3161), .B(n3162), .Z(n3163) );
  XNOR U2247 ( .A(n3164), .B(n3163), .Z(n2231) );
  XNOR U2248 ( .A(n2232), .B(n2231), .Z(n2233) );
  XNOR U2249 ( .A(n2234), .B(n2233), .Z(n1813) );
  XNOR U2250 ( .A(n1814), .B(n1813), .Z(n4441) );
  XOR U2251 ( .A(x[760]), .B(y[760]), .Z(n3170) );
  XOR U2252 ( .A(x[419]), .B(y[419]), .Z(n3167) );
  XNOR U2253 ( .A(x[762]), .B(y[762]), .Z(n3168) );
  XNOR U2254 ( .A(n3167), .B(n3168), .Z(n3169) );
  XOR U2255 ( .A(n3170), .B(n3169), .Z(n2210) );
  XOR U2256 ( .A(x[1358]), .B(y[1358]), .Z(n5559) );
  XOR U2257 ( .A(x[427]), .B(y[427]), .Z(n5556) );
  XNOR U2258 ( .A(x[1360]), .B(y[1360]), .Z(n5557) );
  XNOR U2259 ( .A(n5556), .B(n5557), .Z(n5558) );
  XOR U2260 ( .A(n5559), .B(n5558), .Z(n2208) );
  XOR U2261 ( .A(x[756]), .B(y[756]), .Z(n3158) );
  XOR U2262 ( .A(x[758]), .B(y[758]), .Z(n3155) );
  XNOR U2263 ( .A(x[781]), .B(y[781]), .Z(n3156) );
  XNOR U2264 ( .A(n3155), .B(n3156), .Z(n3157) );
  XNOR U2265 ( .A(n3158), .B(n3157), .Z(n2207) );
  XNOR U2266 ( .A(n2208), .B(n2207), .Z(n2209) );
  XNOR U2267 ( .A(n2210), .B(n2209), .Z(n4452) );
  XOR U2268 ( .A(x[752]), .B(y[752]), .Z(n3146) );
  XOR U2269 ( .A(x[429]), .B(y[429]), .Z(n3143) );
  XNOR U2270 ( .A(x[754]), .B(y[754]), .Z(n3144) );
  XNOR U2271 ( .A(n3143), .B(n3144), .Z(n3145) );
  XOR U2272 ( .A(n3146), .B(n3145), .Z(n1994) );
  XOR U2273 ( .A(x[1882]), .B(y[1882]), .Z(n2582) );
  XOR U2274 ( .A(x[910]), .B(y[910]), .Z(n2579) );
  XNOR U2275 ( .A(x[1884]), .B(y[1884]), .Z(n2580) );
  XNOR U2276 ( .A(n2579), .B(n2580), .Z(n2581) );
  XOR U2277 ( .A(n2582), .B(n2581), .Z(n1992) );
  XOR U2278 ( .A(x[742]), .B(y[742]), .Z(n3152) );
  XOR U2279 ( .A(x[750]), .B(y[750]), .Z(n3149) );
  XNOR U2280 ( .A(x[787]), .B(y[787]), .Z(n3150) );
  XNOR U2281 ( .A(n3149), .B(n3150), .Z(n3151) );
  XNOR U2282 ( .A(n3152), .B(n3151), .Z(n1991) );
  XNOR U2283 ( .A(n1992), .B(n1991), .Z(n1993) );
  XNOR U2284 ( .A(n1994), .B(n1993), .Z(n4453) );
  XOR U2285 ( .A(n4452), .B(n4453), .Z(n4455) );
  XOR U2286 ( .A(x[736]), .B(y[736]), .Z(n3987) );
  XOR U2287 ( .A(x[740]), .B(y[740]), .Z(n3984) );
  XNOR U2288 ( .A(x[1927]), .B(y[1927]), .Z(n3985) );
  XNOR U2289 ( .A(n3984), .B(n3985), .Z(n3986) );
  XOR U2290 ( .A(n3987), .B(n3986), .Z(n1970) );
  XOR U2291 ( .A(x[1350]), .B(y[1350]), .Z(n5547) );
  XOR U2292 ( .A(x[35]), .B(y[35]), .Z(n5544) );
  XNOR U2293 ( .A(x[1352]), .B(y[1352]), .Z(n5545) );
  XNOR U2294 ( .A(n5544), .B(n5545), .Z(n5546) );
  XOR U2295 ( .A(n5547), .B(n5546), .Z(n1968) );
  XOR U2296 ( .A(x[730]), .B(y[730]), .Z(n3975) );
  XOR U2297 ( .A(x[435]), .B(y[435]), .Z(n3972) );
  XNOR U2298 ( .A(x[732]), .B(y[732]), .Z(n3973) );
  XNOR U2299 ( .A(n3972), .B(n3973), .Z(n3974) );
  XNOR U2300 ( .A(n3975), .B(n3974), .Z(n1967) );
  XNOR U2301 ( .A(n1968), .B(n1967), .Z(n1969) );
  XNOR U2302 ( .A(n1970), .B(n1969), .Z(n4454) );
  XNOR U2303 ( .A(n4455), .B(n4454), .Z(n4440) );
  XOR U2304 ( .A(n4441), .B(n4440), .Z(n4442) );
  XNOR U2305 ( .A(n4443), .B(n4442), .Z(n4813) );
  XOR U2306 ( .A(x[726]), .B(y[726]), .Z(n3981) );
  XOR U2307 ( .A(x[728]), .B(y[728]), .Z(n3978) );
  XNOR U2308 ( .A(x[1925]), .B(y[1925]), .Z(n3979) );
  XNOR U2309 ( .A(n3978), .B(n3979), .Z(n3980) );
  XOR U2310 ( .A(n3981), .B(n3980), .Z(n2024) );
  XOR U2311 ( .A(x[1886]), .B(y[1886]), .Z(n101) );
  XOR U2312 ( .A(x[1888]), .B(y[1888]), .Z(n98) );
  XNOR U2313 ( .A(x[1890]), .B(y[1890]), .Z(n99) );
  XNOR U2314 ( .A(n98), .B(n99), .Z(n100) );
  XOR U2315 ( .A(n101), .B(n100), .Z(n2022) );
  XOR U2316 ( .A(x[716]), .B(y[716]), .Z(n3969) );
  XOR U2317 ( .A(x[443]), .B(y[443]), .Z(n3966) );
  XNOR U2318 ( .A(x[724]), .B(y[724]), .Z(n3967) );
  XNOR U2319 ( .A(n3966), .B(n3967), .Z(n3968) );
  XNOR U2320 ( .A(n3969), .B(n3968), .Z(n2021) );
  XNOR U2321 ( .A(n2022), .B(n2021), .Z(n2023) );
  XNOR U2322 ( .A(n2024), .B(n2023), .Z(n4068) );
  XOR U2323 ( .A(x[708]), .B(y[708]), .Z(n3957) );
  XOR U2324 ( .A(x[449]), .B(y[449]), .Z(n3954) );
  XNOR U2325 ( .A(x[710]), .B(y[710]), .Z(n3955) );
  XNOR U2326 ( .A(n3954), .B(n3955), .Z(n3956) );
  XOR U2327 ( .A(n3957), .B(n3956), .Z(n2000) );
  XOR U2328 ( .A(x[1342]), .B(y[1342]), .Z(n6045) );
  XOR U2329 ( .A(x[41]), .B(y[41]), .Z(n6042) );
  XNOR U2330 ( .A(x[1344]), .B(y[1344]), .Z(n6043) );
  XNOR U2331 ( .A(n6042), .B(n6043), .Z(n6044) );
  XOR U2332 ( .A(n6045), .B(n6044), .Z(n1998) );
  XOR U2333 ( .A(x[704]), .B(y[704]), .Z(n3963) );
  XOR U2334 ( .A(x[706]), .B(y[706]), .Z(n3960) );
  XNOR U2335 ( .A(x[801]), .B(y[801]), .Z(n3961) );
  XNOR U2336 ( .A(n3960), .B(n3961), .Z(n3962) );
  XNOR U2337 ( .A(n3963), .B(n3962), .Z(n1997) );
  XNOR U2338 ( .A(n1998), .B(n1997), .Z(n1999) );
  XOR U2339 ( .A(n2000), .B(n1999), .Z(n4069) );
  XNOR U2340 ( .A(n4068), .B(n4069), .Z(n4071) );
  XOR U2341 ( .A(x[696]), .B(y[696]), .Z(n2864) );
  XOR U2342 ( .A(x[455]), .B(y[455]), .Z(n2861) );
  XNOR U2343 ( .A(x[700]), .B(y[700]), .Z(n2862) );
  XNOR U2344 ( .A(n2861), .B(n2862), .Z(n2863) );
  XOR U2345 ( .A(n2864), .B(n2863), .Z(n2054) );
  XOR U2346 ( .A(x[1892]), .B(y[1892]), .Z(n343) );
  XOR U2347 ( .A(x[648]), .B(y[648]), .Z(n340) );
  XNOR U2348 ( .A(x[1894]), .B(y[1894]), .Z(n341) );
  XNOR U2349 ( .A(n340), .B(n341), .Z(n342) );
  XOR U2350 ( .A(n343), .B(n342), .Z(n2052) );
  XOR U2351 ( .A(x[688]), .B(y[688]), .Z(n2852) );
  XOR U2352 ( .A(x[690]), .B(y[690]), .Z(n2849) );
  XNOR U2353 ( .A(x[807]), .B(y[807]), .Z(n2850) );
  XNOR U2354 ( .A(n2849), .B(n2850), .Z(n2851) );
  XNOR U2355 ( .A(n2852), .B(n2851), .Z(n2051) );
  XNOR U2356 ( .A(n2052), .B(n2051), .Z(n2053) );
  XNOR U2357 ( .A(n2054), .B(n2053), .Z(n4070) );
  XOR U2358 ( .A(n4071), .B(n4070), .Z(n4449) );
  XOR U2359 ( .A(x[684]), .B(y[684]), .Z(n2858) );
  XOR U2360 ( .A(x[686]), .B(y[686]), .Z(n2855) );
  XNOR U2361 ( .A(x[1923]), .B(y[1923]), .Z(n2856) );
  XNOR U2362 ( .A(n2855), .B(n2856), .Z(n2857) );
  XOR U2363 ( .A(n2858), .B(n2857), .Z(n2030) );
  XOR U2364 ( .A(x[1334]), .B(y[1334]), .Z(n5151) );
  XOR U2365 ( .A(x[441]), .B(y[441]), .Z(n5148) );
  XNOR U2366 ( .A(x[1336]), .B(y[1336]), .Z(n5149) );
  XNOR U2367 ( .A(n5148), .B(n5149), .Z(n5150) );
  XOR U2368 ( .A(n5151), .B(n5150), .Z(n2028) );
  XOR U2369 ( .A(x[680]), .B(y[680]), .Z(n2678) );
  XOR U2370 ( .A(x[463]), .B(y[463]), .Z(n2675) );
  XNOR U2371 ( .A(x[682]), .B(y[682]), .Z(n2676) );
  XNOR U2372 ( .A(n2675), .B(n2676), .Z(n2677) );
  XNOR U2373 ( .A(n2678), .B(n2677), .Z(n2027) );
  XNOR U2374 ( .A(n2028), .B(n2027), .Z(n2029) );
  XNOR U2375 ( .A(n2030), .B(n2029), .Z(n4008) );
  XOR U2376 ( .A(x[668]), .B(y[668]), .Z(n2672) );
  XOR U2377 ( .A(x[471]), .B(y[471]), .Z(n2669) );
  XNOR U2378 ( .A(x[670]), .B(y[670]), .Z(n2670) );
  XNOR U2379 ( .A(n2669), .B(n2670), .Z(n2671) );
  XOR U2380 ( .A(n2672), .B(n2671), .Z(n2084) );
  XOR U2381 ( .A(x[1896]), .B(y[1896]), .Z(n378) );
  XOR U2382 ( .A(x[652]), .B(y[652]), .Z(n375) );
  XNOR U2383 ( .A(x[1898]), .B(y[1898]), .Z(n376) );
  XNOR U2384 ( .A(n375), .B(n376), .Z(n377) );
  XOR U2385 ( .A(n378), .B(n377), .Z(n2082) );
  XOR U2386 ( .A(x[658]), .B(y[658]), .Z(n2648) );
  XOR U2387 ( .A(x[660]), .B(y[660]), .Z(n2645) );
  XNOR U2388 ( .A(x[821]), .B(y[821]), .Z(n2646) );
  XNOR U2389 ( .A(n2645), .B(n2646), .Z(n2647) );
  XNOR U2390 ( .A(n2648), .B(n2647), .Z(n2081) );
  XNOR U2391 ( .A(n2082), .B(n2081), .Z(n2083) );
  XOR U2392 ( .A(n2084), .B(n2083), .Z(n4009) );
  XNOR U2393 ( .A(n4008), .B(n4009), .Z(n4011) );
  XOR U2394 ( .A(x[650]), .B(y[650]), .Z(n2654) );
  XOR U2395 ( .A(x[483]), .B(y[483]), .Z(n2651) );
  XNOR U2396 ( .A(x[654]), .B(y[654]), .Z(n2652) );
  XNOR U2397 ( .A(n2651), .B(n2652), .Z(n2653) );
  XOR U2398 ( .A(n2654), .B(n2653), .Z(n2060) );
  XOR U2399 ( .A(x[1326]), .B(y[1326]), .Z(n5145) );
  XOR U2400 ( .A(x[447]), .B(y[447]), .Z(n5142) );
  XNOR U2401 ( .A(x[1328]), .B(y[1328]), .Z(n5143) );
  XNOR U2402 ( .A(n5142), .B(n5143), .Z(n5144) );
  XOR U2403 ( .A(n5145), .B(n5144), .Z(n2058) );
  XOR U2404 ( .A(x[642]), .B(y[642]), .Z(n2954) );
  XOR U2405 ( .A(x[646]), .B(y[646]), .Z(n2951) );
  XNOR U2406 ( .A(x[827]), .B(y[827]), .Z(n2952) );
  XNOR U2407 ( .A(n2951), .B(n2952), .Z(n2953) );
  XNOR U2408 ( .A(n2954), .B(n2953), .Z(n2057) );
  XNOR U2409 ( .A(n2058), .B(n2057), .Z(n2059) );
  XNOR U2410 ( .A(n2060), .B(n2059), .Z(n4010) );
  XNOR U2411 ( .A(n4011), .B(n4010), .Z(n4447) );
  XOR U2412 ( .A(x[600]), .B(y[600]), .Z(n1928) );
  XOR U2413 ( .A(x[511]), .B(y[511]), .Z(n1925) );
  XNOR U2414 ( .A(x[602]), .B(y[602]), .Z(n1926) );
  XNOR U2415 ( .A(n1925), .B(n1926), .Z(n1927) );
  XOR U2416 ( .A(n1928), .B(n1927), .Z(n2144) );
  XOR U2417 ( .A(x[1904]), .B(y[1904]), .Z(n197) );
  XOR U2418 ( .A(x[1906]), .B(y[1906]), .Z(n194) );
  XNOR U2419 ( .A(x[1908]), .B(y[1908]), .Z(n195) );
  XNOR U2420 ( .A(n194), .B(n195), .Z(n196) );
  XOR U2421 ( .A(n197), .B(n196), .Z(n2142) );
  XOR U2422 ( .A(x[596]), .B(y[596]), .Z(n1934) );
  XOR U2423 ( .A(x[598]), .B(y[598]), .Z(n1931) );
  XNOR U2424 ( .A(x[847]), .B(y[847]), .Z(n1932) );
  XNOR U2425 ( .A(n1931), .B(n1932), .Z(n1933) );
  XNOR U2426 ( .A(n1934), .B(n1933), .Z(n2141) );
  XNOR U2427 ( .A(n2142), .B(n2141), .Z(n2143) );
  XNOR U2428 ( .A(n2144), .B(n2143), .Z(n4152) );
  XOR U2429 ( .A(x[634]), .B(y[634]), .Z(n2942) );
  XOR U2430 ( .A(x[638]), .B(y[638]), .Z(n2939) );
  XNOR U2431 ( .A(x[1919]), .B(y[1919]), .Z(n2940) );
  XNOR U2432 ( .A(n2939), .B(n2940), .Z(n2941) );
  XOR U2433 ( .A(n2942), .B(n2941), .Z(n2114) );
  XOR U2434 ( .A(x[1900]), .B(y[1900]), .Z(n552) );
  XOR U2435 ( .A(x[656]), .B(y[656]), .Z(n549) );
  XNOR U2436 ( .A(x[1902]), .B(y[1902]), .Z(n550) );
  XNOR U2437 ( .A(n549), .B(n550), .Z(n551) );
  XOR U2438 ( .A(n552), .B(n551), .Z(n2112) );
  XOR U2439 ( .A(x[626]), .B(y[626]), .Z(n2948) );
  XOR U2440 ( .A(x[491]), .B(y[491]), .Z(n2945) );
  XNOR U2441 ( .A(x[630]), .B(y[630]), .Z(n2946) );
  XNOR U2442 ( .A(n2945), .B(n2946), .Z(n2947) );
  XNOR U2443 ( .A(n2948), .B(n2947), .Z(n2111) );
  XNOR U2444 ( .A(n2112), .B(n2111), .Z(n2113) );
  XOR U2445 ( .A(n2114), .B(n2113), .Z(n4153) );
  XNOR U2446 ( .A(n4152), .B(n4153), .Z(n4155) );
  XOR U2447 ( .A(x[622]), .B(y[622]), .Z(n648) );
  XOR U2448 ( .A(x[624]), .B(y[624]), .Z(n645) );
  XNOR U2449 ( .A(x[1917]), .B(y[1917]), .Z(n646) );
  XNOR U2450 ( .A(n645), .B(n646), .Z(n647) );
  XOR U2451 ( .A(n648), .B(n647), .Z(n2090) );
  XOR U2452 ( .A(x[1318]), .B(y[1318]), .Z(n5121) );
  XOR U2453 ( .A(x[57]), .B(y[57]), .Z(n5118) );
  XNOR U2454 ( .A(x[1320]), .B(y[1320]), .Z(n5119) );
  XNOR U2455 ( .A(n5118), .B(n5119), .Z(n5120) );
  XOR U2456 ( .A(n5121), .B(n5120), .Z(n2088) );
  XOR U2457 ( .A(x[610]), .B(y[610]), .Z(n642) );
  XOR U2458 ( .A(x[503]), .B(y[503]), .Z(n639) );
  XNOR U2459 ( .A(x[614]), .B(y[614]), .Z(n640) );
  XNOR U2460 ( .A(n639), .B(n640), .Z(n641) );
  XNOR U2461 ( .A(n642), .B(n641), .Z(n2087) );
  XNOR U2462 ( .A(n2088), .B(n2087), .Z(n2089) );
  XNOR U2463 ( .A(n2090), .B(n2089), .Z(n4154) );
  XNOR U2464 ( .A(n4155), .B(n4154), .Z(n4446) );
  XOR U2465 ( .A(n4447), .B(n4446), .Z(n4448) );
  XOR U2466 ( .A(n4449), .B(n4448), .Z(n4812) );
  XOR U2467 ( .A(n4813), .B(n4812), .Z(n4815) );
  XOR U2468 ( .A(x[554]), .B(y[554]), .Z(n1892) );
  XOR U2469 ( .A(x[556]), .B(y[556]), .Z(n1889) );
  XNOR U2470 ( .A(x[861]), .B(y[861]), .Z(n1890) );
  XNOR U2471 ( .A(n1889), .B(n1890), .Z(n1891) );
  XOR U2472 ( .A(n1892), .B(n1891), .Z(n1922) );
  XOR U2473 ( .A(x[1302]), .B(y[1302]), .Z(n4875) );
  XOR U2474 ( .A(x[461]), .B(y[461]), .Z(n4872) );
  XNOR U2475 ( .A(x[1304]), .B(y[1304]), .Z(n4873) );
  XNOR U2476 ( .A(n4872), .B(n4873), .Z(n4874) );
  XOR U2477 ( .A(n4875), .B(n4874), .Z(n1920) );
  XOR U2478 ( .A(x[542]), .B(y[542]), .Z(n1904) );
  XOR U2479 ( .A(x[544]), .B(y[544]), .Z(n1901) );
  XNOR U2480 ( .A(x[867]), .B(y[867]), .Z(n1902) );
  XNOR U2481 ( .A(n1901), .B(n1902), .Z(n1903) );
  XNOR U2482 ( .A(n1904), .B(n1903), .Z(n1919) );
  XNOR U2483 ( .A(n1920), .B(n1919), .Z(n1921) );
  XNOR U2484 ( .A(n1922), .B(n1921), .Z(n3924) );
  XOR U2485 ( .A(x[592]), .B(y[592]), .Z(n1958) );
  XOR U2486 ( .A(x[594]), .B(y[594]), .Z(n1955) );
  XNOR U2487 ( .A(x[1915]), .B(y[1915]), .Z(n1956) );
  XNOR U2488 ( .A(n1955), .B(n1956), .Z(n1957) );
  XOR U2489 ( .A(n1958), .B(n1957), .Z(n2120) );
  XOR U2490 ( .A(x[1310]), .B(y[1310]), .Z(n4881) );
  XOR U2491 ( .A(x[63]), .B(y[63]), .Z(n4878) );
  XNOR U2492 ( .A(x[1312]), .B(y[1312]), .Z(n4879) );
  XNOR U2493 ( .A(n4878), .B(n4879), .Z(n4880) );
  XOR U2494 ( .A(n4881), .B(n4880), .Z(n2118) );
  XOR U2495 ( .A(x[580]), .B(y[580]), .Z(n1946) );
  XOR U2496 ( .A(x[517]), .B(y[517]), .Z(n1943) );
  XNOR U2497 ( .A(x[584]), .B(y[584]), .Z(n1944) );
  XNOR U2498 ( .A(n1943), .B(n1944), .Z(n1945) );
  XNOR U2499 ( .A(n1946), .B(n1945), .Z(n2117) );
  XNOR U2500 ( .A(n2118), .B(n2117), .Z(n2119) );
  XOR U2501 ( .A(n2120), .B(n2119), .Z(n3925) );
  XNOR U2502 ( .A(n3924), .B(n3925), .Z(n3926) );
  XOR U2503 ( .A(x[576]), .B(y[576]), .Z(n1952) );
  XOR U2504 ( .A(x[578]), .B(y[578]), .Z(n1949) );
  XNOR U2505 ( .A(x[1913]), .B(y[1913]), .Z(n1950) );
  XNOR U2506 ( .A(n1949), .B(n1950), .Z(n1951) );
  XOR U2507 ( .A(n1952), .B(n1951), .Z(n1964) );
  XOR U2508 ( .A(x[1910]), .B(y[1910]), .Z(n534) );
  XOR U2509 ( .A(x[1912]), .B(y[1912]), .Z(n531) );
  XNOR U2510 ( .A(x[1914]), .B(y[1914]), .Z(n532) );
  XNOR U2511 ( .A(n531), .B(n532), .Z(n533) );
  XOR U2512 ( .A(n534), .B(n533), .Z(n1962) );
  XOR U2513 ( .A(x[568]), .B(y[568]), .Z(n1898) );
  XOR U2514 ( .A(x[525]), .B(y[525]), .Z(n1895) );
  XNOR U2515 ( .A(x[574]), .B(y[574]), .Z(n1896) );
  XNOR U2516 ( .A(n1895), .B(n1896), .Z(n1897) );
  XNOR U2517 ( .A(n1898), .B(n1897), .Z(n1961) );
  XNOR U2518 ( .A(n1962), .B(n1961), .Z(n1963) );
  XOR U2519 ( .A(n1964), .B(n1963), .Z(n3927) );
  XNOR U2520 ( .A(n3926), .B(n3927), .Z(n4593) );
  XOR U2521 ( .A(x[486]), .B(y[486]), .Z(n790) );
  XOR U2522 ( .A(x[488]), .B(y[488]), .Z(n788) );
  XOR U2523 ( .A(x[1907]), .B(y[1907]), .Z(n787) );
  XOR U2524 ( .A(n788), .B(n787), .Z(n789) );
  XOR U2525 ( .A(n790), .B(n789), .Z(n934) );
  XOR U2526 ( .A(x[1286]), .B(y[1286]), .Z(n4725) );
  XOR U2527 ( .A(x[79]), .B(y[79]), .Z(n4723) );
  XOR U2528 ( .A(x[1288]), .B(y[1288]), .Z(n4722) );
  XOR U2529 ( .A(n4723), .B(n4722), .Z(n4724) );
  XOR U2530 ( .A(n4725), .B(n4724), .Z(n932) );
  XOR U2531 ( .A(x[482]), .B(y[482]), .Z(n796) );
  XOR U2532 ( .A(x[484]), .B(y[484]), .Z(n794) );
  XOR U2533 ( .A(x[573]), .B(y[573]), .Z(n793) );
  XOR U2534 ( .A(n794), .B(n793), .Z(n795) );
  XNOR U2535 ( .A(n796), .B(n795), .Z(n931) );
  XNOR U2536 ( .A(n932), .B(n931), .Z(n933) );
  XNOR U2537 ( .A(n934), .B(n933), .Z(n4938) );
  XOR U2538 ( .A(x[476]), .B(y[476]), .Z(n820) );
  XOR U2539 ( .A(x[478]), .B(y[478]), .Z(n818) );
  XOR U2540 ( .A(x[1905]), .B(y[1905]), .Z(n817) );
  XOR U2541 ( .A(n818), .B(n817), .Z(n819) );
  XOR U2542 ( .A(n820), .B(n819), .Z(n880) );
  XOR U2543 ( .A(x[1924]), .B(y[1924]), .Z(n3548) );
  XOR U2544 ( .A(x[678]), .B(y[678]), .Z(n3546) );
  XOR U2545 ( .A(x[1926]), .B(y[1926]), .Z(n3545) );
  XOR U2546 ( .A(n3546), .B(n3545), .Z(n3547) );
  XOR U2547 ( .A(n3548), .B(n3547), .Z(n878) );
  XOR U2548 ( .A(x[468]), .B(y[468]), .Z(n808) );
  XOR U2549 ( .A(x[470]), .B(y[470]), .Z(n806) );
  XOR U2550 ( .A(x[579]), .B(y[579]), .Z(n805) );
  XOR U2551 ( .A(n806), .B(n805), .Z(n807) );
  XNOR U2552 ( .A(n808), .B(n807), .Z(n877) );
  XNOR U2553 ( .A(n878), .B(n877), .Z(n879) );
  XOR U2554 ( .A(n880), .B(n879), .Z(n4939) );
  XNOR U2555 ( .A(n4938), .B(n4939), .Z(n4940) );
  XOR U2556 ( .A(x[464]), .B(y[464]), .Z(n814) );
  XOR U2557 ( .A(x[466]), .B(y[466]), .Z(n811) );
  XNOR U2558 ( .A(x[585]), .B(y[585]), .Z(n812) );
  XNOR U2559 ( .A(n811), .B(n812), .Z(n813) );
  XOR U2560 ( .A(n814), .B(n813), .Z(n1462) );
  XOR U2561 ( .A(x[1278]), .B(y[1278]), .Z(n4719) );
  XOR U2562 ( .A(x[85]), .B(y[85]), .Z(n4716) );
  XNOR U2563 ( .A(x[1280]), .B(y[1280]), .Z(n4717) );
  XNOR U2564 ( .A(n4716), .B(n4717), .Z(n4718) );
  XOR U2565 ( .A(n4719), .B(n4718), .Z(n1460) );
  XOR U2566 ( .A(x[460]), .B(y[460]), .Z(n682) );
  XOR U2567 ( .A(x[462]), .B(y[462]), .Z(n679) );
  XNOR U2568 ( .A(x[901]), .B(y[901]), .Z(n680) );
  XNOR U2569 ( .A(n679), .B(n680), .Z(n681) );
  XNOR U2570 ( .A(n682), .B(n681), .Z(n1459) );
  XNOR U2571 ( .A(n1460), .B(n1459), .Z(n1461) );
  XOR U2572 ( .A(n1462), .B(n1461), .Z(n4941) );
  XNOR U2573 ( .A(n4940), .B(n4941), .Z(n4590) );
  XOR U2574 ( .A(x[536]), .B(y[536]), .Z(n1910) );
  XOR U2575 ( .A(x[538]), .B(y[538]), .Z(n1907) );
  XNOR U2576 ( .A(x[1911]), .B(y[1911]), .Z(n1908) );
  XNOR U2577 ( .A(n1907), .B(n1908), .Z(n1909) );
  XOR U2578 ( .A(n1910), .B(n1909), .Z(n778) );
  XOR U2579 ( .A(x[1916]), .B(y[1916]), .Z(n3777) );
  XOR U2580 ( .A(x[936]), .B(y[936]), .Z(n3774) );
  XNOR U2581 ( .A(x[1918]), .B(y[1918]), .Z(n3775) );
  XNOR U2582 ( .A(n3774), .B(n3775), .Z(n3776) );
  XOR U2583 ( .A(n3777), .B(n3776), .Z(n776) );
  XOR U2584 ( .A(x[532]), .B(y[532]), .Z(n754) );
  XOR U2585 ( .A(x[534]), .B(y[534]), .Z(n751) );
  XNOR U2586 ( .A(x[545]), .B(y[545]), .Z(n752) );
  XNOR U2587 ( .A(n751), .B(n752), .Z(n753) );
  XNOR U2588 ( .A(n754), .B(n753), .Z(n775) );
  XNOR U2589 ( .A(n776), .B(n775), .Z(n777) );
  XNOR U2590 ( .A(n778), .B(n777), .Z(n3996) );
  XOR U2591 ( .A(x[528]), .B(y[528]), .Z(n742) );
  XOR U2592 ( .A(x[530]), .B(y[530]), .Z(n739) );
  XNOR U2593 ( .A(x[1909]), .B(y[1909]), .Z(n740) );
  XNOR U2594 ( .A(n739), .B(n740), .Z(n741) );
  XOR U2595 ( .A(n742), .B(n741), .Z(n826) );
  XOR U2596 ( .A(x[1294]), .B(y[1294]), .Z(n4731) );
  XOR U2597 ( .A(x[467]), .B(y[467]), .Z(n4728) );
  XNOR U2598 ( .A(x[1296]), .B(y[1296]), .Z(n4729) );
  XNOR U2599 ( .A(n4728), .B(n4729), .Z(n4730) );
  XOR U2600 ( .A(n4731), .B(n4730), .Z(n824) );
  XOR U2601 ( .A(x[522]), .B(y[522]), .Z(n748) );
  XOR U2602 ( .A(x[526]), .B(y[526]), .Z(n745) );
  XNOR U2603 ( .A(x[553]), .B(y[553]), .Z(n746) );
  XNOR U2604 ( .A(n745), .B(n746), .Z(n747) );
  XNOR U2605 ( .A(n748), .B(n747), .Z(n823) );
  XNOR U2606 ( .A(n824), .B(n823), .Z(n825) );
  XOR U2607 ( .A(n826), .B(n825), .Z(n3997) );
  XNOR U2608 ( .A(n3996), .B(n3997), .Z(n3998) );
  XOR U2609 ( .A(x[514]), .B(y[514]), .Z(n772) );
  XOR U2610 ( .A(x[518]), .B(y[518]), .Z(n770) );
  XOR U2611 ( .A(x[557]), .B(y[557]), .Z(n769) );
  XOR U2612 ( .A(n770), .B(n769), .Z(n771) );
  XOR U2613 ( .A(n772), .B(n771), .Z(n718) );
  XOR U2614 ( .A(x[1920]), .B(y[1920]), .Z(n3699) );
  XOR U2615 ( .A(x[672]), .B(y[672]), .Z(n3697) );
  XOR U2616 ( .A(x[1922]), .B(y[1922]), .Z(n3696) );
  XOR U2617 ( .A(n3697), .B(n3696), .Z(n3698) );
  XOR U2618 ( .A(n3699), .B(n3698), .Z(n716) );
  XOR U2619 ( .A(x[502]), .B(y[502]), .Z(n766) );
  XOR U2620 ( .A(x[506]), .B(y[506]), .Z(n764) );
  XOR U2621 ( .A(x[565]), .B(y[565]), .Z(n763) );
  XOR U2622 ( .A(n764), .B(n763), .Z(n765) );
  XNOR U2623 ( .A(n766), .B(n765), .Z(n715) );
  XNOR U2624 ( .A(n716), .B(n715), .Z(n717) );
  XOR U2625 ( .A(n718), .B(n717), .Z(n3999) );
  XNOR U2626 ( .A(n3998), .B(n3999), .Z(n4591) );
  XOR U2627 ( .A(n4590), .B(n4591), .Z(n4592) );
  XOR U2628 ( .A(n4593), .B(n4592), .Z(n4814) );
  XNOR U2629 ( .A(n4815), .B(n4814), .Z(n4599) );
  XOR U2630 ( .A(x[312]), .B(y[312]), .Z(n922) );
  XOR U2631 ( .A(x[314]), .B(y[314]), .Z(n919) );
  XNOR U2632 ( .A(x[1891]), .B(y[1891]), .Z(n920) );
  XNOR U2633 ( .A(n919), .B(n920), .Z(n921) );
  XOR U2634 ( .A(n922), .B(n921), .Z(n1600) );
  XOR U2635 ( .A(x[1950]), .B(y[1950]), .Z(n5283) );
  XOR U2636 ( .A(x[702]), .B(y[702]), .Z(n5280) );
  XNOR U2637 ( .A(x[1952]), .B(y[1952]), .Z(n5281) );
  XNOR U2638 ( .A(n5280), .B(n5281), .Z(n5282) );
  XOR U2639 ( .A(n5283), .B(n5282), .Z(n1598) );
  XOR U2640 ( .A(x[300]), .B(y[300]), .Z(n2450) );
  XOR U2641 ( .A(x[304]), .B(y[304]), .Z(n2447) );
  XNOR U2642 ( .A(x[1889]), .B(y[1889]), .Z(n2448) );
  XNOR U2643 ( .A(n2447), .B(n2448), .Z(n2449) );
  XNOR U2644 ( .A(n2450), .B(n2449), .Z(n1597) );
  XNOR U2645 ( .A(n1598), .B(n1597), .Z(n1599) );
  XNOR U2646 ( .A(n1600), .B(n1599), .Z(n3948) );
  XOR U2647 ( .A(x[324]), .B(y[324]), .Z(n928) );
  XOR U2648 ( .A(x[328]), .B(y[328]), .Z(n926) );
  XOR U2649 ( .A(x[675]), .B(y[675]), .Z(n925) );
  XOR U2650 ( .A(n926), .B(n925), .Z(n927) );
  XOR U2651 ( .A(n928), .B(n927), .Z(n1856) );
  XOR U2652 ( .A(x[1238]), .B(y[1238]), .Z(n5061) );
  XOR U2653 ( .A(x[501]), .B(y[501]), .Z(n5059) );
  XOR U2654 ( .A(x[1240]), .B(y[1240]), .Z(n5058) );
  XOR U2655 ( .A(n5059), .B(n5058), .Z(n5060) );
  XOR U2656 ( .A(n5061), .B(n5060), .Z(n1854) );
  XOR U2657 ( .A(x[316]), .B(y[316]), .Z(n2564) );
  XOR U2658 ( .A(x[320]), .B(y[320]), .Z(n2562) );
  XOR U2659 ( .A(x[967]), .B(y[967]), .Z(n2561) );
  XOR U2660 ( .A(n2562), .B(n2561), .Z(n2563) );
  XNOR U2661 ( .A(n2564), .B(n2563), .Z(n1853) );
  XNOR U2662 ( .A(n1854), .B(n1853), .Z(n1855) );
  XOR U2663 ( .A(n1856), .B(n1855), .Z(n3949) );
  XNOR U2664 ( .A(n3948), .B(n3949), .Z(n3951) );
  XOR U2665 ( .A(x[290]), .B(y[290]), .Z(n2420) );
  XOR U2666 ( .A(x[292]), .B(y[292]), .Z(n2417) );
  XNOR U2667 ( .A(x[695]), .B(y[695]), .Z(n2418) );
  XNOR U2668 ( .A(n2417), .B(n2418), .Z(n2419) );
  XOR U2669 ( .A(n2420), .B(n2419), .Z(n1660) );
  XOR U2670 ( .A(x[1230]), .B(y[1230]), .Z(n5049) );
  XOR U2671 ( .A(x[507]), .B(y[507]), .Z(n5046) );
  XNOR U2672 ( .A(x[1232]), .B(y[1232]), .Z(n5047) );
  XNOR U2673 ( .A(n5046), .B(n5047), .Z(n5048) );
  XOR U2674 ( .A(n5049), .B(n5048), .Z(n1658) );
  XOR U2675 ( .A(x[286]), .B(y[286]), .Z(n2390) );
  XOR U2676 ( .A(x[288]), .B(y[288]), .Z(n2387) );
  XNOR U2677 ( .A(x[981]), .B(y[981]), .Z(n2388) );
  XNOR U2678 ( .A(n2387), .B(n2388), .Z(n2389) );
  XNOR U2679 ( .A(n2390), .B(n2389), .Z(n1657) );
  XNOR U2680 ( .A(n1658), .B(n1657), .Z(n1659) );
  XNOR U2681 ( .A(n1660), .B(n1659), .Z(n3950) );
  XNOR U2682 ( .A(n3951), .B(n3950), .Z(n4239) );
  XOR U2683 ( .A(x[254]), .B(y[254]), .Z(n2366) );
  XOR U2684 ( .A(x[258]), .B(y[258]), .Z(n2363) );
  XNOR U2685 ( .A(x[717]), .B(y[717]), .Z(n2364) );
  XNOR U2686 ( .A(n2363), .B(n2364), .Z(n2365) );
  XOR U2687 ( .A(n2366), .B(n2365), .Z(n1720) );
  XOR U2688 ( .A(x[1958]), .B(y[1958]), .Z(n3416) );
  XOR U2689 ( .A(x[1960]), .B(y[1960]), .Z(n3413) );
  XNOR U2690 ( .A(x[1962]), .B(y[1962]), .Z(n3414) );
  XNOR U2691 ( .A(n3413), .B(n3414), .Z(n3415) );
  XOR U2692 ( .A(n3416), .B(n3415), .Z(n1718) );
  XOR U2693 ( .A(x[244]), .B(y[244]), .Z(n2780) );
  XOR U2694 ( .A(x[246]), .B(y[246]), .Z(n2777) );
  XNOR U2695 ( .A(x[1001]), .B(y[1001]), .Z(n2778) );
  XNOR U2696 ( .A(n2777), .B(n2778), .Z(n2779) );
  XNOR U2697 ( .A(n2780), .B(n2779), .Z(n1717) );
  XNOR U2698 ( .A(n1718), .B(n1717), .Z(n1719) );
  XNOR U2699 ( .A(n1720), .B(n1719), .Z(n3912) );
  XOR U2700 ( .A(x[226]), .B(y[226]), .Z(n2558) );
  XOR U2701 ( .A(x[228]), .B(y[228]), .Z(n2555) );
  XNOR U2702 ( .A(x[1883]), .B(y[1883]), .Z(n2556) );
  XNOR U2703 ( .A(n2555), .B(n2556), .Z(n2557) );
  XOR U2704 ( .A(n2558), .B(n2557), .Z(n5661) );
  XOR U2705 ( .A(x[1964]), .B(y[1964]), .Z(n5709) );
  XOR U2706 ( .A(x[714]), .B(y[714]), .Z(n5706) );
  XNOR U2707 ( .A(x[1966]), .B(y[1966]), .Z(n5707) );
  XNOR U2708 ( .A(n5706), .B(n5707), .Z(n5708) );
  XOR U2709 ( .A(n5709), .B(n5708), .Z(n5659) );
  XOR U2710 ( .A(x[222]), .B(y[222]), .Z(n2750) );
  XOR U2711 ( .A(x[224]), .B(y[224]), .Z(n2747) );
  XNOR U2712 ( .A(x[737]), .B(y[737]), .Z(n2748) );
  XNOR U2713 ( .A(n2747), .B(n2748), .Z(n2749) );
  XNOR U2714 ( .A(n2750), .B(n2749), .Z(n5658) );
  XNOR U2715 ( .A(n5659), .B(n5658), .Z(n5660) );
  XOR U2716 ( .A(n5661), .B(n5660), .Z(n3913) );
  XNOR U2717 ( .A(n3912), .B(n3913), .Z(n3915) );
  XOR U2718 ( .A(x[198]), .B(y[198]), .Z(n1642) );
  XOR U2719 ( .A(x[200]), .B(y[200]), .Z(n1639) );
  XNOR U2720 ( .A(x[757]), .B(y[757]), .Z(n1640) );
  XNOR U2721 ( .A(n1639), .B(n1640), .Z(n1641) );
  XOR U2722 ( .A(n1642), .B(n1641), .Z(n5505) );
  XOR U2723 ( .A(x[1968]), .B(y[1968]), .Z(n5703) );
  XOR U2724 ( .A(x[718]), .B(y[718]), .Z(n5700) );
  XNOR U2725 ( .A(x[1970]), .B(y[1970]), .Z(n5701) );
  XNOR U2726 ( .A(n5700), .B(n5701), .Z(n5702) );
  XOR U2727 ( .A(n5703), .B(n5702), .Z(n5503) );
  XOR U2728 ( .A(x[192]), .B(y[192]), .Z(n4137) );
  XOR U2729 ( .A(x[196]), .B(y[196]), .Z(n4134) );
  XNOR U2730 ( .A(x[1027]), .B(y[1027]), .Z(n4135) );
  XNOR U2731 ( .A(n4134), .B(n4135), .Z(n4136) );
  XNOR U2732 ( .A(n4137), .B(n4136), .Z(n5502) );
  XNOR U2733 ( .A(n5503), .B(n5502), .Z(n5504) );
  XNOR U2734 ( .A(n5505), .B(n5504), .Z(n3914) );
  XNOR U2735 ( .A(n3915), .B(n3914), .Z(n4237) );
  XOR U2736 ( .A(x[176]), .B(y[176]), .Z(n1060) );
  XOR U2737 ( .A(x[178]), .B(y[178]), .Z(n1057) );
  XNOR U2738 ( .A(x[1877]), .B(y[1877]), .Z(n1058) );
  XNOR U2739 ( .A(n1057), .B(n1058), .Z(n1059) );
  XOR U2740 ( .A(n1060), .B(n1059), .Z(n5967) );
  XOR U2741 ( .A(x[1972]), .B(y[1972]), .Z(n3320) );
  XOR U2742 ( .A(x[722]), .B(y[722]), .Z(n3317) );
  XNOR U2743 ( .A(x[1974]), .B(y[1974]), .Z(n3318) );
  XNOR U2744 ( .A(n3317), .B(n3318), .Z(n3319) );
  XOR U2745 ( .A(n3320), .B(n3319), .Z(n5965) );
  XOR U2746 ( .A(x[172]), .B(y[172]), .Z(n1612) );
  XOR U2747 ( .A(x[174]), .B(y[174]), .Z(n1609) );
  XNOR U2748 ( .A(x[773]), .B(y[773]), .Z(n1610) );
  XNOR U2749 ( .A(n1609), .B(n1610), .Z(n1611) );
  XNOR U2750 ( .A(n1612), .B(n1611), .Z(n5964) );
  XNOR U2751 ( .A(n5965), .B(n5964), .Z(n5966) );
  XNOR U2752 ( .A(n5967), .B(n5966), .Z(n4524) );
  XOR U2753 ( .A(x[164]), .B(y[164]), .Z(n1480) );
  XOR U2754 ( .A(x[166]), .B(y[166]), .Z(n1477) );
  XNOR U2755 ( .A(x[1041]), .B(y[1041]), .Z(n1478) );
  XNOR U2756 ( .A(n1477), .B(n1478), .Z(n1479) );
  XOR U2757 ( .A(n1480), .B(n1479), .Z(n1564) );
  XOR U2758 ( .A(x[1190]), .B(y[1190]), .Z(n916) );
  XOR U2759 ( .A(x[145]), .B(y[145]), .Z(n913) );
  XNOR U2760 ( .A(x[1192]), .B(y[1192]), .Z(n914) );
  XNOR U2761 ( .A(n913), .B(n914), .Z(n915) );
  XOR U2762 ( .A(n916), .B(n915), .Z(n1562) );
  XOR U2763 ( .A(x[156]), .B(y[156]), .Z(n4215) );
  XOR U2764 ( .A(x[158]), .B(y[158]), .Z(n4212) );
  XNOR U2765 ( .A(x[1047]), .B(y[1047]), .Z(n4213) );
  XNOR U2766 ( .A(n4212), .B(n4213), .Z(n4214) );
  XNOR U2767 ( .A(n4215), .B(n4214), .Z(n1561) );
  XNOR U2768 ( .A(n1562), .B(n1561), .Z(n1563) );
  XOR U2769 ( .A(n1564), .B(n1563), .Z(n4525) );
  XNOR U2770 ( .A(n4524), .B(n4525), .Z(n4527) );
  XOR U2771 ( .A(x[152]), .B(y[152]), .Z(n2324) );
  XOR U2772 ( .A(x[154]), .B(y[154]), .Z(n2321) );
  XNOR U2773 ( .A(x[1875]), .B(y[1875]), .Z(n2322) );
  XNOR U2774 ( .A(n2321), .B(n2322), .Z(n2323) );
  XOR U2775 ( .A(n2324), .B(n2323), .Z(n5823) );
  XOR U2776 ( .A(x[1976]), .B(y[1976]), .Z(n5115) );
  XOR U2777 ( .A(x[1978]), .B(y[1978]), .Z(n5112) );
  XNOR U2778 ( .A(x[1980]), .B(y[1980]), .Z(n5113) );
  XNOR U2779 ( .A(n5112), .B(n5113), .Z(n5114) );
  XOR U2780 ( .A(n5115), .B(n5114), .Z(n5821) );
  XOR U2781 ( .A(x[148]), .B(y[148]), .Z(n4479) );
  XOR U2782 ( .A(x[150]), .B(y[150]), .Z(n4476) );
  XNOR U2783 ( .A(x[793]), .B(y[793]), .Z(n4477) );
  XNOR U2784 ( .A(n4476), .B(n4477), .Z(n4478) );
  XNOR U2785 ( .A(n4479), .B(n4478), .Z(n5820) );
  XNOR U2786 ( .A(n5821), .B(n5820), .Z(n5822) );
  XNOR U2787 ( .A(n5823), .B(n5822), .Z(n4526) );
  XNOR U2788 ( .A(n4527), .B(n4526), .Z(n4236) );
  XOR U2789 ( .A(n4237), .B(n4236), .Z(n4238) );
  XNOR U2790 ( .A(n4239), .B(n4238), .Z(n4081) );
  XOR U2791 ( .A(x[446]), .B(y[446]), .Z(n700) );
  XOR U2792 ( .A(x[448]), .B(y[448]), .Z(n697) );
  XNOR U2793 ( .A(x[907]), .B(y[907]), .Z(n698) );
  XNOR U2794 ( .A(n697), .B(n698), .Z(n699) );
  XOR U2795 ( .A(n700), .B(n699), .Z(n1784) );
  XOR U2796 ( .A(x[1928]), .B(y[1928]), .Z(n3434) );
  XOR U2797 ( .A(x[1930]), .B(y[1930]), .Z(n3431) );
  XNOR U2798 ( .A(x[1932]), .B(y[1932]), .Z(n3432) );
  XNOR U2799 ( .A(n3431), .B(n3432), .Z(n3433) );
  XOR U2800 ( .A(n3434), .B(n3433), .Z(n1782) );
  XOR U2801 ( .A(x[432]), .B(y[432]), .Z(n910) );
  XOR U2802 ( .A(x[436]), .B(y[436]), .Z(n907) );
  XNOR U2803 ( .A(x[599]), .B(y[599]), .Z(n908) );
  XNOR U2804 ( .A(n907), .B(n908), .Z(n909) );
  XNOR U2805 ( .A(n910), .B(n909), .Z(n1781) );
  XNOR U2806 ( .A(n1782), .B(n1781), .Z(n1783) );
  XNOR U2807 ( .A(n1784), .B(n1783), .Z(n4806) );
  XOR U2808 ( .A(x[426]), .B(y[426]), .Z(n904) );
  XOR U2809 ( .A(x[428]), .B(y[428]), .Z(n901) );
  XNOR U2810 ( .A(x[1901]), .B(y[1901]), .Z(n902) );
  XNOR U2811 ( .A(n901), .B(n902), .Z(n903) );
  XOR U2812 ( .A(n904), .B(n903), .Z(n1516) );
  XOR U2813 ( .A(x[1270]), .B(y[1270]), .Z(n361) );
  XOR U2814 ( .A(x[481]), .B(y[481]), .Z(n358) );
  XNOR U2815 ( .A(x[1272]), .B(y[1272]), .Z(n359) );
  XNOR U2816 ( .A(n358), .B(n359), .Z(n360) );
  XOR U2817 ( .A(n361), .B(n360), .Z(n1514) );
  XOR U2818 ( .A(x[422]), .B(y[422]), .Z(n2138) );
  XOR U2819 ( .A(x[424]), .B(y[424]), .Z(n2136) );
  XOR U2820 ( .A(x[609]), .B(y[609]), .Z(n2135) );
  XOR U2821 ( .A(n2136), .B(n2135), .Z(n2137) );
  XNOR U2822 ( .A(n2138), .B(n2137), .Z(n1513) );
  XNOR U2823 ( .A(n1514), .B(n1513), .Z(n1515) );
  XOR U2824 ( .A(n1516), .B(n1515), .Z(n4807) );
  XNOR U2825 ( .A(n4806), .B(n4807), .Z(n4808) );
  XOR U2826 ( .A(x[418]), .B(y[418]), .Z(n2132) );
  XOR U2827 ( .A(x[420]), .B(y[420]), .Z(n2130) );
  XOR U2828 ( .A(x[613]), .B(y[613]), .Z(n2129) );
  XOR U2829 ( .A(n2130), .B(n2129), .Z(n2131) );
  XOR U2830 ( .A(n2132), .B(n2131), .Z(n1844) );
  XOR U2831 ( .A(x[1934]), .B(y[1934]), .Z(n3602) );
  XOR U2832 ( .A(x[950]), .B(y[950]), .Z(n3599) );
  XNOR U2833 ( .A(x[1936]), .B(y[1936]), .Z(n3600) );
  XNOR U2834 ( .A(n3599), .B(n3600), .Z(n3601) );
  XOR U2835 ( .A(n3602), .B(n3601), .Z(n1842) );
  XOR U2836 ( .A(x[412]), .B(y[412]), .Z(n2108) );
  XOR U2837 ( .A(x[416]), .B(y[416]), .Z(n2106) );
  XOR U2838 ( .A(x[921]), .B(y[921]), .Z(n2105) );
  XOR U2839 ( .A(n2106), .B(n2105), .Z(n2107) );
  XNOR U2840 ( .A(n2108), .B(n2107), .Z(n1841) );
  XNOR U2841 ( .A(n1842), .B(n1841), .Z(n1843) );
  XOR U2842 ( .A(n1844), .B(n1843), .Z(n4809) );
  XOR U2843 ( .A(n4808), .B(n4809), .Z(n4520) );
  XOR U2844 ( .A(x[406]), .B(y[406]), .Z(n2102) );
  XOR U2845 ( .A(x[410]), .B(y[410]), .Z(n2100) );
  XOR U2846 ( .A(x[619]), .B(y[619]), .Z(n2099) );
  XOR U2847 ( .A(n2100), .B(n2099), .Z(n2101) );
  XOR U2848 ( .A(n2102), .B(n2101), .Z(n1820) );
  XOR U2849 ( .A(x[1262]), .B(y[1262]), .Z(n4971) );
  XOR U2850 ( .A(x[487]), .B(y[487]), .Z(n4968) );
  XNOR U2851 ( .A(x[1264]), .B(y[1264]), .Z(n4969) );
  XNOR U2852 ( .A(n4968), .B(n4969), .Z(n4970) );
  XOR U2853 ( .A(n4971), .B(n4970), .Z(n1818) );
  XOR U2854 ( .A(x[398]), .B(y[398]), .Z(n2072) );
  XOR U2855 ( .A(x[400]), .B(y[400]), .Z(n2069) );
  XNOR U2856 ( .A(x[1899]), .B(y[1899]), .Z(n2070) );
  XNOR U2857 ( .A(n2069), .B(n2070), .Z(n2071) );
  XNOR U2858 ( .A(n2072), .B(n2071), .Z(n1817) );
  XNOR U2859 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U2860 ( .A(n1820), .B(n1819), .Z(n4770) );
  XOR U2861 ( .A(x[386]), .B(y[386]), .Z(n2042) );
  XOR U2862 ( .A(x[390]), .B(y[390]), .Z(n2039) );
  XNOR U2863 ( .A(x[1897]), .B(y[1897]), .Z(n2040) );
  XNOR U2864 ( .A(n2039), .B(n2040), .Z(n2041) );
  XOR U2865 ( .A(n2042), .B(n2041), .Z(n1808) );
  XOR U2866 ( .A(x[1938]), .B(y[1938]), .Z(n3362) );
  XOR U2867 ( .A(x[954]), .B(y[954]), .Z(n3359) );
  XNOR U2868 ( .A(x[1940]), .B(y[1940]), .Z(n3360) );
  XNOR U2869 ( .A(n3359), .B(n3360), .Z(n3361) );
  XOR U2870 ( .A(n3362), .B(n3361), .Z(n1806) );
  XOR U2871 ( .A(x[380]), .B(y[380]), .Z(n2018) );
  XOR U2872 ( .A(x[382]), .B(y[382]), .Z(n2015) );
  XNOR U2873 ( .A(x[635]), .B(y[635]), .Z(n2016) );
  XNOR U2874 ( .A(n2015), .B(n2016), .Z(n2017) );
  XNOR U2875 ( .A(n2018), .B(n2017), .Z(n1805) );
  XNOR U2876 ( .A(n1806), .B(n1805), .Z(n1807) );
  XOR U2877 ( .A(n1808), .B(n1807), .Z(n4771) );
  XNOR U2878 ( .A(n4770), .B(n4771), .Z(n4772) );
  XOR U2879 ( .A(x[376]), .B(y[376]), .Z(n2012) );
  XOR U2880 ( .A(x[378]), .B(y[378]), .Z(n2010) );
  XOR U2881 ( .A(x[639]), .B(y[639]), .Z(n2009) );
  XOR U2882 ( .A(n2010), .B(n2009), .Z(n2011) );
  XOR U2883 ( .A(n2012), .B(n2011), .Z(n1738) );
  XOR U2884 ( .A(x[1254]), .B(y[1254]), .Z(n5067) );
  XOR U2885 ( .A(x[101]), .B(y[101]), .Z(n5065) );
  XOR U2886 ( .A(x[1256]), .B(y[1256]), .Z(n5064) );
  XOR U2887 ( .A(n5065), .B(n5064), .Z(n5066) );
  XOR U2888 ( .A(n5067), .B(n5066), .Z(n1736) );
  XOR U2889 ( .A(x[370]), .B(y[370]), .Z(n1988) );
  XOR U2890 ( .A(x[374]), .B(y[374]), .Z(n1986) );
  XOR U2891 ( .A(x[941]), .B(y[941]), .Z(n1985) );
  XOR U2892 ( .A(n1986), .B(n1985), .Z(n1987) );
  XNOR U2893 ( .A(n1988), .B(n1987), .Z(n1735) );
  XNOR U2894 ( .A(n1736), .B(n1735), .Z(n1737) );
  XOR U2895 ( .A(n1738), .B(n1737), .Z(n4773) );
  XOR U2896 ( .A(n4772), .B(n4773), .Z(n4519) );
  XOR U2897 ( .A(x[362]), .B(y[362]), .Z(n1982) );
  XOR U2898 ( .A(x[366]), .B(y[366]), .Z(n1980) );
  XOR U2899 ( .A(x[649]), .B(y[649]), .Z(n1979) );
  XOR U2900 ( .A(n1980), .B(n1979), .Z(n1981) );
  XOR U2901 ( .A(n1982), .B(n1981), .Z(n1762) );
  XOR U2902 ( .A(x[1942]), .B(y[1942]), .Z(n5997) );
  XOR U2903 ( .A(x[694]), .B(y[694]), .Z(n5995) );
  XOR U2904 ( .A(x[1944]), .B(y[1944]), .Z(n5994) );
  XOR U2905 ( .A(n5995), .B(n5994), .Z(n5996) );
  XOR U2906 ( .A(n5997), .B(n5996), .Z(n1760) );
  XOR U2907 ( .A(x[358]), .B(y[358]), .Z(n2228) );
  XOR U2908 ( .A(x[360]), .B(y[360]), .Z(n2226) );
  XOR U2909 ( .A(x[947]), .B(y[947]), .Z(n2225) );
  XOR U2910 ( .A(n2226), .B(n2225), .Z(n2227) );
  XNOR U2911 ( .A(n2228), .B(n2227), .Z(n1759) );
  XNOR U2912 ( .A(n1760), .B(n1759), .Z(n1761) );
  XNOR U2913 ( .A(n1762), .B(n1761), .Z(n4944) );
  XOR U2914 ( .A(x[350]), .B(y[350]), .Z(n2198) );
  XOR U2915 ( .A(x[352]), .B(y[352]), .Z(n2195) );
  XNOR U2916 ( .A(x[655]), .B(y[655]), .Z(n2196) );
  XNOR U2917 ( .A(n2195), .B(n2196), .Z(n2197) );
  XOR U2918 ( .A(n2198), .B(n2197), .Z(n1606) );
  XOR U2919 ( .A(x[1246]), .B(y[1246]), .Z(n5697) );
  XOR U2920 ( .A(x[107]), .B(y[107]), .Z(n5694) );
  XNOR U2921 ( .A(x[1248]), .B(y[1248]), .Z(n5695) );
  XNOR U2922 ( .A(n5694), .B(n5695), .Z(n5696) );
  XOR U2923 ( .A(n5697), .B(n5696), .Z(n1604) );
  XOR U2924 ( .A(x[338]), .B(y[338]), .Z(n2168) );
  XOR U2925 ( .A(x[340]), .B(y[340]), .Z(n2165) );
  XNOR U2926 ( .A(x[663]), .B(y[663]), .Z(n2166) );
  XNOR U2927 ( .A(n2165), .B(n2166), .Z(n2167) );
  XNOR U2928 ( .A(n2168), .B(n2167), .Z(n1603) );
  XNOR U2929 ( .A(n1604), .B(n1603), .Z(n1605) );
  XOR U2930 ( .A(n1606), .B(n1605), .Z(n4945) );
  XNOR U2931 ( .A(n4944), .B(n4945), .Z(n4946) );
  XOR U2932 ( .A(x[334]), .B(y[334]), .Z(n2162) );
  XOR U2933 ( .A(x[336]), .B(y[336]), .Z(n2160) );
  XOR U2934 ( .A(x[669]), .B(y[669]), .Z(n2159) );
  XOR U2935 ( .A(n2160), .B(n2159), .Z(n2161) );
  XOR U2936 ( .A(n2162), .B(n2161), .Z(n1880) );
  XOR U2937 ( .A(x[1946]), .B(y[1946]), .Z(n3230) );
  XOR U2938 ( .A(x[698]), .B(y[698]), .Z(n3228) );
  XOR U2939 ( .A(x[1948]), .B(y[1948]), .Z(n3227) );
  XOR U2940 ( .A(n3228), .B(n3227), .Z(n3229) );
  XOR U2941 ( .A(n3230), .B(n3229), .Z(n1878) );
  XOR U2942 ( .A(x[330]), .B(y[330]), .Z(n2690) );
  XOR U2943 ( .A(x[332]), .B(y[332]), .Z(n2688) );
  XOR U2944 ( .A(x[961]), .B(y[961]), .Z(n2687) );
  XOR U2945 ( .A(n2688), .B(n2687), .Z(n2689) );
  XNOR U2946 ( .A(n2690), .B(n2689), .Z(n1877) );
  XNOR U2947 ( .A(n1878), .B(n1877), .Z(n1879) );
  XOR U2948 ( .A(n1880), .B(n1879), .Z(n4947) );
  XOR U2949 ( .A(n4946), .B(n4947), .Z(n4518) );
  XNOR U2950 ( .A(n4519), .B(n4518), .Z(n4521) );
  XOR U2951 ( .A(n4520), .B(n4521), .Z(n4080) );
  XOR U2952 ( .A(n4081), .B(n4080), .Z(n4083) );
  XOR U2953 ( .A(x[136]), .B(y[136]), .Z(n3128) );
  XOR U2954 ( .A(x[138]), .B(y[138]), .Z(n3125) );
  XNOR U2955 ( .A(x[805]), .B(y[805]), .Z(n3126) );
  XNOR U2956 ( .A(n3125), .B(n3126), .Z(n3127) );
  XOR U2957 ( .A(n3128), .B(n3127), .Z(n4767) );
  XOR U2958 ( .A(x[1982]), .B(y[1982]), .Z(n5109) );
  XOR U2959 ( .A(x[1984]), .B(y[1984]), .Z(n5106) );
  XNOR U2960 ( .A(x[1986]), .B(y[1986]), .Z(n5107) );
  XNOR U2961 ( .A(n5106), .B(n5107), .Z(n5108) );
  XOR U2962 ( .A(n5109), .B(n5108), .Z(n4765) );
  XOR U2963 ( .A(x[128]), .B(y[128]), .Z(n3212) );
  XOR U2964 ( .A(x[130]), .B(y[130]), .Z(n3209) );
  XNOR U2965 ( .A(x[813]), .B(y[813]), .Z(n3210) );
  XNOR U2966 ( .A(n3209), .B(n3210), .Z(n3211) );
  XNOR U2967 ( .A(n3212), .B(n3211), .Z(n4764) );
  XNOR U2968 ( .A(n4765), .B(n4764), .Z(n4766) );
  XNOR U2969 ( .A(n4767), .B(n4766), .Z(n4230) );
  XOR U2970 ( .A(x[120]), .B(y[120]), .Z(n4497) );
  XOR U2971 ( .A(x[122]), .B(y[122]), .Z(n4494) );
  XNOR U2972 ( .A(x[1871]), .B(y[1871]), .Z(n4495) );
  XNOR U2973 ( .A(n4494), .B(n4495), .Z(n4496) );
  XOR U2974 ( .A(n4497), .B(n4496), .Z(n4695) );
  XOR U2975 ( .A(x[1174]), .B(y[1174]), .Z(n2306) );
  XOR U2976 ( .A(x[541]), .B(y[541]), .Z(n2303) );
  XNOR U2977 ( .A(x[1176]), .B(y[1176]), .Z(n2304) );
  XNOR U2978 ( .A(n2303), .B(n2304), .Z(n2305) );
  XOR U2979 ( .A(n2306), .B(n2305), .Z(n4693) );
  XOR U2980 ( .A(x[116]), .B(y[116]), .Z(n2828) );
  XOR U2981 ( .A(x[118]), .B(y[118]), .Z(n2825) );
  XNOR U2982 ( .A(x[819]), .B(y[819]), .Z(n2826) );
  XNOR U2983 ( .A(n2825), .B(n2826), .Z(n2827) );
  XNOR U2984 ( .A(n2828), .B(n2827), .Z(n4692) );
  XNOR U2985 ( .A(n4693), .B(n4692), .Z(n4694) );
  XOR U2986 ( .A(n4695), .B(n4694), .Z(n4231) );
  XNOR U2987 ( .A(n4230), .B(n4231), .Z(n4232) );
  XOR U2988 ( .A(x[144]), .B(y[144]), .Z(n2552) );
  XOR U2989 ( .A(x[146]), .B(y[146]), .Z(n2549) );
  XNOR U2990 ( .A(x[1873]), .B(y[1873]), .Z(n2550) );
  XNOR U2991 ( .A(n2549), .B(n2550), .Z(n2551) );
  XOR U2992 ( .A(n2552), .B(n2551), .Z(n5493) );
  XOR U2993 ( .A(x[1182]), .B(y[1182]), .Z(n2414) );
  XOR U2994 ( .A(x[151]), .B(y[151]), .Z(n2411) );
  XNOR U2995 ( .A(x[1184]), .B(y[1184]), .Z(n2412) );
  XNOR U2996 ( .A(n2411), .B(n2412), .Z(n2413) );
  XOR U2997 ( .A(n2414), .B(n2413), .Z(n5491) );
  XOR U2998 ( .A(x[140]), .B(y[140]), .Z(n3134) );
  XOR U2999 ( .A(x[142]), .B(y[142]), .Z(n3131) );
  XNOR U3000 ( .A(x[799]), .B(y[799]), .Z(n3132) );
  XNOR U3001 ( .A(n3131), .B(n3132), .Z(n3133) );
  XNOR U3002 ( .A(n3134), .B(n3133), .Z(n5490) );
  XNOR U3003 ( .A(n5491), .B(n5490), .Z(n5492) );
  XOR U3004 ( .A(n5493), .B(n5492), .Z(n4233) );
  XNOR U3005 ( .A(n4232), .B(n4233), .Z(n4833) );
  XOR U3006 ( .A(x[102]), .B(y[102]), .Z(n3680) );
  XOR U3007 ( .A(x[104]), .B(y[104]), .Z(n3677) );
  XNOR U3008 ( .A(x[106]), .B(y[106]), .Z(n3678) );
  XNOR U3009 ( .A(n3677), .B(n3678), .Z(n3679) );
  XOR U3010 ( .A(n3680), .B(n3679), .Z(n5499) );
  XOR U3011 ( .A(x[1166]), .B(y[1166]), .Z(n2768) );
  XOR U3012 ( .A(x[547]), .B(y[547]), .Z(n2765) );
  XNOR U3013 ( .A(x[1168]), .B(y[1168]), .Z(n2766) );
  XNOR U3014 ( .A(n2765), .B(n2766), .Z(n2767) );
  XOR U3015 ( .A(n2768), .B(n2767), .Z(n5497) );
  XOR U3016 ( .A(x[96]), .B(y[96]), .Z(n2498) );
  XOR U3017 ( .A(x[98]), .B(y[98]), .Z(n2495) );
  XNOR U3018 ( .A(x[100]), .B(y[100]), .Z(n2496) );
  XNOR U3019 ( .A(n2495), .B(n2496), .Z(n2497) );
  XNOR U3020 ( .A(n2498), .B(n2497), .Z(n5496) );
  XNOR U3021 ( .A(n5497), .B(n5496), .Z(n5498) );
  XNOR U3022 ( .A(n5499), .B(n5498), .Z(n4170) );
  XOR U3023 ( .A(x[88]), .B(y[88]), .Z(n2594) );
  XOR U3024 ( .A(x[90]), .B(y[90]), .Z(n2591) );
  XNOR U3025 ( .A(x[485]), .B(y[485]), .Z(n2592) );
  XNOR U3026 ( .A(n2591), .B(n2592), .Z(n2593) );
  XOR U3027 ( .A(n2594), .B(n2593), .Z(n5529) );
  XOR U3028 ( .A(x[1992]), .B(y[1992]), .Z(n3464) );
  XOR U3029 ( .A(x[738]), .B(y[738]), .Z(n3461) );
  XNOR U3030 ( .A(x[1994]), .B(y[1994]), .Z(n3462) );
  XNOR U3031 ( .A(n3461), .B(n3462), .Z(n3463) );
  XOR U3032 ( .A(n3464), .B(n3463), .Z(n5527) );
  XOR U3033 ( .A(x[76]), .B(y[76]), .Z(n4053) );
  XOR U3034 ( .A(x[78]), .B(y[78]), .Z(n4050) );
  XNOR U3035 ( .A(x[80]), .B(y[80]), .Z(n4051) );
  XNOR U3036 ( .A(n4050), .B(n4051), .Z(n4052) );
  XNOR U3037 ( .A(n4053), .B(n4052), .Z(n5526) );
  XNOR U3038 ( .A(n5527), .B(n5526), .Z(n5528) );
  XOR U3039 ( .A(n5529), .B(n5528), .Z(n4171) );
  XNOR U3040 ( .A(n4170), .B(n4171), .Z(n4172) );
  XOR U3041 ( .A(x[112]), .B(y[112]), .Z(n4269) );
  XOR U3042 ( .A(x[114]), .B(y[114]), .Z(n4266) );
  XNOR U3043 ( .A(x[1869]), .B(y[1869]), .Z(n4267) );
  XNOR U3044 ( .A(n4266), .B(n4267), .Z(n4268) );
  XOR U3045 ( .A(n4269), .B(n4268), .Z(n4761) );
  XOR U3046 ( .A(x[1988]), .B(y[1988]), .Z(n3470) );
  XOR U3047 ( .A(x[992]), .B(y[992]), .Z(n3467) );
  XNOR U3048 ( .A(x[1990]), .B(y[1990]), .Z(n3468) );
  XNOR U3049 ( .A(n3467), .B(n3468), .Z(n3469) );
  XOR U3050 ( .A(n3470), .B(n3469), .Z(n4759) );
  XOR U3051 ( .A(x[108]), .B(y[108]), .Z(n3686) );
  XOR U3052 ( .A(x[110]), .B(y[110]), .Z(n3683) );
  XNOR U3053 ( .A(x[451]), .B(y[451]), .Z(n3684) );
  XNOR U3054 ( .A(n3683), .B(n3684), .Z(n3685) );
  XNOR U3055 ( .A(n3686), .B(n3685), .Z(n4758) );
  XNOR U3056 ( .A(n4759), .B(n4758), .Z(n4760) );
  XOR U3057 ( .A(n4761), .B(n4760), .Z(n4173) );
  XNOR U3058 ( .A(n4172), .B(n4173), .Z(n4831) );
  XOR U3059 ( .A(x[72]), .B(y[72]), .Z(n2720) );
  XOR U3060 ( .A(x[74]), .B(y[74]), .Z(n2717) );
  XNOR U3061 ( .A(x[513]), .B(y[513]), .Z(n2718) );
  XNOR U3062 ( .A(n2717), .B(n2718), .Z(n2719) );
  XOR U3063 ( .A(n2720), .B(n2719), .Z(n5589) );
  XOR U3064 ( .A(x[1158]), .B(y[1158]), .Z(n3122) );
  XOR U3065 ( .A(x[167]), .B(y[167]), .Z(n3119) );
  XNOR U3066 ( .A(x[1160]), .B(y[1160]), .Z(n3120) );
  XNOR U3067 ( .A(n3119), .B(n3120), .Z(n3121) );
  XOR U3068 ( .A(n3122), .B(n3121), .Z(n5587) );
  XOR U3069 ( .A(x[68]), .B(y[68]), .Z(n4197) );
  XOR U3070 ( .A(x[70]), .B(y[70]), .Z(n4194) );
  XNOR U3071 ( .A(x[519]), .B(y[519]), .Z(n4195) );
  XNOR U3072 ( .A(n4194), .B(n4195), .Z(n4196) );
  XNOR U3073 ( .A(n4197), .B(n4196), .Z(n5586) );
  XNOR U3074 ( .A(n5587), .B(n5586), .Z(n5588) );
  XNOR U3075 ( .A(n5589), .B(n5588), .Z(n4584) );
  XOR U3076 ( .A(x[62]), .B(y[62]), .Z(n2714) );
  XOR U3077 ( .A(x[64]), .B(y[64]), .Z(n2711) );
  XNOR U3078 ( .A(x[66]), .B(y[66]), .Z(n2712) );
  XNOR U3079 ( .A(n2711), .B(n2712), .Z(n2713) );
  XOR U3080 ( .A(n2714), .B(n2713), .Z(n125) );
  XOR U3081 ( .A(x[1996]), .B(y[1996]), .Z(n372) );
  XNOR U3082 ( .A(x[748]), .B(y[748]), .Z(n370) );
  XNOR U3083 ( .A(oglobal[0]), .B(n370), .Z(n371) );
  XOR U3084 ( .A(n372), .B(n371), .Z(n123) );
  XOR U3085 ( .A(x[56]), .B(y[56]), .Z(n113) );
  XOR U3086 ( .A(x[58]), .B(y[58]), .Z(n110) );
  XNOR U3087 ( .A(x[60]), .B(y[60]), .Z(n111) );
  XNOR U3088 ( .A(n110), .B(n111), .Z(n112) );
  XNOR U3089 ( .A(n113), .B(n112), .Z(n122) );
  XNOR U3090 ( .A(n123), .B(n122), .Z(n124) );
  XOR U3091 ( .A(n125), .B(n124), .Z(n4585) );
  XNOR U3092 ( .A(n4584), .B(n4585), .Z(n4586) );
  XOR U3093 ( .A(x[52]), .B(y[52]), .Z(n107) );
  XOR U3094 ( .A(x[54]), .B(y[54]), .Z(n104) );
  XNOR U3095 ( .A(x[549]), .B(y[549]), .Z(n105) );
  XNOR U3096 ( .A(n104), .B(n105), .Z(n106) );
  XOR U3097 ( .A(n107), .B(n106), .Z(n3741) );
  XOR U3098 ( .A(x[1150]), .B(y[1150]), .Z(n2822) );
  XOR U3099 ( .A(x[173]), .B(y[173]), .Z(n2819) );
  XNOR U3100 ( .A(x[1152]), .B(y[1152]), .Z(n2820) );
  XNOR U3101 ( .A(n2819), .B(n2820), .Z(n2821) );
  XOR U3102 ( .A(n2822), .B(n2821), .Z(n3739) );
  XOR U3103 ( .A(x[42]), .B(y[42]), .Z(n179) );
  XOR U3104 ( .A(x[44]), .B(y[44]), .Z(n176) );
  XNOR U3105 ( .A(x[46]), .B(y[46]), .Z(n177) );
  XNOR U3106 ( .A(n176), .B(n177), .Z(n178) );
  XNOR U3107 ( .A(n179), .B(n178), .Z(n3738) );
  XNOR U3108 ( .A(n3739), .B(n3738), .Z(n3740) );
  XOR U3109 ( .A(n3741), .B(n3740), .Z(n4587) );
  XNOR U3110 ( .A(n4586), .B(n4587), .Z(n4830) );
  XOR U3111 ( .A(n4831), .B(n4830), .Z(n4832) );
  XOR U3112 ( .A(n4833), .B(n4832), .Z(n4082) );
  XNOR U3113 ( .A(n4083), .B(n4082), .Z(n4597) );
  XOR U3114 ( .A(x[1189]), .B(y[1189]), .Z(n4059) );
  XOR U3115 ( .A(x[1185]), .B(y[1185]), .Z(n4056) );
  XNOR U3116 ( .A(x[1535]), .B(y[1535]), .Z(n4057) );
  XNOR U3117 ( .A(n4056), .B(n4057), .Z(n4058) );
  XOR U3118 ( .A(n4059), .B(n4058), .Z(n3692) );
  XOR U3119 ( .A(x[1193]), .B(y[1193]), .Z(n4209) );
  XOR U3120 ( .A(x[1191]), .B(y[1191]), .Z(n4206) );
  XNOR U3121 ( .A(x[1835]), .B(y[1835]), .Z(n4207) );
  XNOR U3122 ( .A(n4206), .B(n4207), .Z(n4208) );
  XOR U3123 ( .A(n4209), .B(n4208), .Z(n3690) );
  XOR U3124 ( .A(x[1197]), .B(y[1197]), .Z(n4203) );
  XOR U3125 ( .A(x[1195]), .B(y[1195]), .Z(n4200) );
  XNOR U3126 ( .A(x[1539]), .B(y[1539]), .Z(n4201) );
  XNOR U3127 ( .A(n4200), .B(n4201), .Z(n4202) );
  XNOR U3128 ( .A(n4203), .B(n4202), .Z(n3689) );
  XNOR U3129 ( .A(n3690), .B(n3689), .Z(n3691) );
  XNOR U3130 ( .A(n3692), .B(n3691), .Z(n721) );
  XOR U3131 ( .A(x[1533]), .B(y[1533]), .Z(n1678) );
  XOR U3132 ( .A(x[1525]), .B(y[1525]), .Z(n1675) );
  XNOR U3133 ( .A(x[1529]), .B(y[1529]), .Z(n1676) );
  XNOR U3134 ( .A(n1675), .B(n1676), .Z(n1677) );
  XOR U3135 ( .A(n1678), .B(n1677), .Z(n3380) );
  XOR U3136 ( .A(x[1545]), .B(y[1545]), .Z(n982) );
  XOR U3137 ( .A(x[1537]), .B(y[1537]), .Z(n979) );
  XNOR U3138 ( .A(x[1541]), .B(y[1541]), .Z(n980) );
  XNOR U3139 ( .A(n979), .B(n980), .Z(n981) );
  XOR U3140 ( .A(n982), .B(n981), .Z(n3378) );
  XOR U3141 ( .A(x[1557]), .B(y[1557]), .Z(n976) );
  XOR U3142 ( .A(x[1549]), .B(y[1549]), .Z(n973) );
  XNOR U3143 ( .A(x[1553]), .B(y[1553]), .Z(n974) );
  XNOR U3144 ( .A(n973), .B(n974), .Z(n975) );
  XNOR U3145 ( .A(n976), .B(n975), .Z(n3377) );
  XNOR U3146 ( .A(n3378), .B(n3377), .Z(n3379) );
  XOR U3147 ( .A(n3380), .B(n3379), .Z(n722) );
  XNOR U3148 ( .A(n721), .B(n722), .Z(n724) );
  XOR U3149 ( .A(x[1203]), .B(y[1203]), .Z(n4029) );
  XOR U3150 ( .A(x[1199]), .B(y[1199]), .Z(n4026) );
  XNOR U3151 ( .A(x[1833]), .B(y[1833]), .Z(n4027) );
  XNOR U3152 ( .A(n4026), .B(n4027), .Z(n4028) );
  XOR U3153 ( .A(n4029), .B(n4028), .Z(n2504) );
  XOR U3154 ( .A(x[1209]), .B(y[1209]), .Z(n4017) );
  XOR U3155 ( .A(x[1207]), .B(y[1207]), .Z(n4014) );
  XNOR U3156 ( .A(x[1543]), .B(y[1543]), .Z(n4015) );
  XNOR U3157 ( .A(n4014), .B(n4015), .Z(n4016) );
  XOR U3158 ( .A(n4017), .B(n4016), .Z(n2502) );
  XOR U3159 ( .A(x[1213]), .B(y[1213]), .Z(n4023) );
  XOR U3160 ( .A(x[1211]), .B(y[1211]), .Z(n4020) );
  XNOR U3161 ( .A(x[1831]), .B(y[1831]), .Z(n4021) );
  XNOR U3162 ( .A(n4020), .B(n4021), .Z(n4022) );
  XNOR U3163 ( .A(n4023), .B(n4022), .Z(n2501) );
  XNOR U3164 ( .A(n2502), .B(n2501), .Z(n2503) );
  XNOR U3165 ( .A(n2504), .B(n2503), .Z(n723) );
  XNOR U3166 ( .A(n724), .B(n723), .Z(n946) );
  XOR U3167 ( .A(x[1239]), .B(y[1239]), .Z(n5811) );
  XOR U3168 ( .A(x[1235]), .B(y[1235]), .Z(n5808) );
  XNOR U3169 ( .A(x[1555]), .B(y[1555]), .Z(n5809) );
  XNOR U3170 ( .A(n5808), .B(n5809), .Z(n5810) );
  XOR U3171 ( .A(n5811), .B(n5810), .Z(n119) );
  XOR U3172 ( .A(x[1245]), .B(y[1245]), .Z(n5655) );
  XOR U3173 ( .A(x[1243]), .B(y[1243]), .Z(n5652) );
  XNOR U3174 ( .A(x[1825]), .B(y[1825]), .Z(n5653) );
  XNOR U3175 ( .A(n5652), .B(n5653), .Z(n5654) );
  XOR U3176 ( .A(n5655), .B(n5654), .Z(n117) );
  XOR U3177 ( .A(x[1249]), .B(y[1249]), .Z(n5649) );
  XOR U3178 ( .A(x[1247]), .B(y[1247]), .Z(n5646) );
  XNOR U3179 ( .A(x[1559]), .B(y[1559]), .Z(n5647) );
  XNOR U3180 ( .A(n5646), .B(n5647), .Z(n5648) );
  XNOR U3181 ( .A(n5649), .B(n5648), .Z(n116) );
  XNOR U3182 ( .A(n117), .B(n116), .Z(n118) );
  XNOR U3183 ( .A(n119), .B(n118), .Z(n268) );
  XOR U3184 ( .A(x[1485]), .B(y[1485]), .Z(n1156) );
  XOR U3185 ( .A(x[1477]), .B(y[1477]), .Z(n1153) );
  XNOR U3186 ( .A(x[1481]), .B(y[1481]), .Z(n1154) );
  XNOR U3187 ( .A(n1153), .B(n1154), .Z(n1155) );
  XOR U3188 ( .A(n1156), .B(n1155), .Z(n3452) );
  XOR U3189 ( .A(x[269]), .B(y[269]), .Z(n3440) );
  XOR U3190 ( .A(x[263]), .B(y[263]), .Z(n3437) );
  XNOR U3191 ( .A(x[267]), .B(y[267]), .Z(n3438) );
  XNOR U3192 ( .A(n3437), .B(n3438), .Z(n3439) );
  XOR U3193 ( .A(n3440), .B(n3439), .Z(n3450) );
  XOR U3194 ( .A(x[1497]), .B(y[1497]), .Z(n1144) );
  XOR U3195 ( .A(x[1489]), .B(y[1489]), .Z(n1141) );
  XNOR U3196 ( .A(x[1493]), .B(y[1493]), .Z(n1142) );
  XNOR U3197 ( .A(n1141), .B(n1142), .Z(n1143) );
  XNOR U3198 ( .A(n1144), .B(n1143), .Z(n3449) );
  XNOR U3199 ( .A(n3450), .B(n3449), .Z(n3451) );
  XOR U3200 ( .A(n3452), .B(n3451), .Z(n269) );
  XNOR U3201 ( .A(n268), .B(n269), .Z(n271) );
  XOR U3202 ( .A(x[1253]), .B(y[1253]), .Z(n4263) );
  XOR U3203 ( .A(x[1251]), .B(y[1251]), .Z(n4260) );
  XNOR U3204 ( .A(x[1823]), .B(y[1823]), .Z(n4261) );
  XNOR U3205 ( .A(n4260), .B(n4261), .Z(n4262) );
  XOR U3206 ( .A(n4263), .B(n4262), .Z(n191) );
  XOR U3207 ( .A(x[1261]), .B(y[1261]), .Z(n4251) );
  XOR U3208 ( .A(x[1257]), .B(y[1257]), .Z(n4248) );
  XNOR U3209 ( .A(x[1563]), .B(y[1563]), .Z(n4249) );
  XNOR U3210 ( .A(n4248), .B(n4249), .Z(n4250) );
  XOR U3211 ( .A(n4251), .B(n4250), .Z(n189) );
  XOR U3212 ( .A(x[1265]), .B(y[1265]), .Z(n4257) );
  XOR U3213 ( .A(x[1263]), .B(y[1263]), .Z(n4254) );
  XNOR U3214 ( .A(x[1821]), .B(y[1821]), .Z(n4255) );
  XNOR U3215 ( .A(n4254), .B(n4255), .Z(n4256) );
  XNOR U3216 ( .A(n4257), .B(n4256), .Z(n188) );
  XNOR U3217 ( .A(n189), .B(n188), .Z(n190) );
  XNOR U3218 ( .A(n191), .B(n190), .Z(n270) );
  XNOR U3219 ( .A(n271), .B(n270), .Z(n944) );
  XOR U3220 ( .A(x[1217]), .B(y[1217]), .Z(n4131) );
  XOR U3221 ( .A(x[1215]), .B(y[1215]), .Z(n4128) );
  XNOR U3222 ( .A(x[1547]), .B(y[1547]), .Z(n4129) );
  XNOR U3223 ( .A(n4128), .B(n4129), .Z(n4130) );
  XOR U3224 ( .A(n4131), .B(n4130), .Z(n2600) );
  XOR U3225 ( .A(x[48]), .B(y[48]), .Z(n185) );
  XOR U3226 ( .A(x[50]), .B(y[50]), .Z(n182) );
  XNOR U3227 ( .A(x[555]), .B(y[555]), .Z(n183) );
  XNOR U3228 ( .A(n182), .B(n183), .Z(n184) );
  XOR U3229 ( .A(n185), .B(n184), .Z(n2598) );
  XOR U3230 ( .A(x[1225]), .B(y[1225]), .Z(n4119) );
  XOR U3231 ( .A(x[1221]), .B(y[1221]), .Z(n4116) );
  XNOR U3232 ( .A(x[1829]), .B(y[1829]), .Z(n4117) );
  XNOR U3233 ( .A(n4116), .B(n4117), .Z(n4118) );
  XNOR U3234 ( .A(n4119), .B(n4118), .Z(n2597) );
  XNOR U3235 ( .A(n2598), .B(n2597), .Z(n2599) );
  XNOR U3236 ( .A(n2600), .B(n2599), .Z(n829) );
  XOR U3237 ( .A(x[1509]), .B(y[1509]), .Z(n1150) );
  XOR U3238 ( .A(x[1501]), .B(y[1501]), .Z(n1147) );
  XNOR U3239 ( .A(x[1505]), .B(y[1505]), .Z(n1148) );
  XNOR U3240 ( .A(n1147), .B(n1148), .Z(n1149) );
  XOR U3241 ( .A(n1150), .B(n1149), .Z(n2642) );
  XOR U3242 ( .A(x[285]), .B(y[285]), .Z(n2630) );
  XOR U3243 ( .A(x[281]), .B(y[281]), .Z(n2628) );
  XOR U3244 ( .A(x[917]), .B(y[917]), .Z(n2627) );
  XOR U3245 ( .A(n2628), .B(n2627), .Z(n2629) );
  XOR U3246 ( .A(n2630), .B(n2629), .Z(n2640) );
  XOR U3247 ( .A(x[1521]), .B(y[1521]), .Z(n1684) );
  XOR U3248 ( .A(x[1513]), .B(y[1513]), .Z(n1681) );
  XNOR U3249 ( .A(x[1517]), .B(y[1517]), .Z(n1682) );
  XNOR U3250 ( .A(n1681), .B(n1682), .Z(n1683) );
  XNOR U3251 ( .A(n1684), .B(n1683), .Z(n2639) );
  XNOR U3252 ( .A(n2640), .B(n2639), .Z(n2641) );
  XOR U3253 ( .A(n2642), .B(n2641), .Z(n830) );
  XNOR U3254 ( .A(n829), .B(n830), .Z(n832) );
  XOR U3255 ( .A(x[1229]), .B(y[1229]), .Z(n4125) );
  XOR U3256 ( .A(x[1227]), .B(y[1227]), .Z(n4122) );
  XNOR U3257 ( .A(x[1551]), .B(y[1551]), .Z(n4123) );
  XNOR U3258 ( .A(n4122), .B(n4123), .Z(n4124) );
  XOR U3259 ( .A(n4125), .B(n4124), .Z(n2726) );
  XOR U3260 ( .A(x[36]), .B(y[36]), .Z(n355) );
  XOR U3261 ( .A(x[38]), .B(y[38]), .Z(n352) );
  XNOR U3262 ( .A(x[40]), .B(y[40]), .Z(n353) );
  XNOR U3263 ( .A(n352), .B(n353), .Z(n354) );
  XOR U3264 ( .A(n355), .B(n354), .Z(n2724) );
  XOR U3265 ( .A(x[1233]), .B(y[1233]), .Z(n5817) );
  XOR U3266 ( .A(x[1231]), .B(y[1231]), .Z(n5814) );
  XNOR U3267 ( .A(x[1827]), .B(y[1827]), .Z(n5815) );
  XNOR U3268 ( .A(n5814), .B(n5815), .Z(n5816) );
  XNOR U3269 ( .A(n5817), .B(n5816), .Z(n2723) );
  XNOR U3270 ( .A(n2724), .B(n2723), .Z(n2725) );
  XNOR U3271 ( .A(n2726), .B(n2725), .Z(n831) );
  XNOR U3272 ( .A(n832), .B(n831), .Z(n943) );
  XOR U3273 ( .A(n944), .B(n943), .Z(n945) );
  XNOR U3274 ( .A(n946), .B(n945), .Z(n663) );
  XOR U3275 ( .A(x[1117]), .B(y[1117]), .Z(n3861) );
  XOR U3276 ( .A(x[1113]), .B(y[1113]), .Z(n3858) );
  XNOR U3277 ( .A(x[1507]), .B(y[1507]), .Z(n3859) );
  XNOR U3278 ( .A(n3858), .B(n3859), .Z(n3860) );
  XOR U3279 ( .A(n3861), .B(n3860), .Z(n1366) );
  XOR U3280 ( .A(x[132]), .B(y[132]), .Z(n3218) );
  XOR U3281 ( .A(x[134]), .B(y[134]), .Z(n3215) );
  XNOR U3282 ( .A(x[1061]), .B(y[1061]), .Z(n3216) );
  XNOR U3283 ( .A(n3215), .B(n3216), .Z(n3217) );
  XOR U3284 ( .A(n3218), .B(n3217), .Z(n1364) );
  XOR U3285 ( .A(x[1121]), .B(y[1121]), .Z(n3849) );
  XOR U3286 ( .A(x[1119]), .B(y[1119]), .Z(n3846) );
  XNOR U3287 ( .A(x[1849]), .B(y[1849]), .Z(n3847) );
  XNOR U3288 ( .A(n3846), .B(n3847), .Z(n3848) );
  XNOR U3289 ( .A(n3849), .B(n3848), .Z(n1363) );
  XNOR U3290 ( .A(n1364), .B(n1363), .Z(n1365) );
  XNOR U3291 ( .A(n1366), .B(n1365), .Z(n883) );
  XOR U3292 ( .A(x[1615]), .B(y[1615]), .Z(n1354) );
  XOR U3293 ( .A(x[1611]), .B(y[1611]), .Z(n1351) );
  XNOR U3294 ( .A(x[1613]), .B(y[1613]), .Z(n1352) );
  XNOR U3295 ( .A(n1351), .B(n1352), .Z(n1353) );
  XOR U3296 ( .A(n1354), .B(n1353), .Z(n2684) );
  XOR U3297 ( .A(x[355]), .B(y[355]), .Z(n3260) );
  XOR U3298 ( .A(x[351]), .B(y[351]), .Z(n3257) );
  XNOR U3299 ( .A(x[969]), .B(y[969]), .Z(n3258) );
  XNOR U3300 ( .A(n3257), .B(n3258), .Z(n3259) );
  XOR U3301 ( .A(n3260), .B(n3259), .Z(n2682) );
  XOR U3302 ( .A(x[1621]), .B(y[1621]), .Z(n1048) );
  XOR U3303 ( .A(x[1617]), .B(y[1617]), .Z(n1045) );
  XNOR U3304 ( .A(x[1619]), .B(y[1619]), .Z(n1046) );
  XNOR U3305 ( .A(n1045), .B(n1046), .Z(n1047) );
  XNOR U3306 ( .A(n1048), .B(n1047), .Z(n2681) );
  XNOR U3307 ( .A(n2682), .B(n2681), .Z(n2683) );
  XOR U3308 ( .A(n2684), .B(n2683), .Z(n884) );
  XNOR U3309 ( .A(n883), .B(n884), .Z(n886) );
  XOR U3310 ( .A(x[1125]), .B(y[1125]), .Z(n3855) );
  XOR U3311 ( .A(x[1123]), .B(y[1123]), .Z(n3852) );
  XNOR U3312 ( .A(x[1511]), .B(y[1511]), .Z(n3853) );
  XNOR U3313 ( .A(n3852), .B(n3853), .Z(n3854) );
  XOR U3314 ( .A(n3855), .B(n3854), .Z(n1390) );
  XOR U3315 ( .A(x[124]), .B(y[124]), .Z(n2834) );
  XOR U3316 ( .A(x[126]), .B(y[126]), .Z(n2831) );
  XNOR U3317 ( .A(x[1067]), .B(y[1067]), .Z(n2832) );
  XNOR U3318 ( .A(n2831), .B(n2832), .Z(n2833) );
  XOR U3319 ( .A(n2834), .B(n2833), .Z(n1388) );
  XOR U3320 ( .A(x[1131]), .B(y[1131]), .Z(n4509) );
  XOR U3321 ( .A(x[1127]), .B(y[1127]), .Z(n4506) );
  XNOR U3322 ( .A(x[1847]), .B(y[1847]), .Z(n4507) );
  XNOR U3323 ( .A(n4506), .B(n4507), .Z(n4508) );
  XNOR U3324 ( .A(n4509), .B(n4508), .Z(n1387) );
  XNOR U3325 ( .A(n1388), .B(n1387), .Z(n1389) );
  XNOR U3326 ( .A(n1390), .B(n1389), .Z(n885) );
  XOR U3327 ( .A(n886), .B(n885), .Z(n1329) );
  XOR U3328 ( .A(x[1569]), .B(y[1569]), .Z(n1408) );
  XOR U3329 ( .A(x[1561]), .B(y[1561]), .Z(n1405) );
  XNOR U3330 ( .A(x[1565]), .B(y[1565]), .Z(n1406) );
  XNOR U3331 ( .A(n1405), .B(n1406), .Z(n1407) );
  XOR U3332 ( .A(n1408), .B(n1407), .Z(n3266) );
  XOR U3333 ( .A(x[1581]), .B(y[1581]), .Z(n1396) );
  XOR U3334 ( .A(x[1573]), .B(y[1573]), .Z(n1393) );
  XNOR U3335 ( .A(x[1577]), .B(y[1577]), .Z(n1394) );
  XNOR U3336 ( .A(n1393), .B(n1394), .Z(n1395) );
  XOR U3337 ( .A(n1396), .B(n1395), .Z(n3264) );
  XOR U3338 ( .A(x[1593]), .B(y[1593]), .Z(n1402) );
  XOR U3339 ( .A(x[1585]), .B(y[1585]), .Z(n1399) );
  XNOR U3340 ( .A(x[1589]), .B(y[1589]), .Z(n1400) );
  XNOR U3341 ( .A(n1399), .B(n1400), .Z(n1401) );
  XNOR U3342 ( .A(n1402), .B(n1401), .Z(n3263) );
  XNOR U3343 ( .A(n3264), .B(n3263), .Z(n3265) );
  XNOR U3344 ( .A(n3266), .B(n3265), .Z(n937) );
  XOR U3345 ( .A(x[1177]), .B(y[1177]), .Z(n4407) );
  XOR U3346 ( .A(x[1175]), .B(y[1175]), .Z(n4404) );
  XNOR U3347 ( .A(x[1531]), .B(y[1531]), .Z(n4405) );
  XNOR U3348 ( .A(n4404), .B(n4405), .Z(n4406) );
  XOR U3349 ( .A(n4407), .B(n4406), .Z(n2840) );
  XOR U3350 ( .A(x[82]), .B(y[82]), .Z(n2588) );
  XOR U3351 ( .A(x[84]), .B(y[84]), .Z(n2585) );
  XNOR U3352 ( .A(x[86]), .B(y[86]), .Z(n2586) );
  XNOR U3353 ( .A(n2585), .B(n2586), .Z(n2587) );
  XOR U3354 ( .A(n2588), .B(n2587), .Z(n2838) );
  XOR U3355 ( .A(x[1181]), .B(y[1181]), .Z(n4065) );
  XOR U3356 ( .A(x[1179]), .B(y[1179]), .Z(n4062) );
  XNOR U3357 ( .A(x[1837]), .B(y[1837]), .Z(n4063) );
  XNOR U3358 ( .A(n4062), .B(n4063), .Z(n4064) );
  XNOR U3359 ( .A(n4065), .B(n4064), .Z(n2837) );
  XNOR U3360 ( .A(n2838), .B(n2837), .Z(n2839) );
  XOR U3361 ( .A(n2840), .B(n2839), .Z(n938) );
  XNOR U3362 ( .A(n937), .B(n938), .Z(n940) );
  XOR U3363 ( .A(x[1167]), .B(y[1167]), .Z(n4413) );
  XOR U3364 ( .A(x[1163]), .B(y[1163]), .Z(n4410) );
  XNOR U3365 ( .A(x[1527]), .B(y[1527]), .Z(n4411) );
  XNOR U3366 ( .A(n4410), .B(n4411), .Z(n4412) );
  XOR U3367 ( .A(n4413), .B(n4412), .Z(n3224) );
  XOR U3368 ( .A(x[92]), .B(y[92]), .Z(n2492) );
  XOR U3369 ( .A(x[94]), .B(y[94]), .Z(n2489) );
  XNOR U3370 ( .A(x[477]), .B(y[477]), .Z(n2490) );
  XNOR U3371 ( .A(n2489), .B(n2490), .Z(n2491) );
  XOR U3372 ( .A(n2492), .B(n2491), .Z(n3222) );
  XOR U3373 ( .A(x[1173]), .B(y[1173]), .Z(n4401) );
  XOR U3374 ( .A(x[1171]), .B(y[1171]), .Z(n4398) );
  XNOR U3375 ( .A(x[1839]), .B(y[1839]), .Z(n4399) );
  XNOR U3376 ( .A(n4398), .B(n4399), .Z(n4400) );
  XNOR U3377 ( .A(n4401), .B(n4400), .Z(n3221) );
  XNOR U3378 ( .A(n3222), .B(n3221), .Z(n3223) );
  XNOR U3379 ( .A(n3224), .B(n3223), .Z(n939) );
  XOR U3380 ( .A(n940), .B(n939), .Z(n1328) );
  XOR U3381 ( .A(x[1137]), .B(y[1137]), .Z(n4503) );
  XOR U3382 ( .A(x[1135]), .B(y[1135]), .Z(n4500) );
  XNOR U3383 ( .A(x[1515]), .B(y[1515]), .Z(n4501) );
  XNOR U3384 ( .A(n4500), .B(n4501), .Z(n4502) );
  XOR U3385 ( .A(n4503), .B(n4502), .Z(n1006) );
  XOR U3386 ( .A(x[1141]), .B(y[1141]), .Z(n4281) );
  XOR U3387 ( .A(x[1139]), .B(y[1139]), .Z(n4278) );
  XNOR U3388 ( .A(x[1845]), .B(y[1845]), .Z(n4279) );
  XNOR U3389 ( .A(n4278), .B(n4279), .Z(n4280) );
  XOR U3390 ( .A(n4281), .B(n4280), .Z(n1004) );
  XOR U3391 ( .A(x[1145]), .B(y[1145]), .Z(n4275) );
  XOR U3392 ( .A(x[1143]), .B(y[1143]), .Z(n4272) );
  XNOR U3393 ( .A(x[1519]), .B(y[1519]), .Z(n4273) );
  XNOR U3394 ( .A(n4272), .B(n4273), .Z(n4274) );
  XNOR U3395 ( .A(n4275), .B(n4274), .Z(n1003) );
  XNOR U3396 ( .A(n1004), .B(n1003), .Z(n1005) );
  XNOR U3397 ( .A(n1006), .B(n1005), .Z(n835) );
  XOR U3398 ( .A(x[1603]), .B(y[1603]), .Z(n1360) );
  XOR U3399 ( .A(x[1597]), .B(y[1597]), .Z(n1357) );
  XNOR U3400 ( .A(x[1601]), .B(y[1601]), .Z(n1358) );
  XNOR U3401 ( .A(n1357), .B(n1358), .Z(n1359) );
  XOR U3402 ( .A(n1360), .B(n1359), .Z(n654) );
  XOR U3403 ( .A(x[341]), .B(y[341]), .Z(n3374) );
  XOR U3404 ( .A(x[335]), .B(y[335]), .Z(n3371) );
  XNOR U3405 ( .A(x[339]), .B(y[339]), .Z(n3372) );
  XNOR U3406 ( .A(n3371), .B(n3372), .Z(n3373) );
  XOR U3407 ( .A(n3374), .B(n3373), .Z(n652) );
  XOR U3408 ( .A(x[1609]), .B(y[1609]), .Z(n1348) );
  XOR U3409 ( .A(x[1605]), .B(y[1605]), .Z(n1345) );
  XNOR U3410 ( .A(x[1607]), .B(y[1607]), .Z(n1346) );
  XNOR U3411 ( .A(n1345), .B(n1346), .Z(n1347) );
  XNOR U3412 ( .A(n1348), .B(n1347), .Z(n651) );
  XNOR U3413 ( .A(n652), .B(n651), .Z(n653) );
  XOR U3414 ( .A(n654), .B(n653), .Z(n836) );
  XNOR U3415 ( .A(n835), .B(n836), .Z(n838) );
  XOR U3416 ( .A(x[1153]), .B(y[1153]), .Z(n4365) );
  XOR U3417 ( .A(x[1149]), .B(y[1149]), .Z(n4362) );
  XNOR U3418 ( .A(x[1843]), .B(y[1843]), .Z(n4363) );
  XNOR U3419 ( .A(n4362), .B(n4363), .Z(n4364) );
  XOR U3420 ( .A(n4365), .B(n4364), .Z(n3140) );
  XOR U3421 ( .A(x[1157]), .B(y[1157]), .Z(n4353) );
  XOR U3422 ( .A(x[1155]), .B(y[1155]), .Z(n4350) );
  XNOR U3423 ( .A(x[1523]), .B(y[1523]), .Z(n4351) );
  XNOR U3424 ( .A(n4350), .B(n4351), .Z(n4352) );
  XOR U3425 ( .A(n4353), .B(n4352), .Z(n3138) );
  XOR U3426 ( .A(x[1161]), .B(y[1161]), .Z(n4359) );
  XOR U3427 ( .A(x[1159]), .B(y[1159]), .Z(n4356) );
  XNOR U3428 ( .A(x[1841]), .B(y[1841]), .Z(n4357) );
  XNOR U3429 ( .A(n4356), .B(n4357), .Z(n4358) );
  XNOR U3430 ( .A(n4359), .B(n4358), .Z(n3137) );
  XNOR U3431 ( .A(n3138), .B(n3137), .Z(n3139) );
  XNOR U3432 ( .A(n3140), .B(n3139), .Z(n837) );
  XNOR U3433 ( .A(n838), .B(n837), .Z(n1327) );
  XOR U3434 ( .A(n1328), .B(n1327), .Z(n1330) );
  XOR U3435 ( .A(n1329), .B(n1330), .Z(n662) );
  XOR U3436 ( .A(x[1311]), .B(y[1311]), .Z(n3879) );
  XOR U3437 ( .A(x[1309]), .B(y[1309]), .Z(n3877) );
  XOR U3438 ( .A(x[1587]), .B(y[1587]), .Z(n3876) );
  XOR U3439 ( .A(n3877), .B(n3876), .Z(n3878) );
  XOR U3440 ( .A(n3879), .B(n3878), .Z(n570) );
  XOR U3441 ( .A(x[59]), .B(y[59]), .Z(n209) );
  XOR U3442 ( .A(x[53]), .B(y[53]), .Z(n206) );
  XNOR U3443 ( .A(x[55]), .B(y[55]), .Z(n207) );
  XNOR U3444 ( .A(n206), .B(n207), .Z(n208) );
  XOR U3445 ( .A(n209), .B(n208), .Z(n568) );
  XOR U3446 ( .A(x[1315]), .B(y[1315]), .Z(n3867) );
  XOR U3447 ( .A(x[1313]), .B(y[1313]), .Z(n3865) );
  XOR U3448 ( .A(x[1809]), .B(y[1809]), .Z(n3864) );
  XOR U3449 ( .A(n3865), .B(n3864), .Z(n3866) );
  XNOR U3450 ( .A(n3867), .B(n3866), .Z(n567) );
  XNOR U3451 ( .A(n568), .B(n567), .Z(n569) );
  XNOR U3452 ( .A(n570), .B(n569), .Z(n781) );
  XOR U3453 ( .A(x[1429]), .B(y[1429]), .Z(n4323) );
  XOR U3454 ( .A(x[1425]), .B(y[1425]), .Z(n4320) );
  XNOR U3455 ( .A(x[1427]), .B(y[1427]), .Z(n4321) );
  XNOR U3456 ( .A(n4320), .B(n4321), .Z(n4322) );
  XOR U3457 ( .A(n4323), .B(n4322), .Z(n3494) );
  XOR U3458 ( .A(x[215]), .B(y[215]), .Z(n3560) );
  XOR U3459 ( .A(x[209]), .B(y[209]), .Z(n3557) );
  XNOR U3460 ( .A(x[213]), .B(y[213]), .Z(n3558) );
  XNOR U3461 ( .A(n3557), .B(n3558), .Z(n3559) );
  XOR U3462 ( .A(n3560), .B(n3559), .Z(n3492) );
  XOR U3463 ( .A(x[1435]), .B(y[1435]), .Z(n1312) );
  XOR U3464 ( .A(x[1431]), .B(y[1431]), .Z(n1309) );
  XNOR U3465 ( .A(x[1433]), .B(y[1433]), .Z(n1310) );
  XNOR U3466 ( .A(n1309), .B(n1310), .Z(n1311) );
  XNOR U3467 ( .A(n1312), .B(n1311), .Z(n3491) );
  XNOR U3468 ( .A(n3492), .B(n3491), .Z(n3493) );
  XOR U3469 ( .A(n3494), .B(n3493), .Z(n782) );
  XNOR U3470 ( .A(n781), .B(n782), .Z(n783) );
  XOR U3471 ( .A(x[1417]), .B(y[1417]), .Z(n4329) );
  XOR U3472 ( .A(x[1413]), .B(y[1413]), .Z(n4326) );
  XNOR U3473 ( .A(x[1415]), .B(y[1415]), .Z(n4327) );
  XNOR U3474 ( .A(n4326), .B(n4327), .Z(n4328) );
  XOR U3475 ( .A(n4329), .B(n4328), .Z(n3578) );
  XOR U3476 ( .A(x[197]), .B(y[197]), .Z(n3488) );
  XOR U3477 ( .A(x[193]), .B(y[193]), .Z(n3485) );
  XNOR U3478 ( .A(x[855]), .B(y[855]), .Z(n3486) );
  XNOR U3479 ( .A(n3485), .B(n3486), .Z(n3487) );
  XOR U3480 ( .A(n3488), .B(n3487), .Z(n3576) );
  XOR U3481 ( .A(x[1423]), .B(y[1423]), .Z(n4317) );
  XOR U3482 ( .A(x[1419]), .B(y[1419]), .Z(n4314) );
  XNOR U3483 ( .A(x[1421]), .B(y[1421]), .Z(n4315) );
  XNOR U3484 ( .A(n4314), .B(n4315), .Z(n4316) );
  XNOR U3485 ( .A(n4317), .B(n4316), .Z(n3575) );
  XNOR U3486 ( .A(n3576), .B(n3575), .Z(n3577) );
  XOR U3487 ( .A(n3578), .B(n3577), .Z(n784) );
  XNOR U3488 ( .A(n783), .B(n784), .Z(n5871) );
  XOR U3489 ( .A(x[1335]), .B(y[1335]), .Z(n1269) );
  XOR U3490 ( .A(x[1333]), .B(y[1333]), .Z(n1267) );
  XNOR U3491 ( .A(x[1599]), .B(y[1599]), .Z(n1268) );
  XOR U3492 ( .A(n1267), .B(n1268), .Z(n1270) );
  XNOR U3493 ( .A(n1269), .B(n1270), .Z(n212) );
  XOR U3494 ( .A(x[1331]), .B(y[1331]), .Z(n1275) );
  XOR U3495 ( .A(x[1329]), .B(y[1329]), .Z(n1273) );
  XNOR U3496 ( .A(x[1805]), .B(y[1805]), .Z(n1274) );
  XOR U3497 ( .A(n1273), .B(n1274), .Z(n1276) );
  XOR U3498 ( .A(n1275), .B(n1276), .Z(n213) );
  XNOR U3499 ( .A(n212), .B(n213), .Z(n215) );
  XOR U3500 ( .A(x[1327]), .B(y[1327]), .Z(n3836) );
  XOR U3501 ( .A(x[1325]), .B(y[1325]), .Z(n3834) );
  XNOR U3502 ( .A(x[1595]), .B(y[1595]), .Z(n3835) );
  XOR U3503 ( .A(n3834), .B(n3835), .Z(n3837) );
  XNOR U3504 ( .A(n3836), .B(n3837), .Z(n214) );
  XOR U3505 ( .A(n215), .B(n214), .Z(n736) );
  XOR U3506 ( .A(x[1323]), .B(y[1323]), .Z(n3843) );
  XOR U3507 ( .A(x[1321]), .B(y[1321]), .Z(n3841) );
  XOR U3508 ( .A(x[1807]), .B(y[1807]), .Z(n3840) );
  XOR U3509 ( .A(n3841), .B(n3840), .Z(n3842) );
  XOR U3510 ( .A(n3843), .B(n3842), .Z(n3011) );
  XOR U3511 ( .A(x[71]), .B(y[71]), .Z(n3007) );
  XOR U3512 ( .A(x[69]), .B(y[69]), .Z(n3005) );
  XNOR U3513 ( .A(x[733]), .B(y[733]), .Z(n3006) );
  XOR U3514 ( .A(n3005), .B(n3006), .Z(n3008) );
  XOR U3515 ( .A(n3007), .B(n3008), .Z(n3012) );
  XNOR U3516 ( .A(n3011), .B(n3012), .Z(n3014) );
  XOR U3517 ( .A(x[1319]), .B(y[1319]), .Z(n3873) );
  XOR U3518 ( .A(x[1317]), .B(y[1317]), .Z(n3871) );
  XOR U3519 ( .A(x[1591]), .B(y[1591]), .Z(n3870) );
  XOR U3520 ( .A(n3871), .B(n3870), .Z(n3872) );
  XOR U3521 ( .A(n3873), .B(n3872), .Z(n3013) );
  XOR U3522 ( .A(n3014), .B(n3013), .Z(n734) );
  XOR U3523 ( .A(x[1357]), .B(y[1357]), .Z(n4299) );
  XOR U3524 ( .A(x[1353]), .B(y[1353]), .Z(n4296) );
  XNOR U3525 ( .A(x[1355]), .B(y[1355]), .Z(n4297) );
  XNOR U3526 ( .A(n4296), .B(n4297), .Z(n4298) );
  XOR U3527 ( .A(n4299), .B(n4298), .Z(n3092) );
  XOR U3528 ( .A(x[127]), .B(y[127]), .Z(n438) );
  XOR U3529 ( .A(x[125]), .B(y[125]), .Z(n435) );
  XNOR U3530 ( .A(x[795]), .B(y[795]), .Z(n436) );
  XNOR U3531 ( .A(n435), .B(n436), .Z(n437) );
  XOR U3532 ( .A(n438), .B(n437), .Z(n3090) );
  XOR U3533 ( .A(x[1363]), .B(y[1363]), .Z(n4287) );
  XOR U3534 ( .A(x[1359]), .B(y[1359]), .Z(n4284) );
  XNOR U3535 ( .A(x[1361]), .B(y[1361]), .Z(n4285) );
  XNOR U3536 ( .A(n4284), .B(n4285), .Z(n4286) );
  XNOR U3537 ( .A(n4287), .B(n4286), .Z(n3089) );
  XNOR U3538 ( .A(n3090), .B(n3089), .Z(n3091) );
  XNOR U3539 ( .A(n3092), .B(n3091), .Z(n733) );
  XNOR U3540 ( .A(n734), .B(n733), .Z(n735) );
  XNOR U3541 ( .A(n736), .B(n735), .Z(n5868) );
  XOR U3542 ( .A(x[1339]), .B(y[1339]), .Z(n1186) );
  XOR U3543 ( .A(x[1337]), .B(y[1337]), .Z(n1184) );
  XOR U3544 ( .A(x[1803]), .B(y[1803]), .Z(n1183) );
  XOR U3545 ( .A(n1184), .B(n1183), .Z(n1185) );
  XOR U3546 ( .A(n1186), .B(n1185), .Z(n265) );
  XOR U3547 ( .A(x[1345]), .B(y[1345]), .Z(n1174) );
  XOR U3548 ( .A(x[1341]), .B(y[1341]), .Z(n1172) );
  XOR U3549 ( .A(x[1343]), .B(y[1343]), .Z(n1171) );
  XOR U3550 ( .A(n1172), .B(n1171), .Z(n1173) );
  XOR U3551 ( .A(n1174), .B(n1173), .Z(n263) );
  XOR U3552 ( .A(x[1351]), .B(y[1351]), .Z(n1180) );
  XOR U3553 ( .A(x[1347]), .B(y[1347]), .Z(n1178) );
  XOR U3554 ( .A(x[1349]), .B(y[1349]), .Z(n1177) );
  XOR U3555 ( .A(n1178), .B(n1177), .Z(n1179) );
  XNOR U3556 ( .A(n1180), .B(n1179), .Z(n262) );
  XNOR U3557 ( .A(n263), .B(n262), .Z(n264) );
  XNOR U3558 ( .A(n265), .B(n264), .Z(n5869) );
  XOR U3559 ( .A(n5868), .B(n5869), .Z(n5870) );
  XOR U3560 ( .A(n5871), .B(n5870), .Z(n661) );
  XOR U3561 ( .A(n662), .B(n661), .Z(n664) );
  XOR U3562 ( .A(n663), .B(n664), .Z(n4596) );
  XOR U3563 ( .A(n4597), .B(n4596), .Z(n4598) );
  XOR U3564 ( .A(n4599), .B(n4598), .Z(n3903) );
  XOR U3565 ( .A(x[1775]), .B(y[1775]), .Z(n3074) );
  XOR U3566 ( .A(x[1635]), .B(y[1635]), .Z(n3071) );
  XNOR U3567 ( .A(x[1777]), .B(y[1777]), .Z(n3072) );
  XNOR U3568 ( .A(n3071), .B(n3072), .Z(n3073) );
  XOR U3569 ( .A(n3074), .B(n3073), .Z(n4797) );
  XOR U3570 ( .A(x[411]), .B(y[411]), .Z(n4617) );
  XOR U3571 ( .A(x[407]), .B(y[407]), .Z(n4614) );
  XNOR U3572 ( .A(x[1009]), .B(y[1009]), .Z(n4615) );
  XNOR U3573 ( .A(n4614), .B(n4615), .Z(n4616) );
  XOR U3574 ( .A(n4617), .B(n4616), .Z(n4795) );
  XOR U3575 ( .A(x[1769]), .B(y[1769]), .Z(n3062) );
  XOR U3576 ( .A(x[1637]), .B(y[1637]), .Z(n3059) );
  XNOR U3577 ( .A(x[1773]), .B(y[1773]), .Z(n3060) );
  XNOR U3578 ( .A(n3059), .B(n3060), .Z(n3061) );
  XNOR U3579 ( .A(n3062), .B(n3061), .Z(n4794) );
  XNOR U3580 ( .A(n4795), .B(n4794), .Z(n4796) );
  XNOR U3581 ( .A(n4797), .B(n4796), .Z(n1381) );
  XOR U3582 ( .A(x[1023]), .B(y[1023]), .Z(n4533) );
  XOR U3583 ( .A(x[1019]), .B(y[1019]), .Z(n4530) );
  XNOR U3584 ( .A(x[1475]), .B(y[1475]), .Z(n4531) );
  XNOR U3585 ( .A(n4530), .B(n4531), .Z(n4532) );
  XOR U3586 ( .A(n4533), .B(n4532), .Z(n1096) );
  XOR U3587 ( .A(x[1029]), .B(y[1029]), .Z(n1246) );
  XOR U3588 ( .A(x[1025]), .B(y[1025]), .Z(n1243) );
  XNOR U3589 ( .A(x[1865]), .B(y[1865]), .Z(n1244) );
  XNOR U3590 ( .A(n1243), .B(n1244), .Z(n1245) );
  XOR U3591 ( .A(n1246), .B(n1245), .Z(n1094) );
  XOR U3592 ( .A(x[1037]), .B(y[1037]), .Z(n2756) );
  XOR U3593 ( .A(x[1033]), .B(y[1033]), .Z(n2753) );
  XNOR U3594 ( .A(x[1479]), .B(y[1479]), .Z(n2754) );
  XNOR U3595 ( .A(n2753), .B(n2754), .Z(n2755) );
  XNOR U3596 ( .A(n2756), .B(n2755), .Z(n1093) );
  XNOR U3597 ( .A(n1094), .B(n1093), .Z(n1095) );
  XOR U3598 ( .A(n1096), .B(n1095), .Z(n1382) );
  XNOR U3599 ( .A(n1381), .B(n1382), .Z(n1384) );
  XOR U3600 ( .A(x[1043]), .B(y[1043]), .Z(n4581) );
  XOR U3601 ( .A(x[1039]), .B(y[1039]), .Z(n4578) );
  XNOR U3602 ( .A(x[1863]), .B(y[1863]), .Z(n4579) );
  XNOR U3603 ( .A(n4578), .B(n4579), .Z(n4580) );
  XOR U3604 ( .A(n4581), .B(n4580), .Z(n1294) );
  XOR U3605 ( .A(x[1049]), .B(y[1049]), .Z(n4569) );
  XOR U3606 ( .A(x[1045]), .B(y[1045]), .Z(n4566) );
  XNOR U3607 ( .A(x[1483]), .B(y[1483]), .Z(n4567) );
  XNOR U3608 ( .A(n4566), .B(n4567), .Z(n4568) );
  XOR U3609 ( .A(n4569), .B(n4568), .Z(n1292) );
  XOR U3610 ( .A(x[1055]), .B(y[1055]), .Z(n4575) );
  XOR U3611 ( .A(x[1051]), .B(y[1051]), .Z(n4572) );
  XNOR U3612 ( .A(x[1861]), .B(y[1861]), .Z(n4573) );
  XNOR U3613 ( .A(n4572), .B(n4573), .Z(n4574) );
  XNOR U3614 ( .A(n4575), .B(n4574), .Z(n1291) );
  XNOR U3615 ( .A(n1292), .B(n1291), .Z(n1293) );
  XNOR U3616 ( .A(n1294), .B(n1293), .Z(n1383) );
  XNOR U3617 ( .A(n1384), .B(n1383), .Z(n5673) );
  XOR U3618 ( .A(x[1063]), .B(y[1063]), .Z(n4113) );
  XOR U3619 ( .A(x[1059]), .B(y[1059]), .Z(n4110) );
  XNOR U3620 ( .A(x[1487]), .B(y[1487]), .Z(n4111) );
  XNOR U3621 ( .A(n4110), .B(n4111), .Z(n4112) );
  XOR U3622 ( .A(n4113), .B(n4112), .Z(n1414) );
  XOR U3623 ( .A(x[168]), .B(y[168]), .Z(n1790) );
  XOR U3624 ( .A(x[170]), .B(y[170]), .Z(n1787) );
  XNOR U3625 ( .A(x[777]), .B(y[777]), .Z(n1788) );
  XNOR U3626 ( .A(n1787), .B(n1788), .Z(n1789) );
  XOR U3627 ( .A(n1790), .B(n1789), .Z(n1412) );
  XOR U3628 ( .A(x[1069]), .B(y[1069]), .Z(n4101) );
  XOR U3629 ( .A(x[1065]), .B(y[1065]), .Z(n4098) );
  XNOR U3630 ( .A(x[1859]), .B(y[1859]), .Z(n4099) );
  XNOR U3631 ( .A(n4098), .B(n4099), .Z(n4100) );
  XNOR U3632 ( .A(n4101), .B(n4100), .Z(n1411) );
  XNOR U3633 ( .A(n1412), .B(n1411), .Z(n1413) );
  XNOR U3634 ( .A(n1414), .B(n1413), .Z(n991) );
  XOR U3635 ( .A(x[1787]), .B(y[1787]), .Z(n3759) );
  XOR U3636 ( .A(x[1629]), .B(y[1629]), .Z(n3756) );
  XNOR U3637 ( .A(x[1789]), .B(y[1789]), .Z(n3757) );
  XNOR U3638 ( .A(n3756), .B(n3757), .Z(n3758) );
  XOR U3639 ( .A(n3759), .B(n3758), .Z(n3182) );
  XOR U3640 ( .A(x[1783]), .B(y[1783]), .Z(n3747) );
  XOR U3641 ( .A(x[1631]), .B(y[1631]), .Z(n3744) );
  XNOR U3642 ( .A(x[1785]), .B(y[1785]), .Z(n3745) );
  XNOR U3643 ( .A(n3744), .B(n3745), .Z(n3746) );
  XOR U3644 ( .A(n3747), .B(n3746), .Z(n3180) );
  XOR U3645 ( .A(x[1779]), .B(y[1779]), .Z(n3753) );
  XOR U3646 ( .A(x[1633]), .B(y[1633]), .Z(n3750) );
  XNOR U3647 ( .A(x[1781]), .B(y[1781]), .Z(n3751) );
  XNOR U3648 ( .A(n3750), .B(n3751), .Z(n3752) );
  XNOR U3649 ( .A(n3753), .B(n3752), .Z(n3179) );
  XNOR U3650 ( .A(n3180), .B(n3179), .Z(n3181) );
  XOR U3651 ( .A(n3182), .B(n3181), .Z(n992) );
  XNOR U3652 ( .A(n991), .B(n992), .Z(n994) );
  XOR U3653 ( .A(x[1073]), .B(y[1073]), .Z(n4107) );
  XOR U3654 ( .A(x[1071]), .B(y[1071]), .Z(n4104) );
  XNOR U3655 ( .A(x[1491]), .B(y[1491]), .Z(n4105) );
  XNOR U3656 ( .A(n4104), .B(n4105), .Z(n4106) );
  XOR U3657 ( .A(n4107), .B(n4106), .Z(n988) );
  XOR U3658 ( .A(x[160]), .B(y[160]), .Z(n844) );
  XOR U3659 ( .A(x[162]), .B(y[162]), .Z(n841) );
  XNOR U3660 ( .A(x[785]), .B(y[785]), .Z(n842) );
  XNOR U3661 ( .A(n841), .B(n842), .Z(n843) );
  XOR U3662 ( .A(n844), .B(n843), .Z(n986) );
  XOR U3663 ( .A(x[1081]), .B(y[1081]), .Z(n4227) );
  XOR U3664 ( .A(x[1077]), .B(y[1077]), .Z(n4224) );
  XNOR U3665 ( .A(x[1857]), .B(y[1857]), .Z(n4225) );
  XNOR U3666 ( .A(n4224), .B(n4225), .Z(n4226) );
  XNOR U3667 ( .A(n4227), .B(n4226), .Z(n985) );
  XNOR U3668 ( .A(n986), .B(n985), .Z(n987) );
  XNOR U3669 ( .A(n988), .B(n987), .Z(n993) );
  XNOR U3670 ( .A(n994), .B(n993), .Z(n5671) );
  XOR U3671 ( .A(x[1801]), .B(y[1801]), .Z(n1042) );
  XOR U3672 ( .A(x[1623]), .B(y[1623]), .Z(n1039) );
  XNOR U3673 ( .A(x[1799]), .B(y[1799]), .Z(n1040) );
  XNOR U3674 ( .A(n1039), .B(n1040), .Z(n1041) );
  XOR U3675 ( .A(n1042), .B(n1041), .Z(n2792) );
  XOR U3676 ( .A(x[1795]), .B(y[1795]), .Z(n143) );
  XOR U3677 ( .A(x[1625]), .B(y[1625]), .Z(n140) );
  XNOR U3678 ( .A(x[1797]), .B(y[1797]), .Z(n141) );
  XNOR U3679 ( .A(n140), .B(n141), .Z(n142) );
  XOR U3680 ( .A(n143), .B(n142), .Z(n2790) );
  XOR U3681 ( .A(x[1791]), .B(y[1791]), .Z(n137) );
  XOR U3682 ( .A(x[1627]), .B(y[1627]), .Z(n134) );
  XNOR U3683 ( .A(x[1793]), .B(y[1793]), .Z(n135) );
  XNOR U3684 ( .A(n134), .B(n135), .Z(n136) );
  XNOR U3685 ( .A(n137), .B(n136), .Z(n2789) );
  XNOR U3686 ( .A(n2790), .B(n2789), .Z(n2791) );
  XNOR U3687 ( .A(n2792), .B(n2791), .Z(n955) );
  XOR U3688 ( .A(x[1085]), .B(y[1085]), .Z(n4221) );
  XOR U3689 ( .A(x[1083]), .B(y[1083]), .Z(n4218) );
  XNOR U3690 ( .A(x[1495]), .B(y[1495]), .Z(n4219) );
  XNOR U3691 ( .A(n4218), .B(n4219), .Z(n4220) );
  XOR U3692 ( .A(n4221), .B(n4220), .Z(n1342) );
  XOR U3693 ( .A(x[1089]), .B(y[1089]), .Z(n4491) );
  XOR U3694 ( .A(x[1087]), .B(y[1087]), .Z(n4488) );
  XNOR U3695 ( .A(x[1855]), .B(y[1855]), .Z(n4489) );
  XNOR U3696 ( .A(n4488), .B(n4489), .Z(n4490) );
  XOR U3697 ( .A(n4491), .B(n4490), .Z(n1340) );
  XOR U3698 ( .A(x[1095]), .B(y[1095]), .Z(n4485) );
  XOR U3699 ( .A(x[1091]), .B(y[1091]), .Z(n4482) );
  XNOR U3700 ( .A(x[1499]), .B(y[1499]), .Z(n4483) );
  XNOR U3701 ( .A(n4482), .B(n4483), .Z(n4484) );
  XNOR U3702 ( .A(n4485), .B(n4484), .Z(n1339) );
  XNOR U3703 ( .A(n1340), .B(n1339), .Z(n1341) );
  XOR U3704 ( .A(n1342), .B(n1341), .Z(n956) );
  XNOR U3705 ( .A(n955), .B(n956), .Z(n958) );
  XOR U3706 ( .A(x[1101]), .B(y[1101]), .Z(n4563) );
  XOR U3707 ( .A(x[1099]), .B(y[1099]), .Z(n4560) );
  XNOR U3708 ( .A(x[1853]), .B(y[1853]), .Z(n4561) );
  XNOR U3709 ( .A(n4560), .B(n4561), .Z(n4562) );
  XOR U3710 ( .A(n4563), .B(n4562), .Z(n1540) );
  XOR U3711 ( .A(x[1105]), .B(y[1105]), .Z(n4551) );
  XOR U3712 ( .A(x[1103]), .B(y[1103]), .Z(n4548) );
  XNOR U3713 ( .A(x[1503]), .B(y[1503]), .Z(n4549) );
  XNOR U3714 ( .A(n4548), .B(n4549), .Z(n4550) );
  XOR U3715 ( .A(n4551), .B(n4550), .Z(n1538) );
  XOR U3716 ( .A(x[1109]), .B(y[1109]), .Z(n4557) );
  XOR U3717 ( .A(x[1107]), .B(y[1107]), .Z(n4554) );
  XNOR U3718 ( .A(x[1851]), .B(y[1851]), .Z(n4555) );
  XNOR U3719 ( .A(n4554), .B(n4555), .Z(n4556) );
  XNOR U3720 ( .A(n4557), .B(n4556), .Z(n1537) );
  XNOR U3721 ( .A(n1538), .B(n1537), .Z(n1539) );
  XNOR U3722 ( .A(n1540), .B(n1539), .Z(n957) );
  XNOR U3723 ( .A(n958), .B(n957), .Z(n5670) );
  XOR U3724 ( .A(n5671), .B(n5670), .Z(n5672) );
  XNOR U3725 ( .A(n5673), .B(n5672), .Z(n670) );
  XOR U3726 ( .A(x[713]), .B(y[713]), .Z(n2696) );
  XOR U3727 ( .A(x[709]), .B(y[709]), .Z(n2693) );
  XNOR U3728 ( .A(x[1133]), .B(y[1133]), .Z(n2694) );
  XNOR U3729 ( .A(n2693), .B(n2694), .Z(n2695) );
  XOR U3730 ( .A(n2696), .B(n2695), .Z(n4755) );
  XOR U3731 ( .A(x[354]), .B(y[354]), .Z(n2222) );
  XOR U3732 ( .A(x[356]), .B(y[356]), .Z(n2219) );
  XNOR U3733 ( .A(x[1895]), .B(y[1895]), .Z(n2220) );
  XNOR U3734 ( .A(n2219), .B(n2220), .Z(n2221) );
  XOR U3735 ( .A(n2222), .B(n2221), .Z(n4753) );
  XOR U3736 ( .A(x[729]), .B(y[729]), .Z(n2576) );
  XOR U3737 ( .A(x[715]), .B(y[715]), .Z(n2573) );
  XNOR U3738 ( .A(x[719]), .B(y[719]), .Z(n2574) );
  XNOR U3739 ( .A(n2573), .B(n2574), .Z(n2575) );
  XNOR U3740 ( .A(n2576), .B(n2575), .Z(n4752) );
  XNOR U3741 ( .A(n4753), .B(n4752), .Z(n4754) );
  XNOR U3742 ( .A(n4755), .B(n4754), .Z(n1465) );
  XOR U3743 ( .A(x[743]), .B(y[743]), .Z(n2570) );
  XOR U3744 ( .A(x[735]), .B(y[735]), .Z(n2567) );
  XNOR U3745 ( .A(x[739]), .B(y[739]), .Z(n2568) );
  XNOR U3746 ( .A(n2567), .B(n2568), .Z(n2569) );
  XOR U3747 ( .A(n2570), .B(n2569), .Z(n5583) );
  XOR U3748 ( .A(x[344]), .B(y[344]), .Z(n2192) );
  XOR U3749 ( .A(x[346]), .B(y[346]), .Z(n2189) );
  XNOR U3750 ( .A(x[1893]), .B(y[1893]), .Z(n2190) );
  XNOR U3751 ( .A(n2189), .B(n2190), .Z(n2191) );
  XOR U3752 ( .A(n2192), .B(n2191), .Z(n5581) );
  XOR U3753 ( .A(x[753]), .B(y[753]), .Z(n2480) );
  XOR U3754 ( .A(x[749]), .B(y[749]), .Z(n2477) );
  XNOR U3755 ( .A(x[1147]), .B(y[1147]), .Z(n2478) );
  XNOR U3756 ( .A(n2477), .B(n2478), .Z(n2479) );
  XNOR U3757 ( .A(n2480), .B(n2479), .Z(n5580) );
  XNOR U3758 ( .A(n5581), .B(n5580), .Z(n5582) );
  XOR U3759 ( .A(n5583), .B(n5582), .Z(n1466) );
  XNOR U3760 ( .A(n1465), .B(n1466), .Z(n1468) );
  XOR U3761 ( .A(x[763]), .B(y[763]), .Z(n2468) );
  XOR U3762 ( .A(x[755]), .B(y[755]), .Z(n2465) );
  XNOR U3763 ( .A(x[1151]), .B(y[1151]), .Z(n2466) );
  XNOR U3764 ( .A(n2465), .B(n2466), .Z(n2467) );
  XOR U3765 ( .A(n2468), .B(n2467), .Z(n5667) );
  XOR U3766 ( .A(x[779]), .B(y[779]), .Z(n2474) );
  XOR U3767 ( .A(x[771]), .B(y[771]), .Z(n2471) );
  XNOR U3768 ( .A(x[775]), .B(y[775]), .Z(n2472) );
  XNOR U3769 ( .A(n2471), .B(n2472), .Z(n2473) );
  XOR U3770 ( .A(n2474), .B(n2473), .Z(n5665) );
  XOR U3771 ( .A(x[791]), .B(y[791]), .Z(n3668) );
  XOR U3772 ( .A(x[783]), .B(y[783]), .Z(n3665) );
  XNOR U3773 ( .A(x[789]), .B(y[789]), .Z(n3666) );
  XNOR U3774 ( .A(n3665), .B(n3666), .Z(n3667) );
  XNOR U3775 ( .A(n3668), .B(n3667), .Z(n5664) );
  XNOR U3776 ( .A(n5665), .B(n5664), .Z(n5666) );
  XNOR U3777 ( .A(n5667), .B(n5666), .Z(n1467) );
  XNOR U3778 ( .A(n1468), .B(n1467), .Z(n3933) );
  XOR U3779 ( .A(x[809]), .B(y[809]), .Z(n3656) );
  XOR U3780 ( .A(x[797]), .B(y[797]), .Z(n3653) );
  XNOR U3781 ( .A(x[1165]), .B(y[1165]), .Z(n3654) );
  XNOR U3782 ( .A(n3653), .B(n3654), .Z(n3655) );
  XOR U3783 ( .A(n3656), .B(n3655), .Z(n1054) );
  XOR U3784 ( .A(x[815]), .B(y[815]), .Z(n3662) );
  XOR U3785 ( .A(x[811]), .B(y[811]), .Z(n3659) );
  XNOR U3786 ( .A(x[1169]), .B(y[1169]), .Z(n3660) );
  XNOR U3787 ( .A(n3659), .B(n3660), .Z(n3661) );
  XOR U3788 ( .A(n3662), .B(n3661), .Z(n1052) );
  XOR U3789 ( .A(x[825]), .B(y[825]), .Z(n2816) );
  XOR U3790 ( .A(x[817]), .B(y[817]), .Z(n2813) );
  XNOR U3791 ( .A(x[823]), .B(y[823]), .Z(n2814) );
  XNOR U3792 ( .A(n2813), .B(n2814), .Z(n2815) );
  XNOR U3793 ( .A(n2816), .B(n2815), .Z(n1051) );
  XNOR U3794 ( .A(n1052), .B(n1051), .Z(n1053) );
  XNOR U3795 ( .A(n1054), .B(n1053), .Z(n1417) );
  XOR U3796 ( .A(x[837]), .B(y[837]), .Z(n2810) );
  XOR U3797 ( .A(x[831]), .B(y[831]), .Z(n2807) );
  XNOR U3798 ( .A(x[835]), .B(y[835]), .Z(n2808) );
  XNOR U3799 ( .A(n2807), .B(n2808), .Z(n2809) );
  XOR U3800 ( .A(n2810), .B(n2809), .Z(n1240) );
  XOR U3801 ( .A(x[308]), .B(y[308]), .Z(n2456) );
  XOR U3802 ( .A(x[310]), .B(y[310]), .Z(n2453) );
  XNOR U3803 ( .A(x[683]), .B(y[683]), .Z(n2454) );
  XNOR U3804 ( .A(n2453), .B(n2454), .Z(n2455) );
  XOR U3805 ( .A(n2456), .B(n2455), .Z(n1238) );
  XOR U3806 ( .A(x[843]), .B(y[843]), .Z(n3200) );
  XOR U3807 ( .A(x[839]), .B(y[839]), .Z(n3197) );
  XNOR U3808 ( .A(x[1183]), .B(y[1183]), .Z(n3198) );
  XNOR U3809 ( .A(n3197), .B(n3198), .Z(n3199) );
  XNOR U3810 ( .A(n3200), .B(n3199), .Z(n1237) );
  XNOR U3811 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U3812 ( .A(n1240), .B(n1239), .Z(n1418) );
  XNOR U3813 ( .A(n1417), .B(n1418), .Z(n1420) );
  XOR U3814 ( .A(x[849]), .B(y[849]), .Z(n3194) );
  XOR U3815 ( .A(x[845]), .B(y[845]), .Z(n3191) );
  XNOR U3816 ( .A(x[1187]), .B(y[1187]), .Z(n3192) );
  XNOR U3817 ( .A(n3191), .B(n3192), .Z(n3193) );
  XOR U3818 ( .A(n3194), .B(n3193), .Z(n1318) );
  XOR U3819 ( .A(x[294]), .B(y[294]), .Z(n2426) );
  XOR U3820 ( .A(x[296]), .B(y[296]), .Z(n2423) );
  XNOR U3821 ( .A(x[691]), .B(y[691]), .Z(n2424) );
  XNOR U3822 ( .A(n2423), .B(n2424), .Z(n2425) );
  XOR U3823 ( .A(n2426), .B(n2425), .Z(n1316) );
  XOR U3824 ( .A(x[859]), .B(y[859]), .Z(n3116) );
  XOR U3825 ( .A(x[853]), .B(y[853]), .Z(n3113) );
  XNOR U3826 ( .A(x[857]), .B(y[857]), .Z(n3114) );
  XNOR U3827 ( .A(n3113), .B(n3114), .Z(n3115) );
  XNOR U3828 ( .A(n3116), .B(n3115), .Z(n1315) );
  XNOR U3829 ( .A(n1316), .B(n1315), .Z(n1317) );
  XNOR U3830 ( .A(n1318), .B(n1317), .Z(n1419) );
  XNOR U3831 ( .A(n1420), .B(n1419), .Z(n3931) );
  XOR U3832 ( .A(x[869]), .B(y[869]), .Z(n3104) );
  XOR U3833 ( .A(x[863]), .B(y[863]), .Z(n3101) );
  XNOR U3834 ( .A(x[865]), .B(y[865]), .Z(n3102) );
  XNOR U3835 ( .A(n3101), .B(n3102), .Z(n3103) );
  XOR U3836 ( .A(n3104), .B(n3103), .Z(n5961) );
  XOR U3837 ( .A(x[875]), .B(y[875]), .Z(n3110) );
  XOR U3838 ( .A(x[871]), .B(y[871]), .Z(n3107) );
  XNOR U3839 ( .A(x[1201]), .B(y[1201]), .Z(n3108) );
  XNOR U3840 ( .A(n3107), .B(n3108), .Z(n3109) );
  XOR U3841 ( .A(n3110), .B(n3109), .Z(n5959) );
  XOR U3842 ( .A(x[883]), .B(y[883]), .Z(n2540) );
  XOR U3843 ( .A(x[879]), .B(y[879]), .Z(n2537) );
  XNOR U3844 ( .A(x[1205]), .B(y[1205]), .Z(n2538) );
  XNOR U3845 ( .A(n2537), .B(n2538), .Z(n2539) );
  XNOR U3846 ( .A(n2540), .B(n2539), .Z(n5958) );
  XNOR U3847 ( .A(n5959), .B(n5958), .Z(n5960) );
  XNOR U3848 ( .A(n5961), .B(n5960), .Z(n1369) );
  XOR U3849 ( .A(x[1743]), .B(y[1743]), .Z(n618) );
  XOR U3850 ( .A(x[1667]), .B(y[1667]), .Z(n615) );
  XNOR U3851 ( .A(x[1745]), .B(y[1745]), .Z(n616) );
  XNOR U3852 ( .A(n615), .B(n616), .Z(n617) );
  XOR U3853 ( .A(n618), .B(n617), .Z(n5751) );
  XOR U3854 ( .A(x[509]), .B(y[509]), .Z(n2618) );
  XOR U3855 ( .A(x[505]), .B(y[505]), .Z(n2615) );
  XNOR U3856 ( .A(x[1057]), .B(y[1057]), .Z(n2616) );
  XNOR U3857 ( .A(n2615), .B(n2616), .Z(n2617) );
  XOR U3858 ( .A(n2618), .B(n2617), .Z(n5749) );
  XOR U3859 ( .A(x[1741]), .B(y[1741]), .Z(n606) );
  XOR U3860 ( .A(x[1653]), .B(y[1653]), .Z(n603) );
  XNOR U3861 ( .A(x[1659]), .B(y[1659]), .Z(n604) );
  XNOR U3862 ( .A(n603), .B(n604), .Z(n605) );
  XNOR U3863 ( .A(n606), .B(n605), .Z(n5748) );
  XNOR U3864 ( .A(n5749), .B(n5748), .Z(n5750) );
  XOR U3865 ( .A(n5751), .B(n5750), .Z(n1370) );
  XNOR U3866 ( .A(n1369), .B(n1370), .Z(n1372) );
  XOR U3867 ( .A(x[891]), .B(y[891]), .Z(n2528) );
  XOR U3868 ( .A(x[885]), .B(y[885]), .Z(n2525) );
  XNOR U3869 ( .A(x[889]), .B(y[889]), .Z(n2526) );
  XNOR U3870 ( .A(n2525), .B(n2526), .Z(n2527) );
  XOR U3871 ( .A(n2528), .B(n2527), .Z(n1012) );
  XOR U3872 ( .A(x[903]), .B(y[903]), .Z(n2534) );
  XOR U3873 ( .A(x[893]), .B(y[893]), .Z(n2531) );
  XNOR U3874 ( .A(x[897]), .B(y[897]), .Z(n2532) );
  XNOR U3875 ( .A(n2531), .B(n2532), .Z(n2533) );
  XOR U3876 ( .A(n2534), .B(n2533), .Z(n1010) );
  XOR U3877 ( .A(x[909]), .B(y[909]), .Z(n2522) );
  XOR U3878 ( .A(x[905]), .B(y[905]), .Z(n2519) );
  XNOR U3879 ( .A(x[1219]), .B(y[1219]), .Z(n2520) );
  XNOR U3880 ( .A(n2519), .B(n2520), .Z(n2521) );
  XNOR U3881 ( .A(n2522), .B(n2521), .Z(n1009) );
  XNOR U3882 ( .A(n1010), .B(n1009), .Z(n1011) );
  XNOR U3883 ( .A(n1012), .B(n1011), .Z(n1371) );
  XNOR U3884 ( .A(n1372), .B(n1371), .Z(n3930) );
  XOR U3885 ( .A(n3931), .B(n3930), .Z(n3932) );
  XNOR U3886 ( .A(n3933), .B(n3932), .Z(n668) );
  XOR U3887 ( .A(x[913]), .B(y[913]), .Z(n2516) );
  XOR U3888 ( .A(x[911]), .B(y[911]), .Z(n2513) );
  XNOR U3889 ( .A(x[1223]), .B(y[1223]), .Z(n2514) );
  XNOR U3890 ( .A(n2513), .B(n2514), .Z(n2515) );
  XOR U3891 ( .A(n2516), .B(n2515), .Z(n1000) );
  XOR U3892 ( .A(x[262]), .B(y[262]), .Z(n2312) );
  XOR U3893 ( .A(x[264]), .B(y[264]), .Z(n2309) );
  XNOR U3894 ( .A(x[1885]), .B(y[1885]), .Z(n2310) );
  XNOR U3895 ( .A(n2309), .B(n2310), .Z(n2311) );
  XOR U3896 ( .A(n2312), .B(n2311), .Z(n998) );
  XOR U3897 ( .A(x[925]), .B(y[925]), .Z(n2762) );
  XOR U3898 ( .A(x[915]), .B(y[915]), .Z(n2759) );
  XNOR U3899 ( .A(x[919]), .B(y[919]), .Z(n2760) );
  XNOR U3900 ( .A(n2759), .B(n2760), .Z(n2761) );
  XNOR U3901 ( .A(n2762), .B(n2761), .Z(n997) );
  XNOR U3902 ( .A(n998), .B(n997), .Z(n999) );
  XNOR U3903 ( .A(n1000), .B(n999), .Z(n1375) );
  XOR U3904 ( .A(x[1749]), .B(y[1749]), .Z(n420) );
  XOR U3905 ( .A(x[1665]), .B(y[1665]), .Z(n417) );
  XNOR U3906 ( .A(x[1751]), .B(y[1751]), .Z(n418) );
  XNOR U3907 ( .A(n417), .B(n418), .Z(n419) );
  XOR U3908 ( .A(n420), .B(n419), .Z(n5937) );
  XOR U3909 ( .A(x[1647]), .B(y[1647]), .Z(n408) );
  XOR U3910 ( .A(x[1661]), .B(y[1661]), .Z(n405) );
  XNOR U3911 ( .A(x[1747]), .B(y[1747]), .Z(n406) );
  XNOR U3912 ( .A(n405), .B(n406), .Z(n407) );
  XOR U3913 ( .A(n408), .B(n407), .Z(n5935) );
  XOR U3914 ( .A(x[1651]), .B(y[1651]), .Z(n414) );
  XOR U3915 ( .A(x[1649]), .B(y[1649]), .Z(n411) );
  XNOR U3916 ( .A(x[1663]), .B(y[1663]), .Z(n412) );
  XNOR U3917 ( .A(n411), .B(n412), .Z(n413) );
  XNOR U3918 ( .A(n414), .B(n413), .Z(n5934) );
  XNOR U3919 ( .A(n5935), .B(n5934), .Z(n5936) );
  XOR U3920 ( .A(n5937), .B(n5936), .Z(n1376) );
  XNOR U3921 ( .A(n1375), .B(n1376), .Z(n1377) );
  XOR U3922 ( .A(x[933]), .B(y[933]), .Z(n2732) );
  XOR U3923 ( .A(x[929]), .B(y[929]), .Z(n2729) );
  XNOR U3924 ( .A(x[931]), .B(y[931]), .Z(n2730) );
  XNOR U3925 ( .A(n2729), .B(n2730), .Z(n2731) );
  XOR U3926 ( .A(n2732), .B(n2731), .Z(n1666) );
  XOR U3927 ( .A(x[248]), .B(y[248]), .Z(n2360) );
  XOR U3928 ( .A(x[250]), .B(y[250]), .Z(n2357) );
  XNOR U3929 ( .A(x[723]), .B(y[723]), .Z(n2358) );
  XNOR U3930 ( .A(n2357), .B(n2358), .Z(n2359) );
  XOR U3931 ( .A(n2360), .B(n2359), .Z(n1664) );
  XOR U3932 ( .A(x[937]), .B(y[937]), .Z(n2342) );
  XOR U3933 ( .A(x[935]), .B(y[935]), .Z(n2339) );
  XNOR U3934 ( .A(x[1237]), .B(y[1237]), .Z(n2340) );
  XNOR U3935 ( .A(n2339), .B(n2340), .Z(n2341) );
  XNOR U3936 ( .A(n2342), .B(n2341), .Z(n1663) );
  XNOR U3937 ( .A(n1664), .B(n1663), .Z(n1665) );
  XOR U3938 ( .A(n1666), .B(n1665), .Z(n1378) );
  XNOR U3939 ( .A(n1377), .B(n1378), .Z(n4827) );
  XOR U3940 ( .A(x[997]), .B(y[997]), .Z(n1862) );
  XOR U3941 ( .A(x[993]), .B(y[993]), .Z(n1859) );
  XNOR U3942 ( .A(x[995]), .B(y[995]), .Z(n1860) );
  XNOR U3943 ( .A(n1859), .B(n1860), .Z(n1861) );
  XOR U3944 ( .A(n1862), .B(n1861), .Z(n5973) );
  XOR U3945 ( .A(x[212]), .B(y[212]), .Z(n862) );
  XOR U3946 ( .A(x[214]), .B(y[214]), .Z(n859) );
  XNOR U3947 ( .A(x[745]), .B(y[745]), .Z(n860) );
  XNOR U3948 ( .A(n859), .B(n860), .Z(n861) );
  XOR U3949 ( .A(n862), .B(n861), .Z(n5971) );
  XOR U3950 ( .A(x[1003]), .B(y[1003]), .Z(n1582) );
  XOR U3951 ( .A(x[999]), .B(y[999]), .Z(n1579) );
  XNOR U3952 ( .A(x[1273]), .B(y[1273]), .Z(n1580) );
  XNOR U3953 ( .A(n1579), .B(n1580), .Z(n1581) );
  XNOR U3954 ( .A(n1582), .B(n1581), .Z(n5970) );
  XNOR U3955 ( .A(n5971), .B(n5970), .Z(n5972) );
  XNOR U3956 ( .A(n5973), .B(n5972), .Z(n1285) );
  XOR U3957 ( .A(x[1765]), .B(y[1765]), .Z(n3068) );
  XOR U3958 ( .A(x[1639]), .B(y[1639]), .Z(n3065) );
  XNOR U3959 ( .A(x[1767]), .B(y[1767]), .Z(n3066) );
  XNOR U3960 ( .A(n3065), .B(n3066), .Z(n3067) );
  XOR U3961 ( .A(n3068), .B(n3067), .Z(n5637) );
  XOR U3962 ( .A(x[431]), .B(y[431]), .Z(n3236) );
  XOR U3963 ( .A(x[423]), .B(y[423]), .Z(n3233) );
  XNOR U3964 ( .A(x[425]), .B(y[425]), .Z(n3234) );
  XNOR U3965 ( .A(n3233), .B(n3234), .Z(n3235) );
  XOR U3966 ( .A(n3236), .B(n3235), .Z(n5635) );
  XOR U3967 ( .A(x[1771]), .B(y[1771]), .Z(n2894) );
  XOR U3968 ( .A(x[1641]), .B(y[1641]), .Z(n2891) );
  XNOR U3969 ( .A(x[1763]), .B(y[1763]), .Z(n2892) );
  XNOR U3970 ( .A(n2891), .B(n2892), .Z(n2893) );
  XNOR U3971 ( .A(n2894), .B(n2893), .Z(n5634) );
  XNOR U3972 ( .A(n5635), .B(n5634), .Z(n5636) );
  XOR U3973 ( .A(n5637), .B(n5636), .Z(n1286) );
  XNOR U3974 ( .A(n1285), .B(n1286), .Z(n1287) );
  XOR U3975 ( .A(x[1011]), .B(y[1011]), .Z(n1702) );
  XOR U3976 ( .A(x[1005]), .B(y[1005]), .Z(n1699) );
  XNOR U3977 ( .A(x[1471]), .B(y[1471]), .Z(n1700) );
  XNOR U3978 ( .A(n1699), .B(n1700), .Z(n1701) );
  XOR U3979 ( .A(n1702), .B(n1701), .Z(n5829) );
  XOR U3980 ( .A(x[202]), .B(y[202]), .Z(n1744) );
  XOR U3981 ( .A(x[204]), .B(y[204]), .Z(n1741) );
  XNOR U3982 ( .A(x[1021]), .B(y[1021]), .Z(n1742) );
  XNOR U3983 ( .A(n1741), .B(n1742), .Z(n1743) );
  XOR U3984 ( .A(n1744), .B(n1743), .Z(n5827) );
  XOR U3985 ( .A(x[1017]), .B(y[1017]), .Z(n1546) );
  XOR U3986 ( .A(x[1015]), .B(y[1015]), .Z(n1543) );
  XNOR U3987 ( .A(x[1867]), .B(y[1867]), .Z(n1544) );
  XNOR U3988 ( .A(n1543), .B(n1544), .Z(n1545) );
  XNOR U3989 ( .A(n1546), .B(n1545), .Z(n5826) );
  XNOR U3990 ( .A(n5827), .B(n5826), .Z(n5828) );
  XOR U3991 ( .A(n5829), .B(n5828), .Z(n1288) );
  XNOR U3992 ( .A(n1287), .B(n1288), .Z(n4824) );
  XOR U3993 ( .A(x[949]), .B(y[949]), .Z(n2270) );
  XOR U3994 ( .A(x[943]), .B(y[943]), .Z(n2267) );
  XNOR U3995 ( .A(x[1241]), .B(y[1241]), .Z(n2268) );
  XNOR U3996 ( .A(n2267), .B(n2268), .Z(n2269) );
  XOR U3997 ( .A(n2270), .B(n2269), .Z(n1690) );
  XOR U3998 ( .A(x[955]), .B(y[955]), .Z(n2246) );
  XOR U3999 ( .A(x[951]), .B(y[951]), .Z(n2243) );
  XNOR U4000 ( .A(x[953]), .B(y[953]), .Z(n2244) );
  XNOR U4001 ( .A(n2243), .B(n2244), .Z(n2245) );
  XOR U4002 ( .A(n2246), .B(n2245), .Z(n1688) );
  XOR U4003 ( .A(x[965]), .B(y[965]), .Z(n1426) );
  XOR U4004 ( .A(x[957]), .B(y[957]), .Z(n1423) );
  XNOR U4005 ( .A(x[959]), .B(y[959]), .Z(n1424) );
  XNOR U4006 ( .A(n1423), .B(n1424), .Z(n1425) );
  XNOR U4007 ( .A(n1426), .B(n1425), .Z(n1687) );
  XNOR U4008 ( .A(n1688), .B(n1687), .Z(n1689) );
  XNOR U4009 ( .A(n1690), .B(n1689), .Z(n1279) );
  XOR U4010 ( .A(x[1759]), .B(y[1759]), .Z(n2888) );
  XOR U4011 ( .A(x[1643]), .B(y[1643]), .Z(n2885) );
  XNOR U4012 ( .A(x[1761]), .B(y[1761]), .Z(n2886) );
  XNOR U4013 ( .A(n2885), .B(n2886), .Z(n2887) );
  XOR U4014 ( .A(n2888), .B(n2887), .Z(n5853) );
  XOR U4015 ( .A(x[1757]), .B(y[1757]), .Z(n251) );
  XOR U4016 ( .A(x[1645]), .B(y[1645]), .Z(n248) );
  XNOR U4017 ( .A(x[1671]), .B(y[1671]), .Z(n249) );
  XNOR U4018 ( .A(n248), .B(n249), .Z(n250) );
  XOR U4019 ( .A(n251), .B(n250), .Z(n5851) );
  XOR U4020 ( .A(x[1753]), .B(y[1753]), .Z(n245) );
  XOR U4021 ( .A(x[1669]), .B(y[1669]), .Z(n242) );
  XNOR U4022 ( .A(x[1755]), .B(y[1755]), .Z(n243) );
  XNOR U4023 ( .A(n242), .B(n243), .Z(n244) );
  XNOR U4024 ( .A(n245), .B(n244), .Z(n5850) );
  XNOR U4025 ( .A(n5851), .B(n5850), .Z(n5852) );
  XOR U4026 ( .A(n5853), .B(n5852), .Z(n1280) );
  XNOR U4027 ( .A(n1279), .B(n1280), .Z(n1281) );
  XOR U4028 ( .A(x[973]), .B(y[973]), .Z(n1444) );
  XOR U4029 ( .A(x[971]), .B(y[971]), .Z(n1441) );
  XNOR U4030 ( .A(x[1255]), .B(y[1255]), .Z(n1442) );
  XNOR U4031 ( .A(n1441), .B(n1442), .Z(n1443) );
  XOR U4032 ( .A(n1444), .B(n1443), .Z(n964) );
  XOR U4033 ( .A(x[977]), .B(y[977]), .Z(n4179) );
  XOR U4034 ( .A(x[975]), .B(y[975]), .Z(n4176) );
  XNOR U4035 ( .A(x[1259]), .B(y[1259]), .Z(n4177) );
  XNOR U4036 ( .A(n4176), .B(n4177), .Z(n4178) );
  XOR U4037 ( .A(n4179), .B(n4178), .Z(n962) );
  XOR U4038 ( .A(x[989]), .B(y[989]), .Z(n1826) );
  XOR U4039 ( .A(x[979]), .B(y[979]), .Z(n1823) );
  XNOR U4040 ( .A(x[983]), .B(y[983]), .Z(n1824) );
  XNOR U4041 ( .A(n1823), .B(n1824), .Z(n1825) );
  XNOR U4042 ( .A(n1826), .B(n1825), .Z(n961) );
  XNOR U4043 ( .A(n962), .B(n961), .Z(n963) );
  XOR U4044 ( .A(n964), .B(n963), .Z(n1282) );
  XNOR U4045 ( .A(n1281), .B(n1282), .Z(n4825) );
  XOR U4046 ( .A(n4824), .B(n4825), .Z(n4826) );
  XOR U4047 ( .A(n4827), .B(n4826), .Z(n667) );
  XOR U4048 ( .A(n668), .B(n667), .Z(n669) );
  XOR U4049 ( .A(n670), .B(n669), .Z(n3804) );
  XOR U4050 ( .A(x[1283]), .B(y[1283]), .Z(n4034) );
  XOR U4051 ( .A(x[1281]), .B(y[1281]), .Z(n4032) );
  XNOR U4052 ( .A(x[1817]), .B(y[1817]), .Z(n4033) );
  XOR U4053 ( .A(n4032), .B(n4033), .Z(n4035) );
  XNOR U4054 ( .A(n4034), .B(n4035), .Z(n292) );
  XOR U4055 ( .A(x[7]), .B(y[7]), .Z(n455) );
  XOR U4056 ( .A(x[5]), .B(y[5]), .Z(n453) );
  XNOR U4057 ( .A(x[653]), .B(y[653]), .Z(n454) );
  XOR U4058 ( .A(n453), .B(n454), .Z(n456) );
  XOR U4059 ( .A(n455), .B(n456), .Z(n293) );
  XNOR U4060 ( .A(n292), .B(n293), .Z(n295) );
  XOR U4061 ( .A(x[1279]), .B(y[1279]), .Z(n4466) );
  XOR U4062 ( .A(x[1277]), .B(y[1277]), .Z(n4464) );
  XNOR U4063 ( .A(x[1571]), .B(y[1571]), .Z(n4465) );
  XOR U4064 ( .A(n4464), .B(n4465), .Z(n4467) );
  XNOR U4065 ( .A(n4466), .B(n4467), .Z(n294) );
  XOR U4066 ( .A(n295), .B(n294), .Z(n730) );
  XOR U4067 ( .A(x[1275]), .B(y[1275]), .Z(n4460) );
  XOR U4068 ( .A(x[1271]), .B(y[1271]), .Z(n4458) );
  XNOR U4069 ( .A(x[1819]), .B(y[1819]), .Z(n4459) );
  XOR U4070 ( .A(n4458), .B(n4459), .Z(n4461) );
  XNOR U4071 ( .A(n4460), .B(n4461), .Z(n334) );
  XOR U4072 ( .A(x[2]), .B(y[2]), .Z(n383) );
  XOR U4073 ( .A(x[4]), .B(y[4]), .Z(n381) );
  XNOR U4074 ( .A(x[6]), .B(y[6]), .Z(n382) );
  XOR U4075 ( .A(n381), .B(n382), .Z(n384) );
  XOR U4076 ( .A(n383), .B(n384), .Z(n335) );
  XNOR U4077 ( .A(n334), .B(n335), .Z(n337) );
  XOR U4078 ( .A(x[1269]), .B(y[1269]), .Z(n4472) );
  XOR U4079 ( .A(x[1267]), .B(y[1267]), .Z(n4470) );
  XNOR U4080 ( .A(x[1567]), .B(y[1567]), .Z(n4471) );
  XOR U4081 ( .A(n4470), .B(n4471), .Z(n4473) );
  XNOR U4082 ( .A(n4472), .B(n4473), .Z(n336) );
  XOR U4083 ( .A(n337), .B(n336), .Z(n728) );
  XOR U4084 ( .A(x[1459]), .B(y[1459]), .Z(n1030) );
  XOR U4085 ( .A(x[1455]), .B(y[1455]), .Z(n1027) );
  XNOR U4086 ( .A(x[1457]), .B(y[1457]), .Z(n1028) );
  XNOR U4087 ( .A(n1027), .B(n1028), .Z(n1029) );
  XOR U4088 ( .A(n1030), .B(n1029), .Z(n3350) );
  XOR U4089 ( .A(x[1465]), .B(y[1465]), .Z(n1018) );
  XOR U4090 ( .A(x[1461]), .B(y[1461]), .Z(n1015) );
  XNOR U4091 ( .A(x[1463]), .B(y[1463]), .Z(n1016) );
  XNOR U4092 ( .A(n1015), .B(n1016), .Z(n1017) );
  XOR U4093 ( .A(n1018), .B(n1017), .Z(n3348) );
  XOR U4094 ( .A(x[1473]), .B(y[1473]), .Z(n1024) );
  XOR U4095 ( .A(x[1467]), .B(y[1467]), .Z(n1021) );
  XNOR U4096 ( .A(x[1469]), .B(y[1469]), .Z(n1022) );
  XNOR U4097 ( .A(n1021), .B(n1022), .Z(n1023) );
  XNOR U4098 ( .A(n1024), .B(n1023), .Z(n3347) );
  XNOR U4099 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4100 ( .A(n3350), .B(n3349), .Z(n727) );
  XNOR U4101 ( .A(n728), .B(n727), .Z(n729) );
  XNOR U4102 ( .A(n730), .B(n729), .Z(n1527) );
  XOR U4103 ( .A(x[1287]), .B(y[1287]), .Z(n4041) );
  XOR U4104 ( .A(x[1285]), .B(y[1285]), .Z(n4038) );
  XNOR U4105 ( .A(x[1575]), .B(y[1575]), .Z(n4039) );
  XNOR U4106 ( .A(n4038), .B(n4039), .Z(n4040) );
  XOR U4107 ( .A(n4041), .B(n4040), .Z(n396) );
  XOR U4108 ( .A(x[1291]), .B(y[1291]), .Z(n1090) );
  XOR U4109 ( .A(x[1289]), .B(y[1289]), .Z(n1087) );
  XNOR U4110 ( .A(x[1815]), .B(y[1815]), .Z(n1088) );
  XNOR U4111 ( .A(n1087), .B(n1088), .Z(n1089) );
  XOR U4112 ( .A(n1090), .B(n1089), .Z(n394) );
  XOR U4113 ( .A(x[1295]), .B(y[1295]), .Z(n1084) );
  XOR U4114 ( .A(x[1293]), .B(y[1293]), .Z(n1081) );
  XNOR U4115 ( .A(x[1579]), .B(y[1579]), .Z(n1082) );
  XNOR U4116 ( .A(n1081), .B(n1082), .Z(n1083) );
  XNOR U4117 ( .A(n1084), .B(n1083), .Z(n393) );
  XNOR U4118 ( .A(n394), .B(n393), .Z(n395) );
  XNOR U4119 ( .A(n396), .B(n395), .Z(n673) );
  XOR U4120 ( .A(x[1441]), .B(y[1441]), .Z(n1306) );
  XOR U4121 ( .A(x[1437]), .B(y[1437]), .Z(n1303) );
  XNOR U4122 ( .A(x[1439]), .B(y[1439]), .Z(n1304) );
  XNOR U4123 ( .A(n1303), .B(n1304), .Z(n1305) );
  XOR U4124 ( .A(n1306), .B(n1305), .Z(n3566) );
  XOR U4125 ( .A(x[1447]), .B(y[1447]), .Z(n1120) );
  XOR U4126 ( .A(x[1443]), .B(y[1443]), .Z(n1117) );
  XNOR U4127 ( .A(x[1445]), .B(y[1445]), .Z(n1118) );
  XNOR U4128 ( .A(n1117), .B(n1118), .Z(n1119) );
  XOR U4129 ( .A(n1120), .B(n1119), .Z(n3564) );
  XOR U4130 ( .A(x[1453]), .B(y[1453]), .Z(n1114) );
  XOR U4131 ( .A(x[1449]), .B(y[1449]), .Z(n1111) );
  XNOR U4132 ( .A(x[1451]), .B(y[1451]), .Z(n1112) );
  XNOR U4133 ( .A(n1111), .B(n1112), .Z(n1113) );
  XNOR U4134 ( .A(n1114), .B(n1113), .Z(n3563) );
  XNOR U4135 ( .A(n3564), .B(n3563), .Z(n3565) );
  XOR U4136 ( .A(n3566), .B(n3565), .Z(n674) );
  XNOR U4137 ( .A(n673), .B(n674), .Z(n675) );
  XOR U4138 ( .A(x[1299]), .B(y[1299]), .Z(n1204) );
  XOR U4139 ( .A(x[1297]), .B(y[1297]), .Z(n1201) );
  XNOR U4140 ( .A(x[1813]), .B(y[1813]), .Z(n1202) );
  XNOR U4141 ( .A(n1201), .B(n1202), .Z(n1203) );
  XOR U4142 ( .A(n1204), .B(n1203), .Z(n468) );
  XOR U4143 ( .A(x[1303]), .B(y[1303]), .Z(n1192) );
  XOR U4144 ( .A(x[1301]), .B(y[1301]), .Z(n1189) );
  XNOR U4145 ( .A(x[1583]), .B(y[1583]), .Z(n1190) );
  XNOR U4146 ( .A(n1189), .B(n1190), .Z(n1191) );
  XOR U4147 ( .A(n1192), .B(n1191), .Z(n466) );
  XOR U4148 ( .A(x[1307]), .B(y[1307]), .Z(n1198) );
  XOR U4149 ( .A(x[1305]), .B(y[1305]), .Z(n1195) );
  XNOR U4150 ( .A(x[1811]), .B(y[1811]), .Z(n1196) );
  XNOR U4151 ( .A(n1195), .B(n1196), .Z(n1197) );
  XNOR U4152 ( .A(n1198), .B(n1197), .Z(n465) );
  XNOR U4153 ( .A(n466), .B(n465), .Z(n467) );
  XOR U4154 ( .A(n468), .B(n467), .Z(n676) );
  XNOR U4155 ( .A(n675), .B(n676), .Z(n1525) );
  XOR U4156 ( .A(x[1381]), .B(y[1381]), .Z(n4425) );
  XOR U4157 ( .A(x[1377]), .B(y[1377]), .Z(n4422) );
  XNOR U4158 ( .A(x[1379]), .B(y[1379]), .Z(n4423) );
  XNOR U4159 ( .A(n4422), .B(n4423), .Z(n4424) );
  XOR U4160 ( .A(n4425), .B(n4424), .Z(n3795) );
  XOR U4161 ( .A(x[1387]), .B(y[1387]), .Z(n4395) );
  XOR U4162 ( .A(x[1383]), .B(y[1383]), .Z(n4392) );
  XNOR U4163 ( .A(x[1385]), .B(y[1385]), .Z(n4393) );
  XNOR U4164 ( .A(n4392), .B(n4393), .Z(n4394) );
  XOR U4165 ( .A(n4395), .B(n4394), .Z(n3793) );
  XOR U4166 ( .A(x[1393]), .B(y[1393]), .Z(n4389) );
  XOR U4167 ( .A(x[1389]), .B(y[1389]), .Z(n4386) );
  XNOR U4168 ( .A(x[1391]), .B(y[1391]), .Z(n4387) );
  XNOR U4169 ( .A(n4386), .B(n4387), .Z(n4388) );
  XNOR U4170 ( .A(n4389), .B(n4388), .Z(n3792) );
  XNOR U4171 ( .A(n3793), .B(n3792), .Z(n3794) );
  XNOR U4172 ( .A(n3795), .B(n3794), .Z(n889) );
  XOR U4173 ( .A(x[1399]), .B(y[1399]), .Z(n4347) );
  XOR U4174 ( .A(x[1395]), .B(y[1395]), .Z(n4344) );
  XNOR U4175 ( .A(x[1397]), .B(y[1397]), .Z(n4345) );
  XNOR U4176 ( .A(n4344), .B(n4345), .Z(n4346) );
  XOR U4177 ( .A(n4347), .B(n4346), .Z(n3735) );
  XOR U4178 ( .A(x[1405]), .B(y[1405]), .Z(n4335) );
  XOR U4179 ( .A(x[1401]), .B(y[1401]), .Z(n4332) );
  XNOR U4180 ( .A(x[1403]), .B(y[1403]), .Z(n4333) );
  XNOR U4181 ( .A(n4332), .B(n4333), .Z(n4334) );
  XOR U4182 ( .A(n4335), .B(n4334), .Z(n3733) );
  XOR U4183 ( .A(x[1411]), .B(y[1411]), .Z(n4341) );
  XOR U4184 ( .A(x[1407]), .B(y[1407]), .Z(n4338) );
  XNOR U4185 ( .A(x[1409]), .B(y[1409]), .Z(n4339) );
  XNOR U4186 ( .A(n4338), .B(n4339), .Z(n4340) );
  XNOR U4187 ( .A(n4341), .B(n4340), .Z(n3732) );
  XNOR U4188 ( .A(n3733), .B(n3732), .Z(n3734) );
  XOR U4189 ( .A(n3735), .B(n3734), .Z(n890) );
  XNOR U4190 ( .A(n889), .B(n890), .Z(n891) );
  XOR U4191 ( .A(x[1369]), .B(y[1369]), .Z(n4293) );
  XOR U4192 ( .A(x[1365]), .B(y[1365]), .Z(n4290) );
  XNOR U4193 ( .A(x[1367]), .B(y[1367]), .Z(n4291) );
  XNOR U4194 ( .A(n4290), .B(n4291), .Z(n4292) );
  XOR U4195 ( .A(n4293), .B(n4292), .Z(n3044) );
  XOR U4196 ( .A(x[143]), .B(y[143]), .Z(n3783) );
  XOR U4197 ( .A(x[137]), .B(y[137]), .Z(n3780) );
  XNOR U4198 ( .A(x[141]), .B(y[141]), .Z(n3781) );
  XNOR U4199 ( .A(n3780), .B(n3781), .Z(n3782) );
  XOR U4200 ( .A(n3783), .B(n3782), .Z(n3042) );
  XOR U4201 ( .A(x[1375]), .B(y[1375]), .Z(n4431) );
  XOR U4202 ( .A(x[1371]), .B(y[1371]), .Z(n4428) );
  XNOR U4203 ( .A(x[1373]), .B(y[1373]), .Z(n4429) );
  XNOR U4204 ( .A(n4428), .B(n4429), .Z(n4430) );
  XNOR U4205 ( .A(n4431), .B(n4430), .Z(n3041) );
  XNOR U4206 ( .A(n3042), .B(n3041), .Z(n3043) );
  XOR U4207 ( .A(n3044), .B(n3043), .Z(n892) );
  XOR U4208 ( .A(n891), .B(n892), .Z(n1526) );
  XOR U4209 ( .A(n1525), .B(n1526), .Z(n1528) );
  XOR U4210 ( .A(n1527), .B(n1528), .Z(n3805) );
  XNOR U4211 ( .A(n3804), .B(n3805), .Z(n3807) );
  XOR U4212 ( .A(x[379]), .B(y[379]), .Z(n131) );
  XOR U4213 ( .A(x[377]), .B(y[377]), .Z(n128) );
  XNOR U4214 ( .A(x[985]), .B(y[985]), .Z(n129) );
  XNOR U4215 ( .A(n128), .B(n129), .Z(n130) );
  XOR U4216 ( .A(n131), .B(n130), .Z(n2900) );
  XOR U4217 ( .A(x[385]), .B(y[385]), .Z(n6009) );
  XOR U4218 ( .A(x[383]), .B(y[383]), .Z(n6006) );
  XNOR U4219 ( .A(x[991]), .B(y[991]), .Z(n6007) );
  XNOR U4220 ( .A(n6006), .B(n6007), .Z(n6008) );
  XOR U4221 ( .A(n6009), .B(n6008), .Z(n2898) );
  XOR U4222 ( .A(x[395]), .B(y[395]), .Z(n6003) );
  XOR U4223 ( .A(x[389]), .B(y[389]), .Z(n6000) );
  XNOR U4224 ( .A(x[391]), .B(y[391]), .Z(n6001) );
  XNOR U4225 ( .A(n6000), .B(n6001), .Z(n6002) );
  XNOR U4226 ( .A(n6003), .B(n6002), .Z(n2897) );
  XNOR U4227 ( .A(n2898), .B(n2897), .Z(n2899) );
  XNOR U4228 ( .A(n2900), .B(n2899), .Z(n1765) );
  XOR U4229 ( .A(x[405]), .B(y[405]), .Z(n4623) );
  XOR U4230 ( .A(x[399]), .B(y[399]), .Z(n4620) );
  XNOR U4231 ( .A(x[401]), .B(y[401]), .Z(n4621) );
  XNOR U4232 ( .A(n4620), .B(n4621), .Z(n4622) );
  XOR U4233 ( .A(n4623), .B(n4622), .Z(n3080) );
  XOR U4234 ( .A(x[452]), .B(y[452]), .Z(n688) );
  XOR U4235 ( .A(x[456]), .B(y[456]), .Z(n685) );
  XNOR U4236 ( .A(x[593]), .B(y[593]), .Z(n686) );
  XNOR U4237 ( .A(n685), .B(n686), .Z(n687) );
  XOR U4238 ( .A(n688), .B(n687), .Z(n3078) );
  XOR U4239 ( .A(x[417]), .B(y[417]), .Z(n3242) );
  XOR U4240 ( .A(x[413]), .B(y[413]), .Z(n3239) );
  XNOR U4241 ( .A(x[1013]), .B(y[1013]), .Z(n3240) );
  XNOR U4242 ( .A(n3239), .B(n3240), .Z(n3241) );
  XNOR U4243 ( .A(n3242), .B(n3241), .Z(n3077) );
  XNOR U4244 ( .A(n3078), .B(n3077), .Z(n3079) );
  XOR U4245 ( .A(n3080), .B(n3079), .Z(n1766) );
  XNOR U4246 ( .A(n1765), .B(n1766), .Z(n1768) );
  XOR U4247 ( .A(x[439]), .B(y[439]), .Z(n2882) );
  XOR U4248 ( .A(x[433]), .B(y[433]), .Z(n2879) );
  XNOR U4249 ( .A(x[437]), .B(y[437]), .Z(n2880) );
  XNOR U4250 ( .A(n2879), .B(n2880), .Z(n2881) );
  XOR U4251 ( .A(n2882), .B(n2881), .Z(n3765) );
  XOR U4252 ( .A(x[442]), .B(y[442]), .Z(n706) );
  XOR U4253 ( .A(x[444]), .B(y[444]), .Z(n703) );
  XNOR U4254 ( .A(x[1903]), .B(y[1903]), .Z(n704) );
  XNOR U4255 ( .A(n703), .B(n704), .Z(n705) );
  XOR U4256 ( .A(n706), .B(n705), .Z(n3763) );
  XOR U4257 ( .A(x[453]), .B(y[453]), .Z(n4929) );
  XOR U4258 ( .A(x[445]), .B(y[445]), .Z(n4926) );
  XNOR U4259 ( .A(x[1031]), .B(y[1031]), .Z(n4927) );
  XNOR U4260 ( .A(n4926), .B(n4927), .Z(n4928) );
  XNOR U4261 ( .A(n4929), .B(n4928), .Z(n3762) );
  XNOR U4262 ( .A(n3763), .B(n3762), .Z(n3764) );
  XNOR U4263 ( .A(n3765), .B(n3764), .Z(n1767) );
  XNOR U4264 ( .A(n1768), .B(n1767), .Z(n3945) );
  XOR U4265 ( .A(x[459]), .B(y[459]), .Z(n239) );
  XOR U4266 ( .A(x[457]), .B(y[457]), .Z(n236) );
  XNOR U4267 ( .A(x[1035]), .B(y[1035]), .Z(n237) );
  XNOR U4268 ( .A(n236), .B(n237), .Z(n238) );
  XOR U4269 ( .A(n239), .B(n238), .Z(n149) );
  XOR U4270 ( .A(x[473]), .B(y[473]), .Z(n4923) );
  XOR U4271 ( .A(x[465]), .B(y[465]), .Z(n4920) );
  XNOR U4272 ( .A(x[469]), .B(y[469]), .Z(n4921) );
  XNOR U4273 ( .A(n4920), .B(n4921), .Z(n4922) );
  XOR U4274 ( .A(n4923), .B(n4922), .Z(n147) );
  XOR U4275 ( .A(x[493]), .B(y[493]), .Z(n5295) );
  XOR U4276 ( .A(x[479]), .B(y[479]), .Z(n5292) );
  XNOR U4277 ( .A(x[489]), .B(y[489]), .Z(n5293) );
  XNOR U4278 ( .A(n5292), .B(n5293), .Z(n5294) );
  XNOR U4279 ( .A(n5295), .B(n5294), .Z(n146) );
  XNOR U4280 ( .A(n147), .B(n146), .Z(n148) );
  XNOR U4281 ( .A(n149), .B(n148), .Z(n1729) );
  XOR U4282 ( .A(x[499]), .B(y[499]), .Z(n5289) );
  XOR U4283 ( .A(x[495]), .B(y[495]), .Z(n5286) );
  XNOR U4284 ( .A(x[1053]), .B(y[1053]), .Z(n5287) );
  XNOR U4285 ( .A(n5286), .B(n5287), .Z(n5288) );
  XOR U4286 ( .A(n5289), .B(n5288), .Z(n5535) );
  XOR U4287 ( .A(x[529]), .B(y[529]), .Z(n2612) );
  XOR U4288 ( .A(x[515]), .B(y[515]), .Z(n2609) );
  XNOR U4289 ( .A(x[523]), .B(y[523]), .Z(n2610) );
  XNOR U4290 ( .A(n2609), .B(n2610), .Z(n2611) );
  XOR U4291 ( .A(n2612), .B(n2611), .Z(n5533) );
  XOR U4292 ( .A(x[551]), .B(y[551]), .Z(n510) );
  XOR U4293 ( .A(x[543]), .B(y[543]), .Z(n507) );
  XNOR U4294 ( .A(x[1075]), .B(y[1075]), .Z(n508) );
  XNOR U4295 ( .A(n507), .B(n508), .Z(n509) );
  XNOR U4296 ( .A(n510), .B(n509), .Z(n5532) );
  XNOR U4297 ( .A(n5533), .B(n5532), .Z(n5534) );
  XOR U4298 ( .A(n5535), .B(n5534), .Z(n1730) );
  XNOR U4299 ( .A(n1729), .B(n1730), .Z(n1732) );
  XOR U4300 ( .A(x[563]), .B(y[563]), .Z(n283) );
  XOR U4301 ( .A(x[559]), .B(y[559]), .Z(n280) );
  XNOR U4302 ( .A(x[1079]), .B(y[1079]), .Z(n281) );
  XNOR U4303 ( .A(n280), .B(n281), .Z(n282) );
  XOR U4304 ( .A(n283), .B(n282), .Z(n4701) );
  XOR U4305 ( .A(x[402]), .B(y[402]), .Z(n2078) );
  XOR U4306 ( .A(x[404]), .B(y[404]), .Z(n2075) );
  XNOR U4307 ( .A(x[927]), .B(y[927]), .Z(n2076) );
  XNOR U4308 ( .A(n2075), .B(n2076), .Z(n2077) );
  XOR U4309 ( .A(n2078), .B(n2077), .Z(n4699) );
  XOR U4310 ( .A(x[575]), .B(y[575]), .Z(n2912) );
  XOR U4311 ( .A(x[569]), .B(y[569]), .Z(n2909) );
  XNOR U4312 ( .A(x[571]), .B(y[571]), .Z(n2910) );
  XNOR U4313 ( .A(n2909), .B(n2910), .Z(n2911) );
  XNOR U4314 ( .A(n2912), .B(n2911), .Z(n4698) );
  XNOR U4315 ( .A(n4699), .B(n4698), .Z(n4700) );
  XNOR U4316 ( .A(n4701), .B(n4700), .Z(n1731) );
  XNOR U4317 ( .A(n1732), .B(n1731), .Z(n3943) );
  XOR U4318 ( .A(x[595]), .B(y[595]), .Z(n331) );
  XOR U4319 ( .A(x[577]), .B(y[577]), .Z(n328) );
  XNOR U4320 ( .A(x[589]), .B(y[589]), .Z(n329) );
  XNOR U4321 ( .A(n328), .B(n329), .Z(n330) );
  XOR U4322 ( .A(n331), .B(n330), .Z(n630) );
  XOR U4323 ( .A(x[394]), .B(y[394]), .Z(n2048) );
  XOR U4324 ( .A(x[396]), .B(y[396]), .Z(n2045) );
  XNOR U4325 ( .A(x[629]), .B(y[629]), .Z(n2046) );
  XNOR U4326 ( .A(n2045), .B(n2046), .Z(n2047) );
  XOR U4327 ( .A(n2048), .B(n2047), .Z(n628) );
  XOR U4328 ( .A(x[603]), .B(y[603]), .Z(n325) );
  XOR U4329 ( .A(x[597]), .B(y[597]), .Z(n322) );
  XNOR U4330 ( .A(x[1093]), .B(y[1093]), .Z(n323) );
  XNOR U4331 ( .A(n322), .B(n323), .Z(n324) );
  XNOR U4332 ( .A(n325), .B(n324), .Z(n627) );
  XNOR U4333 ( .A(n628), .B(n627), .Z(n629) );
  XNOR U4334 ( .A(n630), .B(n629), .Z(n1519) );
  XOR U4335 ( .A(x[611]), .B(y[611]), .Z(n167) );
  XOR U4336 ( .A(x[605]), .B(y[605]), .Z(n164) );
  XNOR U4337 ( .A(x[1097]), .B(y[1097]), .Z(n165) );
  XNOR U4338 ( .A(n164), .B(n165), .Z(n166) );
  XOR U4339 ( .A(n167), .B(n166), .Z(n5523) );
  XOR U4340 ( .A(x[643]), .B(y[643]), .Z(n161) );
  XOR U4341 ( .A(x[633]), .B(y[633]), .Z(n158) );
  XNOR U4342 ( .A(x[637]), .B(y[637]), .Z(n159) );
  XNOR U4343 ( .A(n158), .B(n159), .Z(n160) );
  XOR U4344 ( .A(n161), .B(n160), .Z(n5521) );
  XOR U4345 ( .A(x[665]), .B(y[665]), .Z(n95) );
  XOR U4346 ( .A(x[657]), .B(y[657]), .Z(n92) );
  XNOR U4347 ( .A(x[1115]), .B(y[1115]), .Z(n93) );
  XNOR U4348 ( .A(n92), .B(n93), .Z(n94) );
  XNOR U4349 ( .A(n95), .B(n94), .Z(n5520) );
  XNOR U4350 ( .A(n5521), .B(n5520), .Z(n5522) );
  XOR U4351 ( .A(n5523), .B(n5522), .Z(n1520) );
  XNOR U4352 ( .A(n1519), .B(n1520), .Z(n1522) );
  XOR U4353 ( .A(x[677]), .B(y[677]), .Z(n83) );
  XOR U4354 ( .A(x[671]), .B(y[671]), .Z(n80) );
  XNOR U4355 ( .A(x[673]), .B(y[673]), .Z(n81) );
  XNOR U4356 ( .A(n80), .B(n81), .Z(n82) );
  XOR U4357 ( .A(n83), .B(n82), .Z(n4707) );
  XOR U4358 ( .A(x[693]), .B(y[693]), .Z(n89) );
  XOR U4359 ( .A(x[679]), .B(y[679]), .Z(n86) );
  XNOR U4360 ( .A(x[685]), .B(y[685]), .Z(n87) );
  XNOR U4361 ( .A(n86), .B(n87), .Z(n88) );
  XOR U4362 ( .A(n89), .B(n88), .Z(n4705) );
  XOR U4363 ( .A(x[705]), .B(y[705]), .Z(n2702) );
  XOR U4364 ( .A(x[699]), .B(y[699]), .Z(n2699) );
  XNOR U4365 ( .A(x[1129]), .B(y[1129]), .Z(n2700) );
  XNOR U4366 ( .A(n2699), .B(n2700), .Z(n2701) );
  XNOR U4367 ( .A(n2702), .B(n2701), .Z(n4704) );
  XNOR U4368 ( .A(n4705), .B(n4704), .Z(n4706) );
  XNOR U4369 ( .A(n4707), .B(n4706), .Z(n1521) );
  XNOR U4370 ( .A(n1522), .B(n1521), .Z(n3942) );
  XOR U4371 ( .A(n3943), .B(n3942), .Z(n3944) );
  XNOR U4372 ( .A(n3945), .B(n3944), .Z(n952) );
  XOR U4373 ( .A(x[153]), .B(y[153]), .Z(n4419) );
  XOR U4374 ( .A(x[147]), .B(y[147]), .Z(n4416) );
  XNOR U4375 ( .A(x[149]), .B(y[149]), .Z(n4417) );
  XNOR U4376 ( .A(n4416), .B(n4417), .Z(n4418) );
  XOR U4377 ( .A(n4419), .B(n4418), .Z(n576) );
  XOR U4378 ( .A(x[159]), .B(y[159]), .Z(n3729) );
  XOR U4379 ( .A(x[157]), .B(y[157]), .Z(n3726) );
  XNOR U4380 ( .A(x[829]), .B(y[829]), .Z(n3727) );
  XNOR U4381 ( .A(n3726), .B(n3727), .Z(n3728) );
  XOR U4382 ( .A(n3729), .B(n3728), .Z(n574) );
  XOR U4383 ( .A(x[165]), .B(y[165]), .Z(n4383) );
  XOR U4384 ( .A(x[163]), .B(y[163]), .Z(n4380) );
  XNOR U4385 ( .A(x[833]), .B(y[833]), .Z(n4381) );
  XNOR U4386 ( .A(n4380), .B(n4381), .Z(n4382) );
  XNOR U4387 ( .A(n4383), .B(n4382), .Z(n573) );
  XNOR U4388 ( .A(n574), .B(n573), .Z(n575) );
  XNOR U4389 ( .A(n576), .B(n575), .Z(n3822) );
  XOR U4390 ( .A(x[175]), .B(y[175]), .Z(n3723) );
  XOR U4391 ( .A(x[169]), .B(y[169]), .Z(n3720) );
  XNOR U4392 ( .A(x[171]), .B(y[171]), .Z(n3721) );
  XNOR U4393 ( .A(n3720), .B(n3721), .Z(n3722) );
  XOR U4394 ( .A(n3723), .B(n3722), .Z(n582) );
  XOR U4395 ( .A(x[185]), .B(y[185]), .Z(n3711) );
  XOR U4396 ( .A(x[179]), .B(y[179]), .Z(n3708) );
  XNOR U4397 ( .A(x[181]), .B(y[181]), .Z(n3709) );
  XNOR U4398 ( .A(n3708), .B(n3709), .Z(n3710) );
  XOR U4399 ( .A(n3711), .B(n3710), .Z(n580) );
  XOR U4400 ( .A(x[191]), .B(y[191]), .Z(n3705) );
  XOR U4401 ( .A(x[187]), .B(y[187]), .Z(n3702) );
  XNOR U4402 ( .A(x[851]), .B(y[851]), .Z(n3703) );
  XNOR U4403 ( .A(n3702), .B(n3703), .Z(n3704) );
  XNOR U4404 ( .A(n3705), .B(n3704), .Z(n579) );
  XNOR U4405 ( .A(n580), .B(n579), .Z(n581) );
  XOR U4406 ( .A(n582), .B(n581), .Z(n3823) );
  XNOR U4407 ( .A(n3822), .B(n3823), .Z(n3825) );
  XOR U4408 ( .A(x[207]), .B(y[207]), .Z(n3482) );
  XOR U4409 ( .A(x[201]), .B(y[201]), .Z(n3479) );
  XNOR U4410 ( .A(x[203]), .B(y[203]), .Z(n3480) );
  XNOR U4411 ( .A(n3479), .B(n3480), .Z(n3481) );
  XOR U4412 ( .A(n3482), .B(n3481), .Z(n2990) );
  XOR U4413 ( .A(x[558]), .B(y[558]), .Z(n1886) );
  XOR U4414 ( .A(x[531]), .B(y[531]), .Z(n1883) );
  XNOR U4415 ( .A(x[560]), .B(y[560]), .Z(n1884) );
  XNOR U4416 ( .A(n1883), .B(n1884), .Z(n1885) );
  XOR U4417 ( .A(n1886), .B(n1885), .Z(n2988) );
  XOR U4418 ( .A(x[223]), .B(y[223]), .Z(n1300) );
  XOR U4419 ( .A(x[219]), .B(y[219]), .Z(n1297) );
  XNOR U4420 ( .A(x[873]), .B(y[873]), .Z(n1298) );
  XNOR U4421 ( .A(n1297), .B(n1298), .Z(n1299) );
  XNOR U4422 ( .A(n1300), .B(n1299), .Z(n2987) );
  XNOR U4423 ( .A(n2988), .B(n2987), .Z(n2989) );
  XNOR U4424 ( .A(n2990), .B(n2989), .Z(n3824) );
  XNOR U4425 ( .A(n3825), .B(n3824), .Z(n3939) );
  XOR U4426 ( .A(x[373]), .B(y[373]), .Z(n3253) );
  XOR U4427 ( .A(x[367]), .B(y[367]), .Z(n3251) );
  XNOR U4428 ( .A(x[369]), .B(y[369]), .Z(n3252) );
  XOR U4429 ( .A(n3251), .B(n3252), .Z(n3254) );
  XNOR U4430 ( .A(n3253), .B(n3254), .Z(n230) );
  XOR U4431 ( .A(x[363]), .B(y[363]), .Z(n1035) );
  XOR U4432 ( .A(x[357]), .B(y[357]), .Z(n1033) );
  XNOR U4433 ( .A(x[361]), .B(y[361]), .Z(n1034) );
  XOR U4434 ( .A(n1033), .B(n1034), .Z(n1036) );
  XOR U4435 ( .A(n1035), .B(n1036), .Z(n231) );
  XNOR U4436 ( .A(n230), .B(n231), .Z(n233) );
  XOR U4437 ( .A(x[347]), .B(y[347]), .Z(n3367) );
  XOR U4438 ( .A(x[345]), .B(y[345]), .Z(n3365) );
  XNOR U4439 ( .A(x[963]), .B(y[963]), .Z(n3366) );
  XOR U4440 ( .A(n3365), .B(n3366), .Z(n3368) );
  XNOR U4441 ( .A(n3367), .B(n3368), .Z(n232) );
  XOR U4442 ( .A(n233), .B(n232), .Z(n1774) );
  XOR U4443 ( .A(x[311]), .B(y[311]), .Z(n970) );
  XOR U4444 ( .A(x[303]), .B(y[303]), .Z(n967) );
  XNOR U4445 ( .A(x[307]), .B(y[307]), .Z(n968) );
  XNOR U4446 ( .A(n967), .B(n968), .Z(n969) );
  XOR U4447 ( .A(n970), .B(n969), .Z(n624) );
  XOR U4448 ( .A(x[508]), .B(y[508]), .Z(n760) );
  XOR U4449 ( .A(x[510]), .B(y[510]), .Z(n757) );
  XNOR U4450 ( .A(x[881]), .B(y[881]), .Z(n758) );
  XNOR U4451 ( .A(n757), .B(n758), .Z(n759) );
  XOR U4452 ( .A(n760), .B(n759), .Z(n622) );
  XOR U4453 ( .A(x[317]), .B(y[317]), .Z(n3608) );
  XOR U4454 ( .A(x[313]), .B(y[313]), .Z(n3605) );
  XNOR U4455 ( .A(x[939]), .B(y[939]), .Z(n3606) );
  XNOR U4456 ( .A(n3605), .B(n3606), .Z(n3607) );
  XNOR U4457 ( .A(n3608), .B(n3607), .Z(n621) );
  XNOR U4458 ( .A(n622), .B(n621), .Z(n623) );
  XNOR U4459 ( .A(n624), .B(n623), .Z(n1772) );
  XOR U4460 ( .A(x[323]), .B(y[323]), .Z(n3631) );
  XOR U4461 ( .A(x[319]), .B(y[319]), .Z(n3629) );
  XNOR U4462 ( .A(x[945]), .B(y[945]), .Z(n3630) );
  XOR U4463 ( .A(n3629), .B(n3630), .Z(n3632) );
  XOR U4464 ( .A(n3631), .B(n3632), .Z(n425) );
  XOR U4465 ( .A(x[492]), .B(y[492]), .Z(n801) );
  XOR U4466 ( .A(x[498]), .B(y[498]), .Z(n799) );
  XNOR U4467 ( .A(x[887]), .B(y[887]), .Z(n800) );
  XOR U4468 ( .A(n799), .B(n800), .Z(n802) );
  XOR U4469 ( .A(n801), .B(n802), .Z(n424) );
  XOR U4470 ( .A(x[333]), .B(y[333]), .Z(n3626) );
  XOR U4471 ( .A(x[325]), .B(y[325]), .Z(n3623) );
  XNOR U4472 ( .A(x[329]), .B(y[329]), .Z(n3624) );
  XNOR U4473 ( .A(n3623), .B(n3624), .Z(n3625) );
  XNOR U4474 ( .A(n3626), .B(n3625), .Z(n423) );
  XOR U4475 ( .A(n424), .B(n423), .Z(n426) );
  XOR U4476 ( .A(n425), .B(n426), .Z(n1771) );
  XOR U4477 ( .A(n1772), .B(n1771), .Z(n1773) );
  XOR U4478 ( .A(n1774), .B(n1773), .Z(n3937) );
  XOR U4479 ( .A(x[229]), .B(y[229]), .Z(n3554) );
  XOR U4480 ( .A(x[225]), .B(y[225]), .Z(n3551) );
  XNOR U4481 ( .A(x[877]), .B(y[877]), .Z(n3552) );
  XNOR U4482 ( .A(n3551), .B(n3552), .Z(n3553) );
  XOR U4483 ( .A(n3554), .B(n3553), .Z(n498) );
  XOR U4484 ( .A(x[550]), .B(y[550]), .Z(n1916) );
  XOR U4485 ( .A(x[537]), .B(y[537]), .Z(n1913) );
  XNOR U4486 ( .A(x[552]), .B(y[552]), .Z(n1914) );
  XNOR U4487 ( .A(n1913), .B(n1914), .Z(n1915) );
  XOR U4488 ( .A(n1916), .B(n1915), .Z(n496) );
  XOR U4489 ( .A(x[237]), .B(y[237]), .Z(n1108) );
  XOR U4490 ( .A(x[231]), .B(y[231]), .Z(n1105) );
  XNOR U4491 ( .A(x[235]), .B(y[235]), .Z(n1106) );
  XNOR U4492 ( .A(n1105), .B(n1106), .Z(n1107) );
  XNOR U4493 ( .A(n1108), .B(n1107), .Z(n495) );
  XNOR U4494 ( .A(n496), .B(n495), .Z(n497) );
  XNOR U4495 ( .A(n498), .B(n497), .Z(n3882) );
  XOR U4496 ( .A(x[247]), .B(y[247]), .Z(n3344) );
  XOR U4497 ( .A(x[241]), .B(y[241]), .Z(n3341) );
  XNOR U4498 ( .A(x[245]), .B(y[245]), .Z(n3342) );
  XNOR U4499 ( .A(n3341), .B(n3342), .Z(n3343) );
  XOR U4500 ( .A(n3344), .B(n3343), .Z(n2930) );
  XOR U4501 ( .A(x[253]), .B(y[253]), .Z(n3338) );
  XOR U4502 ( .A(x[251]), .B(y[251]), .Z(n3335) );
  XNOR U4503 ( .A(x[895]), .B(y[895]), .Z(n3336) );
  XNOR U4504 ( .A(n3335), .B(n3336), .Z(n3337) );
  XOR U4505 ( .A(n3338), .B(n3337), .Z(n2928) );
  XOR U4506 ( .A(x[259]), .B(y[259]), .Z(n3446) );
  XOR U4507 ( .A(x[257]), .B(y[257]), .Z(n3443) );
  XNOR U4508 ( .A(x[899]), .B(y[899]), .Z(n3444) );
  XNOR U4509 ( .A(n3443), .B(n3444), .Z(n3445) );
  XNOR U4510 ( .A(n3446), .B(n3445), .Z(n2927) );
  XNOR U4511 ( .A(n2928), .B(n2927), .Z(n2929) );
  XOR U4512 ( .A(n2930), .B(n2929), .Z(n3883) );
  XNOR U4513 ( .A(n3882), .B(n3883), .Z(n3885) );
  XOR U4514 ( .A(x[279]), .B(y[279]), .Z(n2636) );
  XOR U4515 ( .A(x[273]), .B(y[273]), .Z(n2633) );
  XNOR U4516 ( .A(x[275]), .B(y[275]), .Z(n2634) );
  XNOR U4517 ( .A(n2633), .B(n2634), .Z(n2635) );
  XOR U4518 ( .A(n2636), .B(n2635), .Z(n528) );
  XOR U4519 ( .A(x[291]), .B(y[291]), .Z(n1672) );
  XOR U4520 ( .A(x[289]), .B(y[289]), .Z(n1669) );
  XNOR U4521 ( .A(x[923]), .B(y[923]), .Z(n1670) );
  XNOR U4522 ( .A(n1669), .B(n1670), .Z(n1671) );
  XOR U4523 ( .A(n1672), .B(n1671), .Z(n526) );
  XOR U4524 ( .A(x[301]), .B(y[301]), .Z(n3614) );
  XOR U4525 ( .A(x[295]), .B(y[295]), .Z(n3611) );
  XNOR U4526 ( .A(x[297]), .B(y[297]), .Z(n3612) );
  XNOR U4527 ( .A(n3611), .B(n3612), .Z(n3613) );
  XNOR U4528 ( .A(n3614), .B(n3613), .Z(n525) );
  XNOR U4529 ( .A(n526), .B(n525), .Z(n527) );
  XNOR U4530 ( .A(n528), .B(n527), .Z(n3884) );
  XNOR U4531 ( .A(n3885), .B(n3884), .Z(n3936) );
  XOR U4532 ( .A(n3937), .B(n3936), .Z(n3938) );
  XNOR U4533 ( .A(n3939), .B(n3938), .Z(n950) );
  XOR U4534 ( .A(x[3]), .B(y[3]), .Z(n461) );
  XOR U4535 ( .A(x[0]), .B(y[0]), .Z(n459) );
  XNOR U4536 ( .A(x[1]), .B(y[1]), .Z(n460) );
  XOR U4537 ( .A(n459), .B(n460), .Z(n462) );
  XNOR U4538 ( .A(n461), .B(n462), .Z(n224) );
  XOR U4539 ( .A(x[8]), .B(y[8]), .Z(n389) );
  XOR U4540 ( .A(x[10]), .B(y[10]), .Z(n387) );
  XNOR U4541 ( .A(x[625]), .B(y[625]), .Z(n388) );
  XOR U4542 ( .A(n387), .B(n388), .Z(n390) );
  XOR U4543 ( .A(n389), .B(n390), .Z(n225) );
  XNOR U4544 ( .A(n224), .B(n225), .Z(n226) );
  XOR U4545 ( .A(x[12]), .B(y[12]), .Z(n306) );
  XOR U4546 ( .A(x[14]), .B(y[14]), .Z(n304) );
  XNOR U4547 ( .A(x[617]), .B(y[617]), .Z(n305) );
  XOR U4548 ( .A(n304), .B(n305), .Z(n307) );
  XOR U4549 ( .A(n306), .B(n307), .Z(n227) );
  XOR U4550 ( .A(n226), .B(n227), .Z(n4514) );
  XOR U4551 ( .A(x[32]), .B(y[32]), .Z(n5805) );
  XOR U4552 ( .A(x[34]), .B(y[34]), .Z(n5802) );
  XNOR U4553 ( .A(x[583]), .B(y[583]), .Z(n5803) );
  XNOR U4554 ( .A(n5802), .B(n5803), .Z(n5804) );
  XOR U4555 ( .A(n5805), .B(n5804), .Z(n3056) );
  XOR U4556 ( .A(x[744]), .B(y[744]), .Z(n319) );
  XOR U4557 ( .A(x[746]), .B(y[746]), .Z(n316) );
  XNOR U4558 ( .A(x[1998]), .B(y[1998]), .Z(n317) );
  XNOR U4559 ( .A(n316), .B(n317), .Z(n318) );
  XOR U4560 ( .A(n319), .B(n318), .Z(n3054) );
  XOR U4561 ( .A(x[28]), .B(y[28]), .Z(n349) );
  XOR U4562 ( .A(x[30]), .B(y[30]), .Z(n346) );
  XNOR U4563 ( .A(x[591]), .B(y[591]), .Z(n347) );
  XNOR U4564 ( .A(n346), .B(n347), .Z(n348) );
  XNOR U4565 ( .A(n349), .B(n348), .Z(n3053) );
  XNOR U4566 ( .A(n3054), .B(n3053), .Z(n3055) );
  XNOR U4567 ( .A(n3056), .B(n3055), .Z(n4513) );
  XOR U4568 ( .A(x[16]), .B(y[16]), .Z(n312) );
  XOR U4569 ( .A(x[18]), .B(y[18]), .Z(n310) );
  XNOR U4570 ( .A(x[20]), .B(y[20]), .Z(n311) );
  XOR U4571 ( .A(n310), .B(n311), .Z(n313) );
  XNOR U4572 ( .A(n312), .B(n313), .Z(n2873) );
  XOR U4573 ( .A(x[1142]), .B(y[1142]), .Z(n2485) );
  XOR U4574 ( .A(x[561]), .B(y[561]), .Z(n2483) );
  XNOR U4575 ( .A(x[1144]), .B(y[1144]), .Z(n2484) );
  XOR U4576 ( .A(n2483), .B(n2484), .Z(n2486) );
  XOR U4577 ( .A(n2485), .B(n2486), .Z(n2874) );
  XNOR U4578 ( .A(n2873), .B(n2874), .Z(n2875) );
  XOR U4579 ( .A(x[22]), .B(y[22]), .Z(n5642) );
  XOR U4580 ( .A(x[24]), .B(y[24]), .Z(n5640) );
  XNOR U4581 ( .A(x[26]), .B(y[26]), .Z(n5641) );
  XOR U4582 ( .A(n5640), .B(n5641), .Z(n5643) );
  XOR U4583 ( .A(n5642), .B(n5643), .Z(n2876) );
  XOR U4584 ( .A(n2875), .B(n2876), .Z(n4512) );
  XOR U4585 ( .A(n4513), .B(n4512), .Z(n4515) );
  XOR U4586 ( .A(n4514), .B(n4515), .Z(n4958) );
  XOR U4587 ( .A(x[81]), .B(y[81]), .Z(n3831) );
  XOR U4588 ( .A(x[75]), .B(y[75]), .Z(n3828) );
  XNOR U4589 ( .A(x[77]), .B(y[77]), .Z(n3829) );
  XNOR U4590 ( .A(n3828), .B(n3829), .Z(n3830) );
  XOR U4591 ( .A(n3831), .B(n3830), .Z(n2906) );
  XOR U4592 ( .A(x[91]), .B(y[91]), .Z(n3002) );
  XOR U4593 ( .A(x[83]), .B(y[83]), .Z(n2999) );
  XNOR U4594 ( .A(x[87]), .B(y[87]), .Z(n3000) );
  XNOR U4595 ( .A(n2999), .B(n3000), .Z(n3001) );
  XOR U4596 ( .A(n3002), .B(n3001), .Z(n2904) );
  XOR U4597 ( .A(x[97]), .B(y[97]), .Z(n1264) );
  XOR U4598 ( .A(x[93]), .B(y[93]), .Z(n1261) );
  XNOR U4599 ( .A(x[759]), .B(y[759]), .Z(n1262) );
  XNOR U4600 ( .A(n1261), .B(n1262), .Z(n1263) );
  XNOR U4601 ( .A(n1264), .B(n1263), .Z(n2903) );
  XNOR U4602 ( .A(n2904), .B(n2903), .Z(n2905) );
  XNOR U4603 ( .A(n2906), .B(n2905), .Z(n4302) );
  XOR U4604 ( .A(x[103]), .B(y[103]), .Z(n546) );
  XOR U4605 ( .A(x[99]), .B(y[99]), .Z(n543) );
  XNOR U4606 ( .A(x[769]), .B(y[769]), .Z(n544) );
  XNOR U4607 ( .A(n543), .B(n544), .Z(n545) );
  XOR U4608 ( .A(n546), .B(n545), .Z(n474) );
  XOR U4609 ( .A(x[616]), .B(y[616]), .Z(n636) );
  XOR U4610 ( .A(x[497]), .B(y[497]), .Z(n633) );
  XNOR U4611 ( .A(x[618]), .B(y[618]), .Z(n634) );
  XNOR U4612 ( .A(n633), .B(n634), .Z(n635) );
  XOR U4613 ( .A(n636), .B(n635), .Z(n472) );
  XOR U4614 ( .A(x[113]), .B(y[113]), .Z(n540) );
  XOR U4615 ( .A(x[105]), .B(y[105]), .Z(n537) );
  XNOR U4616 ( .A(x[109]), .B(y[109]), .Z(n538) );
  XNOR U4617 ( .A(n537), .B(n538), .Z(n539) );
  XNOR U4618 ( .A(n540), .B(n539), .Z(n471) );
  XNOR U4619 ( .A(n472), .B(n471), .Z(n473) );
  XOR U4620 ( .A(n474), .B(n473), .Z(n4303) );
  XNOR U4621 ( .A(n4302), .B(n4303), .Z(n4304) );
  XOR U4622 ( .A(x[121]), .B(y[121]), .Z(n444) );
  XOR U4623 ( .A(x[115]), .B(y[115]), .Z(n441) );
  XNOR U4624 ( .A(x[119]), .B(y[119]), .Z(n442) );
  XNOR U4625 ( .A(n441), .B(n442), .Z(n443) );
  XOR U4626 ( .A(n444), .B(n443), .Z(n2966) );
  XOR U4627 ( .A(x[604]), .B(y[604]), .Z(n1940) );
  XOR U4628 ( .A(x[608]), .B(y[608]), .Z(n1937) );
  XNOR U4629 ( .A(x[841]), .B(y[841]), .Z(n1938) );
  XNOR U4630 ( .A(n1937), .B(n1938), .Z(n1939) );
  XOR U4631 ( .A(n1940), .B(n1939), .Z(n2964) );
  XOR U4632 ( .A(x[135]), .B(y[135]), .Z(n3789) );
  XOR U4633 ( .A(x[131]), .B(y[131]), .Z(n3786) );
  XNOR U4634 ( .A(x[803]), .B(y[803]), .Z(n3787) );
  XNOR U4635 ( .A(n3786), .B(n3787), .Z(n3788) );
  XNOR U4636 ( .A(n3789), .B(n3788), .Z(n2963) );
  XNOR U4637 ( .A(n2964), .B(n2963), .Z(n2965) );
  XOR U4638 ( .A(n2966), .B(n2965), .Z(n4305) );
  XNOR U4639 ( .A(n4304), .B(n4305), .Z(n4956) );
  XOR U4640 ( .A(x[11]), .B(y[11]), .Z(n4046) );
  XOR U4641 ( .A(x[9]), .B(y[9]), .Z(n4044) );
  XNOR U4642 ( .A(x[659]), .B(y[659]), .Z(n4045) );
  XOR U4643 ( .A(n4044), .B(n4045), .Z(n4047) );
  XOR U4644 ( .A(n4046), .B(n4047), .Z(n401) );
  XOR U4645 ( .A(x[674]), .B(y[674]), .Z(n2665) );
  XOR U4646 ( .A(x[676]), .B(y[676]), .Z(n2663) );
  XNOR U4647 ( .A(x[1921]), .B(y[1921]), .Z(n2664) );
  XOR U4648 ( .A(n2663), .B(n2664), .Z(n2666) );
  XOR U4649 ( .A(n2665), .B(n2666), .Z(n400) );
  XOR U4650 ( .A(x[17]), .B(y[17]), .Z(n564) );
  XOR U4651 ( .A(x[13]), .B(y[13]), .Z(n561) );
  XNOR U4652 ( .A(x[15]), .B(y[15]), .Z(n562) );
  XNOR U4653 ( .A(n561), .B(n562), .Z(n563) );
  XNOR U4654 ( .A(n564), .B(n563), .Z(n399) );
  XOR U4655 ( .A(n400), .B(n399), .Z(n402) );
  XOR U4656 ( .A(n401), .B(n402), .Z(n1775) );
  XOR U4657 ( .A(x[27]), .B(y[27]), .Z(n1078) );
  XOR U4658 ( .A(x[21]), .B(y[21]), .Z(n1075) );
  XNOR U4659 ( .A(x[25]), .B(y[25]), .Z(n1076) );
  XNOR U4660 ( .A(n1075), .B(n1076), .Z(n1077) );
  XOR U4661 ( .A(n1078), .B(n1077), .Z(n600) );
  XOR U4662 ( .A(x[664]), .B(y[664]), .Z(n2660) );
  XOR U4663 ( .A(x[475]), .B(y[475]), .Z(n2657) );
  XNOR U4664 ( .A(x[666]), .B(y[666]), .Z(n2658) );
  XNOR U4665 ( .A(n2657), .B(n2658), .Z(n2659) );
  XOR U4666 ( .A(n2660), .B(n2659), .Z(n598) );
  XOR U4667 ( .A(x[33]), .B(y[33]), .Z(n558) );
  XOR U4668 ( .A(x[31]), .B(y[31]), .Z(n555) );
  XNOR U4669 ( .A(x[689]), .B(y[689]), .Z(n556) );
  XNOR U4670 ( .A(n555), .B(n556), .Z(n557) );
  XNOR U4671 ( .A(n558), .B(n557), .Z(n597) );
  XNOR U4672 ( .A(n598), .B(n597), .Z(n599) );
  XOR U4673 ( .A(n600), .B(n599), .Z(n1776) );
  XNOR U4674 ( .A(n1775), .B(n1776), .Z(n1777) );
  XOR U4675 ( .A(x[39]), .B(y[39]), .Z(n3032) );
  XOR U4676 ( .A(x[37]), .B(y[37]), .Z(n3029) );
  XNOR U4677 ( .A(x[697]), .B(y[697]), .Z(n3030) );
  XNOR U4678 ( .A(n3029), .B(n3030), .Z(n3031) );
  XOR U4679 ( .A(n3032), .B(n3031), .Z(n504) );
  XOR U4680 ( .A(x[49]), .B(y[49]), .Z(n3026) );
  XOR U4681 ( .A(x[43]), .B(y[43]), .Z(n3023) );
  XNOR U4682 ( .A(x[47]), .B(y[47]), .Z(n3024) );
  XNOR U4683 ( .A(n3023), .B(n3024), .Z(n3025) );
  XOR U4684 ( .A(n3026), .B(n3025), .Z(n502) );
  XOR U4685 ( .A(x[65]), .B(y[65]), .Z(n203) );
  XOR U4686 ( .A(x[61]), .B(y[61]), .Z(n200) );
  XNOR U4687 ( .A(x[725]), .B(y[725]), .Z(n201) );
  XNOR U4688 ( .A(n200), .B(n201), .Z(n202) );
  XNOR U4689 ( .A(n203), .B(n202), .Z(n501) );
  XNOR U4690 ( .A(n502), .B(n501), .Z(n503) );
  XOR U4691 ( .A(n504), .B(n503), .Z(n1778) );
  XOR U4692 ( .A(n1777), .B(n1778), .Z(n4957) );
  XOR U4693 ( .A(n4956), .B(n4957), .Z(n4959) );
  XNOR U4694 ( .A(n4958), .B(n4959), .Z(n949) );
  XOR U4695 ( .A(n950), .B(n949), .Z(n951) );
  XOR U4696 ( .A(n952), .B(n951), .Z(n3806) );
  XOR U4697 ( .A(n3807), .B(n3806), .Z(n3901) );
  XOR U4698 ( .A(x[1680]), .B(y[1680]), .Z(n5979) );
  XOR U4699 ( .A(x[454]), .B(y[454]), .Z(n5976) );
  XNOR U4700 ( .A(x[1682]), .B(y[1682]), .Z(n5977) );
  XNOR U4701 ( .A(n5976), .B(n5977), .Z(n5978) );
  XOR U4702 ( .A(n5979), .B(n5978), .Z(n5247) );
  XOR U4703 ( .A(x[1824]), .B(y[1824]), .Z(n5553) );
  XOR U4704 ( .A(x[586]), .B(y[586]), .Z(n5550) );
  XNOR U4705 ( .A(x[1826]), .B(y[1826]), .Z(n5551) );
  XNOR U4706 ( .A(n5550), .B(n5551), .Z(n5552) );
  XOR U4707 ( .A(n5553), .B(n5552), .Z(n5245) );
  XOR U4708 ( .A(x[1676]), .B(y[1676]), .Z(n3518) );
  XOR U4709 ( .A(x[450]), .B(y[450]), .Z(n3515) );
  XNOR U4710 ( .A(x[1678]), .B(y[1678]), .Z(n3516) );
  XNOR U4711 ( .A(n3515), .B(n3516), .Z(n3517) );
  XNOR U4712 ( .A(n3518), .B(n3517), .Z(n5244) );
  XNOR U4713 ( .A(n5245), .B(n5244), .Z(n5246) );
  XNOR U4714 ( .A(n5247), .B(n5246), .Z(n5952) );
  XOR U4715 ( .A(x[1655]), .B(y[1655]), .Z(n516) );
  XOR U4716 ( .A(x[1701]), .B(y[1701]), .Z(n514) );
  XOR U4717 ( .A(x[1731]), .B(y[1731]), .Z(n513) );
  XOR U4718 ( .A(n514), .B(n513), .Z(n515) );
  XOR U4719 ( .A(n516), .B(n515), .Z(n4887) );
  XOR U4720 ( .A(x[1673]), .B(y[1673]), .Z(n2924) );
  XOR U4721 ( .A(x[1699]), .B(y[1699]), .Z(n2922) );
  XOR U4722 ( .A(x[1729]), .B(y[1729]), .Z(n2921) );
  XOR U4723 ( .A(n2922), .B(n2921), .Z(n2923) );
  XOR U4724 ( .A(n2924), .B(n2923), .Z(n4885) );
  XOR U4725 ( .A(x[1675]), .B(y[1675]), .Z(n2918) );
  XOR U4726 ( .A(x[1695]), .B(y[1695]), .Z(n2916) );
  XOR U4727 ( .A(x[1727]), .B(y[1727]), .Z(n2915) );
  XOR U4728 ( .A(n2916), .B(n2915), .Z(n2917) );
  XNOR U4729 ( .A(n2918), .B(n2917), .Z(n4884) );
  XNOR U4730 ( .A(n4885), .B(n4884), .Z(n4886) );
  XOR U4731 ( .A(n4887), .B(n4886), .Z(n5953) );
  XNOR U4732 ( .A(n5952), .B(n5953), .Z(n5955) );
  XOR U4733 ( .A(x[1670]), .B(y[1670]), .Z(n3530) );
  XOR U4734 ( .A(x[1672]), .B(y[1672]), .Z(n3528) );
  XOR U4735 ( .A(x[1674]), .B(y[1674]), .Z(n3527) );
  XOR U4736 ( .A(n3528), .B(n3527), .Z(n3529) );
  XOR U4737 ( .A(n3530), .B(n3529), .Z(n5277) );
  XOR U4738 ( .A(x[1828]), .B(y[1828]), .Z(n712) );
  XOR U4739 ( .A(x[590]), .B(y[590]), .Z(n710) );
  XOR U4740 ( .A(x[1830]), .B(y[1830]), .Z(n709) );
  XOR U4741 ( .A(n710), .B(n709), .Z(n711) );
  XOR U4742 ( .A(n712), .B(n711), .Z(n5275) );
  XOR U4743 ( .A(x[1666]), .B(y[1666]), .Z(n3638) );
  XOR U4744 ( .A(x[734]), .B(y[734]), .Z(n3636) );
  XOR U4745 ( .A(x[1668]), .B(y[1668]), .Z(n3635) );
  XOR U4746 ( .A(n3636), .B(n3635), .Z(n3637) );
  XNOR U4747 ( .A(n3638), .B(n3637), .Z(n5274) );
  XNOR U4748 ( .A(n5275), .B(n5274), .Z(n5276) );
  XNOR U4749 ( .A(n5277), .B(n5276), .Z(n5954) );
  XNOR U4750 ( .A(n5955), .B(n5954), .Z(n3909) );
  XOR U4751 ( .A(x[1810]), .B(y[1810]), .Z(n5571) );
  XOR U4752 ( .A(x[854]), .B(y[854]), .Z(n5569) );
  XOR U4753 ( .A(x[1812]), .B(y[1812]), .Z(n5568) );
  XOR U4754 ( .A(n5569), .B(n5568), .Z(n5570) );
  XOR U4755 ( .A(n5571), .B(n5570), .Z(n5487) );
  XOR U4756 ( .A(x[1742]), .B(y[1742]), .Z(n5685) );
  XOR U4757 ( .A(x[1744]), .B(y[1744]), .Z(n5683) );
  XOR U4758 ( .A(x[1746]), .B(y[1746]), .Z(n5682) );
  XOR U4759 ( .A(n5683), .B(n5682), .Z(n5684) );
  XOR U4760 ( .A(n5685), .B(n5684), .Z(n5485) );
  XOR U4761 ( .A(x[1814]), .B(y[1814]), .Z(n5565) );
  XOR U4762 ( .A(x[1816]), .B(y[1816]), .Z(n5563) );
  XOR U4763 ( .A(x[1818]), .B(y[1818]), .Z(n5562) );
  XOR U4764 ( .A(n5563), .B(n5562), .Z(n5564) );
  XNOR U4765 ( .A(n5565), .B(n5564), .Z(n5484) );
  XNOR U4766 ( .A(n5485), .B(n5484), .Z(n5486) );
  XNOR U4767 ( .A(n5487), .B(n5486), .Z(n5946) );
  XOR U4768 ( .A(x[218]), .B(y[218]), .Z(n2288) );
  XOR U4769 ( .A(x[220]), .B(y[220]), .Z(n2285) );
  XNOR U4770 ( .A(x[1881]), .B(y[1881]), .Z(n2286) );
  XNOR U4771 ( .A(n2285), .B(n2286), .Z(n2287) );
  XOR U4772 ( .A(n2288), .B(n2287), .Z(n5595) );
  XOR U4773 ( .A(x[1206]), .B(y[1206]), .Z(n1976) );
  XOR U4774 ( .A(x[521]), .B(y[521]), .Z(n1973) );
  XNOR U4775 ( .A(x[1208]), .B(y[1208]), .Z(n1974) );
  XNOR U4776 ( .A(n1973), .B(n1974), .Z(n1975) );
  XOR U4777 ( .A(n1976), .B(n1975), .Z(n5593) );
  XOR U4778 ( .A(x[206]), .B(y[206]), .Z(n1498) );
  XOR U4779 ( .A(x[208]), .B(y[208]), .Z(n1495) );
  XNOR U4780 ( .A(x[751]), .B(y[751]), .Z(n1496) );
  XNOR U4781 ( .A(n1495), .B(n1496), .Z(n1497) );
  XNOR U4782 ( .A(n1498), .B(n1497), .Z(n5592) );
  XNOR U4783 ( .A(n5593), .B(n5592), .Z(n5594) );
  XOR U4784 ( .A(n5595), .B(n5594), .Z(n5947) );
  XNOR U4785 ( .A(n5946), .B(n5947), .Z(n5949) );
  XOR U4786 ( .A(x[1688]), .B(y[1688]), .Z(n5457) );
  XOR U4787 ( .A(x[1690]), .B(y[1690]), .Z(n5454) );
  XNOR U4788 ( .A(x[1692]), .B(y[1692]), .Z(n5455) );
  XNOR U4789 ( .A(n5454), .B(n5455), .Z(n5456) );
  XOR U4790 ( .A(n5457), .B(n5456), .Z(n5157) );
  XOR U4791 ( .A(x[1820]), .B(y[1820]), .Z(n5391) );
  XOR U4792 ( .A(x[582]), .B(y[582]), .Z(n5389) );
  XOR U4793 ( .A(x[1822]), .B(y[1822]), .Z(n5388) );
  XOR U4794 ( .A(n5389), .B(n5388), .Z(n5390) );
  XOR U4795 ( .A(n5391), .B(n5390), .Z(n5155) );
  XOR U4796 ( .A(x[1684]), .B(y[1684]), .Z(n4683) );
  XOR U4797 ( .A(x[458]), .B(y[458]), .Z(n4680) );
  XNOR U4798 ( .A(x[1686]), .B(y[1686]), .Z(n4681) );
  XNOR U4799 ( .A(n4680), .B(n4681), .Z(n4682) );
  XNOR U4800 ( .A(n4683), .B(n4682), .Z(n5154) );
  XNOR U4801 ( .A(n5155), .B(n5154), .Z(n5156) );
  XNOR U4802 ( .A(n5157), .B(n5156), .Z(n5948) );
  XNOR U4803 ( .A(n5949), .B(n5948), .Z(n3907) );
  XOR U4804 ( .A(x[1662]), .B(y[1662]), .Z(n3596) );
  XOR U4805 ( .A(x[438]), .B(y[438]), .Z(n3593) );
  XNOR U4806 ( .A(x[1664]), .B(y[1664]), .Z(n3594) );
  XNOR U4807 ( .A(n3593), .B(n3594), .Z(n3595) );
  XOR U4808 ( .A(n3596), .B(n3595), .Z(n5271) );
  XOR U4809 ( .A(x[1832]), .B(y[1832]), .Z(n2126) );
  XOR U4810 ( .A(x[1834]), .B(y[1834]), .Z(n2123) );
  XNOR U4811 ( .A(x[1836]), .B(y[1836]), .Z(n2124) );
  XNOR U4812 ( .A(n2123), .B(n2124), .Z(n2125) );
  XOR U4813 ( .A(n2126), .B(n2125), .Z(n5269) );
  XOR U4814 ( .A(x[1658]), .B(y[1658]), .Z(n3590) );
  XOR U4815 ( .A(x[434]), .B(y[434]), .Z(n3587) );
  XNOR U4816 ( .A(x[1660]), .B(y[1660]), .Z(n3588) );
  XNOR U4817 ( .A(n3587), .B(n3588), .Z(n3589) );
  XNOR U4818 ( .A(n3590), .B(n3589), .Z(n5268) );
  XNOR U4819 ( .A(n5269), .B(n5268), .Z(n5270) );
  XNOR U4820 ( .A(n5271), .B(n5270), .Z(n5862) );
  XOR U4821 ( .A(x[184]), .B(y[184]), .Z(n1126) );
  XOR U4822 ( .A(x[188]), .B(y[188]), .Z(n1123) );
  XNOR U4823 ( .A(x[1879]), .B(y[1879]), .Z(n1124) );
  XNOR U4824 ( .A(n1123), .B(n1124), .Z(n1125) );
  XOR U4825 ( .A(n1126), .B(n1125), .Z(n1696) );
  XOR U4826 ( .A(x[1198]), .B(y[1198]), .Z(n2186) );
  XOR U4827 ( .A(x[527]), .B(y[527]), .Z(n2183) );
  XNOR U4828 ( .A(x[1200]), .B(y[1200]), .Z(n2184) );
  XNOR U4829 ( .A(n2183), .B(n2184), .Z(n2185) );
  XOR U4830 ( .A(n2186), .B(n2185), .Z(n1694) );
  XOR U4831 ( .A(x[180]), .B(y[180]), .Z(n1210) );
  XOR U4832 ( .A(x[182]), .B(y[182]), .Z(n1207) );
  XNOR U4833 ( .A(x[765]), .B(y[765]), .Z(n1208) );
  XNOR U4834 ( .A(n1207), .B(n1208), .Z(n1209) );
  XNOR U4835 ( .A(n1210), .B(n1209), .Z(n1693) );
  XNOR U4836 ( .A(n1694), .B(n1693), .Z(n1695) );
  XOR U4837 ( .A(n1696), .B(n1695), .Z(n5863) );
  XNOR U4838 ( .A(n5862), .B(n5863), .Z(n5865) );
  XOR U4839 ( .A(x[1654]), .B(y[1654]), .Z(n3650) );
  XOR U4840 ( .A(x[430]), .B(y[430]), .Z(n3647) );
  XNOR U4841 ( .A(x[1656]), .B(y[1656]), .Z(n3648) );
  XNOR U4842 ( .A(n3647), .B(n3648), .Z(n3649) );
  XOR U4843 ( .A(n3650), .B(n3649), .Z(n6039) );
  XOR U4844 ( .A(x[1838]), .B(y[1838]), .Z(n2066) );
  XOR U4845 ( .A(x[1840]), .B(y[1840]), .Z(n2063) );
  XNOR U4846 ( .A(x[1842]), .B(y[1842]), .Z(n2064) );
  XNOR U4847 ( .A(n2063), .B(n2064), .Z(n2065) );
  XOR U4848 ( .A(n2066), .B(n2065), .Z(n6037) );
  XOR U4849 ( .A(x[1650]), .B(y[1650]), .Z(n3644) );
  XOR U4850 ( .A(x[720]), .B(y[720]), .Z(n3641) );
  XNOR U4851 ( .A(x[1652]), .B(y[1652]), .Z(n3642) );
  XNOR U4852 ( .A(n3641), .B(n3642), .Z(n3643) );
  XNOR U4853 ( .A(n3644), .B(n3643), .Z(n6036) );
  XNOR U4854 ( .A(n6037), .B(n6036), .Z(n6038) );
  XNOR U4855 ( .A(n6039), .B(n6038), .Z(n5864) );
  XNOR U4856 ( .A(n5865), .B(n5864), .Z(n3906) );
  XOR U4857 ( .A(n3907), .B(n3906), .Z(n3908) );
  XNOR U4858 ( .A(n3909), .B(n3908), .Z(n3895) );
  XOR U4859 ( .A(x[1430]), .B(y[1430]), .Z(n874) );
  XOR U4860 ( .A(x[490]), .B(y[490]), .Z(n871) );
  XNOR U4861 ( .A(x[1432]), .B(y[1432]), .Z(n872) );
  XNOR U4862 ( .A(n871), .B(n872), .Z(n873) );
  XOR U4863 ( .A(n874), .B(n873), .Z(n4659) );
  XOR U4864 ( .A(x[1424]), .B(y[1424]), .Z(n1216) );
  XOR U4865 ( .A(x[1426]), .B(y[1426]), .Z(n1213) );
  XNOR U4866 ( .A(x[1428]), .B(y[1428]), .Z(n1214) );
  XNOR U4867 ( .A(n1213), .B(n1214), .Z(n1215) );
  XOR U4868 ( .A(n1216), .B(n1215), .Z(n4657) );
  XOR U4869 ( .A(x[1420]), .B(y[1420]), .Z(n1132) );
  XOR U4870 ( .A(x[216]), .B(y[216]), .Z(n1129) );
  XNOR U4871 ( .A(x[1422]), .B(y[1422]), .Z(n1130) );
  XNOR U4872 ( .A(n1129), .B(n1130), .Z(n1131) );
  XNOR U4873 ( .A(n1132), .B(n1131), .Z(n4656) );
  XNOR U4874 ( .A(n4657), .B(n4656), .Z(n4658) );
  XNOR U4875 ( .A(n4659), .B(n4658), .Z(n1723) );
  XOR U4876 ( .A(x[1416]), .B(y[1416]), .Z(n1222) );
  XOR U4877 ( .A(x[210]), .B(y[210]), .Z(n1219) );
  XNOR U4878 ( .A(x[1418]), .B(y[1418]), .Z(n1220) );
  XNOR U4879 ( .A(n1219), .B(n1220), .Z(n1221) );
  XOR U4880 ( .A(n1222), .B(n1221), .Z(n5943) );
  XOR U4881 ( .A(x[1412]), .B(y[1412]), .Z(n1252) );
  XOR U4882 ( .A(x[472]), .B(y[472]), .Z(n1249) );
  XNOR U4883 ( .A(x[1414]), .B(y[1414]), .Z(n1250) );
  XNOR U4884 ( .A(n1249), .B(n1250), .Z(n1251) );
  XOR U4885 ( .A(n1252), .B(n1251), .Z(n5941) );
  XOR U4886 ( .A(x[1406]), .B(y[1406]), .Z(n856) );
  XOR U4887 ( .A(x[1408]), .B(y[1408]), .Z(n853) );
  XNOR U4888 ( .A(x[1410]), .B(y[1410]), .Z(n854) );
  XNOR U4889 ( .A(n853), .B(n854), .Z(n855) );
  XNOR U4890 ( .A(n856), .B(n855), .Z(n5940) );
  XNOR U4891 ( .A(n5941), .B(n5940), .Z(n5942) );
  XOR U4892 ( .A(n5943), .B(n5942), .Z(n1724) );
  XNOR U4893 ( .A(n1723), .B(n1724), .Z(n1726) );
  XOR U4894 ( .A(x[1396]), .B(y[1396]), .Z(n2336) );
  XOR U4895 ( .A(x[194]), .B(y[194]), .Z(n2333) );
  XNOR U4896 ( .A(x[1398]), .B(y[1398]), .Z(n2334) );
  XNOR U4897 ( .A(n2333), .B(n2334), .Z(n2335) );
  XOR U4898 ( .A(n2336), .B(n2335), .Z(n3308) );
  XOR U4899 ( .A(x[1388]), .B(y[1388]), .Z(n5193) );
  XOR U4900 ( .A(x[186]), .B(y[186]), .Z(n5190) );
  XNOR U4901 ( .A(x[1390]), .B(y[1390]), .Z(n5191) );
  XNOR U4902 ( .A(n5190), .B(n5191), .Z(n5192) );
  XOR U4903 ( .A(n5193), .B(n5192), .Z(n3306) );
  XOR U4904 ( .A(x[1378]), .B(y[1378]), .Z(n5427) );
  XOR U4905 ( .A(x[440]), .B(y[440]), .Z(n5424) );
  XNOR U4906 ( .A(x[1380]), .B(y[1380]), .Z(n5425) );
  XNOR U4907 ( .A(n5424), .B(n5425), .Z(n5426) );
  XNOR U4908 ( .A(n5427), .B(n5426), .Z(n3305) );
  XNOR U4909 ( .A(n3306), .B(n3305), .Z(n3307) );
  XNOR U4910 ( .A(n3308), .B(n3307), .Z(n1725) );
  XOR U4911 ( .A(n1726), .B(n1725), .Z(n4161) );
  XOR U4912 ( .A(x[1370]), .B(y[1370]), .Z(n5397) );
  XOR U4913 ( .A(x[23]), .B(y[23]), .Z(n5394) );
  XNOR U4914 ( .A(x[1372]), .B(y[1372]), .Z(n5395) );
  XNOR U4915 ( .A(n5394), .B(n5395), .Z(n5396) );
  XOR U4916 ( .A(n5397), .B(n5396), .Z(n5859) );
  XOR U4917 ( .A(x[1362]), .B(y[1362]), .Z(n5379) );
  XOR U4918 ( .A(x[29]), .B(y[29]), .Z(n5376) );
  XNOR U4919 ( .A(x[1364]), .B(y[1364]), .Z(n5377) );
  XNOR U4920 ( .A(n5376), .B(n5377), .Z(n5378) );
  XOR U4921 ( .A(n5379), .B(n5378), .Z(n5857) );
  XOR U4922 ( .A(x[1354]), .B(y[1354]), .Z(n5541) );
  XOR U4923 ( .A(x[1356]), .B(y[1356]), .Z(n5538) );
  XNOR U4924 ( .A(x[1999]), .B(y[1999]), .Z(n5539) );
  XNOR U4925 ( .A(n5538), .B(n5539), .Z(n5540) );
  XNOR U4926 ( .A(n5541), .B(n5540), .Z(n5856) );
  XNOR U4927 ( .A(n5857), .B(n5856), .Z(n5858) );
  XNOR U4928 ( .A(n5859), .B(n5858), .Z(n1567) );
  XOR U4929 ( .A(x[1346]), .B(y[1346]), .Z(n6057) );
  XOR U4930 ( .A(x[1348]), .B(y[1348]), .Z(n6054) );
  XNOR U4931 ( .A(x[1997]), .B(y[1997]), .Z(n6055) );
  XNOR U4932 ( .A(n6054), .B(n6055), .Z(n6056) );
  XOR U4933 ( .A(n6057), .B(n6056), .Z(n3410) );
  XOR U4934 ( .A(x[1338]), .B(y[1338]), .Z(n6051) );
  XOR U4935 ( .A(x[45]), .B(y[45]), .Z(n6048) );
  XNOR U4936 ( .A(x[1340]), .B(y[1340]), .Z(n6049) );
  XNOR U4937 ( .A(n6048), .B(n6049), .Z(n6050) );
  XOR U4938 ( .A(n6051), .B(n6050), .Z(n3408) );
  XOR U4939 ( .A(x[1330]), .B(y[1330]), .Z(n5139) );
  XOR U4940 ( .A(x[51]), .B(y[51]), .Z(n5136) );
  XNOR U4941 ( .A(x[1332]), .B(y[1332]), .Z(n5137) );
  XNOR U4942 ( .A(n5136), .B(n5137), .Z(n5138) );
  XNOR U4943 ( .A(n5139), .B(n5138), .Z(n3407) );
  XNOR U4944 ( .A(n3408), .B(n3407), .Z(n3409) );
  XOR U4945 ( .A(n3410), .B(n3409), .Z(n1568) );
  XNOR U4946 ( .A(n1567), .B(n1568), .Z(n1570) );
  XOR U4947 ( .A(x[1322]), .B(y[1322]), .Z(n5133) );
  XOR U4948 ( .A(x[1324]), .B(y[1324]), .Z(n5130) );
  XNOR U4949 ( .A(x[1995]), .B(y[1995]), .Z(n5131) );
  XNOR U4950 ( .A(n5130), .B(n5131), .Z(n5132) );
  XOR U4951 ( .A(n5133), .B(n5132), .Z(n4635) );
  XOR U4952 ( .A(x[1314]), .B(y[1314]), .Z(n5127) );
  XOR U4953 ( .A(x[1316]), .B(y[1316]), .Z(n5124) );
  XNOR U4954 ( .A(x[1993]), .B(y[1993]), .Z(n5125) );
  XNOR U4955 ( .A(n5124), .B(n5125), .Z(n5126) );
  XOR U4956 ( .A(n5127), .B(n5126), .Z(n4633) );
  XOR U4957 ( .A(x[1306]), .B(y[1306]), .Z(n4869) );
  XOR U4958 ( .A(x[67]), .B(y[67]), .Z(n4866) );
  XNOR U4959 ( .A(x[1308]), .B(y[1308]), .Z(n4867) );
  XNOR U4960 ( .A(n4866), .B(n4867), .Z(n4868) );
  XNOR U4961 ( .A(n4869), .B(n4868), .Z(n4632) );
  XNOR U4962 ( .A(n4633), .B(n4632), .Z(n4634) );
  XNOR U4963 ( .A(n4635), .B(n4634), .Z(n1569) );
  XNOR U4964 ( .A(n1570), .B(n1569), .Z(n4159) );
  XOR U4965 ( .A(x[1730]), .B(y[1730]), .Z(n5253) );
  XOR U4966 ( .A(x[500]), .B(y[500]), .Z(n5250) );
  XNOR U4967 ( .A(x[1732]), .B(y[1732]), .Z(n5251) );
  XNOR U4968 ( .A(n5250), .B(n5251), .Z(n5252) );
  XOR U4969 ( .A(n5253), .B(n5252), .Z(n2870) );
  XOR U4970 ( .A(x[1752]), .B(y[1752]), .Z(n5091) );
  XOR U4971 ( .A(x[520]), .B(y[520]), .Z(n5088) );
  XNOR U4972 ( .A(x[1754]), .B(y[1754]), .Z(n5089) );
  XNOR U4973 ( .A(n5088), .B(n5089), .Z(n5090) );
  XOR U4974 ( .A(n5091), .B(n5090), .Z(n2868) );
  XOR U4975 ( .A(x[1760]), .B(y[1760]), .Z(n5175) );
  XOR U4976 ( .A(x[1762]), .B(y[1762]), .Z(n5172) );
  XNOR U4977 ( .A(x[1764]), .B(y[1764]), .Z(n5173) );
  XNOR U4978 ( .A(n5172), .B(n5173), .Z(n5174) );
  XNOR U4979 ( .A(n5175), .B(n5174), .Z(n2867) );
  XNOR U4980 ( .A(n2868), .B(n2867), .Z(n2869) );
  XNOR U4981 ( .A(n2870), .B(n2869), .Z(n5514) );
  XOR U4982 ( .A(x[280]), .B(y[280]), .Z(n2804) );
  XOR U4983 ( .A(x[284]), .B(y[284]), .Z(n2801) );
  XNOR U4984 ( .A(x[703]), .B(y[703]), .Z(n2802) );
  XNOR U4985 ( .A(n2801), .B(n2802), .Z(n2803) );
  XOR U4986 ( .A(n2804), .B(n2803), .Z(n1576) );
  XOR U4987 ( .A(x[1954]), .B(y[1954]), .Z(n3422) );
  XOR U4988 ( .A(x[966]), .B(y[966]), .Z(n3420) );
  XOR U4989 ( .A(x[1956]), .B(y[1956]), .Z(n3419) );
  XOR U4990 ( .A(n3420), .B(n3419), .Z(n3421) );
  XOR U4991 ( .A(n3422), .B(n3421), .Z(n1574) );
  XOR U4992 ( .A(x[274]), .B(y[274]), .Z(n2384) );
  XOR U4993 ( .A(x[278]), .B(y[278]), .Z(n2381) );
  XNOR U4994 ( .A(x[987]), .B(y[987]), .Z(n2382) );
  XNOR U4995 ( .A(n2381), .B(n2382), .Z(n2383) );
  XNOR U4996 ( .A(n2384), .B(n2383), .Z(n1573) );
  XNOR U4997 ( .A(n1574), .B(n1573), .Z(n1575) );
  XOR U4998 ( .A(n1576), .B(n1575), .Z(n5515) );
  XNOR U4999 ( .A(n5514), .B(n5515), .Z(n5517) );
  XOR U5000 ( .A(x[1766]), .B(y[1766]), .Z(n5415) );
  XOR U5001 ( .A(x[1768]), .B(y[1768]), .Z(n5413) );
  XOR U5002 ( .A(x[1770]), .B(y[1770]), .Z(n5412) );
  XOR U5003 ( .A(n5413), .B(n5412), .Z(n5414) );
  XOR U5004 ( .A(n5415), .B(n5414), .Z(n5577) );
  XOR U5005 ( .A(x[1738]), .B(y[1738]), .Z(n5691) );
  XOR U5006 ( .A(x[798]), .B(y[798]), .Z(n5689) );
  XOR U5007 ( .A(x[1740]), .B(y[1740]), .Z(n5688) );
  XOR U5008 ( .A(n5689), .B(n5688), .Z(n5690) );
  XOR U5009 ( .A(n5691), .B(n5690), .Z(n5575) );
  XOR U5010 ( .A(x[1772]), .B(y[1772]), .Z(n5421) );
  XOR U5011 ( .A(x[824]), .B(y[824]), .Z(n5419) );
  XOR U5012 ( .A(x[1774]), .B(y[1774]), .Z(n5418) );
  XOR U5013 ( .A(n5419), .B(n5418), .Z(n5420) );
  XNOR U5014 ( .A(n5421), .B(n5420), .Z(n5574) );
  XNOR U5015 ( .A(n5575), .B(n5574), .Z(n5576) );
  XNOR U5016 ( .A(n5577), .B(n5576), .Z(n5516) );
  XNOR U5017 ( .A(n5517), .B(n5516), .Z(n4158) );
  XOR U5018 ( .A(n4159), .B(n4158), .Z(n4160) );
  XOR U5019 ( .A(n4161), .B(n4160), .Z(n3894) );
  XOR U5020 ( .A(n3895), .B(n3894), .Z(n3897) );
  XOR U5021 ( .A(x[1298]), .B(y[1298]), .Z(n4743) );
  XOR U5022 ( .A(x[73]), .B(y[73]), .Z(n4740) );
  XNOR U5023 ( .A(x[1300]), .B(y[1300]), .Z(n4741) );
  XNOR U5024 ( .A(n4740), .B(n4741), .Z(n4742) );
  XOR U5025 ( .A(n4743), .B(n4742), .Z(n3993) );
  XOR U5026 ( .A(x[1290]), .B(y[1290]), .Z(n4737) );
  XOR U5027 ( .A(x[1292]), .B(y[1292]), .Z(n4734) );
  XNOR U5028 ( .A(x[1991]), .B(y[1991]), .Z(n4735) );
  XNOR U5029 ( .A(n4734), .B(n4735), .Z(n4736) );
  XOR U5030 ( .A(n4737), .B(n4736), .Z(n3991) );
  XOR U5031 ( .A(x[1282]), .B(y[1282]), .Z(n4713) );
  XOR U5032 ( .A(x[1284]), .B(y[1284]), .Z(n4710) );
  XNOR U5033 ( .A(x[1989]), .B(y[1989]), .Z(n4711) );
  XNOR U5034 ( .A(n4710), .B(n4711), .Z(n4712) );
  XNOR U5035 ( .A(n4713), .B(n4712), .Z(n3990) );
  XNOR U5036 ( .A(n3991), .B(n3990), .Z(n3992) );
  XNOR U5037 ( .A(n3993), .B(n3992), .Z(n1333) );
  XOR U5038 ( .A(x[1274]), .B(y[1274]), .Z(n4977) );
  XOR U5039 ( .A(x[89]), .B(y[89]), .Z(n4974) );
  XNOR U5040 ( .A(x[1276]), .B(y[1276]), .Z(n4975) );
  XNOR U5041 ( .A(n4974), .B(n4975), .Z(n4976) );
  XOR U5042 ( .A(n4977), .B(n4976), .Z(n4803) );
  XOR U5043 ( .A(x[1266]), .B(y[1266]), .Z(n4965) );
  XOR U5044 ( .A(x[95]), .B(y[95]), .Z(n4962) );
  XNOR U5045 ( .A(x[1268]), .B(y[1268]), .Z(n4963) );
  XNOR U5046 ( .A(n4962), .B(n4963), .Z(n4964) );
  XOR U5047 ( .A(n4965), .B(n4964), .Z(n4801) );
  XOR U5048 ( .A(x[1258]), .B(y[1258]), .Z(n5103) );
  XOR U5049 ( .A(x[1260]), .B(y[1260]), .Z(n5100) );
  XNOR U5050 ( .A(x[1987]), .B(y[1987]), .Z(n5101) );
  XNOR U5051 ( .A(n5100), .B(n5101), .Z(n5102) );
  XNOR U5052 ( .A(n5103), .B(n5102), .Z(n4800) );
  XNOR U5053 ( .A(n4801), .B(n4800), .Z(n4802) );
  XOR U5054 ( .A(n4803), .B(n4802), .Z(n1334) );
  XNOR U5055 ( .A(n1333), .B(n1334), .Z(n1335) );
  XOR U5056 ( .A(x[1250]), .B(y[1250]), .Z(n5055) );
  XOR U5057 ( .A(x[1252]), .B(y[1252]), .Z(n5052) );
  XNOR U5058 ( .A(x[1985]), .B(y[1985]), .Z(n5053) );
  XNOR U5059 ( .A(n5052), .B(n5053), .Z(n5054) );
  XOR U5060 ( .A(n5055), .B(n5054), .Z(n2960) );
  XOR U5061 ( .A(x[1242]), .B(y[1242]), .Z(n694) );
  XOR U5062 ( .A(x[111]), .B(y[111]), .Z(n691) );
  XNOR U5063 ( .A(x[1244]), .B(y[1244]), .Z(n692) );
  XNOR U5064 ( .A(n691), .B(n692), .Z(n693) );
  XOR U5065 ( .A(n694), .B(n693), .Z(n2958) );
  XOR U5066 ( .A(x[1234]), .B(y[1234]), .Z(n898) );
  XOR U5067 ( .A(x[117]), .B(y[117]), .Z(n895) );
  XNOR U5068 ( .A(x[1236]), .B(y[1236]), .Z(n896) );
  XNOR U5069 ( .A(n895), .B(n896), .Z(n897) );
  XNOR U5070 ( .A(n898), .B(n897), .Z(n2957) );
  XNOR U5071 ( .A(n2958), .B(n2957), .Z(n2959) );
  XOR U5072 ( .A(n2960), .B(n2959), .Z(n1336) );
  XNOR U5073 ( .A(n1335), .B(n1336), .Z(n4167) );
  XOR U5074 ( .A(x[1711]), .B(y[1711]), .Z(n2972) );
  XOR U5075 ( .A(x[1683]), .B(y[1683]), .Z(n2969) );
  XNOR U5076 ( .A(x[1713]), .B(y[1713]), .Z(n2970) );
  XNOR U5077 ( .A(n2969), .B(n2970), .Z(n2971) );
  XOR U5078 ( .A(n2972), .B(n2971), .Z(n5210) );
  XOR U5079 ( .A(x[651]), .B(y[651]), .Z(n594) );
  XOR U5080 ( .A(x[645]), .B(y[645]), .Z(n591) );
  XNOR U5081 ( .A(x[1111]), .B(y[1111]), .Z(n592) );
  XNOR U5082 ( .A(n591), .B(n592), .Z(n593) );
  XOR U5083 ( .A(n594), .B(n593), .Z(n5209) );
  XOR U5084 ( .A(x[1707]), .B(y[1707]), .Z(n588) );
  XOR U5085 ( .A(x[1689]), .B(y[1689]), .Z(n585) );
  XNOR U5086 ( .A(x[1709]), .B(y[1709]), .Z(n586) );
  XNOR U5087 ( .A(n585), .B(n586), .Z(n587) );
  XNOR U5088 ( .A(n588), .B(n587), .Z(n5208) );
  XOR U5089 ( .A(n5209), .B(n5208), .Z(n5211) );
  XOR U5090 ( .A(n5210), .B(n5211), .Z(n5240) );
  XOR U5091 ( .A(x[270]), .B(y[270]), .Z(n3188) );
  XOR U5092 ( .A(x[272]), .B(y[272]), .Z(n3185) );
  XNOR U5093 ( .A(x[1887]), .B(y[1887]), .Z(n3186) );
  XNOR U5094 ( .A(n3185), .B(n3186), .Z(n3187) );
  XOR U5095 ( .A(n3188), .B(n3187), .Z(n1629) );
  XOR U5096 ( .A(x[1222]), .B(y[1222]), .Z(n2096) );
  XOR U5097 ( .A(x[123]), .B(y[123]), .Z(n2093) );
  XNOR U5098 ( .A(x[1224]), .B(y[1224]), .Z(n2094) );
  XNOR U5099 ( .A(n2093), .B(n2094), .Z(n2095) );
  XOR U5100 ( .A(n2096), .B(n2095), .Z(n1628) );
  XOR U5101 ( .A(x[266]), .B(y[266]), .Z(n2318) );
  XOR U5102 ( .A(x[268]), .B(y[268]), .Z(n2315) );
  XNOR U5103 ( .A(x[711]), .B(y[711]), .Z(n2316) );
  XNOR U5104 ( .A(n2315), .B(n2316), .Z(n2317) );
  XNOR U5105 ( .A(n2318), .B(n2317), .Z(n1627) );
  XOR U5106 ( .A(n1628), .B(n1627), .Z(n1630) );
  XOR U5107 ( .A(n1629), .B(n1630), .Z(n5239) );
  XOR U5108 ( .A(x[1756]), .B(y[1756]), .Z(n5198) );
  XOR U5109 ( .A(x[524]), .B(y[524]), .Z(n5196) );
  XNOR U5110 ( .A(x[1758]), .B(y[1758]), .Z(n5197) );
  XOR U5111 ( .A(n5196), .B(n5197), .Z(n5199) );
  XNOR U5112 ( .A(n5198), .B(n5199), .Z(n5238) );
  XOR U5113 ( .A(n5239), .B(n5238), .Z(n5241) );
  XNOR U5114 ( .A(n5240), .B(n5241), .Z(n4165) );
  XOR U5115 ( .A(x[1226]), .B(y[1226]), .Z(n2606) );
  XOR U5116 ( .A(x[1228]), .B(y[1228]), .Z(n2603) );
  XNOR U5117 ( .A(x[1983]), .B(y[1983]), .Z(n2604) );
  XNOR U5118 ( .A(n2603), .B(n2604), .Z(n2605) );
  XOR U5119 ( .A(n2606), .B(n2605), .Z(n3386) );
  XOR U5120 ( .A(x[1218]), .B(y[1218]), .Z(n5037) );
  XOR U5121 ( .A(x[1220]), .B(y[1220]), .Z(n5034) );
  XNOR U5122 ( .A(x[1981]), .B(y[1981]), .Z(n5035) );
  XNOR U5123 ( .A(n5034), .B(n5035), .Z(n5036) );
  XOR U5124 ( .A(n5037), .B(n5036), .Z(n3384) );
  XOR U5125 ( .A(x[1210]), .B(y[1210]), .Z(n5043) );
  XOR U5126 ( .A(x[133]), .B(y[133]), .Z(n5040) );
  XNOR U5127 ( .A(x[1212]), .B(y[1212]), .Z(n5041) );
  XNOR U5128 ( .A(n5040), .B(n5041), .Z(n5042) );
  XNOR U5129 ( .A(n5043), .B(n5042), .Z(n3383) );
  XNOR U5130 ( .A(n3384), .B(n3383), .Z(n3385) );
  XNOR U5131 ( .A(n3386), .B(n3385), .Z(n1531) );
  XOR U5132 ( .A(x[1202]), .B(y[1202]), .Z(n5745) );
  XOR U5133 ( .A(x[139]), .B(y[139]), .Z(n5742) );
  XNOR U5134 ( .A(x[1204]), .B(y[1204]), .Z(n5743) );
  XNOR U5135 ( .A(n5742), .B(n5743), .Z(n5744) );
  XOR U5136 ( .A(n5745), .B(n5744), .Z(n2786) );
  XOR U5137 ( .A(x[1194]), .B(y[1194]), .Z(n5733) );
  XOR U5138 ( .A(x[1196]), .B(y[1196]), .Z(n5730) );
  XNOR U5139 ( .A(x[1979]), .B(y[1979]), .Z(n5731) );
  XNOR U5140 ( .A(n5730), .B(n5731), .Z(n5732) );
  XOR U5141 ( .A(n5733), .B(n5732), .Z(n2784) );
  XOR U5142 ( .A(x[1186]), .B(y[1186]), .Z(n5739) );
  XOR U5143 ( .A(x[1188]), .B(y[1188]), .Z(n5736) );
  XNOR U5144 ( .A(x[1977]), .B(y[1977]), .Z(n5737) );
  XNOR U5145 ( .A(n5736), .B(n5737), .Z(n5738) );
  XNOR U5146 ( .A(n5739), .B(n5738), .Z(n2783) );
  XNOR U5147 ( .A(n2784), .B(n2783), .Z(n2785) );
  XOR U5148 ( .A(n2786), .B(n2785), .Z(n1532) );
  XNOR U5149 ( .A(n1531), .B(n1532), .Z(n1533) );
  XOR U5150 ( .A(x[1178]), .B(y[1178]), .Z(n5907) );
  XOR U5151 ( .A(x[155]), .B(y[155]), .Z(n5904) );
  XNOR U5152 ( .A(x[1180]), .B(y[1180]), .Z(n5905) );
  XNOR U5153 ( .A(n5904), .B(n5905), .Z(n5906) );
  XOR U5154 ( .A(n5907), .B(n5906), .Z(n2798) );
  XOR U5155 ( .A(x[1170]), .B(y[1170]), .Z(n5895) );
  XOR U5156 ( .A(x[161]), .B(y[161]), .Z(n5892) );
  XNOR U5157 ( .A(x[1172]), .B(y[1172]), .Z(n5893) );
  XNOR U5158 ( .A(n5892), .B(n5893), .Z(n5894) );
  XOR U5159 ( .A(n5895), .B(n5894), .Z(n2796) );
  XOR U5160 ( .A(x[1162]), .B(y[1162]), .Z(n5901) );
  XOR U5161 ( .A(x[1164]), .B(y[1164]), .Z(n5898) );
  XNOR U5162 ( .A(x[1975]), .B(y[1975]), .Z(n5899) );
  XNOR U5163 ( .A(n5898), .B(n5899), .Z(n5900) );
  XNOR U5164 ( .A(n5901), .B(n5900), .Z(n2795) );
  XNOR U5165 ( .A(n2796), .B(n2795), .Z(n2797) );
  XOR U5166 ( .A(n2798), .B(n2797), .Z(n1534) );
  XNOR U5167 ( .A(n1533), .B(n1534), .Z(n4164) );
  XOR U5168 ( .A(n4165), .B(n4164), .Z(n4166) );
  XOR U5169 ( .A(n4167), .B(n4166), .Z(n3896) );
  XOR U5170 ( .A(n3897), .B(n3896), .Z(n3801) );
  XOR U5171 ( .A(x[1510]), .B(y[1510]), .Z(n5721) );
  XOR U5172 ( .A(x[298]), .B(y[298]), .Z(n5718) );
  XNOR U5173 ( .A(x[1512]), .B(y[1512]), .Z(n5719) );
  XNOR U5174 ( .A(n5718), .B(n5719), .Z(n5720) );
  XOR U5175 ( .A(n5721), .B(n5720), .Z(n5073) );
  XOR U5176 ( .A(x[1506]), .B(y[1506]), .Z(n2330) );
  XOR U5177 ( .A(x[572]), .B(y[572]), .Z(n2327) );
  XNOR U5178 ( .A(x[1508]), .B(y[1508]), .Z(n2328) );
  XNOR U5179 ( .A(n2327), .B(n2328), .Z(n2329) );
  XOR U5180 ( .A(n2330), .B(n2329), .Z(n5071) );
  XOR U5181 ( .A(x[1502]), .B(y[1502]), .Z(n2294) );
  XOR U5182 ( .A(x[564]), .B(y[564]), .Z(n2291) );
  XNOR U5183 ( .A(x[1504]), .B(y[1504]), .Z(n2292) );
  XNOR U5184 ( .A(n2291), .B(n2292), .Z(n2293) );
  XNOR U5185 ( .A(n2294), .B(n2293), .Z(n5070) );
  XNOR U5186 ( .A(n5071), .B(n5070), .Z(n5072) );
  XNOR U5187 ( .A(n5073), .B(n5072), .Z(n1159) );
  XOR U5188 ( .A(x[1496]), .B(y[1496]), .Z(n2276) );
  XOR U5189 ( .A(x[1498]), .B(y[1498]), .Z(n2273) );
  XNOR U5190 ( .A(x[1500]), .B(y[1500]), .Z(n2274) );
  XNOR U5191 ( .A(n2273), .B(n2274), .Z(n2275) );
  XOR U5192 ( .A(n2276), .B(n2275), .Z(n4893) );
  XOR U5193 ( .A(x[1492]), .B(y[1492]), .Z(n850) );
  XOR U5194 ( .A(x[282]), .B(y[282]), .Z(n847) );
  XNOR U5195 ( .A(x[1494]), .B(y[1494]), .Z(n848) );
  XNOR U5196 ( .A(n847), .B(n848), .Z(n849) );
  XOR U5197 ( .A(n850), .B(n849), .Z(n4891) );
  XOR U5198 ( .A(x[1488]), .B(y[1488]), .Z(n868) );
  XOR U5199 ( .A(x[276]), .B(y[276]), .Z(n865) );
  XNOR U5200 ( .A(x[1490]), .B(y[1490]), .Z(n866) );
  XNOR U5201 ( .A(n865), .B(n866), .Z(n867) );
  XNOR U5202 ( .A(n868), .B(n867), .Z(n4890) );
  XNOR U5203 ( .A(n4891), .B(n4890), .Z(n4892) );
  XOR U5204 ( .A(n4893), .B(n4892), .Z(n1160) );
  XNOR U5205 ( .A(n1159), .B(n1160), .Z(n1162) );
  XOR U5206 ( .A(x[1484]), .B(y[1484]), .Z(n1432) );
  XOR U5207 ( .A(x[548]), .B(y[548]), .Z(n1429) );
  XNOR U5208 ( .A(x[1486]), .B(y[1486]), .Z(n1430) );
  XNOR U5209 ( .A(n1429), .B(n1430), .Z(n1431) );
  XOR U5210 ( .A(n1432), .B(n1431), .Z(n5913) );
  XOR U5211 ( .A(x[1478]), .B(y[1478]), .Z(n1486) );
  XOR U5212 ( .A(x[1480]), .B(y[1480]), .Z(n1483) );
  XNOR U5213 ( .A(x[1482]), .B(y[1482]), .Z(n1484) );
  XNOR U5214 ( .A(n1483), .B(n1484), .Z(n1485) );
  XOR U5215 ( .A(n1486), .B(n1485), .Z(n5911) );
  XOR U5216 ( .A(x[1472]), .B(y[1472]), .Z(n1492) );
  XOR U5217 ( .A(x[1474]), .B(y[1474]), .Z(n1489) );
  XNOR U5218 ( .A(x[1476]), .B(y[1476]), .Z(n1490) );
  XNOR U5219 ( .A(n1489), .B(n1490), .Z(n1491) );
  XNOR U5220 ( .A(n1492), .B(n1491), .Z(n5910) );
  XNOR U5221 ( .A(n5911), .B(n5910), .Z(n5912) );
  XNOR U5222 ( .A(n5913), .B(n5912), .Z(n1161) );
  XNOR U5223 ( .A(n1162), .B(n1161), .Z(n4089) );
  XOR U5224 ( .A(x[1468]), .B(y[1468]), .Z(n1450) );
  XOR U5225 ( .A(x[260]), .B(y[260]), .Z(n1448) );
  XOR U5226 ( .A(x[1470]), .B(y[1470]), .Z(n1447) );
  XOR U5227 ( .A(n1448), .B(n1447), .Z(n1449) );
  XOR U5228 ( .A(n1450), .B(n1449), .Z(n4989) );
  XOR U5229 ( .A(x[1464]), .B(y[1464]), .Z(n1438) );
  XOR U5230 ( .A(x[256]), .B(y[256]), .Z(n1436) );
  XOR U5231 ( .A(x[1466]), .B(y[1466]), .Z(n1435) );
  XOR U5232 ( .A(n1436), .B(n1435), .Z(n1437) );
  XOR U5233 ( .A(n1438), .B(n1437), .Z(n4987) );
  XOR U5234 ( .A(x[1460]), .B(y[1460]), .Z(n1750) );
  XOR U5235 ( .A(x[252]), .B(y[252]), .Z(n1747) );
  XNOR U5236 ( .A(x[1462]), .B(y[1462]), .Z(n1748) );
  XNOR U5237 ( .A(n1747), .B(n1748), .Z(n1749) );
  XNOR U5238 ( .A(n1750), .B(n1749), .Z(n4986) );
  XNOR U5239 ( .A(n4987), .B(n4986), .Z(n4988) );
  XNOR U5240 ( .A(n4989), .B(n4988), .Z(n1231) );
  XOR U5241 ( .A(x[1454]), .B(y[1454]), .Z(n1868) );
  XOR U5242 ( .A(x[1456]), .B(y[1456]), .Z(n1865) );
  XNOR U5243 ( .A(x[1458]), .B(y[1458]), .Z(n1866) );
  XNOR U5244 ( .A(n1865), .B(n1866), .Z(n1867) );
  XOR U5245 ( .A(n1868), .B(n1867), .Z(n5031) );
  XOR U5246 ( .A(x[1450]), .B(y[1450]), .Z(n1588) );
  XOR U5247 ( .A(x[512]), .B(y[512]), .Z(n1585) );
  XNOR U5248 ( .A(x[1452]), .B(y[1452]), .Z(n1586) );
  XNOR U5249 ( .A(n1585), .B(n1586), .Z(n1587) );
  XOR U5250 ( .A(n1588), .B(n1587), .Z(n5029) );
  XOR U5251 ( .A(x[1446]), .B(y[1446]), .Z(n1654) );
  XOR U5252 ( .A(x[240]), .B(y[240]), .Z(n1651) );
  XNOR U5253 ( .A(x[1448]), .B(y[1448]), .Z(n1652) );
  XNOR U5254 ( .A(n1651), .B(n1652), .Z(n1653) );
  XNOR U5255 ( .A(n1654), .B(n1653), .Z(n5028) );
  XNOR U5256 ( .A(n5029), .B(n5028), .Z(n5030) );
  XOR U5257 ( .A(n5031), .B(n5030), .Z(n1232) );
  XNOR U5258 ( .A(n1231), .B(n1232), .Z(n1234) );
  XOR U5259 ( .A(x[1442]), .B(y[1442]), .Z(n1874) );
  XOR U5260 ( .A(x[236]), .B(y[236]), .Z(n1871) );
  XNOR U5261 ( .A(x[1444]), .B(y[1444]), .Z(n1872) );
  XNOR U5262 ( .A(n1871), .B(n1872), .Z(n1873) );
  XOR U5263 ( .A(n1874), .B(n1873), .Z(n5757) );
  XOR U5264 ( .A(x[1438]), .B(y[1438]), .Z(n1552) );
  XOR U5265 ( .A(x[232]), .B(y[232]), .Z(n1549) );
  XNOR U5266 ( .A(x[1440]), .B(y[1440]), .Z(n1550) );
  XNOR U5267 ( .A(n1549), .B(n1550), .Z(n1551) );
  XOR U5268 ( .A(n1552), .B(n1551), .Z(n5755) );
  XOR U5269 ( .A(x[1434]), .B(y[1434]), .Z(n1756) );
  XOR U5270 ( .A(x[494]), .B(y[494]), .Z(n1753) );
  XNOR U5271 ( .A(x[1436]), .B(y[1436]), .Z(n1754) );
  XNOR U5272 ( .A(n1753), .B(n1754), .Z(n1755) );
  XNOR U5273 ( .A(n1756), .B(n1755), .Z(n5754) );
  XNOR U5274 ( .A(n5755), .B(n5754), .Z(n5756) );
  XNOR U5275 ( .A(n5757), .B(n5756), .Z(n1233) );
  XNOR U5276 ( .A(n1234), .B(n1233), .Z(n4087) );
  XOR U5277 ( .A(x[1712]), .B(y[1712]), .Z(n5312) );
  XOR U5278 ( .A(x[1714]), .B(y[1714]), .Z(n5310) );
  XNOR U5279 ( .A(x[1716]), .B(y[1716]), .Z(n5311) );
  XOR U5280 ( .A(n5310), .B(n5311), .Z(n5313) );
  XNOR U5281 ( .A(n5312), .B(n5313), .Z(n6025) );
  XOR U5282 ( .A(x[1748]), .B(y[1748]), .Z(n5097) );
  XOR U5283 ( .A(x[516]), .B(y[516]), .Z(n5094) );
  XNOR U5284 ( .A(x[1750]), .B(y[1750]), .Z(n5095) );
  XNOR U5285 ( .A(n5094), .B(n5095), .Z(n5096) );
  XOR U5286 ( .A(n5097), .B(n5096), .Z(n6024) );
  XOR U5287 ( .A(n6025), .B(n6024), .Z(n6027) );
  XOR U5288 ( .A(x[1726]), .B(y[1726]), .Z(n5792) );
  XOR U5289 ( .A(x[496]), .B(y[496]), .Z(n5790) );
  XNOR U5290 ( .A(x[1728]), .B(y[1728]), .Z(n5791) );
  XOR U5291 ( .A(n5790), .B(n5791), .Z(n5793) );
  XNOR U5292 ( .A(n5792), .B(n5793), .Z(n6026) );
  XOR U5293 ( .A(n6027), .B(n6026), .Z(n5509) );
  XOR U5294 ( .A(x[1685]), .B(y[1685]), .Z(n2977) );
  XOR U5295 ( .A(x[1687]), .B(y[1687]), .Z(n2975) );
  XNOR U5296 ( .A(x[1703]), .B(y[1703]), .Z(n2976) );
  XOR U5297 ( .A(n2975), .B(n2976), .Z(n2978) );
  XNOR U5298 ( .A(n2977), .B(n2978), .Z(n5352) );
  XOR U5299 ( .A(x[631]), .B(y[631]), .Z(n154) );
  XOR U5300 ( .A(x[615]), .B(y[615]), .Z(n152) );
  XNOR U5301 ( .A(x[623]), .B(y[623]), .Z(n153) );
  XOR U5302 ( .A(n152), .B(n153), .Z(n155) );
  XOR U5303 ( .A(n154), .B(n155), .Z(n5353) );
  XNOR U5304 ( .A(n5352), .B(n5353), .Z(n5355) );
  XOR U5305 ( .A(x[1715]), .B(y[1715]), .Z(n2983) );
  XOR U5306 ( .A(x[1681]), .B(y[1681]), .Z(n2981) );
  XNOR U5307 ( .A(x[1717]), .B(y[1717]), .Z(n2982) );
  XOR U5308 ( .A(n2981), .B(n2982), .Z(n2984) );
  XNOR U5309 ( .A(n2983), .B(n2984), .Z(n5354) );
  XNOR U5310 ( .A(n5355), .B(n5354), .Z(n5508) );
  XNOR U5311 ( .A(n5509), .B(n5508), .Z(n5511) );
  XOR U5312 ( .A(x[1776]), .B(y[1776]), .Z(n5343) );
  XOR U5313 ( .A(x[540]), .B(y[540]), .Z(n5340) );
  XNOR U5314 ( .A(x[1778]), .B(y[1778]), .Z(n5341) );
  XNOR U5315 ( .A(n5340), .B(n5341), .Z(n5342) );
  XOR U5316 ( .A(n5343), .B(n5342), .Z(n3536) );
  XOR U5317 ( .A(x[1780]), .B(y[1780]), .Z(n5181) );
  XOR U5318 ( .A(x[546]), .B(y[546]), .Z(n5178) );
  XNOR U5319 ( .A(x[1782]), .B(y[1782]), .Z(n5179) );
  XNOR U5320 ( .A(n5178), .B(n5179), .Z(n5180) );
  XOR U5321 ( .A(n5181), .B(n5180), .Z(n3534) );
  XOR U5322 ( .A(x[1704]), .B(y[1704]), .Z(n4857) );
  XOR U5323 ( .A(x[474]), .B(y[474]), .Z(n4854) );
  XNOR U5324 ( .A(x[1706]), .B(y[1706]), .Z(n4855) );
  XNOR U5325 ( .A(n4854), .B(n4855), .Z(n4856) );
  XNOR U5326 ( .A(n4857), .B(n4856), .Z(n3533) );
  XNOR U5327 ( .A(n3534), .B(n3533), .Z(n3535) );
  XNOR U5328 ( .A(n3536), .B(n3535), .Z(n5510) );
  XNOR U5329 ( .A(n5511), .B(n5510), .Z(n4086) );
  XOR U5330 ( .A(n4087), .B(n4086), .Z(n4088) );
  XNOR U5331 ( .A(n4089), .B(n4088), .Z(n660) );
  XOR U5332 ( .A(x[1646]), .B(y[1646]), .Z(n5715) );
  XOR U5333 ( .A(x[712]), .B(y[712]), .Z(n5712) );
  XNOR U5334 ( .A(x[1648]), .B(y[1648]), .Z(n5713) );
  XNOR U5335 ( .A(n5712), .B(n5713), .Z(n5714) );
  XOR U5336 ( .A(n5715), .B(n5714), .Z(n5763) );
  XOR U5337 ( .A(x[1844]), .B(y[1844]), .Z(n2006) );
  XOR U5338 ( .A(x[880]), .B(y[880]), .Z(n2003) );
  XNOR U5339 ( .A(x[1846]), .B(y[1846]), .Z(n2004) );
  XNOR U5340 ( .A(n2003), .B(n2004), .Z(n2005) );
  XOR U5341 ( .A(n2006), .B(n2005), .Z(n5761) );
  XOR U5342 ( .A(x[1640]), .B(y[1640]), .Z(n5769) );
  XOR U5343 ( .A(x[1642]), .B(y[1642]), .Z(n5766) );
  XNOR U5344 ( .A(x[1644]), .B(y[1644]), .Z(n5767) );
  XNOR U5345 ( .A(n5766), .B(n5767), .Z(n5768) );
  XNOR U5346 ( .A(n5769), .B(n5768), .Z(n5760) );
  XNOR U5347 ( .A(n5761), .B(n5760), .Z(n5762) );
  XNOR U5348 ( .A(n5763), .B(n5762), .Z(n4950) );
  XOR U5349 ( .A(x[1737]), .B(y[1737]), .Z(n612) );
  XOR U5350 ( .A(x[1657]), .B(y[1657]), .Z(n610) );
  XOR U5351 ( .A(x[1739]), .B(y[1739]), .Z(n609) );
  XOR U5352 ( .A(n610), .B(n609), .Z(n611) );
  XOR U5353 ( .A(n612), .B(n611), .Z(n4983) );
  XOR U5354 ( .A(x[539]), .B(y[539]), .Z(n289) );
  XOR U5355 ( .A(x[533]), .B(y[533]), .Z(n286) );
  XNOR U5356 ( .A(x[535]), .B(y[535]), .Z(n287) );
  XNOR U5357 ( .A(n286), .B(n287), .Z(n288) );
  XOR U5358 ( .A(n289), .B(n288), .Z(n4981) );
  XOR U5359 ( .A(x[1733]), .B(y[1733]), .Z(n522) );
  XOR U5360 ( .A(x[1705]), .B(y[1705]), .Z(n520) );
  XOR U5361 ( .A(x[1735]), .B(y[1735]), .Z(n519) );
  XOR U5362 ( .A(n520), .B(n519), .Z(n521) );
  XNOR U5363 ( .A(n522), .B(n521), .Z(n4980) );
  XNOR U5364 ( .A(n4981), .B(n4980), .Z(n4982) );
  XOR U5365 ( .A(n4983), .B(n4982), .Z(n4951) );
  XNOR U5366 ( .A(n4950), .B(n4951), .Z(n4953) );
  XOR U5367 ( .A(x[1636]), .B(y[1636]), .Z(n5787) );
  XOR U5368 ( .A(x[414]), .B(y[414]), .Z(n5784) );
  XNOR U5369 ( .A(x[1638]), .B(y[1638]), .Z(n5785) );
  XNOR U5370 ( .A(n5784), .B(n5785), .Z(n5786) );
  XOR U5371 ( .A(n5787), .B(n5786), .Z(n5229) );
  XOR U5372 ( .A(x[1848]), .B(y[1848]), .Z(n2216) );
  XOR U5373 ( .A(x[606]), .B(y[606]), .Z(n2213) );
  XNOR U5374 ( .A(x[1850]), .B(y[1850]), .Z(n2214) );
  XNOR U5375 ( .A(n2213), .B(n2214), .Z(n2215) );
  XOR U5376 ( .A(n2216), .B(n2215), .Z(n5227) );
  XOR U5377 ( .A(x[1632]), .B(y[1632]), .Z(n3500) );
  XOR U5378 ( .A(x[408]), .B(y[408]), .Z(n3497) );
  XNOR U5379 ( .A(x[1634]), .B(y[1634]), .Z(n3498) );
  XNOR U5380 ( .A(n3497), .B(n3498), .Z(n3499) );
  XNOR U5381 ( .A(n3500), .B(n3499), .Z(n5226) );
  XNOR U5382 ( .A(n5227), .B(n5226), .Z(n5228) );
  XNOR U5383 ( .A(n5229), .B(n5228), .Z(n4952) );
  XNOR U5384 ( .A(n4953), .B(n4952), .Z(n4005) );
  XOR U5385 ( .A(x[1628]), .B(y[1628]), .Z(n5301) );
  XOR U5386 ( .A(x[692]), .B(y[692]), .Z(n5298) );
  XNOR U5387 ( .A(x[1630]), .B(y[1630]), .Z(n5299) );
  XNOR U5388 ( .A(n5298), .B(n5299), .Z(n5300) );
  XOR U5389 ( .A(n5301), .B(n5300), .Z(n5325) );
  XOR U5390 ( .A(x[1852]), .B(y[1852]), .Z(n2156) );
  XOR U5391 ( .A(x[612]), .B(y[612]), .Z(n2153) );
  XNOR U5392 ( .A(x[1854]), .B(y[1854]), .Z(n2154) );
  XNOR U5393 ( .A(n2153), .B(n2154), .Z(n2155) );
  XOR U5394 ( .A(n2156), .B(n2155), .Z(n5323) );
  XOR U5395 ( .A(x[1622]), .B(y[1622]), .Z(n3512) );
  XOR U5396 ( .A(x[1624]), .B(y[1624]), .Z(n3509) );
  XNOR U5397 ( .A(x[1626]), .B(y[1626]), .Z(n3510) );
  XNOR U5398 ( .A(n3509), .B(n3510), .Z(n3511) );
  XNOR U5399 ( .A(n3512), .B(n3511), .Z(n5322) );
  XNOR U5400 ( .A(n5323), .B(n5322), .Z(n5324) );
  XNOR U5401 ( .A(n5325), .B(n5324), .Z(n3918) );
  XOR U5402 ( .A(x[1616]), .B(y[1616]), .Z(n4845) );
  XOR U5403 ( .A(x[1618]), .B(y[1618]), .Z(n4842) );
  XNOR U5404 ( .A(x[1620]), .B(y[1620]), .Z(n4843) );
  XNOR U5405 ( .A(n4842), .B(n4843), .Z(n4844) );
  XOR U5406 ( .A(n4845), .B(n4844), .Z(n5349) );
  XOR U5407 ( .A(x[1612]), .B(y[1612]), .Z(n3506) );
  XOR U5408 ( .A(x[392]), .B(y[392]), .Z(n3503) );
  XNOR U5409 ( .A(x[1614]), .B(y[1614]), .Z(n3504) );
  XNOR U5410 ( .A(n3503), .B(n3504), .Z(n3505) );
  XOR U5411 ( .A(n3506), .B(n3505), .Z(n5347) );
  XOR U5412 ( .A(x[1608]), .B(y[1608]), .Z(n4899) );
  XOR U5413 ( .A(x[388]), .B(y[388]), .Z(n4896) );
  XNOR U5414 ( .A(x[1610]), .B(y[1610]), .Z(n4897) );
  XNOR U5415 ( .A(n4896), .B(n4897), .Z(n4898) );
  XNOR U5416 ( .A(n4899), .B(n4898), .Z(n5346) );
  XNOR U5417 ( .A(n5347), .B(n5346), .Z(n5348) );
  XOR U5418 ( .A(n5349), .B(n5348), .Z(n3919) );
  XNOR U5419 ( .A(n3918), .B(n3919), .Z(n3921) );
  XOR U5420 ( .A(x[1604]), .B(y[1604]), .Z(n5469) );
  XOR U5421 ( .A(x[384]), .B(y[384]), .Z(n5466) );
  XNOR U5422 ( .A(x[1606]), .B(y[1606]), .Z(n5467) );
  XNOR U5423 ( .A(n5466), .B(n5467), .Z(n5468) );
  XOR U5424 ( .A(n5469), .B(n5468), .Z(n6033) );
  XOR U5425 ( .A(x[1598]), .B(y[1598]), .Z(n5187) );
  XOR U5426 ( .A(x[1600]), .B(y[1600]), .Z(n5184) );
  XNOR U5427 ( .A(x[1602]), .B(y[1602]), .Z(n5185) );
  XNOR U5428 ( .A(n5184), .B(n5185), .Z(n5186) );
  XOR U5429 ( .A(n5187), .B(n5186), .Z(n6031) );
  XOR U5430 ( .A(x[1594]), .B(y[1594]), .Z(n5085) );
  XOR U5431 ( .A(x[662]), .B(y[662]), .Z(n5082) );
  XNOR U5432 ( .A(x[1596]), .B(y[1596]), .Z(n5083) );
  XNOR U5433 ( .A(n5082), .B(n5083), .Z(n5084) );
  XNOR U5434 ( .A(n5085), .B(n5084), .Z(n6030) );
  XNOR U5435 ( .A(n6031), .B(n6030), .Z(n6032) );
  XNOR U5436 ( .A(n6033), .B(n6032), .Z(n3920) );
  XNOR U5437 ( .A(n3921), .B(n3920), .Z(n4003) );
  XOR U5438 ( .A(x[1798]), .B(y[1798]), .Z(n5373) );
  XOR U5439 ( .A(x[562]), .B(y[562]), .Z(n5370) );
  XNOR U5440 ( .A(x[1800]), .B(y[1800]), .Z(n5371) );
  XNOR U5441 ( .A(n5370), .B(n5371), .Z(n5372) );
  XOR U5442 ( .A(n5373), .B(n5372), .Z(n4605) );
  XOR U5443 ( .A(x[1722]), .B(y[1722]), .Z(n5799) );
  XOR U5444 ( .A(x[786]), .B(y[786]), .Z(n5796) );
  XNOR U5445 ( .A(x[1724]), .B(y[1724]), .Z(n5797) );
  XNOR U5446 ( .A(n5796), .B(n5797), .Z(n5798) );
  XOR U5447 ( .A(n5799), .B(n5798), .Z(n4603) );
  XOR U5448 ( .A(x[1694]), .B(y[1694]), .Z(n5481) );
  XOR U5449 ( .A(x[1696]), .B(y[1696]), .Z(n5478) );
  XNOR U5450 ( .A(x[1698]), .B(y[1698]), .Z(n5479) );
  XNOR U5451 ( .A(n5478), .B(n5479), .Z(n5480) );
  XNOR U5452 ( .A(n5481), .B(n5480), .Z(n4602) );
  XNOR U5453 ( .A(n4603), .B(n4602), .Z(n4604) );
  XNOR U5454 ( .A(n4605), .B(n4604), .Z(n6018) );
  XOR U5455 ( .A(x[1677]), .B(y[1677]), .Z(n492) );
  XOR U5456 ( .A(x[1693]), .B(y[1693]), .Z(n489) );
  XNOR U5457 ( .A(x[1725]), .B(y[1725]), .Z(n490) );
  XNOR U5458 ( .A(n489), .B(n490), .Z(n491) );
  XOR U5459 ( .A(n492), .B(n491), .Z(n6063) );
  XOR U5460 ( .A(x[1679]), .B(y[1679]), .Z(n480) );
  XOR U5461 ( .A(x[1691]), .B(y[1691]), .Z(n477) );
  XNOR U5462 ( .A(x[1723]), .B(y[1723]), .Z(n478) );
  XNOR U5463 ( .A(n477), .B(n478), .Z(n479) );
  XOR U5464 ( .A(n480), .B(n479), .Z(n6061) );
  XOR U5465 ( .A(x[1719]), .B(y[1719]), .Z(n486) );
  XOR U5466 ( .A(x[1697]), .B(y[1697]), .Z(n483) );
  XNOR U5467 ( .A(x[1721]), .B(y[1721]), .Z(n484) );
  XNOR U5468 ( .A(n483), .B(n484), .Z(n485) );
  XNOR U5469 ( .A(n486), .B(n485), .Z(n6060) );
  XNOR U5470 ( .A(n6061), .B(n6060), .Z(n6062) );
  XOR U5471 ( .A(n6063), .B(n6062), .Z(n6019) );
  XNOR U5472 ( .A(n6018), .B(n6019), .Z(n6021) );
  XOR U5473 ( .A(x[1802]), .B(y[1802]), .Z(n5367) );
  XOR U5474 ( .A(x[566]), .B(y[566]), .Z(n5364) );
  XNOR U5475 ( .A(x[1804]), .B(y[1804]), .Z(n5365) );
  XNOR U5476 ( .A(n5364), .B(n5365), .Z(n5366) );
  XOR U5477 ( .A(n5367), .B(n5366), .Z(n4629) );
  XOR U5478 ( .A(x[1734]), .B(y[1734]), .Z(n5727) );
  XOR U5479 ( .A(x[504]), .B(y[504]), .Z(n5724) );
  XNOR U5480 ( .A(x[1736]), .B(y[1736]), .Z(n5725) );
  XNOR U5481 ( .A(n5724), .B(n5725), .Z(n5726) );
  XOR U5482 ( .A(n5727), .B(n5726), .Z(n4627) );
  XOR U5483 ( .A(x[1806]), .B(y[1806]), .Z(n5385) );
  XOR U5484 ( .A(x[570]), .B(y[570]), .Z(n5382) );
  XNOR U5485 ( .A(x[1808]), .B(y[1808]), .Z(n5383) );
  XNOR U5486 ( .A(n5382), .B(n5383), .Z(n5384) );
  XNOR U5487 ( .A(n5385), .B(n5384), .Z(n4626) );
  XNOR U5488 ( .A(n4627), .B(n4626), .Z(n4628) );
  XNOR U5489 ( .A(n4629), .B(n4628), .Z(n6020) );
  XNOR U5490 ( .A(n6021), .B(n6020), .Z(n4002) );
  XOR U5491 ( .A(n4003), .B(n4002), .Z(n4004) );
  XNOR U5492 ( .A(n4005), .B(n4004), .Z(n658) );
  XOR U5493 ( .A(x[1590]), .B(y[1590]), .Z(n3524) );
  XOR U5494 ( .A(x[372]), .B(y[372]), .Z(n3521) );
  XNOR U5495 ( .A(x[1592]), .B(y[1592]), .Z(n3522) );
  XNOR U5496 ( .A(n3521), .B(n3522), .Z(n3523) );
  XOR U5497 ( .A(n3524), .B(n3523), .Z(n5217) );
  XOR U5498 ( .A(x[1586]), .B(y[1586]), .Z(n5679) );
  XOR U5499 ( .A(x[368]), .B(y[368]), .Z(n5676) );
  XNOR U5500 ( .A(x[1588]), .B(y[1588]), .Z(n5677) );
  XNOR U5501 ( .A(n5676), .B(n5677), .Z(n5678) );
  XOR U5502 ( .A(n5679), .B(n5678), .Z(n5215) );
  XOR U5503 ( .A(x[1582]), .B(y[1582]), .Z(n5991) );
  XOR U5504 ( .A(x[364]), .B(y[364]), .Z(n5988) );
  XNOR U5505 ( .A(x[1584]), .B(y[1584]), .Z(n5989) );
  XNOR U5506 ( .A(n5988), .B(n5989), .Z(n5990) );
  XNOR U5507 ( .A(n5991), .B(n5990), .Z(n5214) );
  XNOR U5508 ( .A(n5215), .B(n5214), .Z(n5216) );
  XNOR U5509 ( .A(n5217), .B(n5216), .Z(n1471) );
  XOR U5510 ( .A(x[1578]), .B(y[1578]), .Z(n5451) );
  XOR U5511 ( .A(x[644]), .B(y[644]), .Z(n5448) );
  XNOR U5512 ( .A(x[1580]), .B(y[1580]), .Z(n5449) );
  XNOR U5513 ( .A(n5448), .B(n5449), .Z(n5450) );
  XOR U5514 ( .A(n5451), .B(n5450), .Z(n5205) );
  XOR U5515 ( .A(x[1574]), .B(y[1574]), .Z(n4671) );
  XOR U5516 ( .A(x[640]), .B(y[640]), .Z(n4668) );
  XNOR U5517 ( .A(x[1576]), .B(y[1576]), .Z(n4669) );
  XNOR U5518 ( .A(n4668), .B(n4669), .Z(n4670) );
  XOR U5519 ( .A(n4671), .B(n4670), .Z(n5203) );
  XOR U5520 ( .A(x[1568]), .B(y[1568]), .Z(n5985) );
  XOR U5521 ( .A(x[1570]), .B(y[1570]), .Z(n5982) );
  XNOR U5522 ( .A(x[1572]), .B(y[1572]), .Z(n5983) );
  XNOR U5523 ( .A(n5982), .B(n5983), .Z(n5984) );
  XNOR U5524 ( .A(n5985), .B(n5984), .Z(n5202) );
  XNOR U5525 ( .A(n5203), .B(n5202), .Z(n5204) );
  XOR U5526 ( .A(n5205), .B(n5204), .Z(n1472) );
  XNOR U5527 ( .A(n1471), .B(n1472), .Z(n1474) );
  XOR U5528 ( .A(x[1564]), .B(y[1564]), .Z(n4677) );
  XOR U5529 ( .A(x[348]), .B(y[348]), .Z(n4674) );
  XNOR U5530 ( .A(x[1566]), .B(y[1566]), .Z(n4675) );
  XNOR U5531 ( .A(n4674), .B(n4675), .Z(n4676) );
  XOR U5532 ( .A(n4677), .B(n4676), .Z(n4749) );
  XOR U5533 ( .A(x[1560]), .B(y[1560]), .Z(n5463) );
  XOR U5534 ( .A(x[342]), .B(y[342]), .Z(n5460) );
  XNOR U5535 ( .A(x[1562]), .B(y[1562]), .Z(n5461) );
  XNOR U5536 ( .A(n5460), .B(n5461), .Z(n5462) );
  XOR U5537 ( .A(n5463), .B(n5462), .Z(n4747) );
  XOR U5538 ( .A(x[1556]), .B(y[1556]), .Z(n5439) );
  XOR U5539 ( .A(x[620]), .B(y[620]), .Z(n5436) );
  XNOR U5540 ( .A(x[1558]), .B(y[1558]), .Z(n5437) );
  XNOR U5541 ( .A(n5436), .B(n5437), .Z(n5438) );
  XNOR U5542 ( .A(n5439), .B(n5438), .Z(n4746) );
  XNOR U5543 ( .A(n4747), .B(n4746), .Z(n4748) );
  XNOR U5544 ( .A(n4749), .B(n4748), .Z(n1473) );
  XOR U5545 ( .A(n1474), .B(n1473), .Z(n4077) );
  XOR U5546 ( .A(x[1550]), .B(y[1550]), .Z(n5445) );
  XOR U5547 ( .A(x[1552]), .B(y[1552]), .Z(n5442) );
  XNOR U5548 ( .A(x[1554]), .B(y[1554]), .Z(n5443) );
  XNOR U5549 ( .A(n5442), .B(n5443), .Z(n5444) );
  XOR U5550 ( .A(n5445), .B(n5444), .Z(n5223) );
  XOR U5551 ( .A(x[1544]), .B(y[1544]), .Z(n367) );
  XOR U5552 ( .A(x[1546]), .B(y[1546]), .Z(n364) );
  XNOR U5553 ( .A(x[1548]), .B(y[1548]), .Z(n365) );
  XNOR U5554 ( .A(n364), .B(n365), .Z(n366) );
  XOR U5555 ( .A(n367), .B(n366), .Z(n5221) );
  XOR U5556 ( .A(x[1540]), .B(y[1540]), .Z(n4911) );
  XOR U5557 ( .A(x[326]), .B(y[326]), .Z(n4908) );
  XNOR U5558 ( .A(x[1542]), .B(y[1542]), .Z(n4909) );
  XNOR U5559 ( .A(n4908), .B(n4909), .Z(n4910) );
  XNOR U5560 ( .A(n4911), .B(n4910), .Z(n5220) );
  XNOR U5561 ( .A(n5221), .B(n5220), .Z(n5222) );
  XNOR U5562 ( .A(n5223), .B(n5222), .Z(n1099) );
  XOR U5563 ( .A(x[1536]), .B(y[1536]), .Z(n4905) );
  XOR U5564 ( .A(x[322]), .B(y[322]), .Z(n4902) );
  XNOR U5565 ( .A(x[1538]), .B(y[1538]), .Z(n4903) );
  XNOR U5566 ( .A(n4902), .B(n4903), .Z(n4904) );
  XOR U5567 ( .A(n4905), .B(n4904), .Z(n5235) );
  XOR U5568 ( .A(x[1532]), .B(y[1532]), .Z(n5265) );
  XOR U5569 ( .A(x[318]), .B(y[318]), .Z(n5262) );
  XNOR U5570 ( .A(x[1534]), .B(y[1534]), .Z(n5263) );
  XNOR U5571 ( .A(n5262), .B(n5263), .Z(n5264) );
  XOR U5572 ( .A(n5265), .B(n5264), .Z(n5233) );
  XOR U5573 ( .A(x[1526]), .B(y[1526]), .Z(n3326) );
  XOR U5574 ( .A(x[1528]), .B(y[1528]), .Z(n3323) );
  XNOR U5575 ( .A(x[1530]), .B(y[1530]), .Z(n3324) );
  XNOR U5576 ( .A(n3323), .B(n3324), .Z(n3325) );
  XNOR U5577 ( .A(n3326), .B(n3325), .Z(n5232) );
  XNOR U5578 ( .A(n5233), .B(n5232), .Z(n5234) );
  XOR U5579 ( .A(n5235), .B(n5234), .Z(n1100) );
  XNOR U5580 ( .A(n1099), .B(n1100), .Z(n1102) );
  XOR U5581 ( .A(x[1522]), .B(y[1522]), .Z(n5259) );
  XOR U5582 ( .A(x[588]), .B(y[588]), .Z(n5256) );
  XNOR U5583 ( .A(x[1524]), .B(y[1524]), .Z(n5257) );
  XNOR U5584 ( .A(n5256), .B(n5257), .Z(n5258) );
  XOR U5585 ( .A(n5259), .B(n5258), .Z(n6069) );
  XOR U5586 ( .A(x[1518]), .B(y[1518]), .Z(n5781) );
  XOR U5587 ( .A(x[306]), .B(y[306]), .Z(n5778) );
  XNOR U5588 ( .A(x[1520]), .B(y[1520]), .Z(n5779) );
  XNOR U5589 ( .A(n5778), .B(n5779), .Z(n5780) );
  XOR U5590 ( .A(n5781), .B(n5780), .Z(n6067) );
  XOR U5591 ( .A(x[1514]), .B(y[1514]), .Z(n5775) );
  XOR U5592 ( .A(x[302]), .B(y[302]), .Z(n5772) );
  XNOR U5593 ( .A(x[1516]), .B(y[1516]), .Z(n5773) );
  XNOR U5594 ( .A(n5772), .B(n5773), .Z(n5774) );
  XNOR U5595 ( .A(n5775), .B(n5774), .Z(n6066) );
  XNOR U5596 ( .A(n6067), .B(n6066), .Z(n6068) );
  XNOR U5597 ( .A(n6069), .B(n6068), .Z(n1101) );
  XNOR U5598 ( .A(n1102), .B(n1101), .Z(n4075) );
  XOR U5599 ( .A(x[230]), .B(y[230]), .Z(n2509) );
  XOR U5600 ( .A(x[234]), .B(y[234]), .Z(n2507) );
  XNOR U5601 ( .A(x[1007]), .B(y[1007]), .Z(n2508) );
  XOR U5602 ( .A(n2507), .B(n2508), .Z(n2510) );
  XNOR U5603 ( .A(n2509), .B(n2510), .Z(n1633) );
  XOR U5604 ( .A(x[1214]), .B(y[1214]), .Z(n2035) );
  XOR U5605 ( .A(x[129]), .B(y[129]), .Z(n2033) );
  XNOR U5606 ( .A(x[1216]), .B(y[1216]), .Z(n2034) );
  XOR U5607 ( .A(n2033), .B(n2034), .Z(n2036) );
  XOR U5608 ( .A(n2035), .B(n2036), .Z(n1634) );
  XNOR U5609 ( .A(n1633), .B(n1634), .Z(n1636) );
  XOR U5610 ( .A(x[238]), .B(y[238]), .Z(n2773) );
  XOR U5611 ( .A(x[242]), .B(y[242]), .Z(n2771) );
  XNOR U5612 ( .A(x[731]), .B(y[731]), .Z(n2772) );
  XOR U5613 ( .A(n2771), .B(n2772), .Z(n2774) );
  XNOR U5614 ( .A(n2773), .B(n2774), .Z(n1635) );
  XOR U5615 ( .A(n1636), .B(n1635), .Z(n5317) );
  XOR U5616 ( .A(x[1784]), .B(y[1784]), .Z(n5408) );
  XOR U5617 ( .A(x[1786]), .B(y[1786]), .Z(n5406) );
  XNOR U5618 ( .A(x[1788]), .B(y[1788]), .Z(n5407) );
  XOR U5619 ( .A(n5406), .B(n5407), .Z(n5409) );
  XOR U5620 ( .A(n5408), .B(n5409), .Z(n4664) );
  XOR U5621 ( .A(x[1708]), .B(y[1708]), .Z(n4850) );
  XOR U5622 ( .A(x[480]), .B(y[480]), .Z(n4848) );
  XNOR U5623 ( .A(x[1710]), .B(y[1710]), .Z(n4849) );
  XOR U5624 ( .A(n4848), .B(n4849), .Z(n4851) );
  XOR U5625 ( .A(n4850), .B(n4851), .Z(n4663) );
  XOR U5626 ( .A(x[1790]), .B(y[1790]), .Z(n5337) );
  XOR U5627 ( .A(x[838]), .B(y[838]), .Z(n5334) );
  XNOR U5628 ( .A(x[1792]), .B(y[1792]), .Z(n5335) );
  XNOR U5629 ( .A(n5334), .B(n5335), .Z(n5336) );
  XNOR U5630 ( .A(n5337), .B(n5336), .Z(n4662) );
  XOR U5631 ( .A(n4663), .B(n4662), .Z(n4665) );
  XOR U5632 ( .A(n4664), .B(n4665), .Z(n5316) );
  XNOR U5633 ( .A(n5317), .B(n5316), .Z(n5319) );
  XOR U5634 ( .A(x[1794]), .B(y[1794]), .Z(n5402) );
  XOR U5635 ( .A(x[842]), .B(y[842]), .Z(n5400) );
  XNOR U5636 ( .A(x[1796]), .B(y[1796]), .Z(n5401) );
  XOR U5637 ( .A(n5400), .B(n5401), .Z(n5403) );
  XOR U5638 ( .A(n5402), .B(n5403), .Z(n4688) );
  XOR U5639 ( .A(x[1718]), .B(y[1718]), .Z(n5306) );
  XOR U5640 ( .A(x[782]), .B(y[782]), .Z(n5304) );
  XNOR U5641 ( .A(x[1720]), .B(y[1720]), .Z(n5305) );
  XOR U5642 ( .A(n5304), .B(n5305), .Z(n5307) );
  XOR U5643 ( .A(n5306), .B(n5307), .Z(n4687) );
  XOR U5644 ( .A(x[1700]), .B(y[1700]), .Z(n5475) );
  XOR U5645 ( .A(x[768]), .B(y[768]), .Z(n5472) );
  XNOR U5646 ( .A(x[1702]), .B(y[1702]), .Z(n5473) );
  XNOR U5647 ( .A(n5472), .B(n5473), .Z(n5474) );
  XNOR U5648 ( .A(n5475), .B(n5474), .Z(n4686) );
  XOR U5649 ( .A(n4687), .B(n4686), .Z(n4689) );
  XOR U5650 ( .A(n4688), .B(n4689), .Z(n5318) );
  XNOR U5651 ( .A(n5319), .B(n5318), .Z(n4074) );
  XOR U5652 ( .A(n4075), .B(n4074), .Z(n4076) );
  XOR U5653 ( .A(n4077), .B(n4076), .Z(n657) );
  XOR U5654 ( .A(n658), .B(n657), .Z(n659) );
  XNOR U5655 ( .A(n660), .B(n659), .Z(n3799) );
  XOR U5656 ( .A(x[920]), .B(y[920]), .Z(n1708) );
  XOR U5657 ( .A(x[922]), .B(y[922]), .Z(n1705) );
  XNOR U5658 ( .A(x[1945]), .B(y[1945]), .Z(n1706) );
  XNOR U5659 ( .A(n1705), .B(n1706), .Z(n1707) );
  XOR U5660 ( .A(n1708), .B(n1707), .Z(n221) );
  XOR U5661 ( .A(x[916]), .B(y[916]), .Z(n1558) );
  XOR U5662 ( .A(x[327]), .B(y[327]), .Z(n1555) );
  XNOR U5663 ( .A(x[918]), .B(y[918]), .Z(n1556) );
  XNOR U5664 ( .A(n1555), .B(n1556), .Z(n1557) );
  XOR U5665 ( .A(n1558), .B(n1557), .Z(n219) );
  XOR U5666 ( .A(x[912]), .B(y[912]), .Z(n1066) );
  XOR U5667 ( .A(x[331]), .B(y[331]), .Z(n1063) );
  XNOR U5668 ( .A(x[914]), .B(y[914]), .Z(n1064) );
  XNOR U5669 ( .A(n1063), .B(n1064), .Z(n1065) );
  XNOR U5670 ( .A(n1066), .B(n1065), .Z(n218) );
  XNOR U5671 ( .A(n219), .B(n218), .Z(n220) );
  XNOR U5672 ( .A(n221), .B(n220), .Z(n4368) );
  XOR U5673 ( .A(x[906]), .B(y[906]), .Z(n4149) );
  XOR U5674 ( .A(x[701]), .B(y[701]), .Z(n4146) );
  XNOR U5675 ( .A(x[908]), .B(y[908]), .Z(n4147) );
  XNOR U5676 ( .A(n4146), .B(n4147), .Z(n4148) );
  XOR U5677 ( .A(n4149), .B(n4148), .Z(n2180) );
  XOR U5678 ( .A(x[902]), .B(y[902]), .Z(n4143) );
  XOR U5679 ( .A(x[337]), .B(y[337]), .Z(n4140) );
  XNOR U5680 ( .A(x[904]), .B(y[904]), .Z(n4141) );
  XNOR U5681 ( .A(n4140), .B(n4141), .Z(n4142) );
  XOR U5682 ( .A(n4143), .B(n4142), .Z(n2178) );
  XOR U5683 ( .A(x[896]), .B(y[896]), .Z(n4539) );
  XOR U5684 ( .A(x[707]), .B(y[707]), .Z(n4536) );
  XNOR U5685 ( .A(x[900]), .B(y[900]), .Z(n4537) );
  XNOR U5686 ( .A(n4536), .B(n4537), .Z(n4538) );
  XNOR U5687 ( .A(n4539), .B(n4538), .Z(n2177) );
  XNOR U5688 ( .A(n2178), .B(n2177), .Z(n2179) );
  XOR U5689 ( .A(n2180), .B(n2179), .Z(n4369) );
  XNOR U5690 ( .A(n4368), .B(n4369), .Z(n4371) );
  XOR U5691 ( .A(x[890]), .B(y[890]), .Z(n1138) );
  XOR U5692 ( .A(x[892]), .B(y[892]), .Z(n1135) );
  XNOR U5693 ( .A(x[1943]), .B(y[1943]), .Z(n1136) );
  XNOR U5694 ( .A(n1135), .B(n1136), .Z(n1137) );
  XOR U5695 ( .A(n1138), .B(n1137), .Z(n5163) );
  XOR U5696 ( .A(x[886]), .B(y[886]), .Z(n1258) );
  XOR U5697 ( .A(x[343]), .B(y[343]), .Z(n1255) );
  XNOR U5698 ( .A(x[888]), .B(y[888]), .Z(n1256) );
  XNOR U5699 ( .A(n1255), .B(n1256), .Z(n1257) );
  XOR U5700 ( .A(n1258), .B(n1257), .Z(n5161) );
  XOR U5701 ( .A(x[882]), .B(y[882]), .Z(n4545) );
  XOR U5702 ( .A(x[884]), .B(y[884]), .Z(n4542) );
  XNOR U5703 ( .A(x[1941]), .B(y[1941]), .Z(n4543) );
  XNOR U5704 ( .A(n4542), .B(n4543), .Z(n4544) );
  XNOR U5705 ( .A(n4545), .B(n4544), .Z(n5160) );
  XNOR U5706 ( .A(n5161), .B(n5160), .Z(n5162) );
  XNOR U5707 ( .A(n5163), .B(n5162), .Z(n4370) );
  XNOR U5708 ( .A(n4371), .B(n4370), .Z(n4821) );
  XOR U5709 ( .A(x[876]), .B(y[876]), .Z(n1072) );
  XOR U5710 ( .A(x[349]), .B(y[349]), .Z(n1070) );
  XOR U5711 ( .A(x[878]), .B(y[878]), .Z(n1069) );
  XOR U5712 ( .A(n1070), .B(n1069), .Z(n1071) );
  XOR U5713 ( .A(n1072), .B(n1071), .Z(n2408) );
  XOR U5714 ( .A(x[872]), .B(y[872]), .Z(n1714) );
  XOR U5715 ( .A(x[353]), .B(y[353]), .Z(n1712) );
  XOR U5716 ( .A(x[874]), .B(y[874]), .Z(n1711) );
  XOR U5717 ( .A(n1712), .B(n1711), .Z(n1713) );
  XOR U5718 ( .A(n1714), .B(n1713), .Z(n2406) );
  XOR U5719 ( .A(x[868]), .B(y[868]), .Z(n1624) );
  XOR U5720 ( .A(x[721]), .B(y[721]), .Z(n1622) );
  XOR U5721 ( .A(x[870]), .B(y[870]), .Z(n1621) );
  XOR U5722 ( .A(n1622), .B(n1621), .Z(n1623) );
  XNOR U5723 ( .A(n1624), .B(n1623), .Z(n2405) );
  XNOR U5724 ( .A(n2406), .B(n2405), .Z(n2407) );
  XNOR U5725 ( .A(n2408), .B(n2407), .Z(n4242) );
  XOR U5726 ( .A(x[864]), .B(y[864]), .Z(n1796) );
  XOR U5727 ( .A(x[359]), .B(y[359]), .Z(n1794) );
  XOR U5728 ( .A(x[866]), .B(y[866]), .Z(n1793) );
  XOR U5729 ( .A(n1794), .B(n1793), .Z(n1795) );
  XOR U5730 ( .A(n1796), .B(n1795), .Z(n2378) );
  XOR U5731 ( .A(x[1856]), .B(y[1856]), .Z(n2444) );
  XOR U5732 ( .A(x[1858]), .B(y[1858]), .Z(n2441) );
  XNOR U5733 ( .A(x[1860]), .B(y[1860]), .Z(n2442) );
  XNOR U5734 ( .A(n2441), .B(n2442), .Z(n2443) );
  XOR U5735 ( .A(n2444), .B(n2443), .Z(n2376) );
  XOR U5736 ( .A(x[860]), .B(y[860]), .Z(n1802) );
  XOR U5737 ( .A(x[727]), .B(y[727]), .Z(n1800) );
  XOR U5738 ( .A(x[862]), .B(y[862]), .Z(n1799) );
  XOR U5739 ( .A(n1800), .B(n1799), .Z(n1801) );
  XNOR U5740 ( .A(n1802), .B(n1801), .Z(n2375) );
  XNOR U5741 ( .A(n2376), .B(n2375), .Z(n2377) );
  XOR U5742 ( .A(n2378), .B(n2377), .Z(n4243) );
  XNOR U5743 ( .A(n4242), .B(n4243), .Z(n4245) );
  XOR U5744 ( .A(x[856]), .B(y[856]), .Z(n4191) );
  XOR U5745 ( .A(x[858]), .B(y[858]), .Z(n4188) );
  XNOR U5746 ( .A(x[1939]), .B(y[1939]), .Z(n4189) );
  XNOR U5747 ( .A(n4188), .B(n4189), .Z(n4190) );
  XOR U5748 ( .A(n4191), .B(n4190), .Z(n2264) );
  XOR U5749 ( .A(x[1400]), .B(y[1400]), .Z(n2282) );
  XOR U5750 ( .A(x[1402]), .B(y[1402]), .Z(n2279) );
  XNOR U5751 ( .A(x[1404]), .B(y[1404]), .Z(n2280) );
  XNOR U5752 ( .A(n2279), .B(n2280), .Z(n2281) );
  XOR U5753 ( .A(n2282), .B(n2281), .Z(n2262) );
  XOR U5754 ( .A(x[850]), .B(y[850]), .Z(n1456) );
  XOR U5755 ( .A(x[365]), .B(y[365]), .Z(n1453) );
  XNOR U5756 ( .A(x[852]), .B(y[852]), .Z(n1454) );
  XNOR U5757 ( .A(n1453), .B(n1454), .Z(n1455) );
  XNOR U5758 ( .A(n1456), .B(n1455), .Z(n2261) );
  XNOR U5759 ( .A(n2262), .B(n2261), .Z(n2263) );
  XNOR U5760 ( .A(n2264), .B(n2263), .Z(n4244) );
  XNOR U5761 ( .A(n4245), .B(n4244), .Z(n4819) );
  XOR U5762 ( .A(x[846]), .B(y[846]), .Z(n2258) );
  XOR U5763 ( .A(x[848]), .B(y[848]), .Z(n2256) );
  XOR U5764 ( .A(x[1937]), .B(y[1937]), .Z(n2255) );
  XOR U5765 ( .A(n2256), .B(n2255), .Z(n2257) );
  XOR U5766 ( .A(n2258), .B(n2257), .Z(n2432) );
  XOR U5767 ( .A(x[1862]), .B(y[1862]), .Z(n2396) );
  XOR U5768 ( .A(x[894]), .B(y[894]), .Z(n2393) );
  XNOR U5769 ( .A(x[1864]), .B(y[1864]), .Z(n2394) );
  XNOR U5770 ( .A(n2393), .B(n2394), .Z(n2395) );
  XOR U5771 ( .A(n2396), .B(n2395), .Z(n2430) );
  XOR U5772 ( .A(x[840]), .B(y[840]), .Z(n2252) );
  XOR U5773 ( .A(x[371]), .B(y[371]), .Z(n2250) );
  XOR U5774 ( .A(x[844]), .B(y[844]), .Z(n2249) );
  XOR U5775 ( .A(n2250), .B(n2249), .Z(n2251) );
  XNOR U5776 ( .A(n2252), .B(n2251), .Z(n2429) );
  XNOR U5777 ( .A(n2430), .B(n2429), .Z(n2431) );
  XNOR U5778 ( .A(n2432), .B(n2431), .Z(n1847) );
  XOR U5779 ( .A(x[834]), .B(y[834]), .Z(n2300) );
  XOR U5780 ( .A(x[375]), .B(y[375]), .Z(n2297) );
  XNOR U5781 ( .A(x[836]), .B(y[836]), .Z(n2298) );
  XNOR U5782 ( .A(n2297), .B(n2298), .Z(n2299) );
  XOR U5783 ( .A(n2300), .B(n2299), .Z(n2462) );
  XOR U5784 ( .A(x[1392]), .B(y[1392]), .Z(n2348) );
  XOR U5785 ( .A(x[190]), .B(y[190]), .Z(n2346) );
  XOR U5786 ( .A(x[1394]), .B(y[1394]), .Z(n2345) );
  XOR U5787 ( .A(n2346), .B(n2345), .Z(n2347) );
  XOR U5788 ( .A(n2348), .B(n2347), .Z(n2460) );
  XOR U5789 ( .A(x[830]), .B(y[830]), .Z(n2354) );
  XOR U5790 ( .A(x[741]), .B(y[741]), .Z(n2352) );
  XOR U5791 ( .A(x[832]), .B(y[832]), .Z(n2351) );
  XOR U5792 ( .A(n2352), .B(n2351), .Z(n2353) );
  XNOR U5793 ( .A(n2354), .B(n2353), .Z(n2459) );
  XNOR U5794 ( .A(n2460), .B(n2459), .Z(n2461) );
  XOR U5795 ( .A(n2462), .B(n2461), .Z(n1848) );
  XNOR U5796 ( .A(n1847), .B(n1848), .Z(n1850) );
  XOR U5797 ( .A(x[826]), .B(y[826]), .Z(n2744) );
  XOR U5798 ( .A(x[381]), .B(y[381]), .Z(n2741) );
  XNOR U5799 ( .A(x[828]), .B(y[828]), .Z(n2742) );
  XNOR U5800 ( .A(n2741), .B(n2742), .Z(n2743) );
  XOR U5801 ( .A(n2744), .B(n2743), .Z(n2240) );
  XOR U5802 ( .A(x[1866]), .B(y[1866]), .Z(n2372) );
  XOR U5803 ( .A(x[898]), .B(y[898]), .Z(n2369) );
  XNOR U5804 ( .A(x[1868]), .B(y[1868]), .Z(n2370) );
  XNOR U5805 ( .A(n2369), .B(n2370), .Z(n2371) );
  XOR U5806 ( .A(n2372), .B(n2371), .Z(n2238) );
  XOR U5807 ( .A(x[820]), .B(y[820]), .Z(n3290) );
  XOR U5808 ( .A(x[747]), .B(y[747]), .Z(n3287) );
  XNOR U5809 ( .A(x[822]), .B(y[822]), .Z(n3288) );
  XNOR U5810 ( .A(n3287), .B(n3288), .Z(n3289) );
  XNOR U5811 ( .A(n3290), .B(n3289), .Z(n2237) );
  XNOR U5812 ( .A(n2238), .B(n2237), .Z(n2239) );
  XNOR U5813 ( .A(n2240), .B(n2239), .Z(n1849) );
  XNOR U5814 ( .A(n1850), .B(n1849), .Z(n4818) );
  XOR U5815 ( .A(n4819), .B(n4818), .Z(n4820) );
  XNOR U5816 ( .A(n4821), .B(n4820), .Z(n3812) );
  XOR U5817 ( .A(x[1154]), .B(y[1154]), .Z(n5889) );
  XOR U5818 ( .A(x[1156]), .B(y[1156]), .Z(n5886) );
  XNOR U5819 ( .A(x[1973]), .B(y[1973]), .Z(n5887) );
  XNOR U5820 ( .A(n5886), .B(n5887), .Z(n5888) );
  XOR U5821 ( .A(n5889), .B(n5888), .Z(n2846) );
  XOR U5822 ( .A(x[1146]), .B(y[1146]), .Z(n5877) );
  XOR U5823 ( .A(x[177]), .B(y[177]), .Z(n5874) );
  XNOR U5824 ( .A(x[1148]), .B(y[1148]), .Z(n5875) );
  XNOR U5825 ( .A(n5874), .B(n5875), .Z(n5876) );
  XOR U5826 ( .A(n5877), .B(n5876), .Z(n2844) );
  XOR U5827 ( .A(x[1138]), .B(y[1138]), .Z(n5883) );
  XOR U5828 ( .A(x[183]), .B(y[183]), .Z(n5880) );
  XNOR U5829 ( .A(x[1140]), .B(y[1140]), .Z(n5881) );
  XNOR U5830 ( .A(n5880), .B(n5881), .Z(n5882) );
  XNOR U5831 ( .A(n5883), .B(n5882), .Z(n2843) );
  XNOR U5832 ( .A(n2844), .B(n2843), .Z(n2845) );
  XNOR U5833 ( .A(n2846), .B(n2845), .Z(n1321) );
  XOR U5834 ( .A(x[1134]), .B(y[1134]), .Z(n2708) );
  XOR U5835 ( .A(x[567]), .B(y[567]), .Z(n2705) );
  XNOR U5836 ( .A(x[1136]), .B(y[1136]), .Z(n2706) );
  XNOR U5837 ( .A(n2705), .B(n2706), .Z(n2707) );
  XOR U5838 ( .A(n2708), .B(n2707), .Z(n3356) );
  XOR U5839 ( .A(x[1130]), .B(y[1130]), .Z(n5931) );
  XOR U5840 ( .A(x[1132]), .B(y[1132]), .Z(n5928) );
  XNOR U5841 ( .A(x[1971]), .B(y[1971]), .Z(n5929) );
  XNOR U5842 ( .A(n5928), .B(n5929), .Z(n5930) );
  XOR U5843 ( .A(n5931), .B(n5930), .Z(n3354) );
  XOR U5844 ( .A(x[1126]), .B(y[1126]), .Z(n173) );
  XOR U5845 ( .A(x[189]), .B(y[189]), .Z(n170) );
  XNOR U5846 ( .A(x[1128]), .B(y[1128]), .Z(n171) );
  XNOR U5847 ( .A(n170), .B(n171), .Z(n172) );
  XNOR U5848 ( .A(n173), .B(n172), .Z(n3353) );
  XNOR U5849 ( .A(n3354), .B(n3353), .Z(n3355) );
  XOR U5850 ( .A(n3356), .B(n3355), .Z(n1322) );
  XNOR U5851 ( .A(n1321), .B(n1322), .Z(n1324) );
  XOR U5852 ( .A(x[1122]), .B(y[1122]), .Z(n5919) );
  XOR U5853 ( .A(x[1124]), .B(y[1124]), .Z(n5916) );
  XNOR U5854 ( .A(x[1969]), .B(y[1969]), .Z(n5917) );
  XNOR U5855 ( .A(n5916), .B(n5917), .Z(n5918) );
  XOR U5856 ( .A(n5919), .B(n5918), .Z(n2936) );
  XOR U5857 ( .A(x[1118]), .B(y[1118]), .Z(n301) );
  XOR U5858 ( .A(x[195]), .B(y[195]), .Z(n298) );
  XNOR U5859 ( .A(x[1120]), .B(y[1120]), .Z(n299) );
  XNOR U5860 ( .A(n298), .B(n299), .Z(n300) );
  XOR U5861 ( .A(n301), .B(n300), .Z(n2934) );
  XOR U5862 ( .A(x[1114]), .B(y[1114]), .Z(n5925) );
  XOR U5863 ( .A(x[199]), .B(y[199]), .Z(n5922) );
  XNOR U5864 ( .A(x[1116]), .B(y[1116]), .Z(n5923) );
  XNOR U5865 ( .A(n5922), .B(n5923), .Z(n5924) );
  XNOR U5866 ( .A(n5925), .B(n5924), .Z(n2933) );
  XNOR U5867 ( .A(n2934), .B(n2933), .Z(n2935) );
  XNOR U5868 ( .A(n2936), .B(n2935), .Z(n1323) );
  XNOR U5869 ( .A(n1324), .B(n1323), .Z(n3891) );
  XOR U5870 ( .A(x[1066]), .B(y[1066]), .Z(n5000) );
  XOR U5871 ( .A(x[1068]), .B(y[1068]), .Z(n4998) );
  XNOR U5872 ( .A(x[1963]), .B(y[1963]), .Z(n4999) );
  XOR U5873 ( .A(n4998), .B(n4999), .Z(n5001) );
  XNOR U5874 ( .A(n5000), .B(n5001), .Z(n3768) );
  XOR U5875 ( .A(x[1070]), .B(y[1070]), .Z(n3475) );
  XOR U5876 ( .A(x[607]), .B(y[607]), .Z(n3473) );
  XNOR U5877 ( .A(x[1072]), .B(y[1072]), .Z(n3474) );
  XOR U5878 ( .A(n3473), .B(n3474), .Z(n3476) );
  XOR U5879 ( .A(n3475), .B(n3476), .Z(n3769) );
  XNOR U5880 ( .A(n3768), .B(n3769), .Z(n3771) );
  XOR U5881 ( .A(x[1074]), .B(y[1074]), .Z(n4994) );
  XOR U5882 ( .A(x[227]), .B(y[227]), .Z(n4992) );
  XNOR U5883 ( .A(x[1076]), .B(y[1076]), .Z(n4993) );
  XOR U5884 ( .A(n4992), .B(n4993), .Z(n4995) );
  XNOR U5885 ( .A(n4994), .B(n4995), .Z(n3770) );
  XOR U5886 ( .A(n3771), .B(n3770), .Z(n4375) );
  XOR U5887 ( .A(x[1062]), .B(y[1062]), .Z(n3332) );
  XOR U5888 ( .A(x[233]), .B(y[233]), .Z(n3329) );
  XNOR U5889 ( .A(x[1064]), .B(y[1064]), .Z(n3330) );
  XNOR U5890 ( .A(n3329), .B(n3330), .Z(n3331) );
  XOR U5891 ( .A(n3332), .B(n3331), .Z(n3050) );
  XOR U5892 ( .A(x[1058]), .B(y[1058]), .Z(n5847) );
  XOR U5893 ( .A(x[1060]), .B(y[1060]), .Z(n5844) );
  XNOR U5894 ( .A(x[1961]), .B(y[1961]), .Z(n5845) );
  XNOR U5895 ( .A(n5844), .B(n5845), .Z(n5846) );
  XOR U5896 ( .A(n5847), .B(n5846), .Z(n3048) );
  XOR U5897 ( .A(x[1054]), .B(y[1054]), .Z(n2624) );
  XOR U5898 ( .A(x[239]), .B(y[239]), .Z(n2621) );
  XNOR U5899 ( .A(x[1056]), .B(y[1056]), .Z(n2622) );
  XNOR U5900 ( .A(n2621), .B(n2622), .Z(n2623) );
  XNOR U5901 ( .A(n2624), .B(n2623), .Z(n3047) );
  XNOR U5902 ( .A(n3048), .B(n3047), .Z(n3049) );
  XNOR U5903 ( .A(n3050), .B(n3049), .Z(n4374) );
  XNOR U5904 ( .A(n4375), .B(n4374), .Z(n4377) );
  XOR U5905 ( .A(x[1050]), .B(y[1050]), .Z(n5835) );
  XOR U5906 ( .A(x[243]), .B(y[243]), .Z(n5832) );
  XNOR U5907 ( .A(x[1052]), .B(y[1052]), .Z(n5833) );
  XNOR U5908 ( .A(n5832), .B(n5833), .Z(n5834) );
  XOR U5909 ( .A(n5835), .B(n5834), .Z(n3038) );
  XOR U5910 ( .A(x[1046]), .B(y[1046]), .Z(n3620) );
  XOR U5911 ( .A(x[621]), .B(y[621]), .Z(n3617) );
  XNOR U5912 ( .A(x[1048]), .B(y[1048]), .Z(n3618) );
  XNOR U5913 ( .A(n3617), .B(n3618), .Z(n3619) );
  XOR U5914 ( .A(n3620), .B(n3619), .Z(n3036) );
  XOR U5915 ( .A(x[1042]), .B(y[1042]), .Z(n5433) );
  XOR U5916 ( .A(x[249]), .B(y[249]), .Z(n5430) );
  XNOR U5917 ( .A(x[1044]), .B(y[1044]), .Z(n5431) );
  XNOR U5918 ( .A(n5430), .B(n5431), .Z(n5432) );
  XNOR U5919 ( .A(n5433), .B(n5432), .Z(n3035) );
  XNOR U5920 ( .A(n3036), .B(n3035), .Z(n3037) );
  XNOR U5921 ( .A(n3038), .B(n3037), .Z(n4376) );
  XNOR U5922 ( .A(n4377), .B(n4376), .Z(n3889) );
  XOR U5923 ( .A(x[1110]), .B(y[1110]), .Z(n450) );
  XOR U5924 ( .A(x[581]), .B(y[581]), .Z(n447) );
  XNOR U5925 ( .A(x[1112]), .B(y[1112]), .Z(n448) );
  XNOR U5926 ( .A(n447), .B(n448), .Z(n449) );
  XOR U5927 ( .A(n450), .B(n449), .Z(n3542) );
  XOR U5928 ( .A(x[1106]), .B(y[1106]), .Z(n5025) );
  XOR U5929 ( .A(x[205]), .B(y[205]), .Z(n5022) );
  XNOR U5930 ( .A(x[1108]), .B(y[1108]), .Z(n5023) );
  XNOR U5931 ( .A(n5022), .B(n5023), .Z(n5024) );
  XOR U5932 ( .A(n5025), .B(n5024), .Z(n3540) );
  XOR U5933 ( .A(x[1102]), .B(y[1102]), .Z(n3020) );
  XOR U5934 ( .A(x[587]), .B(y[587]), .Z(n3017) );
  XNOR U5935 ( .A(x[1104]), .B(y[1104]), .Z(n3018) );
  XNOR U5936 ( .A(n3017), .B(n3018), .Z(n3019) );
  XNOR U5937 ( .A(n3020), .B(n3019), .Z(n3539) );
  XNOR U5938 ( .A(n3540), .B(n3539), .Z(n3541) );
  XNOR U5939 ( .A(n3542), .B(n3541), .Z(n1225) );
  XOR U5940 ( .A(x[1098]), .B(y[1098]), .Z(n5013) );
  XOR U5941 ( .A(x[1100]), .B(y[1100]), .Z(n5010) );
  XNOR U5942 ( .A(x[1967]), .B(y[1967]), .Z(n5011) );
  XNOR U5943 ( .A(n5010), .B(n5011), .Z(n5012) );
  XOR U5944 ( .A(n5013), .B(n5012), .Z(n3584) );
  XOR U5945 ( .A(x[1094]), .B(y[1094]), .Z(n2996) );
  XOR U5946 ( .A(x[211]), .B(y[211]), .Z(n2993) );
  XNOR U5947 ( .A(x[1096]), .B(y[1096]), .Z(n2994) );
  XNOR U5948 ( .A(n2993), .B(n2994), .Z(n2995) );
  XOR U5949 ( .A(n2996), .B(n2995), .Z(n3582) );
  XOR U5950 ( .A(x[1090]), .B(y[1090]), .Z(n5019) );
  XOR U5951 ( .A(x[1092]), .B(y[1092]), .Z(n5016) );
  XNOR U5952 ( .A(x[1965]), .B(y[1965]), .Z(n5017) );
  XNOR U5953 ( .A(n5016), .B(n5017), .Z(n5018) );
  XNOR U5954 ( .A(n5019), .B(n5018), .Z(n3581) );
  XNOR U5955 ( .A(n3582), .B(n3581), .Z(n3583) );
  XOR U5956 ( .A(n3584), .B(n3583), .Z(n1226) );
  XNOR U5957 ( .A(n1225), .B(n1226), .Z(n1228) );
  XOR U5958 ( .A(x[1086]), .B(y[1086]), .Z(n432) );
  XOR U5959 ( .A(x[217]), .B(y[217]), .Z(n429) );
  XNOR U5960 ( .A(x[1088]), .B(y[1088]), .Z(n430) );
  XNOR U5961 ( .A(n429), .B(n430), .Z(n431) );
  XOR U5962 ( .A(n432), .B(n431), .Z(n3572) );
  XOR U5963 ( .A(x[1082]), .B(y[1082]), .Z(n5007) );
  XOR U5964 ( .A(x[221]), .B(y[221]), .Z(n5004) );
  XNOR U5965 ( .A(x[1084]), .B(y[1084]), .Z(n5005) );
  XNOR U5966 ( .A(n5004), .B(n5005), .Z(n5006) );
  XOR U5967 ( .A(n5007), .B(n5006), .Z(n3570) );
  XOR U5968 ( .A(x[1078]), .B(y[1078]), .Z(n3717) );
  XOR U5969 ( .A(x[601]), .B(y[601]), .Z(n3714) );
  XNOR U5970 ( .A(x[1080]), .B(y[1080]), .Z(n3715) );
  XNOR U5971 ( .A(n3714), .B(n3715), .Z(n3716) );
  XNOR U5972 ( .A(n3717), .B(n3716), .Z(n3569) );
  XNOR U5973 ( .A(n3570), .B(n3569), .Z(n3571) );
  XNOR U5974 ( .A(n3572), .B(n3571), .Z(n1227) );
  XNOR U5975 ( .A(n1228), .B(n1227), .Z(n3888) );
  XOR U5976 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U5977 ( .A(n3891), .B(n3890), .Z(n3810) );
  XOR U5978 ( .A(x[1006]), .B(y[1006]), .Z(n4916) );
  XOR U5979 ( .A(x[647]), .B(y[647]), .Z(n4914) );
  XNOR U5980 ( .A(x[1008]), .B(y[1008]), .Z(n4915) );
  XOR U5981 ( .A(n4914), .B(n4915), .Z(n4917) );
  XNOR U5982 ( .A(n4916), .B(n4917), .Z(n259) );
  XOR U5983 ( .A(x[1010]), .B(y[1010]), .Z(n4641) );
  XOR U5984 ( .A(x[271]), .B(y[271]), .Z(n4639) );
  XOR U5985 ( .A(x[1012]), .B(y[1012]), .Z(n4638) );
  XOR U5986 ( .A(n4639), .B(n4638), .Z(n4640) );
  XOR U5987 ( .A(n4641), .B(n4640), .Z(n258) );
  XOR U5988 ( .A(n259), .B(n258), .Z(n261) );
  XOR U5989 ( .A(x[1014]), .B(y[1014]), .Z(n3313) );
  XOR U5990 ( .A(x[641]), .B(y[641]), .Z(n3311) );
  XNOR U5991 ( .A(x[1016]), .B(y[1016]), .Z(n3312) );
  XOR U5992 ( .A(n3311), .B(n3312), .Z(n3314) );
  XNOR U5993 ( .A(n3313), .B(n3314), .Z(n260) );
  XOR U5994 ( .A(n261), .B(n260), .Z(n1166) );
  XOR U5995 ( .A(x[1038]), .B(y[1038]), .Z(n277) );
  XOR U5996 ( .A(x[627]), .B(y[627]), .Z(n274) );
  XNOR U5997 ( .A(x[1040]), .B(y[1040]), .Z(n275) );
  XNOR U5998 ( .A(n274), .B(n275), .Z(n276) );
  XOR U5999 ( .A(n277), .B(n276), .Z(n3098) );
  XOR U6000 ( .A(x[1034]), .B(y[1034]), .Z(n5841) );
  XOR U6001 ( .A(x[1036]), .B(y[1036]), .Z(n5838) );
  XNOR U6002 ( .A(x[1959]), .B(y[1959]), .Z(n5839) );
  XNOR U6003 ( .A(n5838), .B(n5839), .Z(n5840) );
  XOR U6004 ( .A(n5841), .B(n5840), .Z(n3096) );
  XOR U6005 ( .A(x[1030]), .B(y[1030]), .Z(n3248) );
  XOR U6006 ( .A(x[255]), .B(y[255]), .Z(n3245) );
  XNOR U6007 ( .A(x[1032]), .B(y[1032]), .Z(n3246) );
  XNOR U6008 ( .A(n3245), .B(n3246), .Z(n3247) );
  XNOR U6009 ( .A(n3248), .B(n3247), .Z(n3095) );
  XNOR U6010 ( .A(n3096), .B(n3095), .Z(n3097) );
  XNOR U6011 ( .A(n3098), .B(n3097), .Z(n1165) );
  XNOR U6012 ( .A(n1166), .B(n1165), .Z(n1167) );
  XOR U6013 ( .A(x[1026]), .B(y[1026]), .Z(n3458) );
  XOR U6014 ( .A(x[1028]), .B(y[1028]), .Z(n3455) );
  XNOR U6015 ( .A(x[1957]), .B(y[1957]), .Z(n3456) );
  XNOR U6016 ( .A(n3455), .B(n3456), .Z(n3457) );
  XOR U6017 ( .A(n3458), .B(n3457), .Z(n3086) );
  XOR U6018 ( .A(x[1022]), .B(y[1022]), .Z(n4653) );
  XOR U6019 ( .A(x[261]), .B(y[261]), .Z(n4650) );
  XNOR U6020 ( .A(x[1024]), .B(y[1024]), .Z(n4651) );
  XNOR U6021 ( .A(n4650), .B(n4651), .Z(n4652) );
  XOR U6022 ( .A(n4653), .B(n4652), .Z(n3084) );
  XOR U6023 ( .A(x[1018]), .B(y[1018]), .Z(n4611) );
  XOR U6024 ( .A(x[265]), .B(y[265]), .Z(n4608) );
  XNOR U6025 ( .A(x[1020]), .B(y[1020]), .Z(n4609) );
  XNOR U6026 ( .A(n4608), .B(n4609), .Z(n4610) );
  XNOR U6027 ( .A(n4611), .B(n4610), .Z(n3083) );
  XNOR U6028 ( .A(n3084), .B(n3083), .Z(n3085) );
  XOR U6029 ( .A(n3086), .B(n3085), .Z(n1168) );
  XNOR U6030 ( .A(n1167), .B(n1168), .Z(n3819) );
  XOR U6031 ( .A(x[946]), .B(y[946]), .Z(n4185) );
  XOR U6032 ( .A(x[309]), .B(y[309]), .Z(n4182) );
  XNOR U6033 ( .A(x[948]), .B(y[948]), .Z(n4183) );
  XNOR U6034 ( .A(n4182), .B(n4183), .Z(n4184) );
  XOR U6035 ( .A(n4185), .B(n4184), .Z(n4863) );
  XOR U6036 ( .A(x[942]), .B(y[942]), .Z(n1838) );
  XOR U6037 ( .A(x[681]), .B(y[681]), .Z(n1836) );
  XOR U6038 ( .A(x[944]), .B(y[944]), .Z(n1835) );
  XOR U6039 ( .A(n1836), .B(n1835), .Z(n1837) );
  XOR U6040 ( .A(n1838), .B(n1837), .Z(n4861) );
  XOR U6041 ( .A(x[938]), .B(y[938]), .Z(n1832) );
  XOR U6042 ( .A(x[315]), .B(y[315]), .Z(n1830) );
  XOR U6043 ( .A(x[940]), .B(y[940]), .Z(n1829) );
  XOR U6044 ( .A(n1830), .B(n1829), .Z(n1831) );
  XNOR U6045 ( .A(n1832), .B(n1831), .Z(n4860) );
  XNOR U6046 ( .A(n4861), .B(n4860), .Z(n4862) );
  XNOR U6047 ( .A(n4863), .B(n4862), .Z(n4308) );
  XOR U6048 ( .A(x[962]), .B(y[962]), .Z(n2738) );
  XOR U6049 ( .A(x[299]), .B(y[299]), .Z(n2736) );
  XOR U6050 ( .A(x[964]), .B(y[964]), .Z(n2735) );
  XOR U6051 ( .A(n2736), .B(n2735), .Z(n2737) );
  XOR U6052 ( .A(n2738), .B(n2737), .Z(n4839) );
  XOR U6053 ( .A(x[958]), .B(y[958]), .Z(n1510) );
  XOR U6054 ( .A(x[960]), .B(y[960]), .Z(n1507) );
  XNOR U6055 ( .A(x[1949]), .B(y[1949]), .Z(n1508) );
  XNOR U6056 ( .A(n1507), .B(n1508), .Z(n1509) );
  XOR U6057 ( .A(n1510), .B(n1509), .Z(n4837) );
  XOR U6058 ( .A(x[952]), .B(y[952]), .Z(n1504) );
  XOR U6059 ( .A(x[305]), .B(y[305]), .Z(n1501) );
  XNOR U6060 ( .A(x[956]), .B(y[956]), .Z(n1502) );
  XNOR U6061 ( .A(n1501), .B(n1502), .Z(n1503) );
  XNOR U6062 ( .A(n1504), .B(n1503), .Z(n4836) );
  XNOR U6063 ( .A(n4837), .B(n4836), .Z(n4838) );
  XOR U6064 ( .A(n4839), .B(n4838), .Z(n4309) );
  XNOR U6065 ( .A(n4308), .B(n4309), .Z(n4310) );
  XOR U6066 ( .A(x[932]), .B(y[932]), .Z(n1594) );
  XOR U6067 ( .A(x[687]), .B(y[687]), .Z(n1591) );
  XNOR U6068 ( .A(x[934]), .B(y[934]), .Z(n1592) );
  XNOR U6069 ( .A(n1591), .B(n1592), .Z(n1593) );
  XOR U6070 ( .A(n1594), .B(n1593), .Z(n5079) );
  XOR U6071 ( .A(x[928]), .B(y[928]), .Z(n1618) );
  XOR U6072 ( .A(x[930]), .B(y[930]), .Z(n1615) );
  XNOR U6073 ( .A(x[1947]), .B(y[1947]), .Z(n1616) );
  XNOR U6074 ( .A(n1615), .B(n1616), .Z(n1617) );
  XOR U6075 ( .A(n1618), .B(n1617), .Z(n5077) );
  XOR U6076 ( .A(x[924]), .B(y[924]), .Z(n1648) );
  XOR U6077 ( .A(x[321]), .B(y[321]), .Z(n1645) );
  XNOR U6078 ( .A(x[926]), .B(y[926]), .Z(n1646) );
  XNOR U6079 ( .A(n1645), .B(n1646), .Z(n1647) );
  XNOR U6080 ( .A(n1648), .B(n1647), .Z(n5076) );
  XNOR U6081 ( .A(n5077), .B(n5076), .Z(n5078) );
  XOR U6082 ( .A(n5079), .B(n5078), .Z(n4311) );
  XNOR U6083 ( .A(n4310), .B(n4311), .Z(n3816) );
  XOR U6084 ( .A(x[994]), .B(y[994]), .Z(n5631) );
  XOR U6085 ( .A(x[996]), .B(y[996]), .Z(n5629) );
  XOR U6086 ( .A(x[1953]), .B(y[1953]), .Z(n5628) );
  XOR U6087 ( .A(n5629), .B(n5628), .Z(n5630) );
  XOR U6088 ( .A(n5631), .B(n5630), .Z(n255) );
  XOR U6089 ( .A(x[998]), .B(y[998]), .Z(n4647) );
  XOR U6090 ( .A(x[277]), .B(y[277]), .Z(n4645) );
  XOR U6091 ( .A(x[1000]), .B(y[1000]), .Z(n4644) );
  XOR U6092 ( .A(n4645), .B(n4644), .Z(n4646) );
  XOR U6093 ( .A(n4647), .B(n4646), .Z(n254) );
  XOR U6094 ( .A(n255), .B(n254), .Z(n257) );
  XOR U6095 ( .A(x[1002]), .B(y[1002]), .Z(n3428) );
  XOR U6096 ( .A(x[1004]), .B(y[1004]), .Z(n3426) );
  XOR U6097 ( .A(x[1955]), .B(y[1955]), .Z(n3425) );
  XOR U6098 ( .A(n3426), .B(n3425), .Z(n3427) );
  XOR U6099 ( .A(n3428), .B(n3427), .Z(n256) );
  XOR U6100 ( .A(n257), .B(n256), .Z(n4435) );
  XOR U6101 ( .A(x[988]), .B(y[988]), .Z(n5619) );
  XOR U6102 ( .A(x[283]), .B(y[283]), .Z(n5616) );
  XNOR U6103 ( .A(x[990]), .B(y[990]), .Z(n5617) );
  XNOR U6104 ( .A(n5616), .B(n5617), .Z(n5618) );
  XOR U6105 ( .A(n5619), .B(n5618), .Z(n6015) );
  XOR U6106 ( .A(x[984]), .B(y[984]), .Z(n5625) );
  XOR U6107 ( .A(x[287]), .B(y[287]), .Z(n5622) );
  XNOR U6108 ( .A(x[986]), .B(y[986]), .Z(n5623) );
  XNOR U6109 ( .A(n5622), .B(n5623), .Z(n5624) );
  XOR U6110 ( .A(n5625), .B(n5624), .Z(n6013) );
  XOR U6111 ( .A(x[980]), .B(y[980]), .Z(n5613) );
  XOR U6112 ( .A(x[661]), .B(y[661]), .Z(n5610) );
  XNOR U6113 ( .A(x[982]), .B(y[982]), .Z(n5611) );
  XNOR U6114 ( .A(n5610), .B(n5611), .Z(n5612) );
  XNOR U6115 ( .A(n5613), .B(n5612), .Z(n6012) );
  XNOR U6116 ( .A(n6013), .B(n6012), .Z(n6014) );
  XNOR U6117 ( .A(n6015), .B(n6014), .Z(n4434) );
  XNOR U6118 ( .A(n4435), .B(n4434), .Z(n4436) );
  XOR U6119 ( .A(x[976]), .B(y[976]), .Z(n5601) );
  XOR U6120 ( .A(x[293]), .B(y[293]), .Z(n5599) );
  XOR U6121 ( .A(x[978]), .B(y[978]), .Z(n5598) );
  XOR U6122 ( .A(n5599), .B(n5598), .Z(n5600) );
  XOR U6123 ( .A(n5601), .B(n5600), .Z(n4935) );
  XOR U6124 ( .A(x[972]), .B(y[972]), .Z(n5607) );
  XOR U6125 ( .A(x[667]), .B(y[667]), .Z(n5605) );
  XOR U6126 ( .A(x[974]), .B(y[974]), .Z(n5604) );
  XOR U6127 ( .A(n5605), .B(n5604), .Z(n5606) );
  XOR U6128 ( .A(n5607), .B(n5606), .Z(n4933) );
  XOR U6129 ( .A(x[968]), .B(y[968]), .Z(n3302) );
  XOR U6130 ( .A(x[970]), .B(y[970]), .Z(n3300) );
  XOR U6131 ( .A(x[1951]), .B(y[1951]), .Z(n3299) );
  XOR U6132 ( .A(n3300), .B(n3299), .Z(n3301) );
  XNOR U6133 ( .A(n3302), .B(n3301), .Z(n4932) );
  XNOR U6134 ( .A(n4933), .B(n4932), .Z(n4934) );
  XOR U6135 ( .A(n4935), .B(n4934), .Z(n4437) );
  XNOR U6136 ( .A(n4436), .B(n4437), .Z(n3817) );
  XOR U6137 ( .A(n3816), .B(n3817), .Z(n3818) );
  XOR U6138 ( .A(n3819), .B(n3818), .Z(n3811) );
  XOR U6139 ( .A(n3810), .B(n3811), .Z(n3813) );
  XNOR U6140 ( .A(n3812), .B(n3813), .Z(n3798) );
  XOR U6141 ( .A(n3799), .B(n3798), .Z(n3800) );
  XNOR U6142 ( .A(n3801), .B(n3800), .Z(n3900) );
  XNOR U6143 ( .A(n3901), .B(n3900), .Z(n3902) );
  XOR U6144 ( .A(n3903), .B(n3902), .Z(o[0]) );
  NANDN U6145 ( .A(n81), .B(n80), .Z(n85) );
  NAND U6146 ( .A(n83), .B(n82), .Z(n84) );
  AND U6147 ( .A(n85), .B(n84), .Z(n7480) );
  NANDN U6148 ( .A(n87), .B(n86), .Z(n91) );
  NAND U6149 ( .A(n89), .B(n88), .Z(n90) );
  NAND U6150 ( .A(n91), .B(n90), .Z(n7481) );
  XNOR U6151 ( .A(n7480), .B(n7481), .Z(n7483) );
  NANDN U6152 ( .A(n93), .B(n92), .Z(n97) );
  NAND U6153 ( .A(n95), .B(n94), .Z(n96) );
  AND U6154 ( .A(n97), .B(n96), .Z(n7482) );
  XOR U6155 ( .A(n7483), .B(n7482), .Z(n6602) );
  NANDN U6156 ( .A(n99), .B(n98), .Z(n103) );
  NAND U6157 ( .A(n101), .B(n100), .Z(n102) );
  AND U6158 ( .A(n103), .B(n102), .Z(n9009) );
  NANDN U6159 ( .A(n105), .B(n104), .Z(n109) );
  NAND U6160 ( .A(n107), .B(n106), .Z(n108) );
  NAND U6161 ( .A(n109), .B(n108), .Z(n9010) );
  XNOR U6162 ( .A(n9009), .B(n9010), .Z(n9012) );
  NANDN U6163 ( .A(n111), .B(n110), .Z(n115) );
  NAND U6164 ( .A(n113), .B(n112), .Z(n114) );
  AND U6165 ( .A(n115), .B(n114), .Z(n9011) );
  XOR U6166 ( .A(n9012), .B(n9011), .Z(n6601) );
  NANDN U6167 ( .A(n117), .B(n116), .Z(n121) );
  NANDN U6168 ( .A(n119), .B(n118), .Z(n120) );
  AND U6169 ( .A(n121), .B(n120), .Z(n6600) );
  XOR U6170 ( .A(n6601), .B(n6600), .Z(n6603) );
  XOR U6171 ( .A(n6602), .B(n6603), .Z(n7189) );
  NANDN U6172 ( .A(n123), .B(n122), .Z(n127) );
  NANDN U6173 ( .A(n125), .B(n124), .Z(n126) );
  AND U6174 ( .A(n127), .B(n126), .Z(n6913) );
  NANDN U6175 ( .A(n129), .B(n128), .Z(n133) );
  NAND U6176 ( .A(n131), .B(n130), .Z(n132) );
  AND U6177 ( .A(n133), .B(n132), .Z(n8613) );
  NANDN U6178 ( .A(n135), .B(n134), .Z(n139) );
  NAND U6179 ( .A(n137), .B(n136), .Z(n138) );
  NAND U6180 ( .A(n139), .B(n138), .Z(n8614) );
  XNOR U6181 ( .A(n8613), .B(n8614), .Z(n8616) );
  NANDN U6182 ( .A(n141), .B(n140), .Z(n145) );
  NAND U6183 ( .A(n143), .B(n142), .Z(n144) );
  AND U6184 ( .A(n145), .B(n144), .Z(n8615) );
  XOR U6185 ( .A(n8616), .B(n8615), .Z(n6911) );
  NANDN U6186 ( .A(n147), .B(n146), .Z(n151) );
  NANDN U6187 ( .A(n149), .B(n148), .Z(n150) );
  AND U6188 ( .A(n151), .B(n150), .Z(n6910) );
  XNOR U6189 ( .A(n6911), .B(n6910), .Z(n6912) );
  XOR U6190 ( .A(n6913), .B(n6912), .Z(n7187) );
  NANDN U6191 ( .A(n153), .B(n152), .Z(n157) );
  NANDN U6192 ( .A(n155), .B(n154), .Z(n156) );
  AND U6193 ( .A(n157), .B(n156), .Z(n7588) );
  NANDN U6194 ( .A(n159), .B(n158), .Z(n163) );
  NAND U6195 ( .A(n161), .B(n160), .Z(n162) );
  NAND U6196 ( .A(n163), .B(n162), .Z(n7589) );
  XNOR U6197 ( .A(n7588), .B(n7589), .Z(n7591) );
  NANDN U6198 ( .A(n165), .B(n164), .Z(n169) );
  NAND U6199 ( .A(n167), .B(n166), .Z(n168) );
  AND U6200 ( .A(n169), .B(n168), .Z(n7590) );
  XOR U6201 ( .A(n7591), .B(n7590), .Z(n6608) );
  NANDN U6202 ( .A(n171), .B(n170), .Z(n175) );
  NAND U6203 ( .A(n173), .B(n172), .Z(n174) );
  AND U6204 ( .A(n175), .B(n174), .Z(n8337) );
  NANDN U6205 ( .A(n177), .B(n176), .Z(n181) );
  NAND U6206 ( .A(n179), .B(n178), .Z(n180) );
  NAND U6207 ( .A(n181), .B(n180), .Z(n8338) );
  XNOR U6208 ( .A(n8337), .B(n8338), .Z(n8340) );
  NANDN U6209 ( .A(n183), .B(n182), .Z(n187) );
  NAND U6210 ( .A(n185), .B(n184), .Z(n186) );
  AND U6211 ( .A(n187), .B(n186), .Z(n8339) );
  XOR U6212 ( .A(n8340), .B(n8339), .Z(n6607) );
  NANDN U6213 ( .A(n189), .B(n188), .Z(n193) );
  NANDN U6214 ( .A(n191), .B(n190), .Z(n192) );
  AND U6215 ( .A(n193), .B(n192), .Z(n6606) );
  XOR U6216 ( .A(n6607), .B(n6606), .Z(n6609) );
  XNOR U6217 ( .A(n6608), .B(n6609), .Z(n7186) );
  XNOR U6218 ( .A(n7187), .B(n7186), .Z(n7188) );
  XNOR U6219 ( .A(n7189), .B(n7188), .Z(n6117) );
  NANDN U6220 ( .A(n195), .B(n194), .Z(n199) );
  NAND U6221 ( .A(n197), .B(n196), .Z(n198) );
  AND U6222 ( .A(n199), .B(n198), .Z(n6384) );
  NANDN U6223 ( .A(n201), .B(n200), .Z(n205) );
  NAND U6224 ( .A(n203), .B(n202), .Z(n204) );
  NAND U6225 ( .A(n205), .B(n204), .Z(n6385) );
  XNOR U6226 ( .A(n6384), .B(n6385), .Z(n6387) );
  NANDN U6227 ( .A(n207), .B(n206), .Z(n211) );
  NAND U6228 ( .A(n209), .B(n208), .Z(n210) );
  AND U6229 ( .A(n211), .B(n210), .Z(n6386) );
  XOR U6230 ( .A(n6387), .B(n6386), .Z(n7213) );
  NANDN U6231 ( .A(n213), .B(n212), .Z(n217) );
  NAND U6232 ( .A(n215), .B(n214), .Z(n216) );
  AND U6233 ( .A(n217), .B(n216), .Z(n7211) );
  NANDN U6234 ( .A(n219), .B(n218), .Z(n223) );
  NANDN U6235 ( .A(n221), .B(n220), .Z(n222) );
  AND U6236 ( .A(n223), .B(n222), .Z(n7210) );
  XNOR U6237 ( .A(n7211), .B(n7210), .Z(n7212) );
  XNOR U6238 ( .A(n7213), .B(n7212), .Z(n7156) );
  NANDN U6239 ( .A(n225), .B(n224), .Z(n229) );
  NANDN U6240 ( .A(n227), .B(n226), .Z(n228) );
  AND U6241 ( .A(n229), .B(n228), .Z(n7105) );
  NANDN U6242 ( .A(n231), .B(n230), .Z(n235) );
  NAND U6243 ( .A(n233), .B(n232), .Z(n234) );
  AND U6244 ( .A(n235), .B(n234), .Z(n7103) );
  NANDN U6245 ( .A(n237), .B(n236), .Z(n241) );
  NAND U6246 ( .A(n239), .B(n238), .Z(n240) );
  AND U6247 ( .A(n241), .B(n240), .Z(n6372) );
  NANDN U6248 ( .A(n243), .B(n242), .Z(n247) );
  NAND U6249 ( .A(n245), .B(n244), .Z(n246) );
  NAND U6250 ( .A(n247), .B(n246), .Z(n6373) );
  XNOR U6251 ( .A(n6372), .B(n6373), .Z(n6375) );
  NANDN U6252 ( .A(n249), .B(n248), .Z(n253) );
  NAND U6253 ( .A(n251), .B(n250), .Z(n252) );
  AND U6254 ( .A(n253), .B(n252), .Z(n6374) );
  XNOR U6255 ( .A(n6375), .B(n6374), .Z(n7102) );
  XNOR U6256 ( .A(n7103), .B(n7102), .Z(n7104) );
  XOR U6257 ( .A(n7105), .B(n7104), .Z(n7157) );
  XNOR U6258 ( .A(n7156), .B(n7157), .Z(n7159) );
  NANDN U6259 ( .A(n263), .B(n262), .Z(n267) );
  NANDN U6260 ( .A(n265), .B(n264), .Z(n266) );
  AND U6261 ( .A(n267), .B(n266), .Z(n8469) );
  XNOR U6262 ( .A(n8470), .B(n8469), .Z(n8471) );
  XNOR U6263 ( .A(n8472), .B(n8471), .Z(n7158) );
  XNOR U6264 ( .A(n7159), .B(n7158), .Z(n6115) );
  NANDN U6265 ( .A(n269), .B(n268), .Z(n273) );
  NAND U6266 ( .A(n271), .B(n270), .Z(n272) );
  AND U6267 ( .A(n273), .B(n272), .Z(n7162) );
  NANDN U6268 ( .A(n275), .B(n274), .Z(n279) );
  NAND U6269 ( .A(n277), .B(n276), .Z(n278) );
  AND U6270 ( .A(n279), .B(n278), .Z(n7600) );
  NANDN U6271 ( .A(n281), .B(n280), .Z(n285) );
  NAND U6272 ( .A(n283), .B(n282), .Z(n284) );
  NAND U6273 ( .A(n285), .B(n284), .Z(n7601) );
  XNOR U6274 ( .A(n7600), .B(n7601), .Z(n7603) );
  NANDN U6275 ( .A(n287), .B(n286), .Z(n291) );
  NAND U6276 ( .A(n289), .B(n288), .Z(n290) );
  AND U6277 ( .A(n291), .B(n290), .Z(n7602) );
  XOR U6278 ( .A(n7603), .B(n7602), .Z(n8292) );
  NANDN U6279 ( .A(n293), .B(n292), .Z(n297) );
  NAND U6280 ( .A(n295), .B(n294), .Z(n296) );
  AND U6281 ( .A(n297), .B(n296), .Z(n8290) );
  NANDN U6282 ( .A(n299), .B(n298), .Z(n303) );
  NAND U6283 ( .A(n301), .B(n300), .Z(n302) );
  AND U6284 ( .A(n303), .B(n302), .Z(n8703) );
  NANDN U6285 ( .A(n305), .B(n304), .Z(n309) );
  NANDN U6286 ( .A(n307), .B(n306), .Z(n308) );
  NAND U6287 ( .A(n309), .B(n308), .Z(n8704) );
  XNOR U6288 ( .A(n8703), .B(n8704), .Z(n8706) );
  NANDN U6289 ( .A(n311), .B(n310), .Z(n315) );
  NANDN U6290 ( .A(n313), .B(n312), .Z(n314) );
  AND U6291 ( .A(n315), .B(n314), .Z(n8705) );
  XNOR U6292 ( .A(n8706), .B(n8705), .Z(n8289) );
  XNOR U6293 ( .A(n8290), .B(n8289), .Z(n8291) );
  XOR U6294 ( .A(n8292), .B(n8291), .Z(n7163) );
  XNOR U6295 ( .A(n7162), .B(n7163), .Z(n7165) );
  NANDN U6296 ( .A(n317), .B(n316), .Z(n321) );
  NAND U6297 ( .A(n319), .B(n318), .Z(n320) );
  AND U6298 ( .A(n321), .B(n320), .Z(n7606) );
  NANDN U6299 ( .A(n323), .B(n322), .Z(n327) );
  NAND U6300 ( .A(n325), .B(n324), .Z(n326) );
  NAND U6301 ( .A(n327), .B(n326), .Z(n7607) );
  XNOR U6302 ( .A(n7606), .B(n7607), .Z(n7609) );
  NANDN U6303 ( .A(n329), .B(n328), .Z(n333) );
  NAND U6304 ( .A(n331), .B(n330), .Z(n332) );
  AND U6305 ( .A(n333), .B(n332), .Z(n7608) );
  XOR U6306 ( .A(n7609), .B(n7608), .Z(n8286) );
  NANDN U6307 ( .A(n335), .B(n334), .Z(n339) );
  NAND U6308 ( .A(n337), .B(n336), .Z(n338) );
  AND U6309 ( .A(n339), .B(n338), .Z(n8284) );
  NANDN U6310 ( .A(n341), .B(n340), .Z(n345) );
  NAND U6311 ( .A(n343), .B(n342), .Z(n344) );
  AND U6312 ( .A(n345), .B(n344), .Z(n8685) );
  NANDN U6313 ( .A(n347), .B(n346), .Z(n351) );
  NAND U6314 ( .A(n349), .B(n348), .Z(n350) );
  NAND U6315 ( .A(n351), .B(n350), .Z(n8686) );
  XNOR U6316 ( .A(n8685), .B(n8686), .Z(n8688) );
  NANDN U6317 ( .A(n353), .B(n352), .Z(n357) );
  NAND U6318 ( .A(n355), .B(n354), .Z(n356) );
  AND U6319 ( .A(n357), .B(n356), .Z(n8687) );
  XNOR U6320 ( .A(n8688), .B(n8687), .Z(n8283) );
  XNOR U6321 ( .A(n8284), .B(n8283), .Z(n8285) );
  XNOR U6322 ( .A(n8286), .B(n8285), .Z(n7164) );
  XNOR U6323 ( .A(n7165), .B(n7164), .Z(n6114) );
  XOR U6324 ( .A(n6115), .B(n6114), .Z(n6116) );
  XNOR U6325 ( .A(n6117), .B(n6116), .Z(n8640) );
  NANDN U6326 ( .A(n359), .B(n358), .Z(n363) );
  NAND U6327 ( .A(n361), .B(n360), .Z(n362) );
  AND U6328 ( .A(n363), .B(n362), .Z(n7564) );
  NANDN U6329 ( .A(n365), .B(n364), .Z(n369) );
  NAND U6330 ( .A(n367), .B(n366), .Z(n368) );
  NAND U6331 ( .A(n369), .B(n368), .Z(n7565) );
  XNOR U6332 ( .A(n7564), .B(n7565), .Z(n7567) );
  NANDN U6333 ( .A(n370), .B(oglobal[0]), .Z(n374) );
  NAND U6334 ( .A(n372), .B(n371), .Z(n373) );
  AND U6335 ( .A(n374), .B(n373), .Z(n7566) );
  XOR U6336 ( .A(n7567), .B(n7566), .Z(n8789) );
  NANDN U6337 ( .A(n376), .B(n375), .Z(n380) );
  NAND U6338 ( .A(n378), .B(n377), .Z(n379) );
  AND U6339 ( .A(n380), .B(n379), .Z(n8319) );
  NANDN U6340 ( .A(n382), .B(n381), .Z(n386) );
  NANDN U6341 ( .A(n384), .B(n383), .Z(n385) );
  NAND U6342 ( .A(n386), .B(n385), .Z(n8320) );
  XNOR U6343 ( .A(n8319), .B(n8320), .Z(n8322) );
  NANDN U6344 ( .A(n388), .B(n387), .Z(n392) );
  NANDN U6345 ( .A(n390), .B(n389), .Z(n391) );
  AND U6346 ( .A(n392), .B(n391), .Z(n8321) );
  XOR U6347 ( .A(n8322), .B(n8321), .Z(n8788) );
  NANDN U6348 ( .A(n394), .B(n393), .Z(n398) );
  NANDN U6349 ( .A(n396), .B(n395), .Z(n397) );
  AND U6350 ( .A(n398), .B(n397), .Z(n8787) );
  XOR U6351 ( .A(n8788), .B(n8787), .Z(n8790) );
  XOR U6352 ( .A(n8789), .B(n8790), .Z(n7069) );
  NAND U6353 ( .A(n400), .B(n399), .Z(n404) );
  NAND U6354 ( .A(n402), .B(n401), .Z(n403) );
  AND U6355 ( .A(n404), .B(n403), .Z(n7087) );
  NANDN U6356 ( .A(n406), .B(n405), .Z(n410) );
  NAND U6357 ( .A(n408), .B(n407), .Z(n409) );
  AND U6358 ( .A(n410), .B(n409), .Z(n6378) );
  NANDN U6359 ( .A(n412), .B(n411), .Z(n416) );
  NAND U6360 ( .A(n414), .B(n413), .Z(n415) );
  NAND U6361 ( .A(n416), .B(n415), .Z(n6379) );
  XNOR U6362 ( .A(n6378), .B(n6379), .Z(n6381) );
  NANDN U6363 ( .A(n418), .B(n417), .Z(n422) );
  NAND U6364 ( .A(n420), .B(n419), .Z(n421) );
  AND U6365 ( .A(n422), .B(n421), .Z(n6380) );
  XOR U6366 ( .A(n6381), .B(n6380), .Z(n7085) );
  NAND U6367 ( .A(n424), .B(n423), .Z(n428) );
  NAND U6368 ( .A(n426), .B(n425), .Z(n427) );
  AND U6369 ( .A(n428), .B(n427), .Z(n7084) );
  XNOR U6370 ( .A(n7085), .B(n7084), .Z(n7086) );
  XOR U6371 ( .A(n7087), .B(n7086), .Z(n7067) );
  NANDN U6372 ( .A(n430), .B(n429), .Z(n434) );
  NAND U6373 ( .A(n432), .B(n431), .Z(n433) );
  AND U6374 ( .A(n434), .B(n433), .Z(n6360) );
  NANDN U6375 ( .A(n436), .B(n435), .Z(n440) );
  NAND U6376 ( .A(n438), .B(n437), .Z(n439) );
  NAND U6377 ( .A(n440), .B(n439), .Z(n6361) );
  XNOR U6378 ( .A(n6360), .B(n6361), .Z(n6363) );
  NANDN U6379 ( .A(n442), .B(n441), .Z(n446) );
  NAND U6380 ( .A(n444), .B(n443), .Z(n445) );
  AND U6381 ( .A(n446), .B(n445), .Z(n6362) );
  XOR U6382 ( .A(n6363), .B(n6362), .Z(n8783) );
  NANDN U6383 ( .A(n448), .B(n447), .Z(n452) );
  NAND U6384 ( .A(n450), .B(n449), .Z(n451) );
  AND U6385 ( .A(n452), .B(n451), .Z(n8541) );
  NANDN U6386 ( .A(n454), .B(n453), .Z(n458) );
  NANDN U6387 ( .A(n456), .B(n455), .Z(n457) );
  NAND U6388 ( .A(n458), .B(n457), .Z(n8542) );
  XNOR U6389 ( .A(n8541), .B(n8542), .Z(n8544) );
  NANDN U6390 ( .A(n460), .B(n459), .Z(n464) );
  NANDN U6391 ( .A(n462), .B(n461), .Z(n463) );
  AND U6392 ( .A(n464), .B(n463), .Z(n8543) );
  XOR U6393 ( .A(n8544), .B(n8543), .Z(n8782) );
  NANDN U6394 ( .A(n466), .B(n465), .Z(n470) );
  NANDN U6395 ( .A(n468), .B(n467), .Z(n469) );
  AND U6396 ( .A(n470), .B(n469), .Z(n8781) );
  XOR U6397 ( .A(n8782), .B(n8781), .Z(n8784) );
  XNOR U6398 ( .A(n8783), .B(n8784), .Z(n7066) );
  XNOR U6399 ( .A(n7067), .B(n7066), .Z(n7068) );
  XNOR U6400 ( .A(n7069), .B(n7068), .Z(n6141) );
  NANDN U6401 ( .A(n472), .B(n471), .Z(n476) );
  NANDN U6402 ( .A(n474), .B(n473), .Z(n475) );
  AND U6403 ( .A(n476), .B(n475), .Z(n7303) );
  NANDN U6404 ( .A(n478), .B(n477), .Z(n482) );
  NAND U6405 ( .A(n480), .B(n479), .Z(n481) );
  AND U6406 ( .A(n482), .B(n481), .Z(n8877) );
  NANDN U6407 ( .A(n484), .B(n483), .Z(n488) );
  NAND U6408 ( .A(n486), .B(n485), .Z(n487) );
  NAND U6409 ( .A(n488), .B(n487), .Z(n8878) );
  XNOR U6410 ( .A(n8877), .B(n8878), .Z(n8880) );
  NANDN U6411 ( .A(n490), .B(n489), .Z(n494) );
  NAND U6412 ( .A(n492), .B(n491), .Z(n493) );
  AND U6413 ( .A(n494), .B(n493), .Z(n8879) );
  XOR U6414 ( .A(n8880), .B(n8879), .Z(n7301) );
  NANDN U6415 ( .A(n496), .B(n495), .Z(n500) );
  NANDN U6416 ( .A(n498), .B(n497), .Z(n499) );
  AND U6417 ( .A(n500), .B(n499), .Z(n7300) );
  XNOR U6418 ( .A(n7301), .B(n7300), .Z(n7302) );
  XOR U6419 ( .A(n7303), .B(n7302), .Z(n7393) );
  NANDN U6420 ( .A(n502), .B(n501), .Z(n506) );
  NANDN U6421 ( .A(n504), .B(n503), .Z(n505) );
  AND U6422 ( .A(n506), .B(n505), .Z(n7339) );
  NANDN U6423 ( .A(n508), .B(n507), .Z(n512) );
  NAND U6424 ( .A(n510), .B(n509), .Z(n511) );
  AND U6425 ( .A(n512), .B(n511), .Z(n6408) );
  NAND U6426 ( .A(n514), .B(n513), .Z(n518) );
  NAND U6427 ( .A(n516), .B(n515), .Z(n517) );
  NAND U6428 ( .A(n518), .B(n517), .Z(n6409) );
  XNOR U6429 ( .A(n6408), .B(n6409), .Z(n6411) );
  NAND U6430 ( .A(n520), .B(n519), .Z(n524) );
  NAND U6431 ( .A(n522), .B(n521), .Z(n523) );
  AND U6432 ( .A(n524), .B(n523), .Z(n6410) );
  XOR U6433 ( .A(n6411), .B(n6410), .Z(n7337) );
  NANDN U6434 ( .A(n526), .B(n525), .Z(n530) );
  NANDN U6435 ( .A(n528), .B(n527), .Z(n529) );
  AND U6436 ( .A(n530), .B(n529), .Z(n7336) );
  XNOR U6437 ( .A(n7337), .B(n7336), .Z(n7338) );
  XOR U6438 ( .A(n7339), .B(n7338), .Z(n7391) );
  NANDN U6439 ( .A(n532), .B(n531), .Z(n536) );
  NAND U6440 ( .A(n534), .B(n533), .Z(n535) );
  AND U6441 ( .A(n536), .B(n535), .Z(n6432) );
  NANDN U6442 ( .A(n538), .B(n537), .Z(n542) );
  NAND U6443 ( .A(n540), .B(n539), .Z(n541) );
  NAND U6444 ( .A(n542), .B(n541), .Z(n6433) );
  XNOR U6445 ( .A(n6432), .B(n6433), .Z(n6435) );
  NANDN U6446 ( .A(n544), .B(n543), .Z(n548) );
  NAND U6447 ( .A(n546), .B(n545), .Z(n547) );
  AND U6448 ( .A(n548), .B(n547), .Z(n6434) );
  XOR U6449 ( .A(n6435), .B(n6434), .Z(n6572) );
  NANDN U6450 ( .A(n550), .B(n549), .Z(n554) );
  NAND U6451 ( .A(n552), .B(n551), .Z(n553) );
  AND U6452 ( .A(n554), .B(n553), .Z(n8344) );
  NANDN U6453 ( .A(n556), .B(n555), .Z(n560) );
  NAND U6454 ( .A(n558), .B(n557), .Z(n559) );
  AND U6455 ( .A(n560), .B(n559), .Z(n8343) );
  XOR U6456 ( .A(n8344), .B(n8343), .Z(n8346) );
  NANDN U6457 ( .A(n562), .B(n561), .Z(n566) );
  NAND U6458 ( .A(n564), .B(n563), .Z(n565) );
  AND U6459 ( .A(n566), .B(n565), .Z(n8345) );
  XOR U6460 ( .A(n8346), .B(n8345), .Z(n6571) );
  NANDN U6461 ( .A(n568), .B(n567), .Z(n572) );
  NANDN U6462 ( .A(n570), .B(n569), .Z(n571) );
  AND U6463 ( .A(n572), .B(n571), .Z(n6570) );
  XOR U6464 ( .A(n6571), .B(n6570), .Z(n6573) );
  XNOR U6465 ( .A(n6572), .B(n6573), .Z(n7390) );
  XNOR U6466 ( .A(n7391), .B(n7390), .Z(n7392) );
  XNOR U6467 ( .A(n7393), .B(n7392), .Z(n6138) );
  NANDN U6468 ( .A(n574), .B(n573), .Z(n578) );
  NANDN U6469 ( .A(n576), .B(n575), .Z(n577) );
  AND U6470 ( .A(n578), .B(n577), .Z(n7141) );
  NANDN U6471 ( .A(n580), .B(n579), .Z(n584) );
  NANDN U6472 ( .A(n582), .B(n581), .Z(n583) );
  AND U6473 ( .A(n584), .B(n583), .Z(n7138) );
  NANDN U6474 ( .A(n586), .B(n585), .Z(n590) );
  NAND U6475 ( .A(n588), .B(n587), .Z(n589) );
  AND U6476 ( .A(n590), .B(n589), .Z(n8909) );
  NANDN U6477 ( .A(n592), .B(n591), .Z(n596) );
  NAND U6478 ( .A(n594), .B(n593), .Z(n595) );
  AND U6479 ( .A(n596), .B(n595), .Z(n8907) );
  XNOR U6480 ( .A(n8907), .B(oglobal[1]), .Z(n8908) );
  XOR U6481 ( .A(n8909), .B(n8908), .Z(n7139) );
  XNOR U6482 ( .A(n7138), .B(n7139), .Z(n7140) );
  XOR U6483 ( .A(n7141), .B(n7140), .Z(n7881) );
  NANDN U6484 ( .A(n598), .B(n597), .Z(n602) );
  NANDN U6485 ( .A(n600), .B(n599), .Z(n601) );
  AND U6486 ( .A(n602), .B(n601), .Z(n7387) );
  NANDN U6487 ( .A(n604), .B(n603), .Z(n608) );
  NAND U6488 ( .A(n606), .B(n605), .Z(n607) );
  AND U6489 ( .A(n608), .B(n607), .Z(n6396) );
  NAND U6490 ( .A(n610), .B(n609), .Z(n614) );
  NAND U6491 ( .A(n612), .B(n611), .Z(n613) );
  NAND U6492 ( .A(n614), .B(n613), .Z(n6397) );
  XNOR U6493 ( .A(n6396), .B(n6397), .Z(n6399) );
  NANDN U6494 ( .A(n616), .B(n615), .Z(n620) );
  NAND U6495 ( .A(n618), .B(n617), .Z(n619) );
  AND U6496 ( .A(n620), .B(n619), .Z(n6398) );
  XOR U6497 ( .A(n6399), .B(n6398), .Z(n7385) );
  NANDN U6498 ( .A(n622), .B(n621), .Z(n626) );
  NANDN U6499 ( .A(n624), .B(n623), .Z(n625) );
  AND U6500 ( .A(n626), .B(n625), .Z(n7384) );
  XNOR U6501 ( .A(n7385), .B(n7384), .Z(n7386) );
  XOR U6502 ( .A(n7387), .B(n7386), .Z(n7879) );
  NANDN U6503 ( .A(n628), .B(n627), .Z(n632) );
  NANDN U6504 ( .A(n630), .B(n629), .Z(n631) );
  AND U6505 ( .A(n632), .B(n631), .Z(n7333) );
  NANDN U6506 ( .A(n634), .B(n633), .Z(n638) );
  NAND U6507 ( .A(n636), .B(n635), .Z(n637) );
  AND U6508 ( .A(n638), .B(n637), .Z(n6922) );
  NANDN U6509 ( .A(n640), .B(n639), .Z(n644) );
  NAND U6510 ( .A(n642), .B(n641), .Z(n643) );
  NAND U6511 ( .A(n644), .B(n643), .Z(n6923) );
  XNOR U6512 ( .A(n6922), .B(n6923), .Z(n6925) );
  NANDN U6513 ( .A(n646), .B(n645), .Z(n650) );
  NAND U6514 ( .A(n648), .B(n647), .Z(n649) );
  AND U6515 ( .A(n650), .B(n649), .Z(n6924) );
  XOR U6516 ( .A(n6925), .B(n6924), .Z(n7331) );
  NANDN U6517 ( .A(n652), .B(n651), .Z(n656) );
  NANDN U6518 ( .A(n654), .B(n653), .Z(n655) );
  AND U6519 ( .A(n656), .B(n655), .Z(n7330) );
  XNOR U6520 ( .A(n7331), .B(n7330), .Z(n7332) );
  XNOR U6521 ( .A(n7333), .B(n7332), .Z(n7878) );
  XNOR U6522 ( .A(n7879), .B(n7878), .Z(n7880) );
  XNOR U6523 ( .A(n7881), .B(n7880), .Z(n6139) );
  XOR U6524 ( .A(n6138), .B(n6139), .Z(n6140) );
  XNOR U6525 ( .A(n6141), .B(n6140), .Z(n8638) );
  XOR U6526 ( .A(n8638), .B(n8637), .Z(n8639) );
  XNOR U6527 ( .A(n8640), .B(n8639), .Z(n7260) );
  NANDN U6528 ( .A(n662), .B(n661), .Z(n666) );
  NANDN U6529 ( .A(n664), .B(n663), .Z(n665) );
  NAND U6530 ( .A(n666), .B(n665), .Z(n7259) );
  NAND U6531 ( .A(n668), .B(n667), .Z(n672) );
  NAND U6532 ( .A(n670), .B(n669), .Z(n671) );
  NAND U6533 ( .A(n672), .B(n671), .Z(n7258) );
  XOR U6534 ( .A(n7259), .B(n7258), .Z(n7261) );
  XNOR U6535 ( .A(n7260), .B(n7261), .Z(n6662) );
  NANDN U6536 ( .A(n674), .B(n673), .Z(n678) );
  NANDN U6537 ( .A(n676), .B(n675), .Z(n677) );
  AND U6538 ( .A(n678), .B(n677), .Z(n7627) );
  NANDN U6539 ( .A(n680), .B(n679), .Z(n684) );
  NAND U6540 ( .A(n682), .B(n681), .Z(n683) );
  AND U6541 ( .A(n684), .B(n683), .Z(n6693) );
  NANDN U6542 ( .A(n686), .B(n685), .Z(n690) );
  NAND U6543 ( .A(n688), .B(n687), .Z(n689) );
  AND U6544 ( .A(n690), .B(n689), .Z(n6691) );
  NANDN U6545 ( .A(n692), .B(n691), .Z(n696) );
  NAND U6546 ( .A(n694), .B(n693), .Z(n695) );
  AND U6547 ( .A(n696), .B(n695), .Z(n6690) );
  XOR U6548 ( .A(n6691), .B(n6690), .Z(n6692) );
  XOR U6549 ( .A(n6693), .B(n6692), .Z(n6632) );
  NANDN U6550 ( .A(n698), .B(n697), .Z(n702) );
  NAND U6551 ( .A(n700), .B(n699), .Z(n701) );
  AND U6552 ( .A(n702), .B(n701), .Z(n6687) );
  NANDN U6553 ( .A(n704), .B(n703), .Z(n708) );
  NAND U6554 ( .A(n706), .B(n705), .Z(n707) );
  AND U6555 ( .A(n708), .B(n707), .Z(n6685) );
  NAND U6556 ( .A(n710), .B(n709), .Z(n714) );
  NAND U6557 ( .A(n712), .B(n711), .Z(n713) );
  AND U6558 ( .A(n714), .B(n713), .Z(n6684) );
  XOR U6559 ( .A(n6685), .B(n6684), .Z(n6686) );
  XOR U6560 ( .A(n6687), .B(n6686), .Z(n6631) );
  NANDN U6561 ( .A(n716), .B(n715), .Z(n720) );
  NANDN U6562 ( .A(n718), .B(n717), .Z(n719) );
  AND U6563 ( .A(n720), .B(n719), .Z(n6630) );
  XOR U6564 ( .A(n6631), .B(n6630), .Z(n6633) );
  XOR U6565 ( .A(n6632), .B(n6633), .Z(n7625) );
  NANDN U6566 ( .A(n722), .B(n721), .Z(n726) );
  NAND U6567 ( .A(n724), .B(n723), .Z(n725) );
  NAND U6568 ( .A(n726), .B(n725), .Z(n7624) );
  XNOR U6569 ( .A(n7625), .B(n7624), .Z(n7626) );
  XNOR U6570 ( .A(n7627), .B(n7626), .Z(n6219) );
  NANDN U6571 ( .A(n728), .B(n727), .Z(n732) );
  NANDN U6572 ( .A(n730), .B(n729), .Z(n731) );
  AND U6573 ( .A(n732), .B(n731), .Z(n7839) );
  NANDN U6574 ( .A(n734), .B(n733), .Z(n738) );
  NANDN U6575 ( .A(n736), .B(n735), .Z(n737) );
  AND U6576 ( .A(n738), .B(n737), .Z(n7836) );
  NANDN U6577 ( .A(n740), .B(n739), .Z(n744) );
  NAND U6578 ( .A(n742), .B(n741), .Z(n743) );
  AND U6579 ( .A(n744), .B(n743), .Z(n9039) );
  NANDN U6580 ( .A(n746), .B(n745), .Z(n750) );
  NAND U6581 ( .A(n748), .B(n747), .Z(n749) );
  NAND U6582 ( .A(n750), .B(n749), .Z(n9040) );
  XNOR U6583 ( .A(n9039), .B(n9040), .Z(n9042) );
  NANDN U6584 ( .A(n752), .B(n751), .Z(n756) );
  NAND U6585 ( .A(n754), .B(n753), .Z(n755) );
  AND U6586 ( .A(n756), .B(n755), .Z(n9041) );
  XOR U6587 ( .A(n9042), .B(n9041), .Z(n6579) );
  NANDN U6588 ( .A(n758), .B(n757), .Z(n762) );
  NAND U6589 ( .A(n760), .B(n759), .Z(n761) );
  AND U6590 ( .A(n762), .B(n761), .Z(n6757) );
  NAND U6591 ( .A(n764), .B(n763), .Z(n768) );
  NAND U6592 ( .A(n766), .B(n765), .Z(n767) );
  AND U6593 ( .A(n768), .B(n767), .Z(n6756) );
  XOR U6594 ( .A(n6757), .B(n6756), .Z(n6759) );
  NAND U6595 ( .A(n770), .B(n769), .Z(n774) );
  NAND U6596 ( .A(n772), .B(n771), .Z(n773) );
  AND U6597 ( .A(n774), .B(n773), .Z(n6758) );
  XOR U6598 ( .A(n6759), .B(n6758), .Z(n6577) );
  NANDN U6599 ( .A(n776), .B(n775), .Z(n780) );
  NANDN U6600 ( .A(n778), .B(n777), .Z(n779) );
  AND U6601 ( .A(n780), .B(n779), .Z(n6576) );
  XNOR U6602 ( .A(n6577), .B(n6576), .Z(n6578) );
  XOR U6603 ( .A(n6579), .B(n6578), .Z(n7837) );
  XNOR U6604 ( .A(n7836), .B(n7837), .Z(n7838) );
  XOR U6605 ( .A(n7839), .B(n7838), .Z(n6217) );
  NANDN U6606 ( .A(n782), .B(n781), .Z(n786) );
  NANDN U6607 ( .A(n784), .B(n783), .Z(n785) );
  AND U6608 ( .A(n786), .B(n785), .Z(n7621) );
  NAND U6609 ( .A(n788), .B(n787), .Z(n792) );
  NAND U6610 ( .A(n790), .B(n789), .Z(n791) );
  AND U6611 ( .A(n792), .B(n791), .Z(n6750) );
  NAND U6612 ( .A(n794), .B(n793), .Z(n798) );
  NAND U6613 ( .A(n796), .B(n795), .Z(n797) );
  NAND U6614 ( .A(n798), .B(n797), .Z(n6751) );
  XNOR U6615 ( .A(n6750), .B(n6751), .Z(n6753) );
  NANDN U6616 ( .A(n800), .B(n799), .Z(n804) );
  NANDN U6617 ( .A(n802), .B(n801), .Z(n803) );
  AND U6618 ( .A(n804), .B(n803), .Z(n6752) );
  XOR U6619 ( .A(n6753), .B(n6752), .Z(n6344) );
  NAND U6620 ( .A(n806), .B(n805), .Z(n810) );
  NAND U6621 ( .A(n808), .B(n807), .Z(n809) );
  AND U6622 ( .A(n810), .B(n809), .Z(n6744) );
  NANDN U6623 ( .A(n812), .B(n811), .Z(n816) );
  NAND U6624 ( .A(n814), .B(n813), .Z(n815) );
  NAND U6625 ( .A(n816), .B(n815), .Z(n6745) );
  XNOR U6626 ( .A(n6744), .B(n6745), .Z(n6747) );
  NAND U6627 ( .A(n818), .B(n817), .Z(n822) );
  NAND U6628 ( .A(n820), .B(n819), .Z(n821) );
  AND U6629 ( .A(n822), .B(n821), .Z(n6746) );
  XOR U6630 ( .A(n6747), .B(n6746), .Z(n6343) );
  NANDN U6631 ( .A(n824), .B(n823), .Z(n828) );
  NANDN U6632 ( .A(n826), .B(n825), .Z(n827) );
  AND U6633 ( .A(n828), .B(n827), .Z(n6342) );
  XOR U6634 ( .A(n6343), .B(n6342), .Z(n6345) );
  XOR U6635 ( .A(n6344), .B(n6345), .Z(n7619) );
  NANDN U6636 ( .A(n830), .B(n829), .Z(n834) );
  NAND U6637 ( .A(n832), .B(n831), .Z(n833) );
  NAND U6638 ( .A(n834), .B(n833), .Z(n7618) );
  XNOR U6639 ( .A(n7619), .B(n7618), .Z(n7620) );
  XNOR U6640 ( .A(n7621), .B(n7620), .Z(n6216) );
  XNOR U6641 ( .A(n6217), .B(n6216), .Z(n6218) );
  XNOR U6642 ( .A(n6219), .B(n6218), .Z(n9058) );
  NANDN U6643 ( .A(n836), .B(n835), .Z(n840) );
  NAND U6644 ( .A(n838), .B(n837), .Z(n839) );
  AND U6645 ( .A(n840), .B(n839), .Z(n6303) );
  NANDN U6646 ( .A(n842), .B(n841), .Z(n846) );
  NAND U6647 ( .A(n844), .B(n843), .Z(n845) );
  AND U6648 ( .A(n846), .B(n845), .Z(n8913) );
  NANDN U6649 ( .A(n848), .B(n847), .Z(n852) );
  NAND U6650 ( .A(n850), .B(n849), .Z(n851) );
  AND U6651 ( .A(n852), .B(n851), .Z(n8912) );
  XOR U6652 ( .A(n8913), .B(n8912), .Z(n8915) );
  NANDN U6653 ( .A(n854), .B(n853), .Z(n858) );
  NAND U6654 ( .A(n856), .B(n855), .Z(n857) );
  AND U6655 ( .A(n858), .B(n857), .Z(n8914) );
  XOR U6656 ( .A(n8915), .B(n8914), .Z(n6494) );
  NANDN U6657 ( .A(n860), .B(n859), .Z(n864) );
  NAND U6658 ( .A(n862), .B(n861), .Z(n863) );
  AND U6659 ( .A(n864), .B(n863), .Z(n8158) );
  NANDN U6660 ( .A(n866), .B(n865), .Z(n870) );
  NAND U6661 ( .A(n868), .B(n867), .Z(n869) );
  AND U6662 ( .A(n870), .B(n869), .Z(n8157) );
  XOR U6663 ( .A(n8158), .B(n8157), .Z(n8160) );
  NANDN U6664 ( .A(n872), .B(n871), .Z(n876) );
  NAND U6665 ( .A(n874), .B(n873), .Z(n875) );
  AND U6666 ( .A(n876), .B(n875), .Z(n8159) );
  XOR U6667 ( .A(n8160), .B(n8159), .Z(n6493) );
  NANDN U6668 ( .A(n878), .B(n877), .Z(n882) );
  NANDN U6669 ( .A(n880), .B(n879), .Z(n881) );
  AND U6670 ( .A(n882), .B(n881), .Z(n6492) );
  XOR U6671 ( .A(n6493), .B(n6492), .Z(n6495) );
  XOR U6672 ( .A(n6494), .B(n6495), .Z(n6301) );
  NANDN U6673 ( .A(n884), .B(n883), .Z(n888) );
  NAND U6674 ( .A(n886), .B(n885), .Z(n887) );
  NAND U6675 ( .A(n888), .B(n887), .Z(n6300) );
  XNOR U6676 ( .A(n6301), .B(n6300), .Z(n6302) );
  XNOR U6677 ( .A(n6303), .B(n6302), .Z(n6168) );
  NANDN U6678 ( .A(n890), .B(n889), .Z(n894) );
  NANDN U6679 ( .A(n892), .B(n891), .Z(n893) );
  AND U6680 ( .A(n894), .B(n893), .Z(n6315) );
  NANDN U6681 ( .A(n896), .B(n895), .Z(n900) );
  NAND U6682 ( .A(n898), .B(n897), .Z(n899) );
  AND U6683 ( .A(n900), .B(n899), .Z(n8986) );
  NANDN U6684 ( .A(n902), .B(n901), .Z(n906) );
  NAND U6685 ( .A(n904), .B(n903), .Z(n905) );
  AND U6686 ( .A(n906), .B(n905), .Z(n8985) );
  XOR U6687 ( .A(n8986), .B(n8985), .Z(n8988) );
  NANDN U6688 ( .A(n908), .B(n907), .Z(n912) );
  NAND U6689 ( .A(n910), .B(n909), .Z(n911) );
  AND U6690 ( .A(n912), .B(n911), .Z(n8987) );
  XOR U6691 ( .A(n8988), .B(n8987), .Z(n6488) );
  NANDN U6692 ( .A(n914), .B(n913), .Z(n918) );
  NAND U6693 ( .A(n916), .B(n915), .Z(n917) );
  AND U6694 ( .A(n918), .B(n917), .Z(n7867) );
  NANDN U6695 ( .A(n920), .B(n919), .Z(n924) );
  NAND U6696 ( .A(n922), .B(n921), .Z(n923) );
  AND U6697 ( .A(n924), .B(n923), .Z(n7866) );
  XOR U6698 ( .A(n7867), .B(n7866), .Z(n7869) );
  NAND U6699 ( .A(n926), .B(n925), .Z(n930) );
  NAND U6700 ( .A(n928), .B(n927), .Z(n929) );
  AND U6701 ( .A(n930), .B(n929), .Z(n7868) );
  XOR U6702 ( .A(n7869), .B(n7868), .Z(n6487) );
  NANDN U6703 ( .A(n932), .B(n931), .Z(n936) );
  NANDN U6704 ( .A(n934), .B(n933), .Z(n935) );
  AND U6705 ( .A(n936), .B(n935), .Z(n6486) );
  XOR U6706 ( .A(n6487), .B(n6486), .Z(n6489) );
  XOR U6707 ( .A(n6488), .B(n6489), .Z(n6313) );
  NANDN U6708 ( .A(n938), .B(n937), .Z(n942) );
  NAND U6709 ( .A(n940), .B(n939), .Z(n941) );
  NAND U6710 ( .A(n942), .B(n941), .Z(n6312) );
  XNOR U6711 ( .A(n6313), .B(n6312), .Z(n6314) );
  XNOR U6712 ( .A(n6315), .B(n6314), .Z(n6169) );
  XOR U6713 ( .A(n6168), .B(n6169), .Z(n6171) );
  NAND U6714 ( .A(n944), .B(n943), .Z(n948) );
  NAND U6715 ( .A(n946), .B(n945), .Z(n947) );
  AND U6716 ( .A(n948), .B(n947), .Z(n6170) );
  XNOR U6717 ( .A(n6171), .B(n6170), .Z(n9057) );
  XOR U6718 ( .A(n9058), .B(n9057), .Z(n9059) );
  NAND U6719 ( .A(n950), .B(n949), .Z(n954) );
  NAND U6720 ( .A(n952), .B(n951), .Z(n953) );
  AND U6721 ( .A(n954), .B(n953), .Z(n9060) );
  XOR U6722 ( .A(n9059), .B(n9060), .Z(n6661) );
  NANDN U6723 ( .A(n956), .B(n955), .Z(n960) );
  NAND U6724 ( .A(n958), .B(n957), .Z(n959) );
  AND U6725 ( .A(n960), .B(n959), .Z(n7507) );
  NANDN U6726 ( .A(n962), .B(n961), .Z(n966) );
  NANDN U6727 ( .A(n964), .B(n963), .Z(n965) );
  AND U6728 ( .A(n966), .B(n965), .Z(n7033) );
  NANDN U6729 ( .A(n968), .B(n967), .Z(n972) );
  NAND U6730 ( .A(n970), .B(n969), .Z(n971) );
  AND U6731 ( .A(n972), .B(n971), .Z(n8583) );
  NANDN U6732 ( .A(n974), .B(n973), .Z(n978) );
  NAND U6733 ( .A(n976), .B(n975), .Z(n977) );
  NAND U6734 ( .A(n978), .B(n977), .Z(n8584) );
  XNOR U6735 ( .A(n8583), .B(n8584), .Z(n8586) );
  NANDN U6736 ( .A(n980), .B(n979), .Z(n984) );
  NAND U6737 ( .A(n982), .B(n981), .Z(n983) );
  AND U6738 ( .A(n984), .B(n983), .Z(n8585) );
  XOR U6739 ( .A(n8586), .B(n8585), .Z(n7031) );
  NANDN U6740 ( .A(n986), .B(n985), .Z(n990) );
  NANDN U6741 ( .A(n988), .B(n987), .Z(n989) );
  AND U6742 ( .A(n990), .B(n989), .Z(n7030) );
  XNOR U6743 ( .A(n7031), .B(n7030), .Z(n7032) );
  XOR U6744 ( .A(n7033), .B(n7032), .Z(n7505) );
  NANDN U6745 ( .A(n992), .B(n991), .Z(n996) );
  NAND U6746 ( .A(n994), .B(n993), .Z(n995) );
  NAND U6747 ( .A(n996), .B(n995), .Z(n7504) );
  XNOR U6748 ( .A(n7505), .B(n7504), .Z(n7506) );
  XNOR U6749 ( .A(n7507), .B(n7506), .Z(n7060) );
  NANDN U6750 ( .A(n998), .B(n997), .Z(n1002) );
  NANDN U6751 ( .A(n1000), .B(n999), .Z(n1001) );
  AND U6752 ( .A(n1002), .B(n1001), .Z(n7926) );
  NANDN U6753 ( .A(n1004), .B(n1003), .Z(n1008) );
  NANDN U6754 ( .A(n1006), .B(n1005), .Z(n1007) );
  AND U6755 ( .A(n1008), .B(n1007), .Z(n7923) );
  NANDN U6756 ( .A(n1010), .B(n1009), .Z(n1014) );
  NANDN U6757 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U6758 ( .A(n1014), .B(n1013), .Z(n7924) );
  XNOR U6759 ( .A(n7923), .B(n7924), .Z(n7925) );
  XOR U6760 ( .A(n7926), .B(n7925), .Z(n7555) );
  NANDN U6761 ( .A(n1016), .B(n1015), .Z(n1020) );
  NAND U6762 ( .A(n1018), .B(n1017), .Z(n1019) );
  AND U6763 ( .A(n1020), .B(n1019), .Z(n6816) );
  NANDN U6764 ( .A(n1022), .B(n1021), .Z(n1026) );
  NAND U6765 ( .A(n1024), .B(n1023), .Z(n1025) );
  NAND U6766 ( .A(n1026), .B(n1025), .Z(n6817) );
  XNOR U6767 ( .A(n6816), .B(n6817), .Z(n6819) );
  NANDN U6768 ( .A(n1028), .B(n1027), .Z(n1032) );
  NAND U6769 ( .A(n1030), .B(n1029), .Z(n1031) );
  AND U6770 ( .A(n1032), .B(n1031), .Z(n6818) );
  XOR U6771 ( .A(n6819), .B(n6818), .Z(n7404) );
  NANDN U6772 ( .A(n1034), .B(n1033), .Z(n1038) );
  NANDN U6773 ( .A(n1036), .B(n1035), .Z(n1037) );
  AND U6774 ( .A(n1038), .B(n1037), .Z(n8547) );
  NANDN U6775 ( .A(n1040), .B(n1039), .Z(n1044) );
  NAND U6776 ( .A(n1042), .B(n1041), .Z(n1043) );
  NAND U6777 ( .A(n1044), .B(n1043), .Z(n8548) );
  XNOR U6778 ( .A(n8547), .B(n8548), .Z(n8550) );
  NANDN U6779 ( .A(n1046), .B(n1045), .Z(n1050) );
  NAND U6780 ( .A(n1048), .B(n1047), .Z(n1049) );
  AND U6781 ( .A(n1050), .B(n1049), .Z(n8549) );
  XOR U6782 ( .A(n8550), .B(n8549), .Z(n7403) );
  NANDN U6783 ( .A(n1052), .B(n1051), .Z(n1056) );
  NANDN U6784 ( .A(n1054), .B(n1053), .Z(n1055) );
  AND U6785 ( .A(n1056), .B(n1055), .Z(n7402) );
  XOR U6786 ( .A(n7403), .B(n7402), .Z(n7405) );
  XOR U6787 ( .A(n7404), .B(n7405), .Z(n7553) );
  NANDN U6788 ( .A(n1058), .B(n1057), .Z(n1062) );
  NAND U6789 ( .A(n1060), .B(n1059), .Z(n1061) );
  AND U6790 ( .A(n1062), .B(n1061), .Z(n8403) );
  NANDN U6791 ( .A(n1064), .B(n1063), .Z(n1068) );
  NAND U6792 ( .A(n1066), .B(n1065), .Z(n1067) );
  NAND U6793 ( .A(n1068), .B(n1067), .Z(n8404) );
  XNOR U6794 ( .A(n8403), .B(n8404), .Z(n8406) );
  NAND U6795 ( .A(n1070), .B(n1069), .Z(n1074) );
  NAND U6796 ( .A(n1072), .B(n1071), .Z(n1073) );
  AND U6797 ( .A(n1074), .B(n1073), .Z(n8405) );
  XOR U6798 ( .A(n8406), .B(n8405), .Z(n8039) );
  NANDN U6799 ( .A(n1076), .B(n1075), .Z(n1080) );
  NAND U6800 ( .A(n1078), .B(n1077), .Z(n1079) );
  AND U6801 ( .A(n1080), .B(n1079), .Z(n6714) );
  NANDN U6802 ( .A(n1082), .B(n1081), .Z(n1086) );
  NAND U6803 ( .A(n1084), .B(n1083), .Z(n1085) );
  NAND U6804 ( .A(n1086), .B(n1085), .Z(n6715) );
  XNOR U6805 ( .A(n6714), .B(n6715), .Z(n6717) );
  NANDN U6806 ( .A(n1088), .B(n1087), .Z(n1092) );
  NAND U6807 ( .A(n1090), .B(n1089), .Z(n1091) );
  AND U6808 ( .A(n1092), .B(n1091), .Z(n6716) );
  XOR U6809 ( .A(n6717), .B(n6716), .Z(n8038) );
  NANDN U6810 ( .A(n1094), .B(n1093), .Z(n1098) );
  NANDN U6811 ( .A(n1096), .B(n1095), .Z(n1097) );
  AND U6812 ( .A(n1098), .B(n1097), .Z(n8037) );
  XOR U6813 ( .A(n8038), .B(n8037), .Z(n8040) );
  XNOR U6814 ( .A(n8039), .B(n8040), .Z(n7552) );
  XNOR U6815 ( .A(n7553), .B(n7552), .Z(n7554) );
  XOR U6816 ( .A(n7555), .B(n7554), .Z(n7061) );
  XNOR U6817 ( .A(n7060), .B(n7061), .Z(n7063) );
  NANDN U6818 ( .A(n1100), .B(n1099), .Z(n1104) );
  NAND U6819 ( .A(n1102), .B(n1101), .Z(n1103) );
  AND U6820 ( .A(n1104), .B(n1103), .Z(n7561) );
  NANDN U6821 ( .A(n1106), .B(n1105), .Z(n1110) );
  NAND U6822 ( .A(n1108), .B(n1107), .Z(n1109) );
  AND U6823 ( .A(n1110), .B(n1109), .Z(n8733) );
  NANDN U6824 ( .A(n1112), .B(n1111), .Z(n1116) );
  NAND U6825 ( .A(n1114), .B(n1113), .Z(n1115) );
  NAND U6826 ( .A(n1116), .B(n1115), .Z(n8734) );
  XNOR U6827 ( .A(n8733), .B(n8734), .Z(n8736) );
  NANDN U6828 ( .A(n1118), .B(n1117), .Z(n1122) );
  NAND U6829 ( .A(n1120), .B(n1119), .Z(n1121) );
  AND U6830 ( .A(n1122), .B(n1121), .Z(n8735) );
  XOR U6831 ( .A(n8736), .B(n8735), .Z(n7410) );
  NANDN U6832 ( .A(n1124), .B(n1123), .Z(n1128) );
  NAND U6833 ( .A(n1126), .B(n1125), .Z(n1127) );
  AND U6834 ( .A(n1128), .B(n1127), .Z(n8493) );
  NANDN U6835 ( .A(n1130), .B(n1129), .Z(n1134) );
  NAND U6836 ( .A(n1132), .B(n1131), .Z(n1133) );
  NAND U6837 ( .A(n1134), .B(n1133), .Z(n8494) );
  XNOR U6838 ( .A(n8493), .B(n8494), .Z(n8496) );
  NANDN U6839 ( .A(n1136), .B(n1135), .Z(n1140) );
  NAND U6840 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U6841 ( .A(n1140), .B(n1139), .Z(n8495) );
  XOR U6842 ( .A(n8496), .B(n8495), .Z(n7409) );
  NANDN U6843 ( .A(n1142), .B(n1141), .Z(n1146) );
  NAND U6844 ( .A(n1144), .B(n1143), .Z(n1145) );
  AND U6845 ( .A(n1146), .B(n1145), .Z(n6828) );
  NANDN U6846 ( .A(n1148), .B(n1147), .Z(n1152) );
  NAND U6847 ( .A(n1150), .B(n1149), .Z(n1151) );
  NAND U6848 ( .A(n1152), .B(n1151), .Z(n6829) );
  XNOR U6849 ( .A(n6828), .B(n6829), .Z(n6831) );
  NANDN U6850 ( .A(n1154), .B(n1153), .Z(n1158) );
  NAND U6851 ( .A(n1156), .B(n1155), .Z(n1157) );
  AND U6852 ( .A(n1158), .B(n1157), .Z(n6830) );
  XNOR U6853 ( .A(n6831), .B(n6830), .Z(n7408) );
  XOR U6854 ( .A(n7409), .B(n7408), .Z(n7411) );
  XOR U6855 ( .A(n7410), .B(n7411), .Z(n7559) );
  NANDN U6856 ( .A(n1160), .B(n1159), .Z(n1164) );
  NAND U6857 ( .A(n1162), .B(n1161), .Z(n1163) );
  NAND U6858 ( .A(n1164), .B(n1163), .Z(n7558) );
  XNOR U6859 ( .A(n7559), .B(n7558), .Z(n7560) );
  XNOR U6860 ( .A(n7561), .B(n7560), .Z(n7062) );
  XOR U6861 ( .A(n7063), .B(n7062), .Z(n6547) );
  NANDN U6862 ( .A(n1166), .B(n1165), .Z(n1170) );
  NANDN U6863 ( .A(n1168), .B(n1167), .Z(n1169) );
  AND U6864 ( .A(n1170), .B(n1169), .Z(n6327) );
  NAND U6865 ( .A(n1172), .B(n1171), .Z(n1176) );
  NAND U6866 ( .A(n1174), .B(n1173), .Z(n1175) );
  AND U6867 ( .A(n1176), .B(n1175), .Z(n8451) );
  NAND U6868 ( .A(n1178), .B(n1177), .Z(n1182) );
  NAND U6869 ( .A(n1180), .B(n1179), .Z(n1181) );
  NAND U6870 ( .A(n1182), .B(n1181), .Z(n8452) );
  XNOR U6871 ( .A(n8451), .B(n8452), .Z(n8454) );
  NAND U6872 ( .A(n1184), .B(n1183), .Z(n1188) );
  NAND U6873 ( .A(n1186), .B(n1185), .Z(n1187) );
  AND U6874 ( .A(n1188), .B(n1187), .Z(n8453) );
  XOR U6875 ( .A(n8454), .B(n8453), .Z(n7008) );
  NANDN U6876 ( .A(n1190), .B(n1189), .Z(n1194) );
  NAND U6877 ( .A(n1192), .B(n1191), .Z(n1193) );
  AND U6878 ( .A(n1194), .B(n1193), .Z(n8217) );
  NANDN U6879 ( .A(n1196), .B(n1195), .Z(n1200) );
  NAND U6880 ( .A(n1198), .B(n1197), .Z(n1199) );
  NAND U6881 ( .A(n1200), .B(n1199), .Z(n8218) );
  XNOR U6882 ( .A(n8217), .B(n8218), .Z(n8220) );
  NANDN U6883 ( .A(n1202), .B(n1201), .Z(n1206) );
  NAND U6884 ( .A(n1204), .B(n1203), .Z(n1205) );
  AND U6885 ( .A(n1206), .B(n1205), .Z(n8219) );
  XOR U6886 ( .A(n8220), .B(n8219), .Z(n7007) );
  NANDN U6887 ( .A(n1208), .B(n1207), .Z(n1212) );
  NAND U6888 ( .A(n1210), .B(n1209), .Z(n1211) );
  AND U6889 ( .A(n1212), .B(n1211), .Z(n8487) );
  NANDN U6890 ( .A(n1214), .B(n1213), .Z(n1218) );
  NAND U6891 ( .A(n1216), .B(n1215), .Z(n1217) );
  NAND U6892 ( .A(n1218), .B(n1217), .Z(n8488) );
  XNOR U6893 ( .A(n8487), .B(n8488), .Z(n8490) );
  NANDN U6894 ( .A(n1220), .B(n1219), .Z(n1224) );
  NAND U6895 ( .A(n1222), .B(n1221), .Z(n1223) );
  AND U6896 ( .A(n1224), .B(n1223), .Z(n8489) );
  XNOR U6897 ( .A(n8490), .B(n8489), .Z(n7006) );
  XOR U6898 ( .A(n7007), .B(n7006), .Z(n7009) );
  XOR U6899 ( .A(n7008), .B(n7009), .Z(n6325) );
  NANDN U6900 ( .A(n1226), .B(n1225), .Z(n1230) );
  NAND U6901 ( .A(n1228), .B(n1227), .Z(n1229) );
  NAND U6902 ( .A(n1230), .B(n1229), .Z(n6324) );
  XNOR U6903 ( .A(n6325), .B(n6324), .Z(n6326) );
  XNOR U6904 ( .A(n6327), .B(n6326), .Z(n7273) );
  NANDN U6905 ( .A(n1232), .B(n1231), .Z(n1236) );
  NAND U6906 ( .A(n1234), .B(n1233), .Z(n1235) );
  AND U6907 ( .A(n1236), .B(n1235), .Z(n7435) );
  NANDN U6908 ( .A(n1238), .B(n1237), .Z(n1242) );
  NANDN U6909 ( .A(n1240), .B(n1239), .Z(n1241) );
  AND U6910 ( .A(n1242), .B(n1241), .Z(n7893) );
  NANDN U6911 ( .A(n1244), .B(n1243), .Z(n1248) );
  NAND U6912 ( .A(n1246), .B(n1245), .Z(n1247) );
  AND U6913 ( .A(n1248), .B(n1247), .Z(n8475) );
  NANDN U6914 ( .A(n1250), .B(n1249), .Z(n1254) );
  NAND U6915 ( .A(n1252), .B(n1251), .Z(n1253) );
  NAND U6916 ( .A(n1254), .B(n1253), .Z(n8476) );
  XNOR U6917 ( .A(n8475), .B(n8476), .Z(n8478) );
  NANDN U6918 ( .A(n1256), .B(n1255), .Z(n1260) );
  NAND U6919 ( .A(n1258), .B(n1257), .Z(n1259) );
  AND U6920 ( .A(n1260), .B(n1259), .Z(n8477) );
  XOR U6921 ( .A(n8478), .B(n8477), .Z(n7891) );
  NANDN U6922 ( .A(n1262), .B(n1261), .Z(n1266) );
  NAND U6923 ( .A(n1264), .B(n1263), .Z(n1265) );
  AND U6924 ( .A(n1266), .B(n1265), .Z(n8139) );
  NANDN U6925 ( .A(n1268), .B(n1267), .Z(n1272) );
  NANDN U6926 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U6927 ( .A(n1272), .B(n1271), .Z(n8140) );
  XNOR U6928 ( .A(n8139), .B(n8140), .Z(n8142) );
  NANDN U6929 ( .A(n1274), .B(n1273), .Z(n1278) );
  NANDN U6930 ( .A(n1276), .B(n1275), .Z(n1277) );
  AND U6931 ( .A(n1278), .B(n1277), .Z(n8141) );
  XNOR U6932 ( .A(n8142), .B(n8141), .Z(n7890) );
  XNOR U6933 ( .A(n7891), .B(n7890), .Z(n7892) );
  XOR U6934 ( .A(n7893), .B(n7892), .Z(n7433) );
  NANDN U6935 ( .A(n1280), .B(n1279), .Z(n1284) );
  NANDN U6936 ( .A(n1282), .B(n1281), .Z(n1283) );
  NAND U6937 ( .A(n1284), .B(n1283), .Z(n7432) );
  XNOR U6938 ( .A(n7433), .B(n7432), .Z(n7434) );
  XNOR U6939 ( .A(n7435), .B(n7434), .Z(n7270) );
  NANDN U6940 ( .A(n1286), .B(n1285), .Z(n1290) );
  NANDN U6941 ( .A(n1288), .B(n1287), .Z(n1289) );
  AND U6942 ( .A(n1290), .B(n1289), .Z(n7441) );
  NANDN U6943 ( .A(n1292), .B(n1291), .Z(n1296) );
  NANDN U6944 ( .A(n1294), .B(n1293), .Z(n1295) );
  AND U6945 ( .A(n1296), .B(n1295), .Z(n7899) );
  NANDN U6946 ( .A(n1298), .B(n1297), .Z(n1302) );
  NAND U6947 ( .A(n1300), .B(n1299), .Z(n1301) );
  AND U6948 ( .A(n1302), .B(n1301), .Z(n8721) );
  NANDN U6949 ( .A(n1304), .B(n1303), .Z(n1308) );
  NAND U6950 ( .A(n1306), .B(n1305), .Z(n1307) );
  NAND U6951 ( .A(n1308), .B(n1307), .Z(n8722) );
  XNOR U6952 ( .A(n8721), .B(n8722), .Z(n8724) );
  NANDN U6953 ( .A(n1310), .B(n1309), .Z(n1314) );
  NAND U6954 ( .A(n1312), .B(n1311), .Z(n1313) );
  AND U6955 ( .A(n1314), .B(n1313), .Z(n8723) );
  XOR U6956 ( .A(n8724), .B(n8723), .Z(n7897) );
  NANDN U6957 ( .A(n1316), .B(n1315), .Z(n1320) );
  NANDN U6958 ( .A(n1318), .B(n1317), .Z(n1319) );
  AND U6959 ( .A(n1320), .B(n1319), .Z(n7896) );
  XNOR U6960 ( .A(n7897), .B(n7896), .Z(n7898) );
  XOR U6961 ( .A(n7899), .B(n7898), .Z(n7439) );
  NANDN U6962 ( .A(n1322), .B(n1321), .Z(n1326) );
  NAND U6963 ( .A(n1324), .B(n1323), .Z(n1325) );
  NAND U6964 ( .A(n1326), .B(n1325), .Z(n7438) );
  XNOR U6965 ( .A(n7439), .B(n7438), .Z(n7440) );
  XNOR U6966 ( .A(n7441), .B(n7440), .Z(n7271) );
  XOR U6967 ( .A(n7270), .B(n7271), .Z(n7272) );
  XNOR U6968 ( .A(n7273), .B(n7272), .Z(n6546) );
  NANDN U6969 ( .A(n1328), .B(n1327), .Z(n1332) );
  OR U6970 ( .A(n1330), .B(n1329), .Z(n1331) );
  AND U6971 ( .A(n1332), .B(n1331), .Z(n7057) );
  NANDN U6972 ( .A(n1334), .B(n1333), .Z(n1338) );
  NANDN U6973 ( .A(n1336), .B(n1335), .Z(n1337) );
  AND U6974 ( .A(n1338), .B(n1337), .Z(n6242) );
  NANDN U6975 ( .A(n1340), .B(n1339), .Z(n1344) );
  NANDN U6976 ( .A(n1342), .B(n1341), .Z(n1343) );
  AND U6977 ( .A(n1344), .B(n1343), .Z(n7201) );
  NANDN U6978 ( .A(n1346), .B(n1345), .Z(n1350) );
  NAND U6979 ( .A(n1348), .B(n1347), .Z(n1349) );
  AND U6980 ( .A(n1350), .B(n1349), .Z(n6798) );
  NANDN U6981 ( .A(n1352), .B(n1351), .Z(n1356) );
  NAND U6982 ( .A(n1354), .B(n1353), .Z(n1355) );
  NAND U6983 ( .A(n1356), .B(n1355), .Z(n6799) );
  XNOR U6984 ( .A(n6798), .B(n6799), .Z(n6801) );
  NANDN U6985 ( .A(n1358), .B(n1357), .Z(n1362) );
  NAND U6986 ( .A(n1360), .B(n1359), .Z(n1361) );
  AND U6987 ( .A(n1362), .B(n1361), .Z(n6800) );
  XOR U6988 ( .A(n6801), .B(n6800), .Z(n7199) );
  NANDN U6989 ( .A(n1364), .B(n1363), .Z(n1368) );
  NANDN U6990 ( .A(n1366), .B(n1365), .Z(n1367) );
  AND U6991 ( .A(n1368), .B(n1367), .Z(n7198) );
  XNOR U6992 ( .A(n7199), .B(n7198), .Z(n7200) );
  XOR U6993 ( .A(n7201), .B(n7200), .Z(n6241) );
  NANDN U6994 ( .A(n1370), .B(n1369), .Z(n1374) );
  NAND U6995 ( .A(n1372), .B(n1371), .Z(n1373) );
  NAND U6996 ( .A(n1374), .B(n1373), .Z(n6240) );
  XOR U6997 ( .A(n6241), .B(n6240), .Z(n6243) );
  XOR U6998 ( .A(n6242), .B(n6243), .Z(n7055) );
  NANDN U6999 ( .A(n1376), .B(n1375), .Z(n1380) );
  NANDN U7000 ( .A(n1378), .B(n1377), .Z(n1379) );
  AND U7001 ( .A(n1380), .B(n1379), .Z(n6200) );
  NANDN U7002 ( .A(n1382), .B(n1381), .Z(n1386) );
  NAND U7003 ( .A(n1384), .B(n1383), .Z(n1385) );
  AND U7004 ( .A(n1386), .B(n1385), .Z(n6198) );
  NANDN U7005 ( .A(n1388), .B(n1387), .Z(n1392) );
  NANDN U7006 ( .A(n1390), .B(n1389), .Z(n1391) );
  AND U7007 ( .A(n1392), .B(n1391), .Z(n7026) );
  NANDN U7008 ( .A(n1394), .B(n1393), .Z(n1398) );
  NAND U7009 ( .A(n1396), .B(n1395), .Z(n1397) );
  AND U7010 ( .A(n1398), .B(n1397), .Z(n6792) );
  NANDN U7011 ( .A(n1400), .B(n1399), .Z(n1404) );
  NAND U7012 ( .A(n1402), .B(n1401), .Z(n1403) );
  NAND U7013 ( .A(n1404), .B(n1403), .Z(n6793) );
  XNOR U7014 ( .A(n6792), .B(n6793), .Z(n6795) );
  NANDN U7015 ( .A(n1406), .B(n1405), .Z(n1410) );
  NAND U7016 ( .A(n1408), .B(n1407), .Z(n1409) );
  AND U7017 ( .A(n1410), .B(n1409), .Z(n6794) );
  XOR U7018 ( .A(n6795), .B(n6794), .Z(n7025) );
  NANDN U7019 ( .A(n1412), .B(n1411), .Z(n1416) );
  NANDN U7020 ( .A(n1414), .B(n1413), .Z(n1415) );
  AND U7021 ( .A(n1416), .B(n1415), .Z(n7024) );
  XOR U7022 ( .A(n7025), .B(n7024), .Z(n7027) );
  XOR U7023 ( .A(n7026), .B(n7027), .Z(n6199) );
  XOR U7024 ( .A(n6198), .B(n6199), .Z(n6201) );
  XNOR U7025 ( .A(n6200), .B(n6201), .Z(n7054) );
  XNOR U7026 ( .A(n7055), .B(n7054), .Z(n7056) );
  XOR U7027 ( .A(n7057), .B(n7056), .Z(n6549) );
  XOR U7028 ( .A(n6661), .B(n6660), .Z(n6663) );
  XNOR U7029 ( .A(n6662), .B(n6663), .Z(n7236) );
  NANDN U7030 ( .A(n1418), .B(n1417), .Z(n1422) );
  NAND U7031 ( .A(n1420), .B(n1419), .Z(n1421) );
  AND U7032 ( .A(n1422), .B(n1421), .Z(n6134) );
  NANDN U7033 ( .A(n1424), .B(n1423), .Z(n1428) );
  NAND U7034 ( .A(n1426), .B(n1425), .Z(n1427) );
  AND U7035 ( .A(n1428), .B(n1427), .Z(n8193) );
  NANDN U7036 ( .A(n1430), .B(n1429), .Z(n1434) );
  NAND U7037 ( .A(n1432), .B(n1431), .Z(n1433) );
  NAND U7038 ( .A(n1434), .B(n1433), .Z(n8194) );
  XNOR U7039 ( .A(n8193), .B(n8194), .Z(n8196) );
  NAND U7040 ( .A(n1436), .B(n1435), .Z(n1440) );
  NAND U7041 ( .A(n1438), .B(n1437), .Z(n1439) );
  AND U7042 ( .A(n1440), .B(n1439), .Z(n8195) );
  XOR U7043 ( .A(n8196), .B(n8195), .Z(n6428) );
  NANDN U7044 ( .A(n1442), .B(n1441), .Z(n1446) );
  NAND U7045 ( .A(n1444), .B(n1443), .Z(n1445) );
  AND U7046 ( .A(n1446), .B(n1445), .Z(n8163) );
  NAND U7047 ( .A(n1448), .B(n1447), .Z(n1452) );
  NAND U7048 ( .A(n1450), .B(n1449), .Z(n1451) );
  NAND U7049 ( .A(n1452), .B(n1451), .Z(n8164) );
  XNOR U7050 ( .A(n8163), .B(n8164), .Z(n8166) );
  NANDN U7051 ( .A(n1454), .B(n1453), .Z(n1458) );
  NAND U7052 ( .A(n1456), .B(n1455), .Z(n1457) );
  AND U7053 ( .A(n1458), .B(n1457), .Z(n8165) );
  XOR U7054 ( .A(n8166), .B(n8165), .Z(n6427) );
  NANDN U7055 ( .A(n1460), .B(n1459), .Z(n1464) );
  NANDN U7056 ( .A(n1462), .B(n1461), .Z(n1463) );
  AND U7057 ( .A(n1464), .B(n1463), .Z(n6426) );
  XOR U7058 ( .A(n6427), .B(n6426), .Z(n6429) );
  XOR U7059 ( .A(n6428), .B(n6429), .Z(n6133) );
  NANDN U7060 ( .A(n1466), .B(n1465), .Z(n1470) );
  NAND U7061 ( .A(n1468), .B(n1467), .Z(n1469) );
  NAND U7062 ( .A(n1470), .B(n1469), .Z(n6132) );
  XOR U7063 ( .A(n6133), .B(n6132), .Z(n6135) );
  XOR U7064 ( .A(n6134), .B(n6135), .Z(n6086) );
  NANDN U7065 ( .A(n1472), .B(n1471), .Z(n1476) );
  NAND U7066 ( .A(n1474), .B(n1473), .Z(n1475) );
  AND U7067 ( .A(n1476), .B(n1475), .Z(n6122) );
  NANDN U7068 ( .A(n1478), .B(n1477), .Z(n1482) );
  NAND U7069 ( .A(n1480), .B(n1479), .Z(n1481) );
  AND U7070 ( .A(n1482), .B(n1481), .Z(n6871) );
  NANDN U7071 ( .A(n1484), .B(n1483), .Z(n1488) );
  NAND U7072 ( .A(n1486), .B(n1485), .Z(n1487) );
  AND U7073 ( .A(n1488), .B(n1487), .Z(n6870) );
  XOR U7074 ( .A(n6871), .B(n6870), .Z(n6873) );
  NANDN U7075 ( .A(n1490), .B(n1489), .Z(n1494) );
  NAND U7076 ( .A(n1492), .B(n1491), .Z(n1493) );
  AND U7077 ( .A(n1494), .B(n1493), .Z(n6872) );
  XOR U7078 ( .A(n6873), .B(n6872), .Z(n6482) );
  NANDN U7079 ( .A(n1496), .B(n1495), .Z(n1500) );
  NAND U7080 ( .A(n1498), .B(n1497), .Z(n1499) );
  AND U7081 ( .A(n1500), .B(n1499), .Z(n8062) );
  NANDN U7082 ( .A(n1502), .B(n1501), .Z(n1506) );
  NAND U7083 ( .A(n1504), .B(n1503), .Z(n1505) );
  AND U7084 ( .A(n1506), .B(n1505), .Z(n8061) );
  XOR U7085 ( .A(n8062), .B(n8061), .Z(n8064) );
  NANDN U7086 ( .A(n1508), .B(n1507), .Z(n1512) );
  NAND U7087 ( .A(n1510), .B(n1509), .Z(n1511) );
  AND U7088 ( .A(n1512), .B(n1511), .Z(n8063) );
  XOR U7089 ( .A(n8064), .B(n8063), .Z(n6481) );
  NANDN U7090 ( .A(n1514), .B(n1513), .Z(n1518) );
  NANDN U7091 ( .A(n1516), .B(n1515), .Z(n1517) );
  AND U7092 ( .A(n1518), .B(n1517), .Z(n6480) );
  XOR U7093 ( .A(n6481), .B(n6480), .Z(n6483) );
  XOR U7094 ( .A(n6482), .B(n6483), .Z(n6121) );
  NANDN U7095 ( .A(n1520), .B(n1519), .Z(n1524) );
  NAND U7096 ( .A(n1522), .B(n1521), .Z(n1523) );
  NAND U7097 ( .A(n1524), .B(n1523), .Z(n6120) );
  XOR U7098 ( .A(n6121), .B(n6120), .Z(n6123) );
  XOR U7099 ( .A(n6122), .B(n6123), .Z(n6085) );
  NANDN U7100 ( .A(n1526), .B(n1525), .Z(n1530) );
  NANDN U7101 ( .A(n1528), .B(n1527), .Z(n1529) );
  AND U7102 ( .A(n1530), .B(n1529), .Z(n6084) );
  XOR U7103 ( .A(n6085), .B(n6084), .Z(n6087) );
  XNOR U7104 ( .A(n6086), .B(n6087), .Z(n8874) );
  NANDN U7105 ( .A(n1532), .B(n1531), .Z(n1536) );
  NANDN U7106 ( .A(n1534), .B(n1533), .Z(n1535) );
  AND U7107 ( .A(n1536), .B(n1535), .Z(n6237) );
  NANDN U7108 ( .A(n1538), .B(n1537), .Z(n1542) );
  NANDN U7109 ( .A(n1540), .B(n1539), .Z(n1541) );
  AND U7110 ( .A(n1542), .B(n1541), .Z(n7195) );
  NANDN U7111 ( .A(n1544), .B(n1543), .Z(n1548) );
  NAND U7112 ( .A(n1546), .B(n1545), .Z(n1547) );
  AND U7113 ( .A(n1548), .B(n1547), .Z(n8421) );
  NANDN U7114 ( .A(n1550), .B(n1549), .Z(n1554) );
  NAND U7115 ( .A(n1552), .B(n1551), .Z(n1553) );
  NAND U7116 ( .A(n1554), .B(n1553), .Z(n8422) );
  XNOR U7117 ( .A(n8421), .B(n8422), .Z(n8424) );
  NANDN U7118 ( .A(n1556), .B(n1555), .Z(n1560) );
  NAND U7119 ( .A(n1558), .B(n1557), .Z(n1559) );
  AND U7120 ( .A(n1560), .B(n1559), .Z(n8423) );
  XOR U7121 ( .A(n8424), .B(n8423), .Z(n7193) );
  NANDN U7122 ( .A(n1562), .B(n1561), .Z(n1566) );
  NANDN U7123 ( .A(n1564), .B(n1563), .Z(n1565) );
  AND U7124 ( .A(n1566), .B(n1565), .Z(n7192) );
  XNOR U7125 ( .A(n7193), .B(n7192), .Z(n7194) );
  XOR U7126 ( .A(n7195), .B(n7194), .Z(n6235) );
  NANDN U7127 ( .A(n1568), .B(n1567), .Z(n1572) );
  NAND U7128 ( .A(n1570), .B(n1569), .Z(n1571) );
  NAND U7129 ( .A(n1572), .B(n1571), .Z(n6234) );
  XNOR U7130 ( .A(n6235), .B(n6234), .Z(n6236) );
  XNOR U7131 ( .A(n6237), .B(n6236), .Z(n7267) );
  NANDN U7132 ( .A(n1574), .B(n1573), .Z(n1578) );
  NANDN U7133 ( .A(n1576), .B(n1575), .Z(n1577) );
  AND U7134 ( .A(n1578), .B(n1577), .Z(n8256) );
  NANDN U7135 ( .A(n1580), .B(n1579), .Z(n1584) );
  NAND U7136 ( .A(n1582), .B(n1581), .Z(n1583) );
  AND U7137 ( .A(n1584), .B(n1583), .Z(n8386) );
  NANDN U7138 ( .A(n1586), .B(n1585), .Z(n1590) );
  NAND U7139 ( .A(n1588), .B(n1587), .Z(n1589) );
  AND U7140 ( .A(n1590), .B(n1589), .Z(n8385) );
  XOR U7141 ( .A(n8386), .B(n8385), .Z(n8388) );
  NANDN U7142 ( .A(n1592), .B(n1591), .Z(n1596) );
  NAND U7143 ( .A(n1594), .B(n1593), .Z(n1595) );
  AND U7144 ( .A(n1596), .B(n1595), .Z(n8387) );
  XOR U7145 ( .A(n8388), .B(n8387), .Z(n8254) );
  NANDN U7146 ( .A(n1598), .B(n1597), .Z(n1602) );
  NANDN U7147 ( .A(n1600), .B(n1599), .Z(n1601) );
  AND U7148 ( .A(n1602), .B(n1601), .Z(n8253) );
  XNOR U7149 ( .A(n8254), .B(n8253), .Z(n8255) );
  XOR U7150 ( .A(n8256), .B(n8255), .Z(n6159) );
  NANDN U7151 ( .A(n1604), .B(n1603), .Z(n1608) );
  NANDN U7152 ( .A(n1606), .B(n1605), .Z(n1607) );
  AND U7153 ( .A(n1608), .B(n1607), .Z(n7219) );
  NANDN U7154 ( .A(n1610), .B(n1609), .Z(n1614) );
  NAND U7155 ( .A(n1612), .B(n1611), .Z(n1613) );
  AND U7156 ( .A(n1614), .B(n1613), .Z(n8397) );
  NANDN U7157 ( .A(n1616), .B(n1615), .Z(n1620) );
  NAND U7158 ( .A(n1618), .B(n1617), .Z(n1619) );
  NAND U7159 ( .A(n1620), .B(n1619), .Z(n8398) );
  XNOR U7160 ( .A(n8397), .B(n8398), .Z(n8400) );
  NAND U7161 ( .A(n1622), .B(n1621), .Z(n1626) );
  NAND U7162 ( .A(n1624), .B(n1623), .Z(n1625) );
  AND U7163 ( .A(n1626), .B(n1625), .Z(n8399) );
  XOR U7164 ( .A(n8400), .B(n8399), .Z(n7217) );
  NANDN U7165 ( .A(n1628), .B(n1627), .Z(n1632) );
  OR U7166 ( .A(n1630), .B(n1629), .Z(n1631) );
  AND U7167 ( .A(n1632), .B(n1631), .Z(n7216) );
  XNOR U7168 ( .A(n7217), .B(n7216), .Z(n7218) );
  XOR U7169 ( .A(n7219), .B(n7218), .Z(n6157) );
  NANDN U7170 ( .A(n1634), .B(n1633), .Z(n1638) );
  NAND U7171 ( .A(n1636), .B(n1635), .Z(n1637) );
  AND U7172 ( .A(n1638), .B(n1637), .Z(n7170) );
  NANDN U7173 ( .A(n1640), .B(n1639), .Z(n1644) );
  NAND U7174 ( .A(n1642), .B(n1641), .Z(n1643) );
  AND U7175 ( .A(n1644), .B(n1643), .Z(n6876) );
  NANDN U7176 ( .A(n1646), .B(n1645), .Z(n1650) );
  NAND U7177 ( .A(n1648), .B(n1647), .Z(n1649) );
  NAND U7178 ( .A(n1650), .B(n1649), .Z(n6877) );
  XNOR U7179 ( .A(n6876), .B(n6877), .Z(n6879) );
  NANDN U7180 ( .A(n1652), .B(n1651), .Z(n1656) );
  NAND U7181 ( .A(n1654), .B(n1653), .Z(n1655) );
  AND U7182 ( .A(n1656), .B(n1655), .Z(n6878) );
  XOR U7183 ( .A(n6879), .B(n6878), .Z(n7169) );
  NANDN U7184 ( .A(n1658), .B(n1657), .Z(n1662) );
  NANDN U7185 ( .A(n1660), .B(n1659), .Z(n1661) );
  AND U7186 ( .A(n1662), .B(n1661), .Z(n7168) );
  XOR U7187 ( .A(n7169), .B(n7168), .Z(n7171) );
  XNOR U7188 ( .A(n7170), .B(n7171), .Z(n6156) );
  XNOR U7189 ( .A(n6157), .B(n6156), .Z(n6158) );
  XNOR U7190 ( .A(n6159), .B(n6158), .Z(n7265) );
  NANDN U7191 ( .A(n1664), .B(n1663), .Z(n1668) );
  NANDN U7192 ( .A(n1666), .B(n1665), .Z(n1667) );
  AND U7193 ( .A(n1668), .B(n1667), .Z(n7920) );
  NANDN U7194 ( .A(n1670), .B(n1669), .Z(n1674) );
  NAND U7195 ( .A(n1672), .B(n1671), .Z(n1673) );
  AND U7196 ( .A(n1674), .B(n1673), .Z(n8571) );
  NANDN U7197 ( .A(n1676), .B(n1675), .Z(n1680) );
  NAND U7198 ( .A(n1678), .B(n1677), .Z(n1679) );
  NAND U7199 ( .A(n1680), .B(n1679), .Z(n8572) );
  XNOR U7200 ( .A(n8571), .B(n8572), .Z(n8574) );
  NANDN U7201 ( .A(n1682), .B(n1681), .Z(n1686) );
  NAND U7202 ( .A(n1684), .B(n1683), .Z(n1685) );
  AND U7203 ( .A(n1686), .B(n1685), .Z(n8573) );
  XOR U7204 ( .A(n8574), .B(n8573), .Z(n7918) );
  NANDN U7205 ( .A(n1688), .B(n1687), .Z(n1692) );
  NANDN U7206 ( .A(n1690), .B(n1689), .Z(n1691) );
  AND U7207 ( .A(n1692), .B(n1691), .Z(n7917) );
  XNOR U7208 ( .A(n7918), .B(n7917), .Z(n7919) );
  XOR U7209 ( .A(n7920), .B(n7919), .Z(n6153) );
  NANDN U7210 ( .A(n1694), .B(n1693), .Z(n1698) );
  NANDN U7211 ( .A(n1696), .B(n1695), .Z(n1697) );
  AND U7212 ( .A(n1698), .B(n1697), .Z(n7177) );
  NANDN U7213 ( .A(n1700), .B(n1699), .Z(n1704) );
  NAND U7214 ( .A(n1702), .B(n1701), .Z(n1703) );
  AND U7215 ( .A(n1704), .B(n1703), .Z(n8523) );
  NANDN U7216 ( .A(n1706), .B(n1705), .Z(n1710) );
  NAND U7217 ( .A(n1708), .B(n1707), .Z(n1709) );
  NAND U7218 ( .A(n1710), .B(n1709), .Z(n8524) );
  XNOR U7219 ( .A(n8523), .B(n8524), .Z(n8526) );
  NAND U7220 ( .A(n1712), .B(n1711), .Z(n1716) );
  NAND U7221 ( .A(n1714), .B(n1713), .Z(n1715) );
  AND U7222 ( .A(n1716), .B(n1715), .Z(n8525) );
  XOR U7223 ( .A(n8526), .B(n8525), .Z(n7175) );
  NANDN U7224 ( .A(n1718), .B(n1717), .Z(n1722) );
  NANDN U7225 ( .A(n1720), .B(n1719), .Z(n1721) );
  AND U7226 ( .A(n1722), .B(n1721), .Z(n7174) );
  XNOR U7227 ( .A(n7175), .B(n7174), .Z(n7176) );
  XOR U7228 ( .A(n7177), .B(n7176), .Z(n6151) );
  NANDN U7229 ( .A(n1724), .B(n1723), .Z(n1728) );
  NAND U7230 ( .A(n1726), .B(n1725), .Z(n1727) );
  NAND U7231 ( .A(n1728), .B(n1727), .Z(n6150) );
  XNOR U7232 ( .A(n6151), .B(n6150), .Z(n6152) );
  XNOR U7233 ( .A(n6153), .B(n6152), .Z(n7264) );
  XOR U7234 ( .A(n7265), .B(n7264), .Z(n7266) );
  XOR U7235 ( .A(n7267), .B(n7266), .Z(n8872) );
  NANDN U7236 ( .A(n1730), .B(n1729), .Z(n1734) );
  NAND U7237 ( .A(n1732), .B(n1731), .Z(n1733) );
  AND U7238 ( .A(n1734), .B(n1733), .Z(n6099) );
  NANDN U7239 ( .A(n1736), .B(n1735), .Z(n1740) );
  NANDN U7240 ( .A(n1738), .B(n1737), .Z(n1739) );
  AND U7241 ( .A(n1740), .B(n1739), .Z(n6459) );
  NANDN U7242 ( .A(n1742), .B(n1741), .Z(n1746) );
  NAND U7243 ( .A(n1744), .B(n1743), .Z(n1745) );
  AND U7244 ( .A(n1746), .B(n1745), .Z(n8098) );
  NANDN U7245 ( .A(n1748), .B(n1747), .Z(n1752) );
  NAND U7246 ( .A(n1750), .B(n1749), .Z(n1751) );
  AND U7247 ( .A(n1752), .B(n1751), .Z(n8097) );
  XOR U7248 ( .A(n8098), .B(n8097), .Z(n8100) );
  NANDN U7249 ( .A(n1754), .B(n1753), .Z(n1758) );
  NAND U7250 ( .A(n1756), .B(n1755), .Z(n1757) );
  AND U7251 ( .A(n1758), .B(n1757), .Z(n8099) );
  XOR U7252 ( .A(n8100), .B(n8099), .Z(n6457) );
  NANDN U7253 ( .A(n1760), .B(n1759), .Z(n1764) );
  NANDN U7254 ( .A(n1762), .B(n1761), .Z(n1763) );
  AND U7255 ( .A(n1764), .B(n1763), .Z(n6456) );
  XNOR U7256 ( .A(n6457), .B(n6456), .Z(n6458) );
  XOR U7257 ( .A(n6459), .B(n6458), .Z(n6097) );
  NANDN U7258 ( .A(n1766), .B(n1765), .Z(n1770) );
  NAND U7259 ( .A(n1768), .B(n1767), .Z(n1769) );
  NAND U7260 ( .A(n1770), .B(n1769), .Z(n6096) );
  XNOR U7261 ( .A(n6097), .B(n6096), .Z(n6098) );
  XNOR U7262 ( .A(n6099), .B(n6098), .Z(n7278) );
  NANDN U7263 ( .A(n1776), .B(n1775), .Z(n1780) );
  NANDN U7264 ( .A(n1778), .B(n1777), .Z(n1779) );
  AND U7265 ( .A(n1780), .B(n1779), .Z(n7719) );
  NANDN U7266 ( .A(n1782), .B(n1781), .Z(n1786) );
  NANDN U7267 ( .A(n1784), .B(n1783), .Z(n1785) );
  AND U7268 ( .A(n1786), .B(n1785), .Z(n6350) );
  NANDN U7269 ( .A(n1788), .B(n1787), .Z(n1792) );
  NAND U7270 ( .A(n1790), .B(n1789), .Z(n1791) );
  AND U7271 ( .A(n1792), .B(n1791), .Z(n8085) );
  NAND U7272 ( .A(n1794), .B(n1793), .Z(n1798) );
  NAND U7273 ( .A(n1796), .B(n1795), .Z(n1797) );
  NAND U7274 ( .A(n1798), .B(n1797), .Z(n8086) );
  XNOR U7275 ( .A(n8085), .B(n8086), .Z(n8087) );
  NAND U7276 ( .A(n1800), .B(n1799), .Z(n1804) );
  NAND U7277 ( .A(n1802), .B(n1801), .Z(n1803) );
  NAND U7278 ( .A(n1804), .B(n1803), .Z(n8088) );
  XOR U7279 ( .A(n8087), .B(n8088), .Z(n6348) );
  NANDN U7280 ( .A(n1806), .B(n1805), .Z(n1810) );
  NANDN U7281 ( .A(n1808), .B(n1807), .Z(n1809) );
  AND U7282 ( .A(n1810), .B(n1809), .Z(n6349) );
  XOR U7283 ( .A(n6348), .B(n6349), .Z(n6351) );
  XOR U7284 ( .A(n6350), .B(n6351), .Z(n7718) );
  XOR U7285 ( .A(n7719), .B(n7718), .Z(n7720) );
  XNOR U7286 ( .A(n7721), .B(n7720), .Z(n7277) );
  NANDN U7287 ( .A(n1812), .B(n1811), .Z(n1816) );
  NAND U7288 ( .A(n1814), .B(n1813), .Z(n1815) );
  AND U7289 ( .A(n1816), .B(n1815), .Z(n6110) );
  NANDN U7290 ( .A(n1818), .B(n1817), .Z(n1822) );
  NANDN U7291 ( .A(n1820), .B(n1819), .Z(n1821) );
  AND U7292 ( .A(n1822), .B(n1821), .Z(n8939) );
  NANDN U7293 ( .A(n1824), .B(n1823), .Z(n1828) );
  NAND U7294 ( .A(n1826), .B(n1825), .Z(n1827) );
  AND U7295 ( .A(n1828), .B(n1827), .Z(n8079) );
  NAND U7296 ( .A(n1830), .B(n1829), .Z(n1834) );
  NAND U7297 ( .A(n1832), .B(n1831), .Z(n1833) );
  NAND U7298 ( .A(n1834), .B(n1833), .Z(n8080) );
  XNOR U7299 ( .A(n8079), .B(n8080), .Z(n8082) );
  NAND U7300 ( .A(n1836), .B(n1835), .Z(n1840) );
  NAND U7301 ( .A(n1838), .B(n1837), .Z(n1839) );
  AND U7302 ( .A(n1840), .B(n1839), .Z(n8081) );
  XOR U7303 ( .A(n8082), .B(n8081), .Z(n8937) );
  NANDN U7304 ( .A(n1842), .B(n1841), .Z(n1846) );
  NANDN U7305 ( .A(n1844), .B(n1843), .Z(n1845) );
  AND U7306 ( .A(n1846), .B(n1845), .Z(n8936) );
  XNOR U7307 ( .A(n8937), .B(n8936), .Z(n8938) );
  XOR U7308 ( .A(n8939), .B(n8938), .Z(n6109) );
  NANDN U7309 ( .A(n1848), .B(n1847), .Z(n1852) );
  NAND U7310 ( .A(n1850), .B(n1849), .Z(n1851) );
  NAND U7311 ( .A(n1852), .B(n1851), .Z(n6108) );
  XOR U7312 ( .A(n6109), .B(n6108), .Z(n6111) );
  XOR U7313 ( .A(n6110), .B(n6111), .Z(n7276) );
  XNOR U7314 ( .A(n7277), .B(n7276), .Z(n7279) );
  XNOR U7315 ( .A(n7278), .B(n7279), .Z(n8871) );
  XOR U7316 ( .A(n8872), .B(n8871), .Z(n8873) );
  XNOR U7317 ( .A(n8874), .B(n8873), .Z(n7050) );
  NANDN U7318 ( .A(n1854), .B(n1853), .Z(n1858) );
  NANDN U7319 ( .A(n1856), .B(n1855), .Z(n1857) );
  AND U7320 ( .A(n1858), .B(n1857), .Z(n6452) );
  NANDN U7321 ( .A(n1860), .B(n1859), .Z(n1864) );
  NAND U7322 ( .A(n1862), .B(n1861), .Z(n1863) );
  AND U7323 ( .A(n1864), .B(n1863), .Z(n8104) );
  NANDN U7324 ( .A(n1866), .B(n1865), .Z(n1870) );
  NAND U7325 ( .A(n1868), .B(n1867), .Z(n1869) );
  AND U7326 ( .A(n1870), .B(n1869), .Z(n8103) );
  XOR U7327 ( .A(n8104), .B(n8103), .Z(n8106) );
  NANDN U7328 ( .A(n1872), .B(n1871), .Z(n1876) );
  NAND U7329 ( .A(n1874), .B(n1873), .Z(n1875) );
  AND U7330 ( .A(n1876), .B(n1875), .Z(n8105) );
  XOR U7331 ( .A(n8106), .B(n8105), .Z(n6451) );
  NANDN U7332 ( .A(n1878), .B(n1877), .Z(n1882) );
  NANDN U7333 ( .A(n1880), .B(n1879), .Z(n1881) );
  AND U7334 ( .A(n1882), .B(n1881), .Z(n6450) );
  XOR U7335 ( .A(n6451), .B(n6450), .Z(n6453) );
  XNOR U7336 ( .A(n6452), .B(n6453), .Z(n6282) );
  NANDN U7337 ( .A(n1884), .B(n1883), .Z(n1888) );
  NAND U7338 ( .A(n1886), .B(n1885), .Z(n1887) );
  AND U7339 ( .A(n1888), .B(n1887), .Z(n9051) );
  NANDN U7340 ( .A(n1890), .B(n1889), .Z(n1894) );
  NAND U7341 ( .A(n1892), .B(n1891), .Z(n1893) );
  NAND U7342 ( .A(n1894), .B(n1893), .Z(n9052) );
  XNOR U7343 ( .A(n9051), .B(n9052), .Z(n9054) );
  NANDN U7344 ( .A(n1896), .B(n1895), .Z(n1900) );
  NAND U7345 ( .A(n1898), .B(n1897), .Z(n1899) );
  AND U7346 ( .A(n1900), .B(n1899), .Z(n9053) );
  XOR U7347 ( .A(n9054), .B(n9053), .Z(n8604) );
  NANDN U7348 ( .A(n1902), .B(n1901), .Z(n1906) );
  NAND U7349 ( .A(n1904), .B(n1903), .Z(n1905) );
  AND U7350 ( .A(n1906), .B(n1905), .Z(n9045) );
  NANDN U7351 ( .A(n1908), .B(n1907), .Z(n1912) );
  NAND U7352 ( .A(n1910), .B(n1909), .Z(n1911) );
  NAND U7353 ( .A(n1912), .B(n1911), .Z(n9046) );
  XNOR U7354 ( .A(n9045), .B(n9046), .Z(n9048) );
  NANDN U7355 ( .A(n1914), .B(n1913), .Z(n1918) );
  NAND U7356 ( .A(n1916), .B(n1915), .Z(n1917) );
  AND U7357 ( .A(n1918), .B(n1917), .Z(n9047) );
  XOR U7358 ( .A(n9048), .B(n9047), .Z(n8602) );
  NANDN U7359 ( .A(n1920), .B(n1919), .Z(n1924) );
  NANDN U7360 ( .A(n1922), .B(n1921), .Z(n1923) );
  AND U7361 ( .A(n1924), .B(n1923), .Z(n8601) );
  XNOR U7362 ( .A(n8602), .B(n8601), .Z(n8603) );
  XOR U7363 ( .A(n8604), .B(n8603), .Z(n6283) );
  XNOR U7364 ( .A(n6282), .B(n6283), .Z(n6285) );
  NANDN U7365 ( .A(n1926), .B(n1925), .Z(n1930) );
  NAND U7366 ( .A(n1928), .B(n1927), .Z(n1929) );
  AND U7367 ( .A(n1930), .B(n1929), .Z(n6928) );
  NANDN U7368 ( .A(n1932), .B(n1931), .Z(n1936) );
  NAND U7369 ( .A(n1934), .B(n1933), .Z(n1935) );
  NAND U7370 ( .A(n1936), .B(n1935), .Z(n6929) );
  XNOR U7371 ( .A(n6928), .B(n6929), .Z(n6931) );
  NANDN U7372 ( .A(n1938), .B(n1937), .Z(n1942) );
  NAND U7373 ( .A(n1940), .B(n1939), .Z(n1941) );
  AND U7374 ( .A(n1942), .B(n1941), .Z(n6930) );
  XOR U7375 ( .A(n6931), .B(n6930), .Z(n8610) );
  NANDN U7376 ( .A(n1944), .B(n1943), .Z(n1948) );
  NAND U7377 ( .A(n1946), .B(n1945), .Z(n1947) );
  AND U7378 ( .A(n1948), .B(n1947), .Z(n6916) );
  NANDN U7379 ( .A(n1950), .B(n1949), .Z(n1954) );
  NAND U7380 ( .A(n1952), .B(n1951), .Z(n1953) );
  NAND U7381 ( .A(n1954), .B(n1953), .Z(n6917) );
  XNOR U7382 ( .A(n6916), .B(n6917), .Z(n6919) );
  NANDN U7383 ( .A(n1956), .B(n1955), .Z(n1960) );
  NAND U7384 ( .A(n1958), .B(n1957), .Z(n1959) );
  AND U7385 ( .A(n1960), .B(n1959), .Z(n6918) );
  XOR U7386 ( .A(n6919), .B(n6918), .Z(n8608) );
  NANDN U7387 ( .A(n1962), .B(n1961), .Z(n1966) );
  NANDN U7388 ( .A(n1964), .B(n1963), .Z(n1965) );
  AND U7389 ( .A(n1966), .B(n1965), .Z(n8607) );
  XNOR U7390 ( .A(n8608), .B(n8607), .Z(n8609) );
  XNOR U7391 ( .A(n8610), .B(n8609), .Z(n6284) );
  XOR U7392 ( .A(n6285), .B(n6284), .Z(n6183) );
  NANDN U7393 ( .A(n1968), .B(n1967), .Z(n1972) );
  NANDN U7394 ( .A(n1970), .B(n1969), .Z(n1971) );
  AND U7395 ( .A(n1972), .B(n1971), .Z(n8448) );
  NANDN U7396 ( .A(n1974), .B(n1973), .Z(n1978) );
  NAND U7397 ( .A(n1976), .B(n1975), .Z(n1977) );
  AND U7398 ( .A(n1978), .B(n1977), .Z(n7594) );
  NAND U7399 ( .A(n1980), .B(n1979), .Z(n1984) );
  NAND U7400 ( .A(n1982), .B(n1981), .Z(n1983) );
  NAND U7401 ( .A(n1984), .B(n1983), .Z(n7595) );
  XNOR U7402 ( .A(n7594), .B(n7595), .Z(n7597) );
  NAND U7403 ( .A(n1986), .B(n1985), .Z(n1990) );
  NAND U7404 ( .A(n1988), .B(n1987), .Z(n1989) );
  AND U7405 ( .A(n1990), .B(n1989), .Z(n7596) );
  XOR U7406 ( .A(n7597), .B(n7596), .Z(n8446) );
  NANDN U7407 ( .A(n1992), .B(n1991), .Z(n1996) );
  NANDN U7408 ( .A(n1994), .B(n1993), .Z(n1995) );
  AND U7409 ( .A(n1996), .B(n1995), .Z(n8445) );
  XNOR U7410 ( .A(n8446), .B(n8445), .Z(n8447) );
  XOR U7411 ( .A(n8448), .B(n8447), .Z(n7779) );
  NANDN U7412 ( .A(n1998), .B(n1997), .Z(n2002) );
  NANDN U7413 ( .A(n2000), .B(n1999), .Z(n2001) );
  AND U7414 ( .A(n2002), .B(n2001), .Z(n8442) );
  NANDN U7415 ( .A(n2004), .B(n2003), .Z(n2008) );
  NAND U7416 ( .A(n2006), .B(n2005), .Z(n2007) );
  AND U7417 ( .A(n2008), .B(n2007), .Z(n7456) );
  NAND U7418 ( .A(n2010), .B(n2009), .Z(n2014) );
  NAND U7419 ( .A(n2012), .B(n2011), .Z(n2013) );
  NAND U7420 ( .A(n2014), .B(n2013), .Z(n7457) );
  XNOR U7421 ( .A(n7456), .B(n7457), .Z(n7459) );
  NANDN U7422 ( .A(n2016), .B(n2015), .Z(n2020) );
  NAND U7423 ( .A(n2018), .B(n2017), .Z(n2019) );
  AND U7424 ( .A(n2020), .B(n2019), .Z(n7458) );
  XOR U7425 ( .A(n7459), .B(n7458), .Z(n8440) );
  NANDN U7426 ( .A(n2022), .B(n2021), .Z(n2026) );
  NANDN U7427 ( .A(n2024), .B(n2023), .Z(n2025) );
  AND U7428 ( .A(n2026), .B(n2025), .Z(n8439) );
  XNOR U7429 ( .A(n8440), .B(n8439), .Z(n8441) );
  XOR U7430 ( .A(n8442), .B(n8441), .Z(n7777) );
  NANDN U7431 ( .A(n2028), .B(n2027), .Z(n2032) );
  NANDN U7432 ( .A(n2030), .B(n2029), .Z(n2031) );
  AND U7433 ( .A(n2032), .B(n2031), .Z(n8334) );
  NANDN U7434 ( .A(n2034), .B(n2033), .Z(n2038) );
  NANDN U7435 ( .A(n2036), .B(n2035), .Z(n2037) );
  AND U7436 ( .A(n2038), .B(n2037), .Z(n7450) );
  NANDN U7437 ( .A(n2040), .B(n2039), .Z(n2044) );
  NAND U7438 ( .A(n2042), .B(n2041), .Z(n2043) );
  NAND U7439 ( .A(n2044), .B(n2043), .Z(n7451) );
  XNOR U7440 ( .A(n7450), .B(n7451), .Z(n7453) );
  NANDN U7441 ( .A(n2046), .B(n2045), .Z(n2050) );
  NAND U7442 ( .A(n2048), .B(n2047), .Z(n2049) );
  AND U7443 ( .A(n2050), .B(n2049), .Z(n7452) );
  XOR U7444 ( .A(n7453), .B(n7452), .Z(n8332) );
  NANDN U7445 ( .A(n2052), .B(n2051), .Z(n2056) );
  NANDN U7446 ( .A(n2054), .B(n2053), .Z(n2055) );
  AND U7447 ( .A(n2056), .B(n2055), .Z(n8331) );
  XNOR U7448 ( .A(n8332), .B(n8331), .Z(n8333) );
  XNOR U7449 ( .A(n8334), .B(n8333), .Z(n7776) );
  XNOR U7450 ( .A(n7777), .B(n7776), .Z(n7778) );
  XNOR U7451 ( .A(n7779), .B(n7778), .Z(n6180) );
  NANDN U7452 ( .A(n2058), .B(n2057), .Z(n2062) );
  NANDN U7453 ( .A(n2060), .B(n2059), .Z(n2061) );
  AND U7454 ( .A(n2062), .B(n2061), .Z(n6423) );
  NANDN U7455 ( .A(n2064), .B(n2063), .Z(n2068) );
  NAND U7456 ( .A(n2066), .B(n2065), .Z(n2067) );
  AND U7457 ( .A(n2068), .B(n2067), .Z(n7468) );
  NANDN U7458 ( .A(n2070), .B(n2069), .Z(n2074) );
  NAND U7459 ( .A(n2072), .B(n2071), .Z(n2073) );
  NAND U7460 ( .A(n2074), .B(n2073), .Z(n7469) );
  XNOR U7461 ( .A(n7468), .B(n7469), .Z(n7471) );
  NANDN U7462 ( .A(n2076), .B(n2075), .Z(n2080) );
  NAND U7463 ( .A(n2078), .B(n2077), .Z(n2079) );
  AND U7464 ( .A(n2080), .B(n2079), .Z(n7470) );
  XOR U7465 ( .A(n7471), .B(n7470), .Z(n6421) );
  NANDN U7466 ( .A(n2082), .B(n2081), .Z(n2086) );
  NANDN U7467 ( .A(n2084), .B(n2083), .Z(n2085) );
  AND U7468 ( .A(n2086), .B(n2085), .Z(n6420) );
  XNOR U7469 ( .A(n6421), .B(n6420), .Z(n6422) );
  XOR U7470 ( .A(n6423), .B(n6422), .Z(n7845) );
  NANDN U7471 ( .A(n2088), .B(n2087), .Z(n2092) );
  NANDN U7472 ( .A(n2090), .B(n2089), .Z(n2091) );
  AND U7473 ( .A(n2092), .B(n2091), .Z(n8850) );
  NANDN U7474 ( .A(n2094), .B(n2093), .Z(n2098) );
  NAND U7475 ( .A(n2096), .B(n2095), .Z(n2097) );
  AND U7476 ( .A(n2098), .B(n2097), .Z(n8973) );
  NAND U7477 ( .A(n2100), .B(n2099), .Z(n2104) );
  NAND U7478 ( .A(n2102), .B(n2101), .Z(n2103) );
  NAND U7479 ( .A(n2104), .B(n2103), .Z(n8974) );
  XNOR U7480 ( .A(n8973), .B(n8974), .Z(n8976) );
  NAND U7481 ( .A(n2106), .B(n2105), .Z(n2110) );
  NAND U7482 ( .A(n2108), .B(n2107), .Z(n2109) );
  AND U7483 ( .A(n2110), .B(n2109), .Z(n8975) );
  XOR U7484 ( .A(n8976), .B(n8975), .Z(n8848) );
  NANDN U7485 ( .A(n2112), .B(n2111), .Z(n2116) );
  NANDN U7486 ( .A(n2114), .B(n2113), .Z(n2115) );
  AND U7487 ( .A(n2116), .B(n2115), .Z(n8847) );
  XNOR U7488 ( .A(n8848), .B(n8847), .Z(n8849) );
  XOR U7489 ( .A(n8850), .B(n8849), .Z(n7843) );
  NANDN U7490 ( .A(n2118), .B(n2117), .Z(n2122) );
  NANDN U7491 ( .A(n2120), .B(n2119), .Z(n2121) );
  AND U7492 ( .A(n2122), .B(n2121), .Z(n8658) );
  NANDN U7493 ( .A(n2124), .B(n2123), .Z(n2128) );
  NAND U7494 ( .A(n2126), .B(n2125), .Z(n2127) );
  AND U7495 ( .A(n2128), .B(n2127), .Z(n6768) );
  NAND U7496 ( .A(n2130), .B(n2129), .Z(n2134) );
  NAND U7497 ( .A(n2132), .B(n2131), .Z(n2133) );
  NAND U7498 ( .A(n2134), .B(n2133), .Z(n6769) );
  XNOR U7499 ( .A(n6768), .B(n6769), .Z(n6771) );
  NAND U7500 ( .A(n2136), .B(n2135), .Z(n2140) );
  NAND U7501 ( .A(n2138), .B(n2137), .Z(n2139) );
  AND U7502 ( .A(n2140), .B(n2139), .Z(n6770) );
  XOR U7503 ( .A(n6771), .B(n6770), .Z(n8656) );
  NANDN U7504 ( .A(n2142), .B(n2141), .Z(n2146) );
  NANDN U7505 ( .A(n2144), .B(n2143), .Z(n2145) );
  AND U7506 ( .A(n2146), .B(n2145), .Z(n8655) );
  XNOR U7507 ( .A(n8656), .B(n8655), .Z(n8657) );
  XNOR U7508 ( .A(n8658), .B(n8657), .Z(n7842) );
  XNOR U7509 ( .A(n7843), .B(n7842), .Z(n7844) );
  XOR U7510 ( .A(n7845), .B(n7844), .Z(n6181) );
  XNOR U7511 ( .A(n6180), .B(n6181), .Z(n6182) );
  XNOR U7512 ( .A(n6183), .B(n6182), .Z(n8643) );
  NANDN U7513 ( .A(n2148), .B(n2147), .Z(n2152) );
  NANDN U7514 ( .A(n2150), .B(n2149), .Z(n2151) );
  AND U7515 ( .A(n2152), .B(n2151), .Z(n8124) );
  NANDN U7516 ( .A(n2154), .B(n2153), .Z(n2158) );
  NAND U7517 ( .A(n2156), .B(n2155), .Z(n2157) );
  AND U7518 ( .A(n2158), .B(n2157), .Z(n7830) );
  NAND U7519 ( .A(n2160), .B(n2159), .Z(n2164) );
  NAND U7520 ( .A(n2162), .B(n2161), .Z(n2163) );
  NAND U7521 ( .A(n2164), .B(n2163), .Z(n7831) );
  XNOR U7522 ( .A(n7830), .B(n7831), .Z(n7833) );
  NANDN U7523 ( .A(n2166), .B(n2165), .Z(n2170) );
  NAND U7524 ( .A(n2168), .B(n2167), .Z(n2169) );
  AND U7525 ( .A(n2170), .B(n2169), .Z(n7832) );
  XOR U7526 ( .A(n7833), .B(n7832), .Z(n8122) );
  NANDN U7527 ( .A(n2172), .B(n2171), .Z(n2176) );
  NANDN U7528 ( .A(n2174), .B(n2173), .Z(n2175) );
  AND U7529 ( .A(n2176), .B(n2175), .Z(n8121) );
  XNOR U7530 ( .A(n8122), .B(n8121), .Z(n8123) );
  XOR U7531 ( .A(n8124), .B(n8123), .Z(n7773) );
  NANDN U7532 ( .A(n2178), .B(n2177), .Z(n2182) );
  NANDN U7533 ( .A(n2180), .B(n2179), .Z(n2181) );
  AND U7534 ( .A(n2182), .B(n2181), .Z(n6705) );
  NANDN U7535 ( .A(n2184), .B(n2183), .Z(n2188) );
  NAND U7536 ( .A(n2186), .B(n2185), .Z(n2187) );
  AND U7537 ( .A(n2188), .B(n2187), .Z(n7642) );
  NANDN U7538 ( .A(n2190), .B(n2189), .Z(n2194) );
  NAND U7539 ( .A(n2192), .B(n2191), .Z(n2193) );
  NAND U7540 ( .A(n2194), .B(n2193), .Z(n7643) );
  XNOR U7541 ( .A(n7642), .B(n7643), .Z(n7645) );
  NANDN U7542 ( .A(n2196), .B(n2195), .Z(n2200) );
  NAND U7543 ( .A(n2198), .B(n2197), .Z(n2199) );
  AND U7544 ( .A(n2200), .B(n2199), .Z(n7644) );
  XOR U7545 ( .A(n7645), .B(n7644), .Z(n6703) );
  NANDN U7546 ( .A(n2202), .B(n2201), .Z(n2206) );
  NANDN U7547 ( .A(n2204), .B(n2203), .Z(n2205) );
  AND U7548 ( .A(n2206), .B(n2205), .Z(n6702) );
  XNOR U7549 ( .A(n6703), .B(n6702), .Z(n6704) );
  XOR U7550 ( .A(n6705), .B(n6704), .Z(n7771) );
  NANDN U7551 ( .A(n2208), .B(n2207), .Z(n2212) );
  NANDN U7552 ( .A(n2210), .B(n2209), .Z(n2211) );
  AND U7553 ( .A(n2212), .B(n2211), .Z(n8358) );
  NANDN U7554 ( .A(n2214), .B(n2213), .Z(n2218) );
  NAND U7555 ( .A(n2216), .B(n2215), .Z(n2217) );
  AND U7556 ( .A(n2218), .B(n2217), .Z(n7654) );
  NANDN U7557 ( .A(n2220), .B(n2219), .Z(n2224) );
  NAND U7558 ( .A(n2222), .B(n2221), .Z(n2223) );
  NAND U7559 ( .A(n2224), .B(n2223), .Z(n7655) );
  XNOR U7560 ( .A(n7654), .B(n7655), .Z(n7657) );
  NAND U7561 ( .A(n2226), .B(n2225), .Z(n2230) );
  NAND U7562 ( .A(n2228), .B(n2227), .Z(n2229) );
  AND U7563 ( .A(n2230), .B(n2229), .Z(n7656) );
  XOR U7564 ( .A(n7657), .B(n7656), .Z(n8356) );
  NANDN U7565 ( .A(n2232), .B(n2231), .Z(n2236) );
  NANDN U7566 ( .A(n2234), .B(n2233), .Z(n2235) );
  AND U7567 ( .A(n2236), .B(n2235), .Z(n8355) );
  XNOR U7568 ( .A(n8356), .B(n8355), .Z(n8357) );
  XNOR U7569 ( .A(n8358), .B(n8357), .Z(n7770) );
  XNOR U7570 ( .A(n7771), .B(n7770), .Z(n7772) );
  XNOR U7571 ( .A(n7773), .B(n7772), .Z(n6188) );
  NANDN U7572 ( .A(n2238), .B(n2237), .Z(n2242) );
  NANDN U7573 ( .A(n2240), .B(n2239), .Z(n2241) );
  AND U7574 ( .A(n2242), .B(n2241), .Z(n8117) );
  NANDN U7575 ( .A(n2244), .B(n2243), .Z(n2248) );
  NAND U7576 ( .A(n2246), .B(n2245), .Z(n2247) );
  AND U7577 ( .A(n2248), .B(n2247), .Z(n8187) );
  NAND U7578 ( .A(n2250), .B(n2249), .Z(n2254) );
  NAND U7579 ( .A(n2252), .B(n2251), .Z(n2253) );
  NAND U7580 ( .A(n2254), .B(n2253), .Z(n8188) );
  XNOR U7581 ( .A(n8187), .B(n8188), .Z(n8190) );
  NAND U7582 ( .A(n2256), .B(n2255), .Z(n2260) );
  NAND U7583 ( .A(n2258), .B(n2257), .Z(n2259) );
  AND U7584 ( .A(n2260), .B(n2259), .Z(n8189) );
  XOR U7585 ( .A(n8190), .B(n8189), .Z(n8116) );
  NANDN U7586 ( .A(n2262), .B(n2261), .Z(n2266) );
  NANDN U7587 ( .A(n2264), .B(n2263), .Z(n2265) );
  AND U7588 ( .A(n2266), .B(n2265), .Z(n8115) );
  XOR U7589 ( .A(n8116), .B(n8115), .Z(n8118) );
  XNOR U7590 ( .A(n8117), .B(n8118), .Z(n8031) );
  NANDN U7591 ( .A(n2268), .B(n2267), .Z(n2272) );
  NAND U7592 ( .A(n2270), .B(n2269), .Z(n2271) );
  AND U7593 ( .A(n2272), .B(n2271), .Z(n8919) );
  NANDN U7594 ( .A(n2274), .B(n2273), .Z(n2278) );
  NAND U7595 ( .A(n2276), .B(n2275), .Z(n2277) );
  AND U7596 ( .A(n2278), .B(n2277), .Z(n8918) );
  XOR U7597 ( .A(n8919), .B(n8918), .Z(n8921) );
  NANDN U7598 ( .A(n2280), .B(n2279), .Z(n2284) );
  NAND U7599 ( .A(n2282), .B(n2281), .Z(n2283) );
  AND U7600 ( .A(n2284), .B(n2283), .Z(n8920) );
  XOR U7601 ( .A(n8921), .B(n8920), .Z(n6813) );
  NANDN U7602 ( .A(n2286), .B(n2285), .Z(n2290) );
  NAND U7603 ( .A(n2288), .B(n2287), .Z(n2289) );
  AND U7604 ( .A(n2290), .B(n2289), .Z(n8884) );
  NANDN U7605 ( .A(n2292), .B(n2291), .Z(n2296) );
  NAND U7606 ( .A(n2294), .B(n2293), .Z(n2295) );
  AND U7607 ( .A(n2296), .B(n2295), .Z(n8883) );
  XOR U7608 ( .A(n8884), .B(n8883), .Z(n8886) );
  NANDN U7609 ( .A(n2298), .B(n2297), .Z(n2302) );
  NAND U7610 ( .A(n2300), .B(n2299), .Z(n2301) );
  AND U7611 ( .A(n2302), .B(n2301), .Z(n8885) );
  XOR U7612 ( .A(n8886), .B(n8885), .Z(n6811) );
  NANDN U7613 ( .A(n2304), .B(n2303), .Z(n2308) );
  NAND U7614 ( .A(n2306), .B(n2305), .Z(n2307) );
  AND U7615 ( .A(n2308), .B(n2307), .Z(n7612) );
  NANDN U7616 ( .A(n2310), .B(n2309), .Z(n2314) );
  NAND U7617 ( .A(n2312), .B(n2311), .Z(n2313) );
  NAND U7618 ( .A(n2314), .B(n2313), .Z(n7613) );
  XNOR U7619 ( .A(n7612), .B(n7613), .Z(n7615) );
  NANDN U7620 ( .A(n2316), .B(n2315), .Z(n2320) );
  NAND U7621 ( .A(n2318), .B(n2317), .Z(n2319) );
  AND U7622 ( .A(n2320), .B(n2319), .Z(n7614) );
  XNOR U7623 ( .A(n7615), .B(n7614), .Z(n6810) );
  XNOR U7624 ( .A(n6811), .B(n6810), .Z(n6812) );
  XOR U7625 ( .A(n6813), .B(n6812), .Z(n8032) );
  XNOR U7626 ( .A(n8031), .B(n8032), .Z(n8034) );
  NANDN U7627 ( .A(n2322), .B(n2321), .Z(n2326) );
  NAND U7628 ( .A(n2324), .B(n2323), .Z(n2325) );
  AND U7629 ( .A(n2326), .B(n2325), .Z(n6696) );
  NANDN U7630 ( .A(n2328), .B(n2327), .Z(n2332) );
  NAND U7631 ( .A(n2330), .B(n2329), .Z(n2331) );
  NAND U7632 ( .A(n2332), .B(n2331), .Z(n6697) );
  XNOR U7633 ( .A(n6696), .B(n6697), .Z(n6699) );
  NANDN U7634 ( .A(n2334), .B(n2333), .Z(n2338) );
  NAND U7635 ( .A(n2336), .B(n2335), .Z(n2337) );
  AND U7636 ( .A(n2338), .B(n2337), .Z(n6698) );
  XOR U7637 ( .A(n6699), .B(n6698), .Z(n8208) );
  NANDN U7638 ( .A(n2340), .B(n2339), .Z(n2344) );
  NAND U7639 ( .A(n2342), .B(n2341), .Z(n2343) );
  AND U7640 ( .A(n2344), .B(n2343), .Z(n6402) );
  NAND U7641 ( .A(n2346), .B(n2345), .Z(n2350) );
  NAND U7642 ( .A(n2348), .B(n2347), .Z(n2349) );
  NAND U7643 ( .A(n2350), .B(n2349), .Z(n6403) );
  XNOR U7644 ( .A(n6402), .B(n6403), .Z(n6405) );
  NAND U7645 ( .A(n2352), .B(n2351), .Z(n2356) );
  NAND U7646 ( .A(n2354), .B(n2353), .Z(n2355) );
  AND U7647 ( .A(n2356), .B(n2355), .Z(n6404) );
  XOR U7648 ( .A(n6405), .B(n6404), .Z(n8206) );
  NANDN U7649 ( .A(n2358), .B(n2357), .Z(n2362) );
  NAND U7650 ( .A(n2360), .B(n2359), .Z(n2361) );
  AND U7651 ( .A(n2362), .B(n2361), .Z(n7794) );
  NANDN U7652 ( .A(n2364), .B(n2363), .Z(n2368) );
  NAND U7653 ( .A(n2366), .B(n2365), .Z(n2367) );
  NAND U7654 ( .A(n2368), .B(n2367), .Z(n7795) );
  XNOR U7655 ( .A(n7794), .B(n7795), .Z(n7797) );
  NANDN U7656 ( .A(n2370), .B(n2369), .Z(n2374) );
  NAND U7657 ( .A(n2372), .B(n2371), .Z(n2373) );
  AND U7658 ( .A(n2374), .B(n2373), .Z(n7796) );
  XNOR U7659 ( .A(n7797), .B(n7796), .Z(n8205) );
  XNOR U7660 ( .A(n8206), .B(n8205), .Z(n8207) );
  XNOR U7661 ( .A(n8208), .B(n8207), .Z(n8033) );
  XOR U7662 ( .A(n8034), .B(n8033), .Z(n6187) );
  NANDN U7663 ( .A(n2376), .B(n2375), .Z(n2380) );
  NANDN U7664 ( .A(n2378), .B(n2377), .Z(n2379) );
  AND U7665 ( .A(n2380), .B(n2379), .Z(n8568) );
  NANDN U7666 ( .A(n2382), .B(n2381), .Z(n2386) );
  NAND U7667 ( .A(n2384), .B(n2383), .Z(n2385) );
  AND U7668 ( .A(n2386), .B(n2385), .Z(n7807) );
  NANDN U7669 ( .A(n2388), .B(n2387), .Z(n2392) );
  NAND U7670 ( .A(n2390), .B(n2389), .Z(n2391) );
  AND U7671 ( .A(n2392), .B(n2391), .Z(n7806) );
  XOR U7672 ( .A(n7807), .B(n7806), .Z(n7809) );
  NANDN U7673 ( .A(n2394), .B(n2393), .Z(n2398) );
  NAND U7674 ( .A(n2396), .B(n2395), .Z(n2397) );
  AND U7675 ( .A(n2398), .B(n2397), .Z(n7808) );
  XOR U7676 ( .A(n7809), .B(n7808), .Z(n8566) );
  NANDN U7677 ( .A(n2400), .B(n2399), .Z(n2404) );
  NANDN U7678 ( .A(n2402), .B(n2401), .Z(n2403) );
  AND U7679 ( .A(n2404), .B(n2403), .Z(n8565) );
  XNOR U7680 ( .A(n8566), .B(n8565), .Z(n8567) );
  XOR U7681 ( .A(n8568), .B(n8567), .Z(n7980) );
  NANDN U7682 ( .A(n2406), .B(n2405), .Z(n2410) );
  NANDN U7683 ( .A(n2408), .B(n2407), .Z(n2409) );
  AND U7684 ( .A(n2410), .B(n2409), .Z(n8562) );
  NANDN U7685 ( .A(n2412), .B(n2411), .Z(n2416) );
  NAND U7686 ( .A(n2414), .B(n2413), .Z(n2415) );
  AND U7687 ( .A(n2416), .B(n2415), .Z(n7861) );
  NANDN U7688 ( .A(n2418), .B(n2417), .Z(n2422) );
  NAND U7689 ( .A(n2420), .B(n2419), .Z(n2421) );
  AND U7690 ( .A(n2422), .B(n2421), .Z(n7860) );
  XOR U7691 ( .A(n7861), .B(n7860), .Z(n7863) );
  NANDN U7692 ( .A(n2424), .B(n2423), .Z(n2428) );
  NAND U7693 ( .A(n2426), .B(n2425), .Z(n2427) );
  AND U7694 ( .A(n2428), .B(n2427), .Z(n7862) );
  XOR U7695 ( .A(n7863), .B(n7862), .Z(n8560) );
  NANDN U7696 ( .A(n2430), .B(n2429), .Z(n2434) );
  NANDN U7697 ( .A(n2432), .B(n2431), .Z(n2433) );
  AND U7698 ( .A(n2434), .B(n2433), .Z(n8559) );
  XNOR U7699 ( .A(n8560), .B(n8559), .Z(n8561) );
  XOR U7700 ( .A(n8562), .B(n8561), .Z(n7978) );
  NANDN U7701 ( .A(n2436), .B(n2435), .Z(n2440) );
  NANDN U7702 ( .A(n2438), .B(n2437), .Z(n2439) );
  AND U7703 ( .A(n2440), .B(n2439), .Z(n8520) );
  NANDN U7704 ( .A(n2442), .B(n2441), .Z(n2446) );
  NAND U7705 ( .A(n2444), .B(n2443), .Z(n2445) );
  AND U7706 ( .A(n2446), .B(n2445), .Z(n7576) );
  NANDN U7707 ( .A(n2448), .B(n2447), .Z(n2452) );
  NAND U7708 ( .A(n2450), .B(n2449), .Z(n2451) );
  NAND U7709 ( .A(n2452), .B(n2451), .Z(n7577) );
  XNOR U7710 ( .A(n7576), .B(n7577), .Z(n7579) );
  NANDN U7711 ( .A(n2454), .B(n2453), .Z(n2458) );
  NAND U7712 ( .A(n2456), .B(n2455), .Z(n2457) );
  AND U7713 ( .A(n2458), .B(n2457), .Z(n7578) );
  XOR U7714 ( .A(n7579), .B(n7578), .Z(n8518) );
  NANDN U7715 ( .A(n2460), .B(n2459), .Z(n2464) );
  NANDN U7716 ( .A(n2462), .B(n2461), .Z(n2463) );
  AND U7717 ( .A(n2464), .B(n2463), .Z(n8517) );
  XNOR U7718 ( .A(n8518), .B(n8517), .Z(n8519) );
  XNOR U7719 ( .A(n8520), .B(n8519), .Z(n7977) );
  XNOR U7720 ( .A(n7978), .B(n7977), .Z(n7979) );
  XNOR U7721 ( .A(n7980), .B(n7979), .Z(n6186) );
  XOR U7722 ( .A(n6187), .B(n6186), .Z(n6189) );
  XNOR U7723 ( .A(n6188), .B(n6189), .Z(n8644) );
  XOR U7724 ( .A(n8643), .B(n8644), .Z(n8646) );
  NANDN U7725 ( .A(n2466), .B(n2465), .Z(n2470) );
  NAND U7726 ( .A(n2468), .B(n2467), .Z(n2469) );
  AND U7727 ( .A(n2470), .B(n2469), .Z(n7528) );
  NANDN U7728 ( .A(n2472), .B(n2471), .Z(n2476) );
  NAND U7729 ( .A(n2474), .B(n2473), .Z(n2475) );
  NAND U7730 ( .A(n2476), .B(n2475), .Z(n7529) );
  XNOR U7731 ( .A(n7528), .B(n7529), .Z(n7531) );
  NANDN U7732 ( .A(n2478), .B(n2477), .Z(n2482) );
  NAND U7733 ( .A(n2480), .B(n2479), .Z(n2481) );
  AND U7734 ( .A(n2482), .B(n2481), .Z(n7530) );
  XOR U7735 ( .A(n7531), .B(n7530), .Z(n8363) );
  NANDN U7736 ( .A(n2484), .B(n2483), .Z(n2488) );
  NANDN U7737 ( .A(n2486), .B(n2485), .Z(n2487) );
  AND U7738 ( .A(n2488), .B(n2487), .Z(n6612) );
  NANDN U7739 ( .A(n2490), .B(n2489), .Z(n2494) );
  NAND U7740 ( .A(n2492), .B(n2491), .Z(n2493) );
  NAND U7741 ( .A(n2494), .B(n2493), .Z(n6613) );
  XNOR U7742 ( .A(n6612), .B(n6613), .Z(n6615) );
  NANDN U7743 ( .A(n2496), .B(n2495), .Z(n2500) );
  NAND U7744 ( .A(n2498), .B(n2497), .Z(n2499) );
  AND U7745 ( .A(n2500), .B(n2499), .Z(n6614) );
  XOR U7746 ( .A(n6615), .B(n6614), .Z(n8362) );
  NANDN U7747 ( .A(n2502), .B(n2501), .Z(n2506) );
  NANDN U7748 ( .A(n2504), .B(n2503), .Z(n2505) );
  AND U7749 ( .A(n2506), .B(n2505), .Z(n8361) );
  XOR U7750 ( .A(n8362), .B(n8361), .Z(n8364) );
  XOR U7751 ( .A(n8363), .B(n8364), .Z(n8028) );
  NANDN U7752 ( .A(n2508), .B(n2507), .Z(n2512) );
  NANDN U7753 ( .A(n2510), .B(n2509), .Z(n2511) );
  AND U7754 ( .A(n2512), .B(n2511), .Z(n6774) );
  NANDN U7755 ( .A(n2514), .B(n2513), .Z(n2518) );
  NAND U7756 ( .A(n2516), .B(n2515), .Z(n2517) );
  NAND U7757 ( .A(n2518), .B(n2517), .Z(n6775) );
  XNOR U7758 ( .A(n6774), .B(n6775), .Z(n6777) );
  NANDN U7759 ( .A(n2520), .B(n2519), .Z(n2524) );
  NAND U7760 ( .A(n2522), .B(n2521), .Z(n2523) );
  AND U7761 ( .A(n2524), .B(n2523), .Z(n6776) );
  XOR U7762 ( .A(n6777), .B(n6776), .Z(n8813) );
  NANDN U7763 ( .A(n2526), .B(n2525), .Z(n2530) );
  NAND U7764 ( .A(n2528), .B(n2527), .Z(n2529) );
  AND U7765 ( .A(n2530), .B(n2529), .Z(n6444) );
  NANDN U7766 ( .A(n2532), .B(n2531), .Z(n2536) );
  NAND U7767 ( .A(n2534), .B(n2533), .Z(n2535) );
  NAND U7768 ( .A(n2536), .B(n2535), .Z(n6445) );
  XNOR U7769 ( .A(n6444), .B(n6445), .Z(n6447) );
  NANDN U7770 ( .A(n2538), .B(n2537), .Z(n2542) );
  NAND U7771 ( .A(n2540), .B(n2539), .Z(n2541) );
  AND U7772 ( .A(n2542), .B(n2541), .Z(n6446) );
  XOR U7773 ( .A(n6447), .B(n6446), .Z(n8812) );
  NANDN U7774 ( .A(n2544), .B(n2543), .Z(n2548) );
  NAND U7775 ( .A(n2546), .B(n2545), .Z(n2547) );
  AND U7776 ( .A(n2548), .B(n2547), .Z(n7582) );
  NANDN U7777 ( .A(n2550), .B(n2549), .Z(n2554) );
  NAND U7778 ( .A(n2552), .B(n2551), .Z(n2553) );
  NAND U7779 ( .A(n2554), .B(n2553), .Z(n7583) );
  XNOR U7780 ( .A(n7582), .B(n7583), .Z(n7585) );
  NANDN U7781 ( .A(n2556), .B(n2555), .Z(n2560) );
  NAND U7782 ( .A(n2558), .B(n2557), .Z(n2559) );
  AND U7783 ( .A(n2560), .B(n2559), .Z(n7584) );
  XNOR U7784 ( .A(n7585), .B(n7584), .Z(n8811) );
  XOR U7785 ( .A(n8812), .B(n8811), .Z(n8814) );
  XOR U7786 ( .A(n8813), .B(n8814), .Z(n8026) );
  NAND U7787 ( .A(n2562), .B(n2561), .Z(n2566) );
  NAND U7788 ( .A(n2564), .B(n2563), .Z(n2565) );
  AND U7789 ( .A(n2566), .B(n2565), .Z(n7462) );
  NANDN U7790 ( .A(n2568), .B(n2567), .Z(n2572) );
  NAND U7791 ( .A(n2570), .B(n2569), .Z(n2571) );
  NAND U7792 ( .A(n2572), .B(n2571), .Z(n7463) );
  XNOR U7793 ( .A(n7462), .B(n7463), .Z(n7465) );
  NANDN U7794 ( .A(n2574), .B(n2573), .Z(n2578) );
  NAND U7795 ( .A(n2576), .B(n2575), .Z(n2577) );
  AND U7796 ( .A(n2578), .B(n2577), .Z(n7464) );
  XOR U7797 ( .A(n7465), .B(n7464), .Z(n8663) );
  NANDN U7798 ( .A(n2580), .B(n2579), .Z(n2584) );
  NAND U7799 ( .A(n2582), .B(n2581), .Z(n2583) );
  AND U7800 ( .A(n2584), .B(n2583), .Z(n8823) );
  NANDN U7801 ( .A(n2586), .B(n2585), .Z(n2590) );
  NAND U7802 ( .A(n2588), .B(n2587), .Z(n2589) );
  NAND U7803 ( .A(n2590), .B(n2589), .Z(n8824) );
  XNOR U7804 ( .A(n8823), .B(n8824), .Z(n8826) );
  NANDN U7805 ( .A(n2592), .B(n2591), .Z(n2596) );
  NAND U7806 ( .A(n2594), .B(n2593), .Z(n2595) );
  AND U7807 ( .A(n2596), .B(n2595), .Z(n8825) );
  XOR U7808 ( .A(n8826), .B(n8825), .Z(n8662) );
  NANDN U7809 ( .A(n2598), .B(n2597), .Z(n2602) );
  NANDN U7810 ( .A(n2600), .B(n2599), .Z(n2601) );
  AND U7811 ( .A(n2602), .B(n2601), .Z(n8661) );
  XOR U7812 ( .A(n8662), .B(n8661), .Z(n8664) );
  XNOR U7813 ( .A(n8663), .B(n8664), .Z(n8025) );
  XNOR U7814 ( .A(n8026), .B(n8025), .Z(n8027) );
  XNOR U7815 ( .A(n8028), .B(n8027), .Z(n6212) );
  NANDN U7816 ( .A(n2604), .B(n2603), .Z(n2608) );
  NAND U7817 ( .A(n2606), .B(n2605), .Z(n2607) );
  AND U7818 ( .A(n2608), .B(n2607), .Z(n8943) );
  NANDN U7819 ( .A(n2610), .B(n2609), .Z(n2614) );
  NAND U7820 ( .A(n2612), .B(n2611), .Z(n2613) );
  AND U7821 ( .A(n2614), .B(n2613), .Z(n8942) );
  XOR U7822 ( .A(n8943), .B(n8942), .Z(n8945) );
  NANDN U7823 ( .A(n2616), .B(n2615), .Z(n2620) );
  NAND U7824 ( .A(n2618), .B(n2617), .Z(n2619) );
  AND U7825 ( .A(n2620), .B(n2619), .Z(n8944) );
  XOR U7826 ( .A(n8945), .B(n8944), .Z(n9029) );
  NANDN U7827 ( .A(n2622), .B(n2621), .Z(n2626) );
  NAND U7828 ( .A(n2624), .B(n2623), .Z(n2625) );
  AND U7829 ( .A(n2626), .B(n2625), .Z(n6505) );
  NAND U7830 ( .A(n2628), .B(n2627), .Z(n2632) );
  NAND U7831 ( .A(n2630), .B(n2629), .Z(n2631) );
  AND U7832 ( .A(n2632), .B(n2631), .Z(n6504) );
  XOR U7833 ( .A(n6505), .B(n6504), .Z(n6507) );
  NANDN U7834 ( .A(n2634), .B(n2633), .Z(n2638) );
  NAND U7835 ( .A(n2636), .B(n2635), .Z(n2637) );
  AND U7836 ( .A(n2638), .B(n2637), .Z(n6506) );
  XOR U7837 ( .A(n6507), .B(n6506), .Z(n9028) );
  NANDN U7838 ( .A(n2640), .B(n2639), .Z(n2644) );
  NANDN U7839 ( .A(n2642), .B(n2641), .Z(n2643) );
  AND U7840 ( .A(n2644), .B(n2643), .Z(n9027) );
  XOR U7841 ( .A(n9028), .B(n9027), .Z(n9030) );
  XOR U7842 ( .A(n9029), .B(n9030), .Z(n7938) );
  NANDN U7843 ( .A(n2646), .B(n2645), .Z(n2650) );
  NAND U7844 ( .A(n2648), .B(n2647), .Z(n2649) );
  AND U7845 ( .A(n2650), .B(n2649), .Z(n7540) );
  NANDN U7846 ( .A(n2652), .B(n2651), .Z(n2656) );
  NAND U7847 ( .A(n2654), .B(n2653), .Z(n2655) );
  NAND U7848 ( .A(n2656), .B(n2655), .Z(n7541) );
  XNOR U7849 ( .A(n7540), .B(n7541), .Z(n7543) );
  NANDN U7850 ( .A(n2658), .B(n2657), .Z(n2662) );
  NAND U7851 ( .A(n2660), .B(n2659), .Z(n2661) );
  AND U7852 ( .A(n2662), .B(n2661), .Z(n7542) );
  XOR U7853 ( .A(n7543), .B(n7542), .Z(n7296) );
  NANDN U7854 ( .A(n2664), .B(n2663), .Z(n2668) );
  NANDN U7855 ( .A(n2666), .B(n2665), .Z(n2667) );
  AND U7856 ( .A(n2668), .B(n2667), .Z(n7546) );
  NANDN U7857 ( .A(n2670), .B(n2669), .Z(n2674) );
  NAND U7858 ( .A(n2672), .B(n2671), .Z(n2673) );
  NAND U7859 ( .A(n2674), .B(n2673), .Z(n7547) );
  XNOR U7860 ( .A(n7546), .B(n7547), .Z(n7549) );
  NANDN U7861 ( .A(n2676), .B(n2675), .Z(n2680) );
  NAND U7862 ( .A(n2678), .B(n2677), .Z(n2679) );
  AND U7863 ( .A(n2680), .B(n2679), .Z(n7548) );
  XOR U7864 ( .A(n7549), .B(n7548), .Z(n7295) );
  NANDN U7865 ( .A(n2682), .B(n2681), .Z(n2686) );
  NANDN U7866 ( .A(n2684), .B(n2683), .Z(n2685) );
  AND U7867 ( .A(n2686), .B(n2685), .Z(n7294) );
  XOR U7868 ( .A(n7295), .B(n7294), .Z(n7297) );
  XOR U7869 ( .A(n7296), .B(n7297), .Z(n7936) );
  NAND U7870 ( .A(n2688), .B(n2687), .Z(n2692) );
  NAND U7871 ( .A(n2690), .B(n2689), .Z(n2691) );
  AND U7872 ( .A(n2692), .B(n2691), .Z(n7486) );
  NANDN U7873 ( .A(n2694), .B(n2693), .Z(n2698) );
  NAND U7874 ( .A(n2696), .B(n2695), .Z(n2697) );
  NAND U7875 ( .A(n2698), .B(n2697), .Z(n7487) );
  XNOR U7876 ( .A(n7486), .B(n7487), .Z(n7489) );
  NANDN U7877 ( .A(n2700), .B(n2699), .Z(n2704) );
  NAND U7878 ( .A(n2702), .B(n2701), .Z(n2703) );
  AND U7879 ( .A(n2704), .B(n2703), .Z(n7488) );
  XOR U7880 ( .A(n7489), .B(n7488), .Z(n8999) );
  NANDN U7881 ( .A(n2706), .B(n2705), .Z(n2710) );
  NAND U7882 ( .A(n2708), .B(n2707), .Z(n2709) );
  AND U7883 ( .A(n2710), .B(n2709), .Z(n6726) );
  NANDN U7884 ( .A(n2712), .B(n2711), .Z(n2716) );
  NAND U7885 ( .A(n2714), .B(n2713), .Z(n2715) );
  NAND U7886 ( .A(n2716), .B(n2715), .Z(n6727) );
  XNOR U7887 ( .A(n6726), .B(n6727), .Z(n6729) );
  NANDN U7888 ( .A(n2718), .B(n2717), .Z(n2722) );
  NAND U7889 ( .A(n2720), .B(n2719), .Z(n2721) );
  AND U7890 ( .A(n2722), .B(n2721), .Z(n6728) );
  XOR U7891 ( .A(n6729), .B(n6728), .Z(n8998) );
  NANDN U7892 ( .A(n2724), .B(n2723), .Z(n2728) );
  NANDN U7893 ( .A(n2726), .B(n2725), .Z(n2727) );
  AND U7894 ( .A(n2728), .B(n2727), .Z(n8997) );
  XOR U7895 ( .A(n8998), .B(n8997), .Z(n9000) );
  XNOR U7896 ( .A(n8999), .B(n9000), .Z(n7935) );
  XNOR U7897 ( .A(n7936), .B(n7935), .Z(n7937) );
  XNOR U7898 ( .A(n7938), .B(n7937), .Z(n6210) );
  NANDN U7899 ( .A(n2730), .B(n2729), .Z(n2734) );
  NAND U7900 ( .A(n2732), .B(n2731), .Z(n2733) );
  AND U7901 ( .A(n2734), .B(n2733), .Z(n6516) );
  NAND U7902 ( .A(n2736), .B(n2735), .Z(n2740) );
  NAND U7903 ( .A(n2738), .B(n2737), .Z(n2739) );
  NAND U7904 ( .A(n2740), .B(n2739), .Z(n6517) );
  XNOR U7905 ( .A(n6516), .B(n6517), .Z(n6519) );
  NANDN U7906 ( .A(n2742), .B(n2741), .Z(n2746) );
  NAND U7907 ( .A(n2744), .B(n2743), .Z(n2745) );
  AND U7908 ( .A(n2746), .B(n2745), .Z(n6518) );
  XOR U7909 ( .A(n6519), .B(n6518), .Z(n8213) );
  NANDN U7910 ( .A(n2748), .B(n2747), .Z(n2752) );
  NAND U7911 ( .A(n2750), .B(n2749), .Z(n2751) );
  AND U7912 ( .A(n2752), .B(n2751), .Z(n8979) );
  NANDN U7913 ( .A(n2754), .B(n2753), .Z(n2758) );
  NAND U7914 ( .A(n2756), .B(n2755), .Z(n2757) );
  NAND U7915 ( .A(n2758), .B(n2757), .Z(n8980) );
  XNOR U7916 ( .A(n8979), .B(n8980), .Z(n8982) );
  NANDN U7917 ( .A(n2760), .B(n2759), .Z(n2764) );
  NAND U7918 ( .A(n2762), .B(n2761), .Z(n2763) );
  AND U7919 ( .A(n2764), .B(n2763), .Z(n8981) );
  XOR U7920 ( .A(n8982), .B(n8981), .Z(n8212) );
  NANDN U7921 ( .A(n2766), .B(n2765), .Z(n2770) );
  NAND U7922 ( .A(n2768), .B(n2767), .Z(n2769) );
  AND U7923 ( .A(n2770), .B(n2769), .Z(n7444) );
  NANDN U7924 ( .A(n2772), .B(n2771), .Z(n2776) );
  NANDN U7925 ( .A(n2774), .B(n2773), .Z(n2775) );
  NAND U7926 ( .A(n2776), .B(n2775), .Z(n7445) );
  XNOR U7927 ( .A(n7444), .B(n7445), .Z(n7447) );
  NANDN U7928 ( .A(n2778), .B(n2777), .Z(n2782) );
  NAND U7929 ( .A(n2780), .B(n2779), .Z(n2781) );
  AND U7930 ( .A(n2782), .B(n2781), .Z(n7446) );
  XNOR U7931 ( .A(n7447), .B(n7446), .Z(n8211) );
  XOR U7932 ( .A(n8212), .B(n8211), .Z(n8214) );
  XOR U7933 ( .A(n8213), .B(n8214), .Z(n6979) );
  NANDN U7934 ( .A(n2784), .B(n2783), .Z(n2788) );
  NANDN U7935 ( .A(n2786), .B(n2785), .Z(n2787) );
  AND U7936 ( .A(n2788), .B(n2787), .Z(n7291) );
  NANDN U7937 ( .A(n2790), .B(n2789), .Z(n2794) );
  NANDN U7938 ( .A(n2792), .B(n2791), .Z(n2793) );
  AND U7939 ( .A(n2794), .B(n2793), .Z(n7288) );
  NANDN U7940 ( .A(n2796), .B(n2795), .Z(n2800) );
  NANDN U7941 ( .A(n2798), .B(n2797), .Z(n2799) );
  NAND U7942 ( .A(n2800), .B(n2799), .Z(n7289) );
  XNOR U7943 ( .A(n7288), .B(n7289), .Z(n7290) );
  XOR U7944 ( .A(n7291), .B(n7290), .Z(n6977) );
  NANDN U7945 ( .A(n2802), .B(n2801), .Z(n2806) );
  NAND U7946 ( .A(n2804), .B(n2803), .Z(n2805) );
  AND U7947 ( .A(n2806), .B(n2805), .Z(n7722) );
  NANDN U7948 ( .A(n2808), .B(n2807), .Z(n2812) );
  NAND U7949 ( .A(n2810), .B(n2809), .Z(n2811) );
  NAND U7950 ( .A(n2812), .B(n2811), .Z(n7723) );
  XNOR U7951 ( .A(n7722), .B(n7723), .Z(n7725) );
  NANDN U7952 ( .A(n2814), .B(n2813), .Z(n2818) );
  NAND U7953 ( .A(n2816), .B(n2815), .Z(n2817) );
  AND U7954 ( .A(n2818), .B(n2817), .Z(n7724) );
  XOR U7955 ( .A(n7725), .B(n7724), .Z(n9005) );
  NANDN U7956 ( .A(n2820), .B(n2819), .Z(n2824) );
  NAND U7957 ( .A(n2822), .B(n2821), .Z(n2823) );
  AND U7958 ( .A(n2824), .B(n2823), .Z(n6468) );
  NANDN U7959 ( .A(n2826), .B(n2825), .Z(n2830) );
  NAND U7960 ( .A(n2828), .B(n2827), .Z(n2829) );
  NAND U7961 ( .A(n2830), .B(n2829), .Z(n6469) );
  XNOR U7962 ( .A(n6468), .B(n6469), .Z(n6471) );
  NANDN U7963 ( .A(n2832), .B(n2831), .Z(n2836) );
  NAND U7964 ( .A(n2834), .B(n2833), .Z(n2835) );
  AND U7965 ( .A(n2836), .B(n2835), .Z(n6470) );
  XOR U7966 ( .A(n6471), .B(n6470), .Z(n9004) );
  NANDN U7967 ( .A(n2838), .B(n2837), .Z(n2842) );
  NANDN U7968 ( .A(n2840), .B(n2839), .Z(n2841) );
  AND U7969 ( .A(n2842), .B(n2841), .Z(n9003) );
  XOR U7970 ( .A(n9004), .B(n9003), .Z(n9006) );
  XNOR U7971 ( .A(n9005), .B(n9006), .Z(n6976) );
  XNOR U7972 ( .A(n6977), .B(n6976), .Z(n6978) );
  XOR U7973 ( .A(n6979), .B(n6978), .Z(n6211) );
  XOR U7974 ( .A(n6210), .B(n6211), .Z(n6213) );
  XNOR U7975 ( .A(n6212), .B(n6213), .Z(n8645) );
  XNOR U7976 ( .A(n8646), .B(n8645), .Z(n7049) );
  NANDN U7977 ( .A(n2844), .B(n2843), .Z(n2848) );
  NANDN U7978 ( .A(n2846), .B(n2845), .Z(n2847) );
  AND U7979 ( .A(n2848), .B(n2847), .Z(n7368) );
  NANDN U7980 ( .A(n2850), .B(n2849), .Z(n2854) );
  NAND U7981 ( .A(n2852), .B(n2851), .Z(n2853) );
  AND U7982 ( .A(n2854), .B(n2853), .Z(n8763) );
  NANDN U7983 ( .A(n2856), .B(n2855), .Z(n2860) );
  NAND U7984 ( .A(n2858), .B(n2857), .Z(n2859) );
  NAND U7985 ( .A(n2860), .B(n2859), .Z(n8764) );
  XNOR U7986 ( .A(n8763), .B(n8764), .Z(n8766) );
  NANDN U7987 ( .A(n2862), .B(n2861), .Z(n2866) );
  NAND U7988 ( .A(n2864), .B(n2863), .Z(n2865) );
  AND U7989 ( .A(n2866), .B(n2865), .Z(n8765) );
  XOR U7990 ( .A(n8766), .B(n8765), .Z(n7367) );
  NANDN U7991 ( .A(n2868), .B(n2867), .Z(n2872) );
  NANDN U7992 ( .A(n2870), .B(n2869), .Z(n2871) );
  AND U7993 ( .A(n2872), .B(n2871), .Z(n7366) );
  XOR U7994 ( .A(n7367), .B(n7366), .Z(n7369) );
  XNOR U7995 ( .A(n7368), .B(n7369), .Z(n6288) );
  NANDN U7996 ( .A(n2874), .B(n2873), .Z(n2878) );
  NANDN U7997 ( .A(n2876), .B(n2875), .Z(n2877) );
  AND U7998 ( .A(n2878), .B(n2877), .Z(n7345) );
  NANDN U7999 ( .A(n2880), .B(n2879), .Z(n2884) );
  NAND U8000 ( .A(n2882), .B(n2881), .Z(n2883) );
  AND U8001 ( .A(n2884), .B(n2883), .Z(n7688) );
  NANDN U8002 ( .A(n2886), .B(n2885), .Z(n2890) );
  NAND U8003 ( .A(n2888), .B(n2887), .Z(n2889) );
  NAND U8004 ( .A(n2890), .B(n2889), .Z(n7689) );
  XNOR U8005 ( .A(n7688), .B(n7689), .Z(n7691) );
  NANDN U8006 ( .A(n2892), .B(n2891), .Z(n2896) );
  NAND U8007 ( .A(n2894), .B(n2893), .Z(n2895) );
  AND U8008 ( .A(n2896), .B(n2895), .Z(n7690) );
  XOR U8009 ( .A(n7691), .B(n7690), .Z(n7343) );
  NANDN U8010 ( .A(n2898), .B(n2897), .Z(n2902) );
  NANDN U8011 ( .A(n2900), .B(n2899), .Z(n2901) );
  AND U8012 ( .A(n2902), .B(n2901), .Z(n7342) );
  XNOR U8013 ( .A(n7343), .B(n7342), .Z(n7344) );
  XOR U8014 ( .A(n7345), .B(n7344), .Z(n6289) );
  XNOR U8015 ( .A(n6288), .B(n6289), .Z(n6291) );
  NANDN U8016 ( .A(n2904), .B(n2903), .Z(n2908) );
  NANDN U8017 ( .A(n2906), .B(n2905), .Z(n2907) );
  AND U8018 ( .A(n2908), .B(n2907), .Z(n7320) );
  NANDN U8019 ( .A(n2910), .B(n2909), .Z(n2914) );
  NAND U8020 ( .A(n2912), .B(n2911), .Z(n2913) );
  AND U8021 ( .A(n2914), .B(n2913), .Z(n6366) );
  NAND U8022 ( .A(n2916), .B(n2915), .Z(n2920) );
  NAND U8023 ( .A(n2918), .B(n2917), .Z(n2919) );
  NAND U8024 ( .A(n2920), .B(n2919), .Z(n6367) );
  XNOR U8025 ( .A(n6366), .B(n6367), .Z(n6369) );
  NAND U8026 ( .A(n2922), .B(n2921), .Z(n2926) );
  NAND U8027 ( .A(n2924), .B(n2923), .Z(n2925) );
  AND U8028 ( .A(n2926), .B(n2925), .Z(n6368) );
  XOR U8029 ( .A(n6369), .B(n6368), .Z(n7319) );
  NANDN U8030 ( .A(n2928), .B(n2927), .Z(n2932) );
  NANDN U8031 ( .A(n2930), .B(n2929), .Z(n2931) );
  AND U8032 ( .A(n2932), .B(n2931), .Z(n7318) );
  XOR U8033 ( .A(n7319), .B(n7318), .Z(n7321) );
  XNOR U8034 ( .A(n7320), .B(n7321), .Z(n6290) );
  XOR U8035 ( .A(n6291), .B(n6290), .Z(n7110) );
  NANDN U8036 ( .A(n2934), .B(n2933), .Z(n2938) );
  NANDN U8037 ( .A(n2936), .B(n2935), .Z(n2937) );
  AND U8038 ( .A(n2938), .B(n2937), .Z(n7350) );
  NANDN U8039 ( .A(n2940), .B(n2939), .Z(n2944) );
  NAND U8040 ( .A(n2942), .B(n2941), .Z(n2943) );
  AND U8041 ( .A(n2944), .B(n2943), .Z(n7534) );
  NANDN U8042 ( .A(n2946), .B(n2945), .Z(n2950) );
  NAND U8043 ( .A(n2948), .B(n2947), .Z(n2949) );
  NAND U8044 ( .A(n2950), .B(n2949), .Z(n7535) );
  XNOR U8045 ( .A(n7534), .B(n7535), .Z(n7537) );
  NANDN U8046 ( .A(n2952), .B(n2951), .Z(n2956) );
  NAND U8047 ( .A(n2954), .B(n2953), .Z(n2955) );
  AND U8048 ( .A(n2956), .B(n2955), .Z(n7536) );
  XOR U8049 ( .A(n7537), .B(n7536), .Z(n7349) );
  NANDN U8050 ( .A(n2958), .B(n2957), .Z(n2962) );
  NANDN U8051 ( .A(n2960), .B(n2959), .Z(n2961) );
  AND U8052 ( .A(n2962), .B(n2961), .Z(n7348) );
  XOR U8053 ( .A(n7349), .B(n7348), .Z(n7351) );
  XNOR U8054 ( .A(n7350), .B(n7351), .Z(n7498) );
  NANDN U8055 ( .A(n2964), .B(n2963), .Z(n2968) );
  NANDN U8056 ( .A(n2966), .B(n2965), .Z(n2967) );
  AND U8057 ( .A(n2968), .B(n2967), .Z(n7146) );
  NANDN U8058 ( .A(n2970), .B(n2969), .Z(n2974) );
  NAND U8059 ( .A(n2972), .B(n2971), .Z(n2973) );
  AND U8060 ( .A(n2974), .B(n2973), .Z(n8889) );
  NANDN U8061 ( .A(n2976), .B(n2975), .Z(n2980) );
  NANDN U8062 ( .A(n2978), .B(n2977), .Z(n2979) );
  NAND U8063 ( .A(n2980), .B(n2979), .Z(n8890) );
  XNOR U8064 ( .A(n8889), .B(n8890), .Z(n8892) );
  NANDN U8065 ( .A(n2982), .B(n2981), .Z(n2986) );
  NANDN U8066 ( .A(n2984), .B(n2983), .Z(n2985) );
  AND U8067 ( .A(n2986), .B(n2985), .Z(n8891) );
  XOR U8068 ( .A(n8892), .B(n8891), .Z(n7145) );
  NANDN U8069 ( .A(n2988), .B(n2987), .Z(n2992) );
  NANDN U8070 ( .A(n2990), .B(n2989), .Z(n2991) );
  AND U8071 ( .A(n2992), .B(n2991), .Z(n7144) );
  XOR U8072 ( .A(n7145), .B(n7144), .Z(n7147) );
  XOR U8073 ( .A(n7146), .B(n7147), .Z(n7499) );
  XNOR U8074 ( .A(n7498), .B(n7499), .Z(n7501) );
  NANDN U8075 ( .A(n2994), .B(n2993), .Z(n2998) );
  NAND U8076 ( .A(n2996), .B(n2995), .Z(n2997) );
  AND U8077 ( .A(n2998), .B(n2997), .Z(n6438) );
  NANDN U8078 ( .A(n3000), .B(n2999), .Z(n3004) );
  NAND U8079 ( .A(n3002), .B(n3001), .Z(n3003) );
  NAND U8080 ( .A(n3004), .B(n3003), .Z(n6439) );
  XNOR U8081 ( .A(n6438), .B(n6439), .Z(n6441) );
  NANDN U8082 ( .A(n3006), .B(n3005), .Z(n3010) );
  NANDN U8083 ( .A(n3008), .B(n3007), .Z(n3009) );
  AND U8084 ( .A(n3010), .B(n3009), .Z(n6440) );
  XOR U8085 ( .A(n6441), .B(n6440), .Z(n6639) );
  NANDN U8086 ( .A(n3012), .B(n3011), .Z(n3016) );
  NAND U8087 ( .A(n3014), .B(n3013), .Z(n3015) );
  AND U8088 ( .A(n3016), .B(n3015), .Z(n6637) );
  NANDN U8089 ( .A(n3018), .B(n3017), .Z(n3022) );
  NAND U8090 ( .A(n3020), .B(n3019), .Z(n3021) );
  AND U8091 ( .A(n3022), .B(n3021), .Z(n7700) );
  NANDN U8092 ( .A(n3024), .B(n3023), .Z(n3028) );
  NAND U8093 ( .A(n3026), .B(n3025), .Z(n3027) );
  NAND U8094 ( .A(n3028), .B(n3027), .Z(n7701) );
  XNOR U8095 ( .A(n7700), .B(n7701), .Z(n7703) );
  NANDN U8096 ( .A(n3030), .B(n3029), .Z(n3034) );
  NAND U8097 ( .A(n3032), .B(n3031), .Z(n3033) );
  AND U8098 ( .A(n3034), .B(n3033), .Z(n7702) );
  XNOR U8099 ( .A(n7703), .B(n7702), .Z(n6636) );
  XNOR U8100 ( .A(n6637), .B(n6636), .Z(n6638) );
  XNOR U8101 ( .A(n6639), .B(n6638), .Z(n7500) );
  XOR U8102 ( .A(n7501), .B(n7500), .Z(n7109) );
  NANDN U8103 ( .A(n3036), .B(n3035), .Z(n3040) );
  NANDN U8104 ( .A(n3038), .B(n3037), .Z(n3039) );
  AND U8105 ( .A(n3040), .B(n3039), .Z(n7075) );
  NANDN U8106 ( .A(n3042), .B(n3041), .Z(n3046) );
  NANDN U8107 ( .A(n3044), .B(n3043), .Z(n3045) );
  AND U8108 ( .A(n3046), .B(n3045), .Z(n7073) );
  NANDN U8109 ( .A(n3048), .B(n3047), .Z(n3052) );
  NANDN U8110 ( .A(n3050), .B(n3049), .Z(n3051) );
  AND U8111 ( .A(n3052), .B(n3051), .Z(n7072) );
  XOR U8112 ( .A(n7073), .B(n7072), .Z(n7074) );
  XOR U8113 ( .A(n7075), .B(n7074), .Z(n7755) );
  NANDN U8114 ( .A(n3054), .B(n3053), .Z(n3058) );
  NANDN U8115 ( .A(n3056), .B(n3055), .Z(n3057) );
  AND U8116 ( .A(n3058), .B(n3057), .Z(n7381) );
  NANDN U8117 ( .A(n3060), .B(n3059), .Z(n3064) );
  NAND U8118 ( .A(n3062), .B(n3061), .Z(n3063) );
  AND U8119 ( .A(n3064), .B(n3063), .Z(n7676) );
  NANDN U8120 ( .A(n3066), .B(n3065), .Z(n3070) );
  NAND U8121 ( .A(n3068), .B(n3067), .Z(n3069) );
  NAND U8122 ( .A(n3070), .B(n3069), .Z(n7677) );
  XNOR U8123 ( .A(n7676), .B(n7677), .Z(n7679) );
  NANDN U8124 ( .A(n3072), .B(n3071), .Z(n3076) );
  NAND U8125 ( .A(n3074), .B(n3073), .Z(n3075) );
  AND U8126 ( .A(n3076), .B(n3075), .Z(n7678) );
  XOR U8127 ( .A(n7679), .B(n7678), .Z(n7379) );
  NANDN U8128 ( .A(n3078), .B(n3077), .Z(n3082) );
  NANDN U8129 ( .A(n3080), .B(n3079), .Z(n3081) );
  AND U8130 ( .A(n3082), .B(n3081), .Z(n7378) );
  XNOR U8131 ( .A(n7379), .B(n7378), .Z(n7380) );
  XOR U8132 ( .A(n7381), .B(n7380), .Z(n7753) );
  NANDN U8133 ( .A(n3084), .B(n3083), .Z(n3088) );
  NANDN U8134 ( .A(n3086), .B(n3085), .Z(n3087) );
  AND U8135 ( .A(n3088), .B(n3087), .Z(n7081) );
  NANDN U8136 ( .A(n3090), .B(n3089), .Z(n3094) );
  NANDN U8137 ( .A(n3092), .B(n3091), .Z(n3093) );
  AND U8138 ( .A(n3094), .B(n3093), .Z(n7079) );
  NANDN U8139 ( .A(n3096), .B(n3095), .Z(n3100) );
  NANDN U8140 ( .A(n3098), .B(n3097), .Z(n3099) );
  AND U8141 ( .A(n3100), .B(n3099), .Z(n7078) );
  XOR U8142 ( .A(n7079), .B(n7078), .Z(n7080) );
  XNOR U8143 ( .A(n7081), .B(n7080), .Z(n7752) );
  XNOR U8144 ( .A(n7753), .B(n7752), .Z(n7754) );
  XNOR U8145 ( .A(n7755), .B(n7754), .Z(n7108) );
  XOR U8146 ( .A(n7109), .B(n7108), .Z(n7111) );
  XOR U8147 ( .A(n7110), .B(n7111), .Z(n6553) );
  NANDN U8148 ( .A(n3102), .B(n3101), .Z(n3106) );
  NAND U8149 ( .A(n3104), .B(n3103), .Z(n3105) );
  AND U8150 ( .A(n3106), .B(n3105), .Z(n6780) );
  NANDN U8151 ( .A(n3108), .B(n3107), .Z(n3112) );
  NAND U8152 ( .A(n3110), .B(n3109), .Z(n3111) );
  NAND U8153 ( .A(n3112), .B(n3111), .Z(n6781) );
  XNOR U8154 ( .A(n6780), .B(n6781), .Z(n6783) );
  NANDN U8155 ( .A(n3114), .B(n3113), .Z(n3118) );
  NAND U8156 ( .A(n3116), .B(n3115), .Z(n3117) );
  AND U8157 ( .A(n3118), .B(n3117), .Z(n6782) );
  XOR U8158 ( .A(n6783), .B(n6782), .Z(n6711) );
  NANDN U8159 ( .A(n3120), .B(n3119), .Z(n3124) );
  NAND U8160 ( .A(n3122), .B(n3121), .Z(n3123) );
  AND U8161 ( .A(n3124), .B(n3123), .Z(n7492) );
  NANDN U8162 ( .A(n3126), .B(n3125), .Z(n3130) );
  NAND U8163 ( .A(n3128), .B(n3127), .Z(n3129) );
  NAND U8164 ( .A(n3130), .B(n3129), .Z(n7493) );
  XNOR U8165 ( .A(n7492), .B(n7493), .Z(n7495) );
  NANDN U8166 ( .A(n3132), .B(n3131), .Z(n3136) );
  NAND U8167 ( .A(n3134), .B(n3133), .Z(n3135) );
  AND U8168 ( .A(n3136), .B(n3135), .Z(n7494) );
  XOR U8169 ( .A(n7495), .B(n7494), .Z(n6709) );
  NANDN U8170 ( .A(n3138), .B(n3137), .Z(n3142) );
  NANDN U8171 ( .A(n3140), .B(n3139), .Z(n3141) );
  AND U8172 ( .A(n3142), .B(n3141), .Z(n6708) );
  XNOR U8173 ( .A(n6709), .B(n6708), .Z(n6710) );
  XNOR U8174 ( .A(n6711), .B(n6710), .Z(n6970) );
  NANDN U8175 ( .A(n3144), .B(n3143), .Z(n3148) );
  NAND U8176 ( .A(n3146), .B(n3145), .Z(n3147) );
  AND U8177 ( .A(n3148), .B(n3147), .Z(n8745) );
  NANDN U8178 ( .A(n3150), .B(n3149), .Z(n3154) );
  NAND U8179 ( .A(n3152), .B(n3151), .Z(n3153) );
  NAND U8180 ( .A(n3154), .B(n3153), .Z(n8746) );
  XNOR U8181 ( .A(n8745), .B(n8746), .Z(n8748) );
  NANDN U8182 ( .A(n3156), .B(n3155), .Z(n3160) );
  NAND U8183 ( .A(n3158), .B(n3157), .Z(n3159) );
  AND U8184 ( .A(n3160), .B(n3159), .Z(n8747) );
  XOR U8185 ( .A(n8748), .B(n8747), .Z(n7153) );
  NANDN U8186 ( .A(n3162), .B(n3161), .Z(n3166) );
  NAND U8187 ( .A(n3164), .B(n3163), .Z(n3165) );
  AND U8188 ( .A(n3166), .B(n3165), .Z(n8757) );
  NANDN U8189 ( .A(n3168), .B(n3167), .Z(n3172) );
  NAND U8190 ( .A(n3170), .B(n3169), .Z(n3171) );
  NAND U8191 ( .A(n3172), .B(n3171), .Z(n8758) );
  XNOR U8192 ( .A(n8757), .B(n8758), .Z(n8760) );
  NANDN U8193 ( .A(n3174), .B(n3173), .Z(n3178) );
  NAND U8194 ( .A(n3176), .B(n3175), .Z(n3177) );
  AND U8195 ( .A(n3178), .B(n3177), .Z(n8759) );
  XOR U8196 ( .A(n8760), .B(n8759), .Z(n7151) );
  NANDN U8197 ( .A(n3180), .B(n3179), .Z(n3184) );
  NANDN U8198 ( .A(n3182), .B(n3181), .Z(n3183) );
  AND U8199 ( .A(n3184), .B(n3183), .Z(n7150) );
  XNOR U8200 ( .A(n7151), .B(n7150), .Z(n7152) );
  XOR U8201 ( .A(n7153), .B(n7152), .Z(n6971) );
  XNOR U8202 ( .A(n6970), .B(n6971), .Z(n6973) );
  NANDN U8203 ( .A(n3186), .B(n3185), .Z(n3190) );
  NAND U8204 ( .A(n3188), .B(n3187), .Z(n3189) );
  AND U8205 ( .A(n3190), .B(n3189), .Z(n7734) );
  NANDN U8206 ( .A(n3192), .B(n3191), .Z(n3196) );
  NAND U8207 ( .A(n3194), .B(n3193), .Z(n3195) );
  NAND U8208 ( .A(n3196), .B(n3195), .Z(n7735) );
  XNOR U8209 ( .A(n7734), .B(n7735), .Z(n7737) );
  NANDN U8210 ( .A(n3198), .B(n3197), .Z(n3202) );
  NAND U8211 ( .A(n3200), .B(n3199), .Z(n3201) );
  AND U8212 ( .A(n3202), .B(n3201), .Z(n7736) );
  XOR U8213 ( .A(n7737), .B(n7736), .Z(n8820) );
  NAND U8214 ( .A(n3204), .B(n3203), .Z(n3208) );
  NAND U8215 ( .A(n3206), .B(n3205), .Z(n3207) );
  AND U8216 ( .A(n3208), .B(n3207), .Z(n6648) );
  NANDN U8217 ( .A(n3210), .B(n3209), .Z(n3214) );
  NAND U8218 ( .A(n3212), .B(n3211), .Z(n3213) );
  NAND U8219 ( .A(n3214), .B(n3213), .Z(n6649) );
  XNOR U8220 ( .A(n6648), .B(n6649), .Z(n6651) );
  NANDN U8221 ( .A(n3216), .B(n3215), .Z(n3220) );
  NAND U8222 ( .A(n3218), .B(n3217), .Z(n3219) );
  AND U8223 ( .A(n3220), .B(n3219), .Z(n6650) );
  XOR U8224 ( .A(n6651), .B(n6650), .Z(n8818) );
  NANDN U8225 ( .A(n3222), .B(n3221), .Z(n3226) );
  NANDN U8226 ( .A(n3224), .B(n3223), .Z(n3225) );
  AND U8227 ( .A(n3226), .B(n3225), .Z(n8817) );
  XNOR U8228 ( .A(n8818), .B(n8817), .Z(n8819) );
  XNOR U8229 ( .A(n8820), .B(n8819), .Z(n6972) );
  XOR U8230 ( .A(n6973), .B(n6972), .Z(n6092) );
  NAND U8231 ( .A(n3228), .B(n3227), .Z(n3232) );
  NAND U8232 ( .A(n3230), .B(n3229), .Z(n3231) );
  AND U8233 ( .A(n3232), .B(n3231), .Z(n8949) );
  NANDN U8234 ( .A(n3234), .B(n3233), .Z(n3238) );
  NAND U8235 ( .A(n3236), .B(n3235), .Z(n3237) );
  AND U8236 ( .A(n3238), .B(n3237), .Z(n8948) );
  XOR U8237 ( .A(n8949), .B(n8948), .Z(n8951) );
  NANDN U8238 ( .A(n3240), .B(n3239), .Z(n3244) );
  NAND U8239 ( .A(n3242), .B(n3241), .Z(n3243) );
  AND U8240 ( .A(n3244), .B(n3243), .Z(n8950) );
  XOR U8241 ( .A(n8951), .B(n8950), .Z(n9035) );
  NANDN U8242 ( .A(n3246), .B(n3245), .Z(n3250) );
  NAND U8243 ( .A(n3248), .B(n3247), .Z(n3249) );
  AND U8244 ( .A(n3250), .B(n3249), .Z(n7475) );
  NANDN U8245 ( .A(n3252), .B(n3251), .Z(n3256) );
  NANDN U8246 ( .A(n3254), .B(n3253), .Z(n3255) );
  AND U8247 ( .A(n3256), .B(n3255), .Z(n7474) );
  XOR U8248 ( .A(n7475), .B(n7474), .Z(n7477) );
  NANDN U8249 ( .A(n3258), .B(n3257), .Z(n3262) );
  NAND U8250 ( .A(n3260), .B(n3259), .Z(n3261) );
  AND U8251 ( .A(n3262), .B(n3261), .Z(n7476) );
  XOR U8252 ( .A(n7477), .B(n7476), .Z(n9034) );
  NANDN U8253 ( .A(n3264), .B(n3263), .Z(n3268) );
  NANDN U8254 ( .A(n3266), .B(n3265), .Z(n3267) );
  AND U8255 ( .A(n3268), .B(n3267), .Z(n9033) );
  XOR U8256 ( .A(n9034), .B(n9033), .Z(n9036) );
  XOR U8257 ( .A(n9035), .B(n9036), .Z(n7887) );
  NANDN U8258 ( .A(n3270), .B(n3269), .Z(n3274) );
  NAND U8259 ( .A(n3272), .B(n3271), .Z(n3273) );
  AND U8260 ( .A(n3274), .B(n3273), .Z(n6846) );
  NANDN U8261 ( .A(n3276), .B(n3275), .Z(n3280) );
  NAND U8262 ( .A(n3278), .B(n3277), .Z(n3279) );
  NAND U8263 ( .A(n3280), .B(n3279), .Z(n6847) );
  XNOR U8264 ( .A(n6846), .B(n6847), .Z(n6849) );
  NAND U8265 ( .A(n3282), .B(n3281), .Z(n3286) );
  NAND U8266 ( .A(n3284), .B(n3283), .Z(n3285) );
  AND U8267 ( .A(n3286), .B(n3285), .Z(n6848) );
  XOR U8268 ( .A(n6849), .B(n6848), .Z(n7326) );
  NANDN U8269 ( .A(n3288), .B(n3287), .Z(n3292) );
  NAND U8270 ( .A(n3290), .B(n3289), .Z(n3291) );
  AND U8271 ( .A(n3292), .B(n3291), .Z(n6840) );
  NAND U8272 ( .A(n3294), .B(n3293), .Z(n3298) );
  NAND U8273 ( .A(n3296), .B(n3295), .Z(n3297) );
  NAND U8274 ( .A(n3298), .B(n3297), .Z(n6841) );
  XNOR U8275 ( .A(n6840), .B(n6841), .Z(n6843) );
  NAND U8276 ( .A(n3300), .B(n3299), .Z(n3304) );
  NAND U8277 ( .A(n3302), .B(n3301), .Z(n3303) );
  AND U8278 ( .A(n3304), .B(n3303), .Z(n6842) );
  XOR U8279 ( .A(n6843), .B(n6842), .Z(n7325) );
  NANDN U8280 ( .A(n3306), .B(n3305), .Z(n3310) );
  NANDN U8281 ( .A(n3308), .B(n3307), .Z(n3309) );
  AND U8282 ( .A(n3310), .B(n3309), .Z(n7324) );
  XOR U8283 ( .A(n7325), .B(n7324), .Z(n7327) );
  XOR U8284 ( .A(n7326), .B(n7327), .Z(n7885) );
  NANDN U8285 ( .A(n3312), .B(n3311), .Z(n3316) );
  NANDN U8286 ( .A(n3314), .B(n3313), .Z(n3315) );
  AND U8287 ( .A(n3316), .B(n3315), .Z(n7648) );
  NANDN U8288 ( .A(n3318), .B(n3317), .Z(n3322) );
  NAND U8289 ( .A(n3320), .B(n3319), .Z(n3321) );
  NAND U8290 ( .A(n3322), .B(n3321), .Z(n7649) );
  XNOR U8291 ( .A(n7648), .B(n7649), .Z(n7651) );
  NANDN U8292 ( .A(n3324), .B(n3323), .Z(n3328) );
  NAND U8293 ( .A(n3326), .B(n3325), .Z(n3327) );
  AND U8294 ( .A(n3328), .B(n3327), .Z(n7650) );
  XOR U8295 ( .A(n7651), .B(n7650), .Z(n6740) );
  NANDN U8296 ( .A(n3330), .B(n3329), .Z(n3334) );
  NAND U8297 ( .A(n3332), .B(n3331), .Z(n3333) );
  AND U8298 ( .A(n3334), .B(n3333), .Z(n8924) );
  NANDN U8299 ( .A(n3336), .B(n3335), .Z(n3340) );
  NAND U8300 ( .A(n3338), .B(n3337), .Z(n3339) );
  NAND U8301 ( .A(n3340), .B(n3339), .Z(n8925) );
  XNOR U8302 ( .A(n8924), .B(n8925), .Z(n8927) );
  NANDN U8303 ( .A(n3342), .B(n3341), .Z(n3346) );
  NAND U8304 ( .A(n3344), .B(n3343), .Z(n3345) );
  AND U8305 ( .A(n3346), .B(n3345), .Z(n8926) );
  XOR U8306 ( .A(n8927), .B(n8926), .Z(n6739) );
  NANDN U8307 ( .A(n3348), .B(n3347), .Z(n3352) );
  NANDN U8308 ( .A(n3350), .B(n3349), .Z(n3351) );
  AND U8309 ( .A(n3352), .B(n3351), .Z(n6738) );
  XOR U8310 ( .A(n6739), .B(n6738), .Z(n6741) );
  XNOR U8311 ( .A(n6740), .B(n6741), .Z(n7884) );
  XNOR U8312 ( .A(n7885), .B(n7884), .Z(n7886) );
  XNOR U8313 ( .A(n7887), .B(n7886), .Z(n6090) );
  NANDN U8314 ( .A(n3354), .B(n3353), .Z(n3358) );
  NANDN U8315 ( .A(n3356), .B(n3355), .Z(n3357) );
  AND U8316 ( .A(n3358), .B(n3357), .Z(n8742) );
  NANDN U8317 ( .A(n3360), .B(n3359), .Z(n3364) );
  NAND U8318 ( .A(n3362), .B(n3361), .Z(n3363) );
  AND U8319 ( .A(n3364), .B(n3363), .Z(n8859) );
  NANDN U8320 ( .A(n3366), .B(n3365), .Z(n3370) );
  NANDN U8321 ( .A(n3368), .B(n3367), .Z(n3369) );
  NAND U8322 ( .A(n3370), .B(n3369), .Z(n8860) );
  XNOR U8323 ( .A(n8859), .B(n8860), .Z(n8862) );
  NANDN U8324 ( .A(n3372), .B(n3371), .Z(n3376) );
  NAND U8325 ( .A(n3374), .B(n3373), .Z(n3375) );
  AND U8326 ( .A(n3376), .B(n3375), .Z(n8861) );
  XOR U8327 ( .A(n8862), .B(n8861), .Z(n8740) );
  NANDN U8328 ( .A(n3378), .B(n3377), .Z(n3382) );
  NANDN U8329 ( .A(n3380), .B(n3379), .Z(n3381) );
  AND U8330 ( .A(n3382), .B(n3381), .Z(n8739) );
  XNOR U8331 ( .A(n8740), .B(n8739), .Z(n8741) );
  XOR U8332 ( .A(n8742), .B(n8741), .Z(n7003) );
  NANDN U8333 ( .A(n3384), .B(n3383), .Z(n3388) );
  NANDN U8334 ( .A(n3386), .B(n3385), .Z(n3387) );
  AND U8335 ( .A(n3388), .B(n3387), .Z(n7309) );
  NANDN U8336 ( .A(n3390), .B(n3389), .Z(n3394) );
  NAND U8337 ( .A(n3392), .B(n3391), .Z(n3393) );
  AND U8338 ( .A(n3394), .B(n3393), .Z(n8751) );
  NANDN U8339 ( .A(n3396), .B(n3395), .Z(n3400) );
  NAND U8340 ( .A(n3398), .B(n3397), .Z(n3399) );
  NAND U8341 ( .A(n3400), .B(n3399), .Z(n8752) );
  XNOR U8342 ( .A(n8751), .B(n8752), .Z(n8754) );
  NAND U8343 ( .A(n3402), .B(n3401), .Z(n3406) );
  NAND U8344 ( .A(n3404), .B(n3403), .Z(n3405) );
  AND U8345 ( .A(n3406), .B(n3405), .Z(n8753) );
  XOR U8346 ( .A(n8754), .B(n8753), .Z(n7307) );
  NANDN U8347 ( .A(n3408), .B(n3407), .Z(n3412) );
  NANDN U8348 ( .A(n3410), .B(n3409), .Z(n3411) );
  AND U8349 ( .A(n3412), .B(n3411), .Z(n7306) );
  XNOR U8350 ( .A(n7307), .B(n7306), .Z(n7308) );
  XOR U8351 ( .A(n7309), .B(n7308), .Z(n7001) );
  NANDN U8352 ( .A(n3414), .B(n3413), .Z(n3418) );
  NAND U8353 ( .A(n3416), .B(n3415), .Z(n3417) );
  AND U8354 ( .A(n3418), .B(n3417), .Z(n7782) );
  NAND U8355 ( .A(n3420), .B(n3419), .Z(n3424) );
  NAND U8356 ( .A(n3422), .B(n3421), .Z(n3423) );
  NAND U8357 ( .A(n3424), .B(n3423), .Z(n7783) );
  XNOR U8358 ( .A(n7782), .B(n7783), .Z(n7785) );
  NAND U8359 ( .A(n3426), .B(n3425), .Z(n3430) );
  NAND U8360 ( .A(n3428), .B(n3427), .Z(n3429) );
  AND U8361 ( .A(n3430), .B(n3429), .Z(n7784) );
  XOR U8362 ( .A(n7785), .B(n7784), .Z(n7092) );
  NANDN U8363 ( .A(n3432), .B(n3431), .Z(n3436) );
  NAND U8364 ( .A(n3434), .B(n3433), .Z(n3435) );
  AND U8365 ( .A(n3436), .B(n3435), .Z(n6540) );
  NANDN U8366 ( .A(n3438), .B(n3437), .Z(n3442) );
  NAND U8367 ( .A(n3440), .B(n3439), .Z(n3441) );
  NAND U8368 ( .A(n3442), .B(n3441), .Z(n6541) );
  XNOR U8369 ( .A(n6540), .B(n6541), .Z(n6543) );
  NANDN U8370 ( .A(n3444), .B(n3443), .Z(n3448) );
  NAND U8371 ( .A(n3446), .B(n3445), .Z(n3447) );
  AND U8372 ( .A(n3448), .B(n3447), .Z(n6542) );
  XOR U8373 ( .A(n6543), .B(n6542), .Z(n7091) );
  NANDN U8374 ( .A(n3450), .B(n3449), .Z(n3454) );
  NANDN U8375 ( .A(n3452), .B(n3451), .Z(n3453) );
  AND U8376 ( .A(n3454), .B(n3453), .Z(n7090) );
  XOR U8377 ( .A(n7091), .B(n7090), .Z(n7093) );
  XNOR U8378 ( .A(n7092), .B(n7093), .Z(n7000) );
  XNOR U8379 ( .A(n7001), .B(n7000), .Z(n7002) );
  XOR U8380 ( .A(n7003), .B(n7002), .Z(n6091) );
  XOR U8381 ( .A(n6090), .B(n6091), .Z(n6093) );
  XNOR U8382 ( .A(n6092), .B(n6093), .Z(n6552) );
  NANDN U8383 ( .A(n3456), .B(n3455), .Z(n3460) );
  NAND U8384 ( .A(n3458), .B(n3457), .Z(n3459) );
  AND U8385 ( .A(n3460), .B(n3459), .Z(n7824) );
  NANDN U8386 ( .A(n3462), .B(n3461), .Z(n3466) );
  NAND U8387 ( .A(n3464), .B(n3463), .Z(n3465) );
  NAND U8388 ( .A(n3466), .B(n3465), .Z(n7825) );
  XNOR U8389 ( .A(n7824), .B(n7825), .Z(n7827) );
  NANDN U8390 ( .A(n3468), .B(n3467), .Z(n3472) );
  NAND U8391 ( .A(n3470), .B(n3469), .Z(n3471) );
  AND U8392 ( .A(n3472), .B(n3471), .Z(n7826) );
  XOR U8393 ( .A(n7827), .B(n7826), .Z(n8177) );
  NANDN U8394 ( .A(n3474), .B(n3473), .Z(n3478) );
  NANDN U8395 ( .A(n3476), .B(n3475), .Z(n3477) );
  AND U8396 ( .A(n3478), .B(n3477), .Z(n6510) );
  NANDN U8397 ( .A(n3480), .B(n3479), .Z(n3484) );
  NAND U8398 ( .A(n3482), .B(n3481), .Z(n3483) );
  NAND U8399 ( .A(n3484), .B(n3483), .Z(n6511) );
  XNOR U8400 ( .A(n6510), .B(n6511), .Z(n6513) );
  NANDN U8401 ( .A(n3486), .B(n3485), .Z(n3490) );
  NAND U8402 ( .A(n3488), .B(n3487), .Z(n3489) );
  AND U8403 ( .A(n3490), .B(n3489), .Z(n6512) );
  XOR U8404 ( .A(n6513), .B(n6512), .Z(n8176) );
  NANDN U8405 ( .A(n3492), .B(n3491), .Z(n3496) );
  NANDN U8406 ( .A(n3494), .B(n3493), .Z(n3495) );
  AND U8407 ( .A(n3496), .B(n3495), .Z(n8175) );
  XOR U8408 ( .A(n8176), .B(n8175), .Z(n8178) );
  XOR U8409 ( .A(n8177), .B(n8178), .Z(n7398) );
  NANDN U8410 ( .A(n3498), .B(n3497), .Z(n3502) );
  NAND U8411 ( .A(n3500), .B(n3499), .Z(n3501) );
  AND U8412 ( .A(n3502), .B(n3501), .Z(n7682) );
  NANDN U8413 ( .A(n3504), .B(n3503), .Z(n3508) );
  NAND U8414 ( .A(n3506), .B(n3505), .Z(n3507) );
  NAND U8415 ( .A(n3508), .B(n3507), .Z(n7683) );
  XNOR U8416 ( .A(n7682), .B(n7683), .Z(n7685) );
  NANDN U8417 ( .A(n3510), .B(n3509), .Z(n3514) );
  NAND U8418 ( .A(n3512), .B(n3511), .Z(n3513) );
  AND U8419 ( .A(n3514), .B(n3513), .Z(n7684) );
  XOR U8420 ( .A(n7685), .B(n7684), .Z(n8897) );
  NANDN U8421 ( .A(n3516), .B(n3515), .Z(n3520) );
  NAND U8422 ( .A(n3518), .B(n3517), .Z(n3519) );
  AND U8423 ( .A(n3520), .B(n3519), .Z(n8535) );
  NANDN U8424 ( .A(n3522), .B(n3521), .Z(n3526) );
  NAND U8425 ( .A(n3524), .B(n3523), .Z(n3525) );
  NAND U8426 ( .A(n3526), .B(n3525), .Z(n8536) );
  XNOR U8427 ( .A(n8535), .B(n8536), .Z(n8538) );
  NAND U8428 ( .A(n3528), .B(n3527), .Z(n3532) );
  NAND U8429 ( .A(n3530), .B(n3529), .Z(n3531) );
  AND U8430 ( .A(n3532), .B(n3531), .Z(n8537) );
  XOR U8431 ( .A(n8538), .B(n8537), .Z(n8896) );
  NANDN U8432 ( .A(n3534), .B(n3533), .Z(n3538) );
  NANDN U8433 ( .A(n3536), .B(n3535), .Z(n3537) );
  AND U8434 ( .A(n3538), .B(n3537), .Z(n8895) );
  XOR U8435 ( .A(n8896), .B(n8895), .Z(n8898) );
  XOR U8436 ( .A(n8897), .B(n8898), .Z(n7397) );
  NANDN U8437 ( .A(n3540), .B(n3539), .Z(n3544) );
  NANDN U8438 ( .A(n3542), .B(n3541), .Z(n3543) );
  AND U8439 ( .A(n3544), .B(n3543), .Z(n8202) );
  NAND U8440 ( .A(n3546), .B(n3545), .Z(n3550) );
  NAND U8441 ( .A(n3548), .B(n3547), .Z(n3549) );
  AND U8442 ( .A(n3550), .B(n3549), .Z(n6528) );
  NANDN U8443 ( .A(n3552), .B(n3551), .Z(n3556) );
  NAND U8444 ( .A(n3554), .B(n3553), .Z(n3555) );
  NAND U8445 ( .A(n3556), .B(n3555), .Z(n6529) );
  XNOR U8446 ( .A(n6528), .B(n6529), .Z(n6531) );
  NANDN U8447 ( .A(n3558), .B(n3557), .Z(n3562) );
  NAND U8448 ( .A(n3560), .B(n3559), .Z(n3561) );
  AND U8449 ( .A(n3562), .B(n3561), .Z(n6530) );
  XOR U8450 ( .A(n6531), .B(n6530), .Z(n8200) );
  NANDN U8451 ( .A(n3564), .B(n3563), .Z(n3568) );
  NANDN U8452 ( .A(n3566), .B(n3565), .Z(n3567) );
  AND U8453 ( .A(n3568), .B(n3567), .Z(n8199) );
  XNOR U8454 ( .A(n8200), .B(n8199), .Z(n8201) );
  XNOR U8455 ( .A(n8202), .B(n8201), .Z(n7396) );
  XOR U8456 ( .A(n7397), .B(n7396), .Z(n7399) );
  XNOR U8457 ( .A(n7398), .B(n7399), .Z(n6147) );
  NANDN U8458 ( .A(n3570), .B(n3569), .Z(n3574) );
  NANDN U8459 ( .A(n3572), .B(n3571), .Z(n3573) );
  AND U8460 ( .A(n3574), .B(n3573), .Z(n8148) );
  NANDN U8461 ( .A(n3576), .B(n3575), .Z(n3580) );
  NANDN U8462 ( .A(n3578), .B(n3577), .Z(n3579) );
  AND U8463 ( .A(n3580), .B(n3579), .Z(n8145) );
  NANDN U8464 ( .A(n3582), .B(n3581), .Z(n3586) );
  NANDN U8465 ( .A(n3584), .B(n3583), .Z(n3585) );
  NAND U8466 ( .A(n3586), .B(n3585), .Z(n8146) );
  XNOR U8467 ( .A(n8145), .B(n8146), .Z(n8147) );
  XNOR U8468 ( .A(n8148), .B(n8147), .Z(n7916) );
  NANDN U8469 ( .A(n3588), .B(n3587), .Z(n3592) );
  NAND U8470 ( .A(n3590), .B(n3589), .Z(n3591) );
  AND U8471 ( .A(n3592), .B(n3591), .Z(n8903) );
  NANDN U8472 ( .A(n3594), .B(n3593), .Z(n3598) );
  NAND U8473 ( .A(n3596), .B(n3595), .Z(n3597) );
  AND U8474 ( .A(n3598), .B(n3597), .Z(n8902) );
  NANDN U8475 ( .A(n3600), .B(n3599), .Z(n3604) );
  NAND U8476 ( .A(n3602), .B(n3601), .Z(n3603) );
  AND U8477 ( .A(n3604), .B(n3603), .Z(n8529) );
  NANDN U8478 ( .A(n3606), .B(n3605), .Z(n3610) );
  NAND U8479 ( .A(n3608), .B(n3607), .Z(n3609) );
  NAND U8480 ( .A(n3610), .B(n3609), .Z(n8530) );
  XNOR U8481 ( .A(n8529), .B(n8530), .Z(n8532) );
  NANDN U8482 ( .A(n3612), .B(n3611), .Z(n3616) );
  NAND U8483 ( .A(n3614), .B(n3613), .Z(n3615) );
  AND U8484 ( .A(n3616), .B(n3615), .Z(n8531) );
  XNOR U8485 ( .A(n8532), .B(n8531), .Z(n8901) );
  XOR U8486 ( .A(n8902), .B(n8901), .Z(n8904) );
  XOR U8487 ( .A(n8903), .B(n8904), .Z(n8933) );
  NANDN U8488 ( .A(n3618), .B(n3617), .Z(n3622) );
  NAND U8489 ( .A(n3620), .B(n3619), .Z(n3621) );
  AND U8490 ( .A(n3622), .B(n3621), .Z(n8241) );
  NANDN U8491 ( .A(n3624), .B(n3623), .Z(n3628) );
  NAND U8492 ( .A(n3626), .B(n3625), .Z(n3627) );
  NAND U8493 ( .A(n3628), .B(n3627), .Z(n8242) );
  XNOR U8494 ( .A(n8241), .B(n8242), .Z(n8243) );
  NANDN U8495 ( .A(n3630), .B(n3629), .Z(n3634) );
  NANDN U8496 ( .A(n3632), .B(n3631), .Z(n3633) );
  NAND U8497 ( .A(n3634), .B(n3633), .Z(n8244) );
  XNOR U8498 ( .A(n8243), .B(n8244), .Z(n8930) );
  NAND U8499 ( .A(n3636), .B(n3635), .Z(n3640) );
  NAND U8500 ( .A(n3638), .B(n3637), .Z(n3639) );
  AND U8501 ( .A(n3640), .B(n3639), .Z(n7712) );
  NANDN U8502 ( .A(n3642), .B(n3641), .Z(n3646) );
  NAND U8503 ( .A(n3644), .B(n3643), .Z(n3645) );
  NAND U8504 ( .A(n3646), .B(n3645), .Z(n7713) );
  XNOR U8505 ( .A(n7712), .B(n7713), .Z(n7714) );
  NANDN U8506 ( .A(n3648), .B(n3647), .Z(n3652) );
  NAND U8507 ( .A(n3650), .B(n3649), .Z(n3651) );
  NAND U8508 ( .A(n3652), .B(n3651), .Z(n7715) );
  XOR U8509 ( .A(n7714), .B(n7715), .Z(n8931) );
  XNOR U8510 ( .A(n8930), .B(n8931), .Z(n8932) );
  XOR U8511 ( .A(n8933), .B(n8932), .Z(n7914) );
  NANDN U8512 ( .A(n3654), .B(n3653), .Z(n3658) );
  NAND U8513 ( .A(n3656), .B(n3655), .Z(n3657) );
  AND U8514 ( .A(n3658), .B(n3657), .Z(n7522) );
  NANDN U8515 ( .A(n3660), .B(n3659), .Z(n3664) );
  NAND U8516 ( .A(n3662), .B(n3661), .Z(n3663) );
  NAND U8517 ( .A(n3664), .B(n3663), .Z(n7523) );
  XNOR U8518 ( .A(n7522), .B(n7523), .Z(n7525) );
  NANDN U8519 ( .A(n3666), .B(n3665), .Z(n3670) );
  NAND U8520 ( .A(n3668), .B(n3667), .Z(n3669) );
  AND U8521 ( .A(n3670), .B(n3669), .Z(n7524) );
  XOR U8522 ( .A(n7525), .B(n7524), .Z(n8843) );
  NANDN U8523 ( .A(n3672), .B(n3671), .Z(n3676) );
  NAND U8524 ( .A(n3674), .B(n3673), .Z(n3675) );
  AND U8525 ( .A(n3676), .B(n3675), .Z(n7812) );
  NANDN U8526 ( .A(n3678), .B(n3677), .Z(n3682) );
  NAND U8527 ( .A(n3680), .B(n3679), .Z(n3681) );
  NAND U8528 ( .A(n3682), .B(n3681), .Z(n7813) );
  XNOR U8529 ( .A(n7812), .B(n7813), .Z(n7815) );
  NANDN U8530 ( .A(n3684), .B(n3683), .Z(n3688) );
  NAND U8531 ( .A(n3686), .B(n3685), .Z(n3687) );
  AND U8532 ( .A(n3688), .B(n3687), .Z(n7814) );
  XOR U8533 ( .A(n7815), .B(n7814), .Z(n8842) );
  NANDN U8534 ( .A(n3690), .B(n3689), .Z(n3694) );
  NANDN U8535 ( .A(n3692), .B(n3691), .Z(n3693) );
  AND U8536 ( .A(n3694), .B(n3693), .Z(n8841) );
  XOR U8537 ( .A(n8842), .B(n8841), .Z(n8844) );
  XOR U8538 ( .A(n8843), .B(n8844), .Z(n7915) );
  XOR U8539 ( .A(n7914), .B(n7915), .Z(n3695) );
  XNOR U8540 ( .A(n7916), .B(n3695), .Z(n6144) );
  NAND U8541 ( .A(n3697), .B(n3696), .Z(n3701) );
  NAND U8542 ( .A(n3699), .B(n3698), .Z(n3700) );
  AND U8543 ( .A(n3701), .B(n3700), .Z(n6534) );
  NANDN U8544 ( .A(n3703), .B(n3702), .Z(n3707) );
  NAND U8545 ( .A(n3705), .B(n3704), .Z(n3706) );
  NAND U8546 ( .A(n3707), .B(n3706), .Z(n6535) );
  XNOR U8547 ( .A(n6534), .B(n6535), .Z(n6537) );
  NANDN U8548 ( .A(n3709), .B(n3708), .Z(n3713) );
  NAND U8549 ( .A(n3711), .B(n3710), .Z(n3712) );
  AND U8550 ( .A(n3713), .B(n3712), .Z(n6536) );
  XOR U8551 ( .A(n6537), .B(n6536), .Z(n8172) );
  NANDN U8552 ( .A(n3715), .B(n3714), .Z(n3719) );
  NAND U8553 ( .A(n3717), .B(n3716), .Z(n3718) );
  AND U8554 ( .A(n3719), .B(n3718), .Z(n6354) );
  NANDN U8555 ( .A(n3721), .B(n3720), .Z(n3725) );
  NAND U8556 ( .A(n3723), .B(n3722), .Z(n3724) );
  NAND U8557 ( .A(n3725), .B(n3724), .Z(n6355) );
  XNOR U8558 ( .A(n6354), .B(n6355), .Z(n6357) );
  NANDN U8559 ( .A(n3727), .B(n3726), .Z(n3731) );
  NAND U8560 ( .A(n3729), .B(n3728), .Z(n3730) );
  AND U8561 ( .A(n3731), .B(n3730), .Z(n6356) );
  XOR U8562 ( .A(n6357), .B(n6356), .Z(n8170) );
  NANDN U8563 ( .A(n3733), .B(n3732), .Z(n3737) );
  NANDN U8564 ( .A(n3735), .B(n3734), .Z(n3736) );
  AND U8565 ( .A(n3737), .B(n3736), .Z(n8169) );
  XNOR U8566 ( .A(n8170), .B(n8169), .Z(n8171) );
  XNOR U8567 ( .A(n8172), .B(n8171), .Z(n7908) );
  NANDN U8568 ( .A(n3739), .B(n3738), .Z(n3743) );
  NANDN U8569 ( .A(n3741), .B(n3740), .Z(n3742) );
  AND U8570 ( .A(n3743), .B(n3742), .Z(n6906) );
  NANDN U8571 ( .A(n3745), .B(n3744), .Z(n3749) );
  NAND U8572 ( .A(n3747), .B(n3746), .Z(n3748) );
  AND U8573 ( .A(n3749), .B(n3748), .Z(n8625) );
  NANDN U8574 ( .A(n3751), .B(n3750), .Z(n3755) );
  NAND U8575 ( .A(n3753), .B(n3752), .Z(n3754) );
  NAND U8576 ( .A(n3755), .B(n3754), .Z(n8626) );
  XNOR U8577 ( .A(n8625), .B(n8626), .Z(n8628) );
  NANDN U8578 ( .A(n3757), .B(n3756), .Z(n3761) );
  NAND U8579 ( .A(n3759), .B(n3758), .Z(n3760) );
  AND U8580 ( .A(n3761), .B(n3760), .Z(n8627) );
  XOR U8581 ( .A(n8628), .B(n8627), .Z(n6905) );
  NANDN U8582 ( .A(n3763), .B(n3762), .Z(n3767) );
  NANDN U8583 ( .A(n3765), .B(n3764), .Z(n3766) );
  AND U8584 ( .A(n3767), .B(n3766), .Z(n6904) );
  XOR U8585 ( .A(n6905), .B(n6904), .Z(n6907) );
  XOR U8586 ( .A(n6906), .B(n6907), .Z(n7909) );
  XNOR U8587 ( .A(n7908), .B(n7909), .Z(n7910) );
  NANDN U8588 ( .A(n3769), .B(n3768), .Z(n3773) );
  NAND U8589 ( .A(n3771), .B(n3770), .Z(n3772) );
  AND U8590 ( .A(n3773), .B(n3772), .Z(n7099) );
  NANDN U8591 ( .A(n3775), .B(n3774), .Z(n3779) );
  NAND U8592 ( .A(n3777), .B(n3776), .Z(n3778) );
  AND U8593 ( .A(n3779), .B(n3778), .Z(n7706) );
  NANDN U8594 ( .A(n3781), .B(n3780), .Z(n3785) );
  NAND U8595 ( .A(n3783), .B(n3782), .Z(n3784) );
  NAND U8596 ( .A(n3785), .B(n3784), .Z(n7707) );
  XNOR U8597 ( .A(n7706), .B(n7707), .Z(n7709) );
  NANDN U8598 ( .A(n3787), .B(n3786), .Z(n3791) );
  NAND U8599 ( .A(n3789), .B(n3788), .Z(n3790) );
  AND U8600 ( .A(n3791), .B(n3790), .Z(n7708) );
  XOR U8601 ( .A(n7709), .B(n7708), .Z(n7097) );
  NANDN U8602 ( .A(n3793), .B(n3792), .Z(n3797) );
  NANDN U8603 ( .A(n3795), .B(n3794), .Z(n3796) );
  AND U8604 ( .A(n3797), .B(n3796), .Z(n7096) );
  XNOR U8605 ( .A(n7097), .B(n7096), .Z(n7098) );
  XOR U8606 ( .A(n7099), .B(n7098), .Z(n7911) );
  XNOR U8607 ( .A(n7910), .B(n7911), .Z(n6145) );
  XOR U8608 ( .A(n6144), .B(n6145), .Z(n6146) );
  XOR U8609 ( .A(n6147), .B(n6146), .Z(n6554) );
  XOR U8610 ( .A(n6555), .B(n6554), .Z(n7048) );
  XOR U8611 ( .A(n7049), .B(n7048), .Z(n7051) );
  XNOR U8612 ( .A(n7050), .B(n7051), .Z(n7234) );
  NAND U8613 ( .A(n3799), .B(n3798), .Z(n3803) );
  NANDN U8614 ( .A(n3801), .B(n3800), .Z(n3802) );
  AND U8615 ( .A(n3803), .B(n3802), .Z(n7249) );
  NANDN U8616 ( .A(n3805), .B(n3804), .Z(n3809) );
  NAND U8617 ( .A(n3807), .B(n3806), .Z(n3808) );
  NAND U8618 ( .A(n3809), .B(n3808), .Z(n7247) );
  NAND U8619 ( .A(n3811), .B(n3810), .Z(n3815) );
  NAND U8620 ( .A(n3813), .B(n3812), .Z(n3814) );
  AND U8621 ( .A(n3815), .B(n3814), .Z(n6175) );
  NAND U8622 ( .A(n3817), .B(n3816), .Z(n3821) );
  NAND U8623 ( .A(n3819), .B(n3818), .Z(n3820) );
  AND U8624 ( .A(n3821), .B(n3820), .Z(n6897) );
  NANDN U8625 ( .A(n3823), .B(n3822), .Z(n3827) );
  NAND U8626 ( .A(n3825), .B(n3824), .Z(n3826) );
  AND U8627 ( .A(n3827), .B(n3826), .Z(n6332) );
  NANDN U8628 ( .A(n3829), .B(n3828), .Z(n3833) );
  NAND U8629 ( .A(n3831), .B(n3830), .Z(n3832) );
  AND U8630 ( .A(n3833), .B(n3832), .Z(n8127) );
  NANDN U8631 ( .A(n3835), .B(n3834), .Z(n3839) );
  NANDN U8632 ( .A(n3837), .B(n3836), .Z(n3838) );
  NAND U8633 ( .A(n3839), .B(n3838), .Z(n8128) );
  XNOR U8634 ( .A(n8127), .B(n8128), .Z(n8130) );
  NAND U8635 ( .A(n3841), .B(n3840), .Z(n3845) );
  NAND U8636 ( .A(n3843), .B(n3842), .Z(n3844) );
  AND U8637 ( .A(n3845), .B(n3844), .Z(n8129) );
  XOR U8638 ( .A(n8130), .B(n8129), .Z(n6984) );
  NANDN U8639 ( .A(n3847), .B(n3846), .Z(n3851) );
  NAND U8640 ( .A(n3849), .B(n3848), .Z(n3850) );
  AND U8641 ( .A(n3851), .B(n3850), .Z(n6594) );
  NANDN U8642 ( .A(n3853), .B(n3852), .Z(n3857) );
  NAND U8643 ( .A(n3855), .B(n3854), .Z(n3856) );
  NAND U8644 ( .A(n3857), .B(n3856), .Z(n6595) );
  XNOR U8645 ( .A(n6594), .B(n6595), .Z(n6597) );
  NANDN U8646 ( .A(n3859), .B(n3858), .Z(n3863) );
  NAND U8647 ( .A(n3861), .B(n3860), .Z(n3862) );
  AND U8648 ( .A(n3863), .B(n3862), .Z(n6596) );
  XOR U8649 ( .A(n6597), .B(n6596), .Z(n6983) );
  NAND U8650 ( .A(n3865), .B(n3864), .Z(n3869) );
  NAND U8651 ( .A(n3867), .B(n3866), .Z(n3868) );
  AND U8652 ( .A(n3869), .B(n3868), .Z(n8229) );
  NAND U8653 ( .A(n3871), .B(n3870), .Z(n3875) );
  NAND U8654 ( .A(n3873), .B(n3872), .Z(n3874) );
  NAND U8655 ( .A(n3875), .B(n3874), .Z(n8230) );
  XNOR U8656 ( .A(n8229), .B(n8230), .Z(n8232) );
  NAND U8657 ( .A(n3877), .B(n3876), .Z(n3881) );
  NAND U8658 ( .A(n3879), .B(n3878), .Z(n3880) );
  AND U8659 ( .A(n3881), .B(n3880), .Z(n8231) );
  XNOR U8660 ( .A(n8232), .B(n8231), .Z(n6982) );
  XOR U8661 ( .A(n6983), .B(n6982), .Z(n6985) );
  XOR U8662 ( .A(n6984), .B(n6985), .Z(n6331) );
  NANDN U8663 ( .A(n3883), .B(n3882), .Z(n3887) );
  NAND U8664 ( .A(n3885), .B(n3884), .Z(n3886) );
  NAND U8665 ( .A(n3887), .B(n3886), .Z(n6330) );
  XOR U8666 ( .A(n6331), .B(n6330), .Z(n6333) );
  XNOR U8667 ( .A(n6332), .B(n6333), .Z(n6895) );
  NAND U8668 ( .A(n3889), .B(n3888), .Z(n3893) );
  NAND U8669 ( .A(n3891), .B(n3890), .Z(n3892) );
  NAND U8670 ( .A(n3893), .B(n3892), .Z(n6894) );
  XOR U8671 ( .A(n6895), .B(n6894), .Z(n6896) );
  XOR U8672 ( .A(n6897), .B(n6896), .Z(n6174) );
  XOR U8673 ( .A(n6175), .B(n6174), .Z(n6177) );
  NAND U8674 ( .A(n3895), .B(n3894), .Z(n3899) );
  NAND U8675 ( .A(n3897), .B(n3896), .Z(n3898) );
  AND U8676 ( .A(n3899), .B(n3898), .Z(n6176) );
  XNOR U8677 ( .A(n6177), .B(n6176), .Z(n7246) );
  XOR U8678 ( .A(n7247), .B(n7246), .Z(n7248) );
  XOR U8679 ( .A(n7249), .B(n7248), .Z(n7235) );
  XOR U8680 ( .A(n7234), .B(n7235), .Z(n7237) );
  XOR U8681 ( .A(n7236), .B(n7237), .Z(n7228) );
  NANDN U8682 ( .A(n3901), .B(n3900), .Z(n3905) );
  NAND U8683 ( .A(n3903), .B(n3902), .Z(n3904) );
  NAND U8684 ( .A(n3905), .B(n3904), .Z(n7229) );
  XNOR U8685 ( .A(n7228), .B(n7229), .Z(n7231) );
  NAND U8686 ( .A(n3907), .B(n3906), .Z(n3911) );
  NAND U8687 ( .A(n3909), .B(n3908), .Z(n3910) );
  AND U8688 ( .A(n3911), .B(n3910), .Z(n7758) );
  NANDN U8689 ( .A(n3913), .B(n3912), .Z(n3917) );
  NAND U8690 ( .A(n3915), .B(n3914), .Z(n3916) );
  AND U8691 ( .A(n3917), .B(n3916), .Z(n6207) );
  NANDN U8692 ( .A(n3919), .B(n3918), .Z(n3923) );
  NAND U8693 ( .A(n3921), .B(n3920), .Z(n3922) );
  AND U8694 ( .A(n3923), .B(n3922), .Z(n6205) );
  NANDN U8695 ( .A(n3925), .B(n3924), .Z(n3929) );
  NANDN U8696 ( .A(n3927), .B(n3926), .Z(n3928) );
  NAND U8697 ( .A(n3929), .B(n3928), .Z(n6204) );
  XNOR U8698 ( .A(n6205), .B(n6204), .Z(n6206) );
  XNOR U8699 ( .A(n6207), .B(n6206), .Z(n7759) );
  XOR U8700 ( .A(n7758), .B(n7759), .Z(n7761) );
  NAND U8701 ( .A(n3931), .B(n3930), .Z(n3935) );
  NAND U8702 ( .A(n3933), .B(n3932), .Z(n3934) );
  AND U8703 ( .A(n3935), .B(n3934), .Z(n7760) );
  XNOR U8704 ( .A(n7761), .B(n7760), .Z(n6073) );
  NAND U8705 ( .A(n3937), .B(n3936), .Z(n3941) );
  NAND U8706 ( .A(n3939), .B(n3938), .Z(n3940) );
  NAND U8707 ( .A(n3941), .B(n3940), .Z(n8634) );
  NAND U8708 ( .A(n3943), .B(n3942), .Z(n3947) );
  NAND U8709 ( .A(n3945), .B(n3944), .Z(n3946) );
  NAND U8710 ( .A(n3947), .B(n3946), .Z(n8632) );
  NANDN U8711 ( .A(n3949), .B(n3948), .Z(n3953) );
  NAND U8712 ( .A(n3951), .B(n3950), .Z(n3952) );
  AND U8713 ( .A(n3953), .B(n3952), .Z(n6224) );
  NANDN U8714 ( .A(n3955), .B(n3954), .Z(n3959) );
  NAND U8715 ( .A(n3957), .B(n3956), .Z(n3958) );
  AND U8716 ( .A(n3959), .B(n3958), .Z(n8769) );
  NANDN U8717 ( .A(n3961), .B(n3960), .Z(n3965) );
  NAND U8718 ( .A(n3963), .B(n3962), .Z(n3964) );
  NAND U8719 ( .A(n3965), .B(n3964), .Z(n8770) );
  XNOR U8720 ( .A(n8769), .B(n8770), .Z(n8772) );
  NANDN U8721 ( .A(n3967), .B(n3966), .Z(n3971) );
  NAND U8722 ( .A(n3969), .B(n3968), .Z(n3970) );
  AND U8723 ( .A(n3971), .B(n3970), .Z(n8771) );
  XOR U8724 ( .A(n8772), .B(n8771), .Z(n7284) );
  NANDN U8725 ( .A(n3973), .B(n3972), .Z(n3977) );
  NAND U8726 ( .A(n3975), .B(n3974), .Z(n3976) );
  AND U8727 ( .A(n3977), .B(n3976), .Z(n8775) );
  NANDN U8728 ( .A(n3979), .B(n3978), .Z(n3983) );
  NAND U8729 ( .A(n3981), .B(n3980), .Z(n3982) );
  NAND U8730 ( .A(n3983), .B(n3982), .Z(n8776) );
  XNOR U8731 ( .A(n8775), .B(n8776), .Z(n8778) );
  NANDN U8732 ( .A(n3985), .B(n3984), .Z(n3989) );
  NAND U8733 ( .A(n3987), .B(n3986), .Z(n3988) );
  AND U8734 ( .A(n3989), .B(n3988), .Z(n8777) );
  XOR U8735 ( .A(n8778), .B(n8777), .Z(n7283) );
  NANDN U8736 ( .A(n3991), .B(n3990), .Z(n3995) );
  NANDN U8737 ( .A(n3993), .B(n3992), .Z(n3994) );
  AND U8738 ( .A(n3995), .B(n3994), .Z(n7282) );
  XOR U8739 ( .A(n7283), .B(n7282), .Z(n7285) );
  XOR U8740 ( .A(n7284), .B(n7285), .Z(n6223) );
  NANDN U8741 ( .A(n3997), .B(n3996), .Z(n4001) );
  NANDN U8742 ( .A(n3999), .B(n3998), .Z(n4000) );
  NAND U8743 ( .A(n4001), .B(n4000), .Z(n6222) );
  XOR U8744 ( .A(n6223), .B(n6222), .Z(n6225) );
  XNOR U8745 ( .A(n6224), .B(n6225), .Z(n8631) );
  XOR U8746 ( .A(n8632), .B(n8631), .Z(n8633) );
  XOR U8747 ( .A(n8634), .B(n8633), .Z(n6072) );
  XOR U8748 ( .A(n6073), .B(n6072), .Z(n6075) );
  NAND U8749 ( .A(n4003), .B(n4002), .Z(n4007) );
  NAND U8750 ( .A(n4005), .B(n4004), .Z(n4006) );
  NAND U8751 ( .A(n4007), .B(n4006), .Z(n7429) );
  NANDN U8752 ( .A(n4009), .B(n4008), .Z(n4013) );
  NAND U8753 ( .A(n4011), .B(n4010), .Z(n4012) );
  AND U8754 ( .A(n4013), .B(n4012), .Z(n6194) );
  NANDN U8755 ( .A(n4015), .B(n4014), .Z(n4019) );
  NAND U8756 ( .A(n4017), .B(n4016), .Z(n4018) );
  AND U8757 ( .A(n4019), .B(n4018), .Z(n8368) );
  NANDN U8758 ( .A(n4021), .B(n4020), .Z(n4025) );
  NAND U8759 ( .A(n4023), .B(n4022), .Z(n4024) );
  AND U8760 ( .A(n4025), .B(n4024), .Z(n8367) );
  XOR U8761 ( .A(n8368), .B(n8367), .Z(n8370) );
  NANDN U8762 ( .A(n4027), .B(n4026), .Z(n4031) );
  NAND U8763 ( .A(n4029), .B(n4028), .Z(n4030) );
  AND U8764 ( .A(n4031), .B(n4030), .Z(n8369) );
  XOR U8765 ( .A(n8370), .B(n8369), .Z(n8009) );
  NANDN U8766 ( .A(n4033), .B(n4032), .Z(n4037) );
  NANDN U8767 ( .A(n4035), .B(n4034), .Z(n4036) );
  AND U8768 ( .A(n4037), .B(n4036), .Z(n8832) );
  NANDN U8769 ( .A(n4039), .B(n4038), .Z(n4043) );
  NAND U8770 ( .A(n4041), .B(n4040), .Z(n4042) );
  AND U8771 ( .A(n4043), .B(n4042), .Z(n8830) );
  NANDN U8772 ( .A(n4045), .B(n4044), .Z(n4049) );
  NANDN U8773 ( .A(n4047), .B(n4046), .Z(n4048) );
  AND U8774 ( .A(n4049), .B(n4048), .Z(n8829) );
  XOR U8775 ( .A(n8830), .B(n8829), .Z(n8831) );
  XOR U8776 ( .A(n8832), .B(n8831), .Z(n8008) );
  NANDN U8777 ( .A(n4051), .B(n4050), .Z(n4055) );
  NAND U8778 ( .A(n4053), .B(n4052), .Z(n4054) );
  AND U8779 ( .A(n4055), .B(n4054), .Z(n8308) );
  NANDN U8780 ( .A(n4057), .B(n4056), .Z(n4061) );
  NAND U8781 ( .A(n4059), .B(n4058), .Z(n4060) );
  AND U8782 ( .A(n4061), .B(n4060), .Z(n8307) );
  XOR U8783 ( .A(n8308), .B(n8307), .Z(n8310) );
  NANDN U8784 ( .A(n4063), .B(n4062), .Z(n4067) );
  NAND U8785 ( .A(n4065), .B(n4064), .Z(n4066) );
  AND U8786 ( .A(n4067), .B(n4066), .Z(n8309) );
  XNOR U8787 ( .A(n8310), .B(n8309), .Z(n8007) );
  XOR U8788 ( .A(n8008), .B(n8007), .Z(n8010) );
  XOR U8789 ( .A(n8009), .B(n8010), .Z(n6193) );
  NANDN U8790 ( .A(n4069), .B(n4068), .Z(n4073) );
  NAND U8791 ( .A(n4071), .B(n4070), .Z(n4072) );
  NAND U8792 ( .A(n4073), .B(n4072), .Z(n6192) );
  XOR U8793 ( .A(n6193), .B(n6192), .Z(n6195) );
  XNOR U8794 ( .A(n6194), .B(n6195), .Z(n7427) );
  NAND U8795 ( .A(n4075), .B(n4074), .Z(n4079) );
  NANDN U8796 ( .A(n4077), .B(n4076), .Z(n4078) );
  NAND U8797 ( .A(n4079), .B(n4078), .Z(n7426) );
  XOR U8798 ( .A(n7427), .B(n7426), .Z(n7428) );
  XOR U8799 ( .A(n7429), .B(n7428), .Z(n6074) );
  XOR U8800 ( .A(n6075), .B(n6074), .Z(n7255) );
  NAND U8801 ( .A(n4081), .B(n4080), .Z(n4085) );
  NAND U8802 ( .A(n4083), .B(n4082), .Z(n4084) );
  NAND U8803 ( .A(n4085), .B(n4084), .Z(n6081) );
  NAND U8804 ( .A(n4087), .B(n4086), .Z(n4091) );
  NAND U8805 ( .A(n4089), .B(n4088), .Z(n4090) );
  NAND U8806 ( .A(n4091), .B(n4090), .Z(n7663) );
  NANDN U8807 ( .A(n4093), .B(n4092), .Z(n4097) );
  NAND U8808 ( .A(n4095), .B(n4094), .Z(n4096) );
  AND U8809 ( .A(n4097), .B(n4096), .Z(n6254) );
  NANDN U8810 ( .A(n4099), .B(n4098), .Z(n4103) );
  NAND U8811 ( .A(n4101), .B(n4100), .Z(n4102) );
  AND U8812 ( .A(n4103), .B(n4102), .Z(n8260) );
  NANDN U8813 ( .A(n4105), .B(n4104), .Z(n4109) );
  NAND U8814 ( .A(n4107), .B(n4106), .Z(n4108) );
  AND U8815 ( .A(n4109), .B(n4108), .Z(n8259) );
  XOR U8816 ( .A(n8260), .B(n8259), .Z(n8262) );
  NANDN U8817 ( .A(n4111), .B(n4110), .Z(n4115) );
  NAND U8818 ( .A(n4113), .B(n4112), .Z(n4114) );
  AND U8819 ( .A(n4115), .B(n4114), .Z(n8261) );
  XOR U8820 ( .A(n8262), .B(n8261), .Z(n8003) );
  NANDN U8821 ( .A(n4117), .B(n4116), .Z(n4121) );
  NAND U8822 ( .A(n4119), .B(n4118), .Z(n4120) );
  AND U8823 ( .A(n4121), .B(n4120), .Z(n8374) );
  NANDN U8824 ( .A(n4123), .B(n4122), .Z(n4127) );
  NAND U8825 ( .A(n4125), .B(n4124), .Z(n4126) );
  AND U8826 ( .A(n4127), .B(n4126), .Z(n8373) );
  XOR U8827 ( .A(n8374), .B(n8373), .Z(n8376) );
  NANDN U8828 ( .A(n4129), .B(n4128), .Z(n4133) );
  NAND U8829 ( .A(n4131), .B(n4130), .Z(n4132) );
  AND U8830 ( .A(n4133), .B(n4132), .Z(n8375) );
  XOR U8831 ( .A(n8376), .B(n8375), .Z(n8002) );
  NANDN U8832 ( .A(n4135), .B(n4134), .Z(n4139) );
  NAND U8833 ( .A(n4137), .B(n4136), .Z(n4138) );
  AND U8834 ( .A(n4139), .B(n4138), .Z(n8434) );
  NANDN U8835 ( .A(n4141), .B(n4140), .Z(n4145) );
  NAND U8836 ( .A(n4143), .B(n4142), .Z(n4144) );
  AND U8837 ( .A(n4145), .B(n4144), .Z(n8433) );
  XOR U8838 ( .A(n8434), .B(n8433), .Z(n8436) );
  NANDN U8839 ( .A(n4147), .B(n4146), .Z(n4151) );
  NAND U8840 ( .A(n4149), .B(n4148), .Z(n4150) );
  AND U8841 ( .A(n4151), .B(n4150), .Z(n8435) );
  XNOR U8842 ( .A(n8436), .B(n8435), .Z(n8001) );
  XOR U8843 ( .A(n8002), .B(n8001), .Z(n8004) );
  XOR U8844 ( .A(n8003), .B(n8004), .Z(n6253) );
  NANDN U8845 ( .A(n4153), .B(n4152), .Z(n4157) );
  NAND U8846 ( .A(n4155), .B(n4154), .Z(n4156) );
  NAND U8847 ( .A(n4157), .B(n4156), .Z(n6252) );
  XOR U8848 ( .A(n6253), .B(n6252), .Z(n6255) );
  XNOR U8849 ( .A(n6254), .B(n6255), .Z(n7661) );
  NAND U8850 ( .A(n4159), .B(n4158), .Z(n4163) );
  NANDN U8851 ( .A(n4161), .B(n4160), .Z(n4162) );
  NAND U8852 ( .A(n4163), .B(n4162), .Z(n7660) );
  XOR U8853 ( .A(n7661), .B(n7660), .Z(n7662) );
  XNOR U8854 ( .A(n7663), .B(n7662), .Z(n6078) );
  NAND U8855 ( .A(n4165), .B(n4164), .Z(n4169) );
  NAND U8856 ( .A(n4167), .B(n4166), .Z(n4168) );
  NAND U8857 ( .A(n4169), .B(n4168), .Z(n7767) );
  NANDN U8858 ( .A(n4171), .B(n4170), .Z(n4175) );
  NANDN U8859 ( .A(n4173), .B(n4172), .Z(n4174) );
  AND U8860 ( .A(n4175), .B(n4174), .Z(n6267) );
  NANDN U8861 ( .A(n4177), .B(n4176), .Z(n4181) );
  NAND U8862 ( .A(n4179), .B(n4178), .Z(n4180) );
  AND U8863 ( .A(n4181), .B(n4180), .Z(n8067) );
  NANDN U8864 ( .A(n4183), .B(n4182), .Z(n4187) );
  NAND U8865 ( .A(n4185), .B(n4184), .Z(n4186) );
  NAND U8866 ( .A(n4187), .B(n4186), .Z(n8068) );
  XNOR U8867 ( .A(n8067), .B(n8068), .Z(n8070) );
  NANDN U8868 ( .A(n4189), .B(n4188), .Z(n4193) );
  NAND U8869 ( .A(n4191), .B(n4190), .Z(n4192) );
  AND U8870 ( .A(n4193), .B(n4192), .Z(n8069) );
  XOR U8871 ( .A(n8070), .B(n8069), .Z(n7949) );
  NANDN U8872 ( .A(n4195), .B(n4194), .Z(n4199) );
  NAND U8873 ( .A(n4197), .B(n4196), .Z(n4198) );
  AND U8874 ( .A(n4199), .B(n4198), .Z(n8668) );
  NANDN U8875 ( .A(n4201), .B(n4200), .Z(n4205) );
  NAND U8876 ( .A(n4203), .B(n4202), .Z(n4204) );
  AND U8877 ( .A(n4205), .B(n4204), .Z(n8667) );
  XOR U8878 ( .A(n8668), .B(n8667), .Z(n8670) );
  NANDN U8879 ( .A(n4207), .B(n4206), .Z(n4211) );
  NAND U8880 ( .A(n4209), .B(n4208), .Z(n4210) );
  AND U8881 ( .A(n4211), .B(n4210), .Z(n8669) );
  XOR U8882 ( .A(n8670), .B(n8669), .Z(n7948) );
  NANDN U8883 ( .A(n4213), .B(n4212), .Z(n4217) );
  NAND U8884 ( .A(n4215), .B(n4214), .Z(n4216) );
  AND U8885 ( .A(n4217), .B(n4216), .Z(n8271) );
  NANDN U8886 ( .A(n4219), .B(n4218), .Z(n4223) );
  NAND U8887 ( .A(n4221), .B(n4220), .Z(n4222) );
  NAND U8888 ( .A(n4223), .B(n4222), .Z(n8272) );
  XNOR U8889 ( .A(n8271), .B(n8272), .Z(n8274) );
  NANDN U8890 ( .A(n4225), .B(n4224), .Z(n4229) );
  NAND U8891 ( .A(n4227), .B(n4226), .Z(n4228) );
  AND U8892 ( .A(n4229), .B(n4228), .Z(n8273) );
  XNOR U8893 ( .A(n8274), .B(n8273), .Z(n7947) );
  XOR U8894 ( .A(n7948), .B(n7947), .Z(n7950) );
  XOR U8895 ( .A(n7949), .B(n7950), .Z(n6265) );
  NANDN U8896 ( .A(n4231), .B(n4230), .Z(n4235) );
  NANDN U8897 ( .A(n4233), .B(n4232), .Z(n4234) );
  NAND U8898 ( .A(n4235), .B(n4234), .Z(n6264) );
  XNOR U8899 ( .A(n6265), .B(n6264), .Z(n6266) );
  XNOR U8900 ( .A(n6267), .B(n6266), .Z(n7764) );
  NAND U8901 ( .A(n4237), .B(n4236), .Z(n4241) );
  NAND U8902 ( .A(n4239), .B(n4238), .Z(n4240) );
  AND U8903 ( .A(n4241), .B(n4240), .Z(n7765) );
  XOR U8904 ( .A(n7764), .B(n7765), .Z(n7766) );
  XOR U8905 ( .A(n7767), .B(n7766), .Z(n6079) );
  XOR U8906 ( .A(n6078), .B(n6079), .Z(n6080) );
  XNOR U8907 ( .A(n6081), .B(n6080), .Z(n7253) );
  NANDN U8908 ( .A(n4243), .B(n4242), .Z(n4247) );
  NAND U8909 ( .A(n4245), .B(n4244), .Z(n4246) );
  AND U8910 ( .A(n4247), .B(n4246), .Z(n6248) );
  NANDN U8911 ( .A(n4249), .B(n4248), .Z(n4253) );
  NAND U8912 ( .A(n4251), .B(n4250), .Z(n4252) );
  AND U8913 ( .A(n4253), .B(n4252), .Z(n6624) );
  NANDN U8914 ( .A(n4255), .B(n4254), .Z(n4259) );
  NAND U8915 ( .A(n4257), .B(n4256), .Z(n4258) );
  NAND U8916 ( .A(n4259), .B(n4258), .Z(n6625) );
  XNOR U8917 ( .A(n6624), .B(n6625), .Z(n6627) );
  NANDN U8918 ( .A(n4261), .B(n4260), .Z(n4265) );
  NAND U8919 ( .A(n4263), .B(n4262), .Z(n4264) );
  AND U8920 ( .A(n4265), .B(n4264), .Z(n6626) );
  XOR U8921 ( .A(n6627), .B(n6626), .Z(n7967) );
  NANDN U8922 ( .A(n4267), .B(n4266), .Z(n4271) );
  NAND U8923 ( .A(n4269), .B(n4268), .Z(n4270) );
  AND U8924 ( .A(n4271), .B(n4270), .Z(n8793) );
  NANDN U8925 ( .A(n4273), .B(n4272), .Z(n4277) );
  NAND U8926 ( .A(n4275), .B(n4274), .Z(n4276) );
  NAND U8927 ( .A(n4277), .B(n4276), .Z(n8794) );
  XNOR U8928 ( .A(n8793), .B(n8794), .Z(n8796) );
  NANDN U8929 ( .A(n4279), .B(n4278), .Z(n4283) );
  NAND U8930 ( .A(n4281), .B(n4280), .Z(n4282) );
  AND U8931 ( .A(n4283), .B(n4282), .Z(n8795) );
  XOR U8932 ( .A(n8796), .B(n8795), .Z(n7966) );
  NANDN U8933 ( .A(n4285), .B(n4284), .Z(n4289) );
  NAND U8934 ( .A(n4287), .B(n4286), .Z(n4288) );
  AND U8935 ( .A(n4289), .B(n4288), .Z(n8457) );
  NANDN U8936 ( .A(n4291), .B(n4290), .Z(n4295) );
  NAND U8937 ( .A(n4293), .B(n4292), .Z(n4294) );
  NAND U8938 ( .A(n4295), .B(n4294), .Z(n8458) );
  XNOR U8939 ( .A(n8457), .B(n8458), .Z(n8460) );
  NANDN U8940 ( .A(n4297), .B(n4296), .Z(n4301) );
  NAND U8941 ( .A(n4299), .B(n4298), .Z(n4300) );
  AND U8942 ( .A(n4301), .B(n4300), .Z(n8459) );
  XNOR U8943 ( .A(n8460), .B(n8459), .Z(n7965) );
  XOR U8944 ( .A(n7966), .B(n7965), .Z(n7968) );
  XOR U8945 ( .A(n7967), .B(n7968), .Z(n6247) );
  NANDN U8946 ( .A(n4303), .B(n4302), .Z(n4307) );
  NANDN U8947 ( .A(n4305), .B(n4304), .Z(n4306) );
  NAND U8948 ( .A(n4307), .B(n4306), .Z(n6246) );
  XOR U8949 ( .A(n6247), .B(n6246), .Z(n6249) );
  XOR U8950 ( .A(n6248), .B(n6249), .Z(n7116) );
  NANDN U8951 ( .A(n4309), .B(n4308), .Z(n4313) );
  NANDN U8952 ( .A(n4311), .B(n4310), .Z(n4312) );
  AND U8953 ( .A(n4313), .B(n4312), .Z(n6272) );
  NANDN U8954 ( .A(n4315), .B(n4314), .Z(n4319) );
  NAND U8955 ( .A(n4317), .B(n4316), .Z(n4318) );
  AND U8956 ( .A(n4319), .B(n4318), .Z(n8715) );
  NANDN U8957 ( .A(n4321), .B(n4320), .Z(n4325) );
  NAND U8958 ( .A(n4323), .B(n4322), .Z(n4324) );
  NAND U8959 ( .A(n4325), .B(n4324), .Z(n8716) );
  XNOR U8960 ( .A(n8715), .B(n8716), .Z(n8718) );
  NANDN U8961 ( .A(n4327), .B(n4326), .Z(n4331) );
  NAND U8962 ( .A(n4329), .B(n4328), .Z(n4330) );
  AND U8963 ( .A(n4331), .B(n4330), .Z(n8717) );
  XOR U8964 ( .A(n8718), .B(n8717), .Z(n7961) );
  NANDN U8965 ( .A(n4333), .B(n4332), .Z(n4337) );
  NAND U8966 ( .A(n4335), .B(n4334), .Z(n4336) );
  AND U8967 ( .A(n4337), .B(n4336), .Z(n8691) );
  NANDN U8968 ( .A(n4339), .B(n4338), .Z(n4343) );
  NAND U8969 ( .A(n4341), .B(n4340), .Z(n4342) );
  NAND U8970 ( .A(n4343), .B(n4342), .Z(n8692) );
  XNOR U8971 ( .A(n8691), .B(n8692), .Z(n8694) );
  NANDN U8972 ( .A(n4345), .B(n4344), .Z(n4349) );
  NAND U8973 ( .A(n4347), .B(n4346), .Z(n4348) );
  AND U8974 ( .A(n4349), .B(n4348), .Z(n8693) );
  XOR U8975 ( .A(n8694), .B(n8693), .Z(n7960) );
  NANDN U8976 ( .A(n4351), .B(n4350), .Z(n4355) );
  NAND U8977 ( .A(n4353), .B(n4352), .Z(n4354) );
  AND U8978 ( .A(n4355), .B(n4354), .Z(n8805) );
  NANDN U8979 ( .A(n4357), .B(n4356), .Z(n4361) );
  NAND U8980 ( .A(n4359), .B(n4358), .Z(n4360) );
  NAND U8981 ( .A(n4361), .B(n4360), .Z(n8806) );
  XNOR U8982 ( .A(n8805), .B(n8806), .Z(n8808) );
  NANDN U8983 ( .A(n4363), .B(n4362), .Z(n4367) );
  NAND U8984 ( .A(n4365), .B(n4364), .Z(n4366) );
  AND U8985 ( .A(n4367), .B(n4366), .Z(n8807) );
  XNOR U8986 ( .A(n8808), .B(n8807), .Z(n7959) );
  XOR U8987 ( .A(n7960), .B(n7959), .Z(n7962) );
  XOR U8988 ( .A(n7961), .B(n7962), .Z(n6271) );
  NANDN U8989 ( .A(n4369), .B(n4368), .Z(n4373) );
  NAND U8990 ( .A(n4371), .B(n4370), .Z(n4372) );
  NAND U8991 ( .A(n4373), .B(n4372), .Z(n6270) );
  XOR U8992 ( .A(n6271), .B(n6270), .Z(n6273) );
  XOR U8993 ( .A(n6272), .B(n6273), .Z(n7115) );
  NANDN U8994 ( .A(n4375), .B(n4374), .Z(n4379) );
  NAND U8995 ( .A(n4377), .B(n4376), .Z(n4378) );
  AND U8996 ( .A(n4379), .B(n4378), .Z(n6320) );
  NANDN U8997 ( .A(n4381), .B(n4380), .Z(n4385) );
  NAND U8998 ( .A(n4383), .B(n4382), .Z(n4384) );
  AND U8999 ( .A(n4385), .B(n4384), .Z(n8313) );
  NANDN U9000 ( .A(n4387), .B(n4386), .Z(n4391) );
  NAND U9001 ( .A(n4389), .B(n4388), .Z(n4390) );
  NAND U9002 ( .A(n4391), .B(n4390), .Z(n8314) );
  XNOR U9003 ( .A(n8313), .B(n8314), .Z(n8316) );
  NANDN U9004 ( .A(n4393), .B(n4392), .Z(n4397) );
  NAND U9005 ( .A(n4395), .B(n4394), .Z(n4396) );
  AND U9006 ( .A(n4397), .B(n4396), .Z(n8315) );
  XOR U9007 ( .A(n8316), .B(n8315), .Z(n7014) );
  NANDN U9008 ( .A(n4399), .B(n4398), .Z(n4403) );
  NAND U9009 ( .A(n4401), .B(n4400), .Z(n4402) );
  AND U9010 ( .A(n4403), .B(n4402), .Z(n8295) );
  NANDN U9011 ( .A(n4405), .B(n4404), .Z(n4409) );
  NAND U9012 ( .A(n4407), .B(n4406), .Z(n4408) );
  NAND U9013 ( .A(n4409), .B(n4408), .Z(n8296) );
  XNOR U9014 ( .A(n8295), .B(n8296), .Z(n8298) );
  NANDN U9015 ( .A(n4411), .B(n4410), .Z(n4415) );
  NAND U9016 ( .A(n4413), .B(n4412), .Z(n4414) );
  AND U9017 ( .A(n4415), .B(n4414), .Z(n8297) );
  XOR U9018 ( .A(n8298), .B(n8297), .Z(n7013) );
  NANDN U9019 ( .A(n4417), .B(n4416), .Z(n4421) );
  NAND U9020 ( .A(n4419), .B(n4418), .Z(n4420) );
  AND U9021 ( .A(n4421), .B(n4420), .Z(n8235) );
  NANDN U9022 ( .A(n4423), .B(n4422), .Z(n4427) );
  NAND U9023 ( .A(n4425), .B(n4424), .Z(n4426) );
  NAND U9024 ( .A(n4427), .B(n4426), .Z(n8236) );
  XNOR U9025 ( .A(n8235), .B(n8236), .Z(n8238) );
  NANDN U9026 ( .A(n4429), .B(n4428), .Z(n4433) );
  NAND U9027 ( .A(n4431), .B(n4430), .Z(n4432) );
  AND U9028 ( .A(n4433), .B(n4432), .Z(n8237) );
  XNOR U9029 ( .A(n8238), .B(n8237), .Z(n7012) );
  XOR U9030 ( .A(n7013), .B(n7012), .Z(n7015) );
  XOR U9031 ( .A(n7014), .B(n7015), .Z(n6319) );
  NANDN U9032 ( .A(n4435), .B(n4434), .Z(n4439) );
  NANDN U9033 ( .A(n4437), .B(n4436), .Z(n4438) );
  NAND U9034 ( .A(n4439), .B(n4438), .Z(n6318) );
  XOR U9035 ( .A(n6319), .B(n6318), .Z(n6321) );
  XNOR U9036 ( .A(n6320), .B(n6321), .Z(n7114) );
  XOR U9037 ( .A(n7115), .B(n7114), .Z(n7117) );
  XOR U9038 ( .A(n7116), .B(n7117), .Z(n6955) );
  NAND U9039 ( .A(n4441), .B(n4440), .Z(n4445) );
  NAND U9040 ( .A(n4443), .B(n4442), .Z(n4444) );
  NAND U9041 ( .A(n4445), .B(n4444), .Z(n6967) );
  NAND U9042 ( .A(n4447), .B(n4446), .Z(n4451) );
  NANDN U9043 ( .A(n4449), .B(n4448), .Z(n4450) );
  NAND U9044 ( .A(n4451), .B(n4450), .Z(n6965) );
  NAND U9045 ( .A(n4453), .B(n4452), .Z(n4457) );
  NAND U9046 ( .A(n4455), .B(n4454), .Z(n4456) );
  AND U9047 ( .A(n4457), .B(n4456), .Z(n6277) );
  NANDN U9048 ( .A(n4459), .B(n4458), .Z(n4463) );
  NANDN U9049 ( .A(n4461), .B(n4460), .Z(n4462) );
  AND U9050 ( .A(n4463), .B(n4462), .Z(n9021) );
  NANDN U9051 ( .A(n4465), .B(n4464), .Z(n4469) );
  NANDN U9052 ( .A(n4467), .B(n4466), .Z(n4468) );
  NAND U9053 ( .A(n4469), .B(n4468), .Z(n9022) );
  XNOR U9054 ( .A(n9021), .B(n9022), .Z(n9024) );
  NANDN U9055 ( .A(n4471), .B(n4470), .Z(n4475) );
  NANDN U9056 ( .A(n4473), .B(n4472), .Z(n4474) );
  AND U9057 ( .A(n4475), .B(n4474), .Z(n9023) );
  XOR U9058 ( .A(n9024), .B(n9023), .Z(n6990) );
  NANDN U9059 ( .A(n4477), .B(n4476), .Z(n4481) );
  NAND U9060 ( .A(n4479), .B(n4478), .Z(n4480) );
  AND U9061 ( .A(n4481), .B(n4480), .Z(n6642) );
  NANDN U9062 ( .A(n4483), .B(n4482), .Z(n4487) );
  NAND U9063 ( .A(n4485), .B(n4484), .Z(n4486) );
  NAND U9064 ( .A(n4487), .B(n4486), .Z(n6643) );
  XNOR U9065 ( .A(n6642), .B(n6643), .Z(n6645) );
  NANDN U9066 ( .A(n4489), .B(n4488), .Z(n4493) );
  NAND U9067 ( .A(n4491), .B(n4490), .Z(n4492) );
  AND U9068 ( .A(n4493), .B(n4492), .Z(n6644) );
  XOR U9069 ( .A(n6645), .B(n6644), .Z(n6989) );
  NANDN U9070 ( .A(n4495), .B(n4494), .Z(n4499) );
  NAND U9071 ( .A(n4497), .B(n4496), .Z(n4498) );
  AND U9072 ( .A(n4499), .B(n4498), .Z(n6462) );
  NANDN U9073 ( .A(n4501), .B(n4500), .Z(n4505) );
  NAND U9074 ( .A(n4503), .B(n4502), .Z(n4504) );
  NAND U9075 ( .A(n4505), .B(n4504), .Z(n6463) );
  XNOR U9076 ( .A(n6462), .B(n6463), .Z(n6465) );
  NANDN U9077 ( .A(n4507), .B(n4506), .Z(n4511) );
  NAND U9078 ( .A(n4509), .B(n4508), .Z(n4510) );
  AND U9079 ( .A(n4511), .B(n4510), .Z(n6464) );
  XNOR U9080 ( .A(n6465), .B(n6464), .Z(n6988) );
  XOR U9081 ( .A(n6989), .B(n6988), .Z(n6991) );
  XOR U9082 ( .A(n6990), .B(n6991), .Z(n6276) );
  XOR U9083 ( .A(n6277), .B(n6276), .Z(n6279) );
  NAND U9084 ( .A(n4513), .B(n4512), .Z(n4517) );
  NAND U9085 ( .A(n4515), .B(n4514), .Z(n4516) );
  AND U9086 ( .A(n4517), .B(n4516), .Z(n6278) );
  XOR U9087 ( .A(n6279), .B(n6278), .Z(n6964) );
  XOR U9088 ( .A(n6965), .B(n6964), .Z(n6966) );
  XNOR U9089 ( .A(n6967), .B(n6966), .Z(n6953) );
  NAND U9090 ( .A(n4519), .B(n4518), .Z(n4523) );
  NANDN U9091 ( .A(n4521), .B(n4520), .Z(n4522) );
  AND U9092 ( .A(n4523), .B(n4522), .Z(n8022) );
  NANDN U9093 ( .A(n4525), .B(n4524), .Z(n4529) );
  NAND U9094 ( .A(n4527), .B(n4526), .Z(n4528) );
  AND U9095 ( .A(n4529), .B(n4528), .Z(n6260) );
  NANDN U9096 ( .A(n4531), .B(n4530), .Z(n4535) );
  NAND U9097 ( .A(n4533), .B(n4532), .Z(n4534) );
  AND U9098 ( .A(n4535), .B(n4534), .Z(n8410) );
  NANDN U9099 ( .A(n4537), .B(n4536), .Z(n4541) );
  NAND U9100 ( .A(n4539), .B(n4538), .Z(n4540) );
  AND U9101 ( .A(n4541), .B(n4540), .Z(n8409) );
  XOR U9102 ( .A(n8410), .B(n8409), .Z(n8412) );
  NANDN U9103 ( .A(n4543), .B(n4542), .Z(n4547) );
  NAND U9104 ( .A(n4545), .B(n4544), .Z(n4546) );
  AND U9105 ( .A(n4547), .B(n4546), .Z(n8411) );
  XOR U9106 ( .A(n8412), .B(n8411), .Z(n7943) );
  NANDN U9107 ( .A(n4549), .B(n4548), .Z(n4553) );
  NAND U9108 ( .A(n4551), .B(n4550), .Z(n4552) );
  AND U9109 ( .A(n4553), .B(n4552), .Z(n6582) );
  NANDN U9110 ( .A(n4555), .B(n4554), .Z(n4559) );
  NAND U9111 ( .A(n4557), .B(n4556), .Z(n4558) );
  NAND U9112 ( .A(n4559), .B(n4558), .Z(n6583) );
  XNOR U9113 ( .A(n6582), .B(n6583), .Z(n6585) );
  NANDN U9114 ( .A(n4561), .B(n4560), .Z(n4565) );
  NAND U9115 ( .A(n4563), .B(n4562), .Z(n4564) );
  AND U9116 ( .A(n4565), .B(n4564), .Z(n6584) );
  XOR U9117 ( .A(n6585), .B(n6584), .Z(n7942) );
  NANDN U9118 ( .A(n4567), .B(n4566), .Z(n4571) );
  NAND U9119 ( .A(n4569), .B(n4568), .Z(n4570) );
  AND U9120 ( .A(n4571), .B(n4570), .Z(n8505) );
  NANDN U9121 ( .A(n4573), .B(n4572), .Z(n4577) );
  NAND U9122 ( .A(n4575), .B(n4574), .Z(n4576) );
  NAND U9123 ( .A(n4577), .B(n4576), .Z(n8506) );
  XNOR U9124 ( .A(n8505), .B(n8506), .Z(n8508) );
  NANDN U9125 ( .A(n4579), .B(n4578), .Z(n4583) );
  NAND U9126 ( .A(n4581), .B(n4580), .Z(n4582) );
  AND U9127 ( .A(n4583), .B(n4582), .Z(n8507) );
  XNOR U9128 ( .A(n8508), .B(n8507), .Z(n7941) );
  XOR U9129 ( .A(n7942), .B(n7941), .Z(n7944) );
  XOR U9130 ( .A(n7943), .B(n7944), .Z(n6259) );
  NANDN U9131 ( .A(n4585), .B(n4584), .Z(n4589) );
  NANDN U9132 ( .A(n4587), .B(n4586), .Z(n4588) );
  NAND U9133 ( .A(n4589), .B(n4588), .Z(n6258) );
  XOR U9134 ( .A(n6259), .B(n6258), .Z(n6261) );
  XNOR U9135 ( .A(n6260), .B(n6261), .Z(n8020) );
  NAND U9136 ( .A(n4591), .B(n4590), .Z(n4595) );
  NAND U9137 ( .A(n4593), .B(n4592), .Z(n4594) );
  AND U9138 ( .A(n4595), .B(n4594), .Z(n8019) );
  XOR U9139 ( .A(n8020), .B(n8019), .Z(n8021) );
  XOR U9140 ( .A(n8022), .B(n8021), .Z(n6952) );
  XOR U9141 ( .A(n6953), .B(n6952), .Z(n6954) );
  XOR U9142 ( .A(n6955), .B(n6954), .Z(n7252) );
  XOR U9143 ( .A(n7253), .B(n7252), .Z(n7254) );
  XNOR U9144 ( .A(n7255), .B(n7254), .Z(n7243) );
  NAND U9145 ( .A(n4597), .B(n4596), .Z(n4601) );
  NAND U9146 ( .A(n4599), .B(n4598), .Z(n4600) );
  AND U9147 ( .A(n4601), .B(n4600), .Z(n7241) );
  NANDN U9148 ( .A(n4603), .B(n4602), .Z(n4607) );
  NANDN U9149 ( .A(n4605), .B(n4604), .Z(n4606) );
  AND U9150 ( .A(n4607), .B(n4606), .Z(n7697) );
  NANDN U9151 ( .A(n4609), .B(n4608), .Z(n4613) );
  NAND U9152 ( .A(n4611), .B(n4610), .Z(n4612) );
  AND U9153 ( .A(n4613), .B(n4612), .Z(n7516) );
  NANDN U9154 ( .A(n4615), .B(n4614), .Z(n4619) );
  NAND U9155 ( .A(n4617), .B(n4616), .Z(n4618) );
  NAND U9156 ( .A(n4619), .B(n4618), .Z(n7517) );
  XNOR U9157 ( .A(n7516), .B(n7517), .Z(n7519) );
  NANDN U9158 ( .A(n4621), .B(n4620), .Z(n4625) );
  NAND U9159 ( .A(n4623), .B(n4622), .Z(n4624) );
  AND U9160 ( .A(n4625), .B(n4624), .Z(n7518) );
  XOR U9161 ( .A(n7519), .B(n7518), .Z(n7695) );
  NANDN U9162 ( .A(n4627), .B(n4626), .Z(n4631) );
  NANDN U9163 ( .A(n4629), .B(n4628), .Z(n4630) );
  AND U9164 ( .A(n4631), .B(n4630), .Z(n7694) );
  XNOR U9165 ( .A(n7695), .B(n7694), .Z(n7696) );
  XOR U9166 ( .A(n7697), .B(n7696), .Z(n6105) );
  NANDN U9167 ( .A(n4633), .B(n4632), .Z(n4637) );
  NANDN U9168 ( .A(n4635), .B(n4634), .Z(n4636) );
  AND U9169 ( .A(n4637), .B(n4636), .Z(n7363) );
  NAND U9170 ( .A(n4639), .B(n4638), .Z(n4643) );
  NAND U9171 ( .A(n4641), .B(n4640), .Z(n4642) );
  AND U9172 ( .A(n4643), .B(n4642), .Z(n6864) );
  NAND U9173 ( .A(n4645), .B(n4644), .Z(n4649) );
  NAND U9174 ( .A(n4647), .B(n4646), .Z(n4648) );
  NAND U9175 ( .A(n4649), .B(n4648), .Z(n6865) );
  XNOR U9176 ( .A(n6864), .B(n6865), .Z(n6867) );
  NANDN U9177 ( .A(n4651), .B(n4650), .Z(n4655) );
  NAND U9178 ( .A(n4653), .B(n4652), .Z(n4654) );
  AND U9179 ( .A(n4655), .B(n4654), .Z(n6866) );
  XOR U9180 ( .A(n6867), .B(n6866), .Z(n7361) );
  NANDN U9181 ( .A(n4657), .B(n4656), .Z(n4661) );
  NANDN U9182 ( .A(n4659), .B(n4658), .Z(n4660) );
  AND U9183 ( .A(n4661), .B(n4660), .Z(n7360) );
  XNOR U9184 ( .A(n7361), .B(n7360), .Z(n7362) );
  XOR U9185 ( .A(n7363), .B(n7362), .Z(n6103) );
  NAND U9186 ( .A(n4663), .B(n4662), .Z(n4667) );
  NAND U9187 ( .A(n4665), .B(n4664), .Z(n4666) );
  AND U9188 ( .A(n4667), .B(n4666), .Z(n6525) );
  NANDN U9189 ( .A(n4669), .B(n4668), .Z(n4673) );
  NAND U9190 ( .A(n4671), .B(n4670), .Z(n4672) );
  AND U9191 ( .A(n4673), .B(n4672), .Z(n8553) );
  NANDN U9192 ( .A(n4675), .B(n4674), .Z(n4679) );
  NAND U9193 ( .A(n4677), .B(n4676), .Z(n4678) );
  NAND U9194 ( .A(n4679), .B(n4678), .Z(n8554) );
  XNOR U9195 ( .A(n8553), .B(n8554), .Z(n8556) );
  NANDN U9196 ( .A(n4681), .B(n4680), .Z(n4685) );
  NAND U9197 ( .A(n4683), .B(n4682), .Z(n4684) );
  AND U9198 ( .A(n4685), .B(n4684), .Z(n8555) );
  XOR U9199 ( .A(n8556), .B(n8555), .Z(n6523) );
  NAND U9200 ( .A(n4687), .B(n4686), .Z(n4691) );
  NAND U9201 ( .A(n4689), .B(n4688), .Z(n4690) );
  AND U9202 ( .A(n4691), .B(n4690), .Z(n6522) );
  XNOR U9203 ( .A(n6523), .B(n6522), .Z(n6524) );
  XNOR U9204 ( .A(n6525), .B(n6524), .Z(n6102) );
  XNOR U9205 ( .A(n6103), .B(n6102), .Z(n6104) );
  XNOR U9206 ( .A(n6105), .B(n6104), .Z(n6567) );
  NANDN U9207 ( .A(n4693), .B(n4692), .Z(n4697) );
  NANDN U9208 ( .A(n4695), .B(n4694), .Z(n4696) );
  AND U9209 ( .A(n4697), .B(n4696), .Z(n6948) );
  NANDN U9210 ( .A(n4699), .B(n4698), .Z(n4703) );
  NANDN U9211 ( .A(n4701), .B(n4700), .Z(n4702) );
  AND U9212 ( .A(n4703), .B(n4702), .Z(n6946) );
  NANDN U9213 ( .A(n4705), .B(n4704), .Z(n4709) );
  NANDN U9214 ( .A(n4707), .B(n4706), .Z(n4708) );
  NAND U9215 ( .A(n4709), .B(n4708), .Z(n6947) );
  XOR U9216 ( .A(n6946), .B(n6947), .Z(n6949) );
  XNOR U9217 ( .A(n6948), .B(n6949), .Z(n6336) );
  NANDN U9218 ( .A(n4711), .B(n4710), .Z(n4715) );
  NAND U9219 ( .A(n4713), .B(n4712), .Z(n4714) );
  AND U9220 ( .A(n4715), .B(n4714), .Z(n8499) );
  NANDN U9221 ( .A(n4717), .B(n4716), .Z(n4721) );
  NAND U9222 ( .A(n4719), .B(n4718), .Z(n4720) );
  NAND U9223 ( .A(n4721), .B(n4720), .Z(n8500) );
  XNOR U9224 ( .A(n8499), .B(n8500), .Z(n8502) );
  NAND U9225 ( .A(n4723), .B(n4722), .Z(n4727) );
  NAND U9226 ( .A(n4725), .B(n4724), .Z(n4726) );
  AND U9227 ( .A(n4727), .B(n4726), .Z(n8501) );
  XOR U9228 ( .A(n8502), .B(n8501), .Z(n7417) );
  NANDN U9229 ( .A(n4729), .B(n4728), .Z(n4733) );
  NAND U9230 ( .A(n4731), .B(n4730), .Z(n4732) );
  AND U9231 ( .A(n4733), .B(n4732), .Z(n8265) );
  NANDN U9232 ( .A(n4735), .B(n4734), .Z(n4739) );
  NAND U9233 ( .A(n4737), .B(n4736), .Z(n4738) );
  NAND U9234 ( .A(n4739), .B(n4738), .Z(n8266) );
  XNOR U9235 ( .A(n8265), .B(n8266), .Z(n8268) );
  NANDN U9236 ( .A(n4741), .B(n4740), .Z(n4745) );
  NAND U9237 ( .A(n4743), .B(n4742), .Z(n4744) );
  AND U9238 ( .A(n4745), .B(n4744), .Z(n8267) );
  XOR U9239 ( .A(n8268), .B(n8267), .Z(n7415) );
  NANDN U9240 ( .A(n4747), .B(n4746), .Z(n4751) );
  NANDN U9241 ( .A(n4749), .B(n4748), .Z(n4750) );
  AND U9242 ( .A(n4751), .B(n4750), .Z(n7414) );
  XNOR U9243 ( .A(n7415), .B(n7414), .Z(n7416) );
  XOR U9244 ( .A(n7417), .B(n7416), .Z(n6337) );
  XNOR U9245 ( .A(n6336), .B(n6337), .Z(n6339) );
  NANDN U9246 ( .A(n4753), .B(n4752), .Z(n4757) );
  NANDN U9247 ( .A(n4755), .B(n4754), .Z(n4756) );
  AND U9248 ( .A(n4757), .B(n4756), .Z(n6936) );
  NANDN U9249 ( .A(n4759), .B(n4758), .Z(n4763) );
  NANDN U9250 ( .A(n4761), .B(n4760), .Z(n4762) );
  AND U9251 ( .A(n4763), .B(n4762), .Z(n6934) );
  NANDN U9252 ( .A(n4765), .B(n4764), .Z(n4769) );
  NANDN U9253 ( .A(n4767), .B(n4766), .Z(n4768) );
  NAND U9254 ( .A(n4769), .B(n4768), .Z(n6935) );
  XOR U9255 ( .A(n6934), .B(n6935), .Z(n6937) );
  XNOR U9256 ( .A(n6936), .B(n6937), .Z(n6338) );
  XNOR U9257 ( .A(n6339), .B(n6338), .Z(n6565) );
  NANDN U9258 ( .A(n4771), .B(n4770), .Z(n4775) );
  NANDN U9259 ( .A(n4773), .B(n4772), .Z(n4774) );
  AND U9260 ( .A(n4775), .B(n4774), .Z(n8514) );
  NANDN U9261 ( .A(n4777), .B(n4776), .Z(n4781) );
  NAND U9262 ( .A(n4779), .B(n4778), .Z(n4780) );
  AND U9263 ( .A(n4781), .B(n4780), .Z(n6834) );
  NANDN U9264 ( .A(n4783), .B(n4782), .Z(n4787) );
  NAND U9265 ( .A(n4785), .B(n4784), .Z(n4786) );
  NAND U9266 ( .A(n4787), .B(n4786), .Z(n6835) );
  XNOR U9267 ( .A(n6834), .B(n6835), .Z(n6837) );
  NANDN U9268 ( .A(n4789), .B(n4788), .Z(n4793) );
  NAND U9269 ( .A(n4791), .B(n4790), .Z(n4792) );
  AND U9270 ( .A(n4793), .B(n4792), .Z(n6836) );
  XOR U9271 ( .A(n6837), .B(n6836), .Z(n7314) );
  NANDN U9272 ( .A(n4795), .B(n4794), .Z(n4799) );
  NANDN U9273 ( .A(n4797), .B(n4796), .Z(n4798) );
  AND U9274 ( .A(n4799), .B(n4798), .Z(n7312) );
  NANDN U9275 ( .A(n4801), .B(n4800), .Z(n4805) );
  NANDN U9276 ( .A(n4803), .B(n4802), .Z(n4804) );
  NAND U9277 ( .A(n4805), .B(n4804), .Z(n7313) );
  XOR U9278 ( .A(n7312), .B(n7313), .Z(n7315) );
  XOR U9279 ( .A(n7314), .B(n7315), .Z(n8512) );
  NANDN U9280 ( .A(n4807), .B(n4806), .Z(n4811) );
  NANDN U9281 ( .A(n4809), .B(n4808), .Z(n4810) );
  NAND U9282 ( .A(n4811), .B(n4810), .Z(n8511) );
  XNOR U9283 ( .A(n8512), .B(n8511), .Z(n8513) );
  XNOR U9284 ( .A(n8514), .B(n8513), .Z(n6564) );
  XOR U9285 ( .A(n6565), .B(n6564), .Z(n6566) );
  XNOR U9286 ( .A(n6567), .B(n6566), .Z(n6959) );
  NAND U9287 ( .A(n4813), .B(n4812), .Z(n4817) );
  NAND U9288 ( .A(n4815), .B(n4814), .Z(n4816) );
  AND U9289 ( .A(n4817), .B(n4816), .Z(n6958) );
  XOR U9290 ( .A(n6959), .B(n6958), .Z(n6961) );
  NAND U9291 ( .A(n4819), .B(n4818), .Z(n4823) );
  NAND U9292 ( .A(n4821), .B(n4820), .Z(n4822) );
  NAND U9293 ( .A(n4823), .B(n4822), .Z(n6891) );
  NAND U9294 ( .A(n4825), .B(n4824), .Z(n4829) );
  NAND U9295 ( .A(n4827), .B(n4826), .Z(n4828) );
  AND U9296 ( .A(n4829), .B(n4828), .Z(n6888) );
  NAND U9297 ( .A(n4831), .B(n4830), .Z(n4835) );
  NAND U9298 ( .A(n4833), .B(n4832), .Z(n4834) );
  AND U9299 ( .A(n4835), .B(n4834), .Z(n6889) );
  XOR U9300 ( .A(n6888), .B(n6889), .Z(n6890) );
  XOR U9301 ( .A(n6891), .B(n6890), .Z(n6960) );
  XNOR U9302 ( .A(n6961), .B(n6960), .Z(n7423) );
  NANDN U9303 ( .A(n4837), .B(n4836), .Z(n4841) );
  NANDN U9304 ( .A(n4839), .B(n4838), .Z(n4840) );
  AND U9305 ( .A(n4841), .B(n4840), .Z(n7955) );
  NANDN U9306 ( .A(n4843), .B(n4842), .Z(n4847) );
  NAND U9307 ( .A(n4845), .B(n4844), .Z(n4846) );
  AND U9308 ( .A(n4847), .B(n4846), .Z(n8727) );
  NANDN U9309 ( .A(n4849), .B(n4848), .Z(n4853) );
  NANDN U9310 ( .A(n4851), .B(n4850), .Z(n4852) );
  NAND U9311 ( .A(n4853), .B(n4852), .Z(n8728) );
  XNOR U9312 ( .A(n8727), .B(n8728), .Z(n8730) );
  NANDN U9313 ( .A(n4855), .B(n4854), .Z(n4859) );
  NAND U9314 ( .A(n4857), .B(n4856), .Z(n4858) );
  AND U9315 ( .A(n4859), .B(n4858), .Z(n8729) );
  XOR U9316 ( .A(n8730), .B(n8729), .Z(n7954) );
  NANDN U9317 ( .A(n4861), .B(n4860), .Z(n4865) );
  NANDN U9318 ( .A(n4863), .B(n4862), .Z(n4864) );
  AND U9319 ( .A(n4865), .B(n4864), .Z(n7953) );
  XOR U9320 ( .A(n7954), .B(n7953), .Z(n7956) );
  XNOR U9321 ( .A(n7955), .B(n7956), .Z(n6498) );
  NANDN U9322 ( .A(n4867), .B(n4866), .Z(n4871) );
  NAND U9323 ( .A(n4869), .B(n4868), .Z(n4870) );
  AND U9324 ( .A(n4871), .B(n4870), .Z(n6654) );
  NANDN U9325 ( .A(n4873), .B(n4872), .Z(n4877) );
  NAND U9326 ( .A(n4875), .B(n4874), .Z(n4876) );
  NAND U9327 ( .A(n4877), .B(n4876), .Z(n6655) );
  XNOR U9328 ( .A(n6654), .B(n6655), .Z(n6657) );
  NANDN U9329 ( .A(n4879), .B(n4878), .Z(n4883) );
  NAND U9330 ( .A(n4881), .B(n4880), .Z(n4882) );
  AND U9331 ( .A(n4883), .B(n4882), .Z(n6656) );
  XOR U9332 ( .A(n6657), .B(n6656), .Z(n7743) );
  NANDN U9333 ( .A(n4885), .B(n4884), .Z(n4889) );
  NANDN U9334 ( .A(n4887), .B(n4886), .Z(n4888) );
  AND U9335 ( .A(n4889), .B(n4888), .Z(n7740) );
  NANDN U9336 ( .A(n4891), .B(n4890), .Z(n4895) );
  NANDN U9337 ( .A(n4893), .B(n4892), .Z(n4894) );
  NAND U9338 ( .A(n4895), .B(n4894), .Z(n7741) );
  XNOR U9339 ( .A(n7740), .B(n7741), .Z(n7742) );
  XOR U9340 ( .A(n7743), .B(n7742), .Z(n6499) );
  XNOR U9341 ( .A(n6498), .B(n6499), .Z(n6500) );
  NANDN U9342 ( .A(n4897), .B(n4896), .Z(n4901) );
  NAND U9343 ( .A(n4899), .B(n4898), .Z(n4900) );
  AND U9344 ( .A(n4901), .B(n4900), .Z(n6823) );
  NANDN U9345 ( .A(n4903), .B(n4902), .Z(n4907) );
  NAND U9346 ( .A(n4905), .B(n4904), .Z(n4906) );
  AND U9347 ( .A(n4907), .B(n4906), .Z(n6822) );
  XOR U9348 ( .A(n6823), .B(n6822), .Z(n6825) );
  NANDN U9349 ( .A(n4909), .B(n4908), .Z(n4913) );
  NAND U9350 ( .A(n4911), .B(n4910), .Z(n4912) );
  AND U9351 ( .A(n4913), .B(n4912), .Z(n6824) );
  XOR U9352 ( .A(n6825), .B(n6824), .Z(n7639) );
  NANDN U9353 ( .A(n4915), .B(n4914), .Z(n4919) );
  NANDN U9354 ( .A(n4917), .B(n4916), .Z(n4918) );
  AND U9355 ( .A(n4919), .B(n4918), .Z(n7789) );
  NANDN U9356 ( .A(n4921), .B(n4920), .Z(n4925) );
  NAND U9357 ( .A(n4923), .B(n4922), .Z(n4924) );
  AND U9358 ( .A(n4925), .B(n4924), .Z(n7788) );
  XOR U9359 ( .A(n7789), .B(n7788), .Z(n7791) );
  NANDN U9360 ( .A(n4927), .B(n4926), .Z(n4931) );
  NAND U9361 ( .A(n4929), .B(n4928), .Z(n4930) );
  AND U9362 ( .A(n4931), .B(n4930), .Z(n7790) );
  XOR U9363 ( .A(n7791), .B(n7790), .Z(n7637) );
  NANDN U9364 ( .A(n4933), .B(n4932), .Z(n4937) );
  NANDN U9365 ( .A(n4935), .B(n4934), .Z(n4936) );
  AND U9366 ( .A(n4937), .B(n4936), .Z(n7636) );
  XNOR U9367 ( .A(n7637), .B(n7636), .Z(n7638) );
  XOR U9368 ( .A(n7639), .B(n7638), .Z(n6501) );
  XNOR U9369 ( .A(n6500), .B(n6501), .Z(n8280) );
  NANDN U9370 ( .A(n4939), .B(n4938), .Z(n4943) );
  NANDN U9371 ( .A(n4941), .B(n4940), .Z(n4942) );
  AND U9372 ( .A(n4943), .B(n4942), .Z(n6230) );
  NANDN U9373 ( .A(n4945), .B(n4944), .Z(n4949) );
  NANDN U9374 ( .A(n4947), .B(n4946), .Z(n4948) );
  AND U9375 ( .A(n4949), .B(n4948), .Z(n6229) );
  NANDN U9376 ( .A(n4951), .B(n4950), .Z(n4955) );
  NAND U9377 ( .A(n4953), .B(n4952), .Z(n4954) );
  NAND U9378 ( .A(n4955), .B(n4954), .Z(n6228) );
  XOR U9379 ( .A(n6229), .B(n6228), .Z(n6231) );
  XOR U9380 ( .A(n6230), .B(n6231), .Z(n8278) );
  NANDN U9381 ( .A(n4957), .B(n4956), .Z(n4961) );
  NANDN U9382 ( .A(n4959), .B(n4958), .Z(n4960) );
  AND U9383 ( .A(n4961), .B(n4960), .Z(n8277) );
  XNOR U9384 ( .A(n8278), .B(n8277), .Z(n8279) );
  XNOR U9385 ( .A(n8280), .B(n8279), .Z(n7045) );
  NANDN U9386 ( .A(n4963), .B(n4962), .Z(n4967) );
  NAND U9387 ( .A(n4965), .B(n4964), .Z(n4966) );
  AND U9388 ( .A(n4967), .B(n4966), .Z(n8482) );
  NANDN U9389 ( .A(n4969), .B(n4968), .Z(n4973) );
  NAND U9390 ( .A(n4971), .B(n4970), .Z(n4972) );
  AND U9391 ( .A(n4973), .B(n4972), .Z(n8481) );
  XOR U9392 ( .A(n8482), .B(n8481), .Z(n8484) );
  NANDN U9393 ( .A(n4975), .B(n4974), .Z(n4979) );
  NAND U9394 ( .A(n4977), .B(n4976), .Z(n4978) );
  AND U9395 ( .A(n4979), .B(n4978), .Z(n8483) );
  XOR U9396 ( .A(n8484), .B(n8483), .Z(n7749) );
  NANDN U9397 ( .A(n4981), .B(n4980), .Z(n4985) );
  NANDN U9398 ( .A(n4983), .B(n4982), .Z(n4984) );
  AND U9399 ( .A(n4985), .B(n4984), .Z(n7746) );
  NANDN U9400 ( .A(n4987), .B(n4986), .Z(n4991) );
  NANDN U9401 ( .A(n4989), .B(n4988), .Z(n4990) );
  NAND U9402 ( .A(n4991), .B(n4990), .Z(n7747) );
  XNOR U9403 ( .A(n7746), .B(n7747), .Z(n7748) );
  XNOR U9404 ( .A(n7749), .B(n7748), .Z(n8595) );
  NANDN U9405 ( .A(n4993), .B(n4992), .Z(n4997) );
  NANDN U9406 ( .A(n4995), .B(n4994), .Z(n4996) );
  AND U9407 ( .A(n4997), .B(n4996), .Z(n8151) );
  NANDN U9408 ( .A(n4999), .B(n4998), .Z(n5003) );
  NANDN U9409 ( .A(n5001), .B(n5000), .Z(n5002) );
  NAND U9410 ( .A(n5003), .B(n5002), .Z(n8152) );
  XNOR U9411 ( .A(n8151), .B(n8152), .Z(n8154) );
  NANDN U9412 ( .A(n5005), .B(n5004), .Z(n5009) );
  NAND U9413 ( .A(n5007), .B(n5006), .Z(n5008) );
  AND U9414 ( .A(n5009), .B(n5008), .Z(n8153) );
  XOR U9415 ( .A(n8154), .B(n8153), .Z(n7225) );
  NANDN U9416 ( .A(n5011), .B(n5010), .Z(n5015) );
  NAND U9417 ( .A(n5013), .B(n5012), .Z(n5014) );
  AND U9418 ( .A(n5015), .B(n5014), .Z(n6882) );
  NANDN U9419 ( .A(n5017), .B(n5016), .Z(n5021) );
  NAND U9420 ( .A(n5019), .B(n5018), .Z(n5020) );
  NAND U9421 ( .A(n5021), .B(n5020), .Z(n6883) );
  XNOR U9422 ( .A(n6882), .B(n6883), .Z(n6885) );
  NANDN U9423 ( .A(n5023), .B(n5022), .Z(n5027) );
  NAND U9424 ( .A(n5025), .B(n5024), .Z(n5026) );
  AND U9425 ( .A(n5027), .B(n5026), .Z(n6884) );
  XOR U9426 ( .A(n6885), .B(n6884), .Z(n7223) );
  NANDN U9427 ( .A(n5029), .B(n5028), .Z(n5033) );
  NANDN U9428 ( .A(n5031), .B(n5030), .Z(n5032) );
  AND U9429 ( .A(n5033), .B(n5032), .Z(n7222) );
  XNOR U9430 ( .A(n7223), .B(n7222), .Z(n7224) );
  XOR U9431 ( .A(n7225), .B(n7224), .Z(n8596) );
  XNOR U9432 ( .A(n8595), .B(n8596), .Z(n8598) );
  NANDN U9433 ( .A(n5035), .B(n5034), .Z(n5039) );
  NAND U9434 ( .A(n5037), .B(n5036), .Z(n5038) );
  AND U9435 ( .A(n5039), .B(n5038), .Z(n8427) );
  NANDN U9436 ( .A(n5041), .B(n5040), .Z(n5045) );
  NAND U9437 ( .A(n5043), .B(n5042), .Z(n5044) );
  NAND U9438 ( .A(n5045), .B(n5044), .Z(n8428) );
  XNOR U9439 ( .A(n8427), .B(n8428), .Z(n8430) );
  NANDN U9440 ( .A(n5047), .B(n5046), .Z(n5051) );
  NAND U9441 ( .A(n5049), .B(n5048), .Z(n5050) );
  AND U9442 ( .A(n5051), .B(n5050), .Z(n8429) );
  XOR U9443 ( .A(n8430), .B(n8429), .Z(n7932) );
  NANDN U9444 ( .A(n5053), .B(n5052), .Z(n5057) );
  NAND U9445 ( .A(n5055), .B(n5054), .Z(n5056) );
  AND U9446 ( .A(n5057), .B(n5056), .Z(n8415) );
  NAND U9447 ( .A(n5059), .B(n5058), .Z(n5063) );
  NAND U9448 ( .A(n5061), .B(n5060), .Z(n5062) );
  NAND U9449 ( .A(n5063), .B(n5062), .Z(n8416) );
  XNOR U9450 ( .A(n8415), .B(n8416), .Z(n8418) );
  NAND U9451 ( .A(n5065), .B(n5064), .Z(n5069) );
  NAND U9452 ( .A(n5067), .B(n5066), .Z(n5068) );
  AND U9453 ( .A(n5069), .B(n5068), .Z(n8417) );
  XOR U9454 ( .A(n8418), .B(n8417), .Z(n7930) );
  NANDN U9455 ( .A(n5071), .B(n5070), .Z(n5075) );
  NANDN U9456 ( .A(n5073), .B(n5072), .Z(n5074) );
  AND U9457 ( .A(n5075), .B(n5074), .Z(n7929) );
  XNOR U9458 ( .A(n7930), .B(n7929), .Z(n7931) );
  XNOR U9459 ( .A(n7932), .B(n7931), .Z(n8597) );
  XOR U9460 ( .A(n8598), .B(n8597), .Z(n6667) );
  NANDN U9461 ( .A(n5077), .B(n5076), .Z(n5081) );
  NANDN U9462 ( .A(n5079), .B(n5078), .Z(n5080) );
  AND U9463 ( .A(n5081), .B(n5080), .Z(n7973) );
  NANDN U9464 ( .A(n5083), .B(n5082), .Z(n5087) );
  NAND U9465 ( .A(n5085), .B(n5084), .Z(n5086) );
  AND U9466 ( .A(n5087), .B(n5086), .Z(n8133) );
  NANDN U9467 ( .A(n5089), .B(n5088), .Z(n5093) );
  NAND U9468 ( .A(n5091), .B(n5090), .Z(n5092) );
  NAND U9469 ( .A(n5093), .B(n5092), .Z(n8134) );
  XNOR U9470 ( .A(n8133), .B(n8134), .Z(n8136) );
  NANDN U9471 ( .A(n5095), .B(n5094), .Z(n5099) );
  NAND U9472 ( .A(n5097), .B(n5096), .Z(n5098) );
  AND U9473 ( .A(n5099), .B(n5098), .Z(n8135) );
  XOR U9474 ( .A(n8136), .B(n8135), .Z(n7972) );
  NANDN U9475 ( .A(n5101), .B(n5100), .Z(n5105) );
  NAND U9476 ( .A(n5103), .B(n5102), .Z(n5104) );
  AND U9477 ( .A(n5105), .B(n5104), .Z(n7818) );
  NANDN U9478 ( .A(n5107), .B(n5106), .Z(n5111) );
  NAND U9479 ( .A(n5109), .B(n5108), .Z(n5110) );
  NAND U9480 ( .A(n5111), .B(n5110), .Z(n7819) );
  XNOR U9481 ( .A(n7818), .B(n7819), .Z(n7821) );
  NANDN U9482 ( .A(n5113), .B(n5112), .Z(n5117) );
  NAND U9483 ( .A(n5115), .B(n5114), .Z(n5116) );
  AND U9484 ( .A(n5117), .B(n5116), .Z(n7820) );
  XNOR U9485 ( .A(n7821), .B(n7820), .Z(n7971) );
  XOR U9486 ( .A(n7972), .B(n7971), .Z(n7974) );
  XNOR U9487 ( .A(n7973), .B(n7974), .Z(n7126) );
  NANDN U9488 ( .A(n5119), .B(n5118), .Z(n5123) );
  NAND U9489 ( .A(n5121), .B(n5120), .Z(n5122) );
  AND U9490 ( .A(n5123), .B(n5122), .Z(n6589) );
  NANDN U9491 ( .A(n5125), .B(n5124), .Z(n5129) );
  NAND U9492 ( .A(n5127), .B(n5126), .Z(n5128) );
  AND U9493 ( .A(n5129), .B(n5128), .Z(n6588) );
  XOR U9494 ( .A(n6589), .B(n6588), .Z(n6591) );
  NANDN U9495 ( .A(n5131), .B(n5130), .Z(n5135) );
  NAND U9496 ( .A(n5133), .B(n5132), .Z(n5134) );
  AND U9497 ( .A(n5135), .B(n5134), .Z(n6590) );
  XOR U9498 ( .A(n6591), .B(n6590), .Z(n6675) );
  NANDN U9499 ( .A(n5137), .B(n5136), .Z(n5141) );
  NAND U9500 ( .A(n5139), .B(n5138), .Z(n5140) );
  AND U9501 ( .A(n5141), .B(n5140), .Z(n6474) );
  NANDN U9502 ( .A(n5143), .B(n5142), .Z(n5147) );
  NAND U9503 ( .A(n5145), .B(n5144), .Z(n5146) );
  NAND U9504 ( .A(n5147), .B(n5146), .Z(n6475) );
  XNOR U9505 ( .A(n6474), .B(n6475), .Z(n6477) );
  NANDN U9506 ( .A(n5149), .B(n5148), .Z(n5153) );
  NAND U9507 ( .A(n5151), .B(n5150), .Z(n5152) );
  AND U9508 ( .A(n5153), .B(n5152), .Z(n6476) );
  XOR U9509 ( .A(n6477), .B(n6476), .Z(n6673) );
  NANDN U9510 ( .A(n5155), .B(n5154), .Z(n5159) );
  NANDN U9511 ( .A(n5157), .B(n5156), .Z(n5158) );
  AND U9512 ( .A(n5159), .B(n5158), .Z(n6672) );
  XNOR U9513 ( .A(n6673), .B(n6672), .Z(n6674) );
  XOR U9514 ( .A(n6675), .B(n6674), .Z(n7127) );
  XNOR U9515 ( .A(n7126), .B(n7127), .Z(n7129) );
  NANDN U9516 ( .A(n5161), .B(n5160), .Z(n5165) );
  NANDN U9517 ( .A(n5163), .B(n5162), .Z(n5164) );
  AND U9518 ( .A(n5165), .B(n5164), .Z(n7020) );
  NAND U9519 ( .A(n5167), .B(n5166), .Z(n5171) );
  NAND U9520 ( .A(n5169), .B(n5168), .Z(n5170) );
  AND U9521 ( .A(n5171), .B(n5170), .Z(n6720) );
  NANDN U9522 ( .A(n5173), .B(n5172), .Z(n5177) );
  NAND U9523 ( .A(n5175), .B(n5174), .Z(n5176) );
  NAND U9524 ( .A(n5177), .B(n5176), .Z(n6721) );
  XNOR U9525 ( .A(n6720), .B(n6721), .Z(n6723) );
  NANDN U9526 ( .A(n5179), .B(n5178), .Z(n5183) );
  NAND U9527 ( .A(n5181), .B(n5180), .Z(n5182) );
  AND U9528 ( .A(n5183), .B(n5182), .Z(n6722) );
  XOR U9529 ( .A(n6723), .B(n6722), .Z(n7019) );
  NANDN U9530 ( .A(n5185), .B(n5184), .Z(n5189) );
  NAND U9531 ( .A(n5187), .B(n5186), .Z(n5188) );
  AND U9532 ( .A(n5189), .B(n5188), .Z(n8223) );
  NANDN U9533 ( .A(n5191), .B(n5190), .Z(n5195) );
  NAND U9534 ( .A(n5193), .B(n5192), .Z(n5194) );
  NAND U9535 ( .A(n5195), .B(n5194), .Z(n8224) );
  XNOR U9536 ( .A(n8223), .B(n8224), .Z(n8226) );
  NANDN U9537 ( .A(n5197), .B(n5196), .Z(n5201) );
  NANDN U9538 ( .A(n5199), .B(n5198), .Z(n5200) );
  AND U9539 ( .A(n5201), .B(n5200), .Z(n8225) );
  XNOR U9540 ( .A(n8226), .B(n8225), .Z(n7018) );
  XOR U9541 ( .A(n7019), .B(n7018), .Z(n7021) );
  XNOR U9542 ( .A(n7020), .B(n7021), .Z(n7128) );
  XNOR U9543 ( .A(n7129), .B(n7128), .Z(n6666) );
  XNOR U9544 ( .A(n6667), .B(n6666), .Z(n6668) );
  NANDN U9545 ( .A(n5203), .B(n5202), .Z(n5207) );
  NANDN U9546 ( .A(n5205), .B(n5204), .Z(n5206) );
  AND U9547 ( .A(n5207), .B(n5206), .Z(n8970) );
  NANDN U9548 ( .A(n5209), .B(n5208), .Z(n5213) );
  OR U9549 ( .A(n5211), .B(n5210), .Z(n5212) );
  AND U9550 ( .A(n5213), .B(n5212), .Z(n8967) );
  NANDN U9551 ( .A(n5215), .B(n5214), .Z(n5219) );
  NANDN U9552 ( .A(n5217), .B(n5216), .Z(n5218) );
  NAND U9553 ( .A(n5219), .B(n5218), .Z(n8968) );
  XNOR U9554 ( .A(n8967), .B(n8968), .Z(n8969) );
  XOR U9555 ( .A(n8970), .B(n8969), .Z(n7135) );
  NANDN U9556 ( .A(n5221), .B(n5220), .Z(n5225) );
  NANDN U9557 ( .A(n5223), .B(n5222), .Z(n5224) );
  AND U9558 ( .A(n5225), .B(n5224), .Z(n8994) );
  NANDN U9559 ( .A(n5227), .B(n5226), .Z(n5231) );
  NANDN U9560 ( .A(n5229), .B(n5228), .Z(n5230) );
  AND U9561 ( .A(n5231), .B(n5230), .Z(n8991) );
  NANDN U9562 ( .A(n5233), .B(n5232), .Z(n5237) );
  NANDN U9563 ( .A(n5235), .B(n5234), .Z(n5236) );
  NAND U9564 ( .A(n5237), .B(n5236), .Z(n8992) );
  XNOR U9565 ( .A(n8991), .B(n8992), .Z(n8993) );
  XOR U9566 ( .A(n8994), .B(n8993), .Z(n7133) );
  NANDN U9567 ( .A(n5239), .B(n5238), .Z(n5243) );
  OR U9568 ( .A(n5241), .B(n5240), .Z(n5242) );
  AND U9569 ( .A(n5243), .B(n5242), .Z(n7132) );
  XNOR U9570 ( .A(n7133), .B(n7132), .Z(n7134) );
  XOR U9571 ( .A(n7135), .B(n7134), .Z(n6669) );
  XNOR U9572 ( .A(n6668), .B(n6669), .Z(n7042) );
  NANDN U9573 ( .A(n5245), .B(n5244), .Z(n5249) );
  NANDN U9574 ( .A(n5247), .B(n5246), .Z(n5248) );
  AND U9575 ( .A(n5249), .B(n5248), .Z(n7857) );
  NANDN U9576 ( .A(n5251), .B(n5250), .Z(n5255) );
  NAND U9577 ( .A(n5253), .B(n5252), .Z(n5254) );
  AND U9578 ( .A(n5255), .B(n5254), .Z(n8325) );
  NANDN U9579 ( .A(n5257), .B(n5256), .Z(n5261) );
  NAND U9580 ( .A(n5259), .B(n5258), .Z(n5260) );
  NAND U9581 ( .A(n5261), .B(n5260), .Z(n8326) );
  XNOR U9582 ( .A(n8325), .B(n8326), .Z(n8328) );
  NANDN U9583 ( .A(n5263), .B(n5262), .Z(n5267) );
  NAND U9584 ( .A(n5265), .B(n5264), .Z(n5266) );
  AND U9585 ( .A(n5267), .B(n5266), .Z(n8327) );
  XOR U9586 ( .A(n8328), .B(n8327), .Z(n7855) );
  NANDN U9587 ( .A(n5269), .B(n5268), .Z(n5273) );
  NANDN U9588 ( .A(n5271), .B(n5270), .Z(n5272) );
  AND U9589 ( .A(n5273), .B(n5272), .Z(n7854) );
  XNOR U9590 ( .A(n7855), .B(n7854), .Z(n7856) );
  XOR U9591 ( .A(n7857), .B(n7856), .Z(n6297) );
  NANDN U9592 ( .A(n5275), .B(n5274), .Z(n5279) );
  NANDN U9593 ( .A(n5277), .B(n5276), .Z(n5278) );
  AND U9594 ( .A(n5279), .B(n5278), .Z(n7633) );
  NANDN U9595 ( .A(n5281), .B(n5280), .Z(n5285) );
  NAND U9596 ( .A(n5283), .B(n5282), .Z(n5284) );
  AND U9597 ( .A(n5285), .B(n5284), .Z(n7729) );
  NANDN U9598 ( .A(n5287), .B(n5286), .Z(n5291) );
  NAND U9599 ( .A(n5289), .B(n5288), .Z(n5290) );
  AND U9600 ( .A(n5291), .B(n5290), .Z(n7728) );
  XOR U9601 ( .A(n7729), .B(n7728), .Z(n7731) );
  NANDN U9602 ( .A(n5293), .B(n5292), .Z(n5297) );
  NAND U9603 ( .A(n5295), .B(n5294), .Z(n5296) );
  AND U9604 ( .A(n5297), .B(n5296), .Z(n7730) );
  XOR U9605 ( .A(n7731), .B(n7730), .Z(n7631) );
  NANDN U9606 ( .A(n5299), .B(n5298), .Z(n5303) );
  NAND U9607 ( .A(n5301), .B(n5300), .Z(n5302) );
  AND U9608 ( .A(n5303), .B(n5302), .Z(n8710) );
  NANDN U9609 ( .A(n5305), .B(n5304), .Z(n5309) );
  NANDN U9610 ( .A(n5307), .B(n5306), .Z(n5308) );
  AND U9611 ( .A(n5309), .B(n5308), .Z(n8709) );
  XOR U9612 ( .A(n8710), .B(n8709), .Z(n8712) );
  NANDN U9613 ( .A(n5311), .B(n5310), .Z(n5315) );
  NANDN U9614 ( .A(n5313), .B(n5312), .Z(n5314) );
  AND U9615 ( .A(n5315), .B(n5314), .Z(n8711) );
  XNOR U9616 ( .A(n8712), .B(n8711), .Z(n7630) );
  XNOR U9617 ( .A(n7631), .B(n7630), .Z(n7632) );
  XOR U9618 ( .A(n7633), .B(n7632), .Z(n6295) );
  NANDN U9619 ( .A(n5317), .B(n5316), .Z(n5321) );
  NAND U9620 ( .A(n5319), .B(n5318), .Z(n5320) );
  NAND U9621 ( .A(n5321), .B(n5320), .Z(n6294) );
  XNOR U9622 ( .A(n6295), .B(n6294), .Z(n6296) );
  XNOR U9623 ( .A(n6297), .B(n6296), .Z(n8057) );
  NANDN U9624 ( .A(n5323), .B(n5322), .Z(n5327) );
  NANDN U9625 ( .A(n5325), .B(n5324), .Z(n5326) );
  AND U9626 ( .A(n5327), .B(n5326), .Z(n7904) );
  NANDN U9627 ( .A(n5329), .B(n5328), .Z(n5333) );
  NAND U9628 ( .A(n5331), .B(n5330), .Z(n5332) );
  AND U9629 ( .A(n5333), .B(n5332), .Z(n9015) );
  NANDN U9630 ( .A(n5335), .B(n5334), .Z(n5339) );
  NAND U9631 ( .A(n5337), .B(n5336), .Z(n5338) );
  NAND U9632 ( .A(n5339), .B(n5338), .Z(n9016) );
  XNOR U9633 ( .A(n9015), .B(n9016), .Z(n9018) );
  NANDN U9634 ( .A(n5341), .B(n5340), .Z(n5345) );
  NAND U9635 ( .A(n5343), .B(n5342), .Z(n5344) );
  AND U9636 ( .A(n5345), .B(n5344), .Z(n9017) );
  XOR U9637 ( .A(n9018), .B(n9017), .Z(n7903) );
  NANDN U9638 ( .A(n5347), .B(n5346), .Z(n5351) );
  NANDN U9639 ( .A(n5349), .B(n5348), .Z(n5350) );
  AND U9640 ( .A(n5351), .B(n5350), .Z(n7902) );
  XOR U9641 ( .A(n7903), .B(n7902), .Z(n7905) );
  XNOR U9642 ( .A(n7904), .B(n7905), .Z(n6901) );
  NANDN U9643 ( .A(n5353), .B(n5352), .Z(n5357) );
  NAND U9644 ( .A(n5355), .B(n5354), .Z(n5356) );
  NAND U9645 ( .A(n5357), .B(n5356), .Z(n6787) );
  NANDN U9646 ( .A(n5359), .B(n5358), .Z(n5363) );
  NAND U9647 ( .A(n5361), .B(n5360), .Z(n5362) );
  AND U9648 ( .A(n5363), .B(n5362), .Z(n8865) );
  NANDN U9649 ( .A(n5365), .B(n5364), .Z(n5369) );
  NAND U9650 ( .A(n5367), .B(n5366), .Z(n5368) );
  NAND U9651 ( .A(n5369), .B(n5368), .Z(n8866) );
  XNOR U9652 ( .A(n8865), .B(n8866), .Z(n8868) );
  NANDN U9653 ( .A(n5371), .B(n5370), .Z(n5375) );
  NAND U9654 ( .A(n5373), .B(n5372), .Z(n5374) );
  AND U9655 ( .A(n5375), .B(n5374), .Z(n8867) );
  XNOR U9656 ( .A(n8868), .B(n8867), .Z(n6786) );
  XOR U9657 ( .A(n6787), .B(n6786), .Z(n6789) );
  NANDN U9658 ( .A(n5377), .B(n5376), .Z(n5381) );
  NAND U9659 ( .A(n5379), .B(n5378), .Z(n5380) );
  AND U9660 ( .A(n5381), .B(n5380), .Z(n8379) );
  NANDN U9661 ( .A(n5383), .B(n5382), .Z(n5387) );
  NAND U9662 ( .A(n5385), .B(n5384), .Z(n5386) );
  NAND U9663 ( .A(n5387), .B(n5386), .Z(n8380) );
  XNOR U9664 ( .A(n8379), .B(n8380), .Z(n8381) );
  NAND U9665 ( .A(n5389), .B(n5388), .Z(n5393) );
  NAND U9666 ( .A(n5391), .B(n5390), .Z(n5392) );
  NAND U9667 ( .A(n5393), .B(n5392), .Z(n8382) );
  XOR U9668 ( .A(n8381), .B(n8382), .Z(n6788) );
  XOR U9669 ( .A(n6789), .B(n6788), .Z(n6900) );
  XOR U9670 ( .A(n6901), .B(n6900), .Z(n6903) );
  NANDN U9671 ( .A(n5395), .B(n5394), .Z(n5399) );
  NAND U9672 ( .A(n5397), .B(n5396), .Z(n5398) );
  AND U9673 ( .A(n5399), .B(n5398), .Z(n6619) );
  NANDN U9674 ( .A(n5401), .B(n5400), .Z(n5405) );
  NANDN U9675 ( .A(n5403), .B(n5402), .Z(n5404) );
  AND U9676 ( .A(n5405), .B(n5404), .Z(n6618) );
  XOR U9677 ( .A(n6619), .B(n6618), .Z(n6621) );
  NANDN U9678 ( .A(n5407), .B(n5406), .Z(n5411) );
  NANDN U9679 ( .A(n5409), .B(n5408), .Z(n5410) );
  AND U9680 ( .A(n5411), .B(n5410), .Z(n6620) );
  XOR U9681 ( .A(n6621), .B(n6620), .Z(n7513) );
  NAND U9682 ( .A(n5413), .B(n5412), .Z(n5417) );
  NAND U9683 ( .A(n5415), .B(n5414), .Z(n5416) );
  AND U9684 ( .A(n5417), .B(n5416), .Z(n8838) );
  NAND U9685 ( .A(n5419), .B(n5418), .Z(n5423) );
  NAND U9686 ( .A(n5421), .B(n5420), .Z(n5422) );
  AND U9687 ( .A(n5423), .B(n5422), .Z(n8836) );
  NANDN U9688 ( .A(n5425), .B(n5424), .Z(n5429) );
  NAND U9689 ( .A(n5427), .B(n5426), .Z(n5428) );
  AND U9690 ( .A(n5429), .B(n5428), .Z(n8835) );
  XOR U9691 ( .A(n8836), .B(n8835), .Z(n8837) );
  XOR U9692 ( .A(n8838), .B(n8837), .Z(n7511) );
  NANDN U9693 ( .A(n5431), .B(n5430), .Z(n5435) );
  NAND U9694 ( .A(n5433), .B(n5432), .Z(n5434) );
  AND U9695 ( .A(n5435), .B(n5434), .Z(n7570) );
  NANDN U9696 ( .A(n5437), .B(n5436), .Z(n5441) );
  NAND U9697 ( .A(n5439), .B(n5438), .Z(n5440) );
  NAND U9698 ( .A(n5441), .B(n5440), .Z(n7571) );
  XNOR U9699 ( .A(n7570), .B(n7571), .Z(n7573) );
  NANDN U9700 ( .A(n5443), .B(n5442), .Z(n5447) );
  NAND U9701 ( .A(n5445), .B(n5444), .Z(n5446) );
  AND U9702 ( .A(n5447), .B(n5446), .Z(n7572) );
  XNOR U9703 ( .A(n7573), .B(n7572), .Z(n7510) );
  XNOR U9704 ( .A(n7511), .B(n7510), .Z(n7512) );
  XNOR U9705 ( .A(n7513), .B(n7512), .Z(n6902) );
  XOR U9706 ( .A(n6903), .B(n6902), .Z(n8056) );
  NANDN U9707 ( .A(n5449), .B(n5448), .Z(n5453) );
  NAND U9708 ( .A(n5451), .B(n5450), .Z(n5452) );
  AND U9709 ( .A(n5453), .B(n5452), .Z(n6804) );
  NANDN U9710 ( .A(n5455), .B(n5454), .Z(n5459) );
  NAND U9711 ( .A(n5457), .B(n5456), .Z(n5458) );
  NAND U9712 ( .A(n5459), .B(n5458), .Z(n6805) );
  XNOR U9713 ( .A(n6804), .B(n6805), .Z(n6807) );
  NANDN U9714 ( .A(n5461), .B(n5460), .Z(n5465) );
  NAND U9715 ( .A(n5463), .B(n5462), .Z(n5464) );
  AND U9716 ( .A(n5465), .B(n5464), .Z(n6806) );
  XOR U9717 ( .A(n6807), .B(n6806), .Z(n8015) );
  NANDN U9718 ( .A(n5467), .B(n5466), .Z(n5471) );
  NAND U9719 ( .A(n5469), .B(n5468), .Z(n5470) );
  AND U9720 ( .A(n5471), .B(n5470), .Z(n8577) );
  NANDN U9721 ( .A(n5473), .B(n5472), .Z(n5477) );
  NAND U9722 ( .A(n5475), .B(n5474), .Z(n5476) );
  NAND U9723 ( .A(n5477), .B(n5476), .Z(n8578) );
  XNOR U9724 ( .A(n8577), .B(n8578), .Z(n8580) );
  NANDN U9725 ( .A(n5479), .B(n5478), .Z(n5483) );
  NAND U9726 ( .A(n5481), .B(n5480), .Z(n5482) );
  AND U9727 ( .A(n5483), .B(n5482), .Z(n8579) );
  XOR U9728 ( .A(n8580), .B(n8579), .Z(n8014) );
  NANDN U9729 ( .A(n5485), .B(n5484), .Z(n5489) );
  NANDN U9730 ( .A(n5487), .B(n5486), .Z(n5488) );
  AND U9731 ( .A(n5489), .B(n5488), .Z(n8013) );
  XOR U9732 ( .A(n8014), .B(n8013), .Z(n8016) );
  XOR U9733 ( .A(n8015), .B(n8016), .Z(n6417) );
  NANDN U9734 ( .A(n5491), .B(n5490), .Z(n5495) );
  NANDN U9735 ( .A(n5493), .B(n5492), .Z(n5494) );
  AND U9736 ( .A(n5495), .B(n5494), .Z(n7992) );
  NANDN U9737 ( .A(n5497), .B(n5496), .Z(n5501) );
  NANDN U9738 ( .A(n5499), .B(n5498), .Z(n5500) );
  AND U9739 ( .A(n5501), .B(n5500), .Z(n7989) );
  NANDN U9740 ( .A(n5503), .B(n5502), .Z(n5507) );
  NANDN U9741 ( .A(n5505), .B(n5504), .Z(n5506) );
  NAND U9742 ( .A(n5507), .B(n5506), .Z(n7990) );
  XNOR U9743 ( .A(n7989), .B(n7990), .Z(n7991) );
  XOR U9744 ( .A(n7992), .B(n7991), .Z(n6415) );
  NANDN U9745 ( .A(n5509), .B(n5508), .Z(n5513) );
  NAND U9746 ( .A(n5511), .B(n5510), .Z(n5512) );
  NAND U9747 ( .A(n5513), .B(n5512), .Z(n6414) );
  XNOR U9748 ( .A(n6415), .B(n6414), .Z(n6416) );
  XNOR U9749 ( .A(n6417), .B(n6416), .Z(n8055) );
  XOR U9750 ( .A(n8056), .B(n8055), .Z(n8058) );
  XNOR U9751 ( .A(n8057), .B(n8058), .Z(n7043) );
  XOR U9752 ( .A(n7042), .B(n7043), .Z(n7044) );
  XOR U9753 ( .A(n7045), .B(n7044), .Z(n7421) );
  NANDN U9754 ( .A(n5515), .B(n5514), .Z(n5519) );
  NAND U9755 ( .A(n5517), .B(n5516), .Z(n5518) );
  AND U9756 ( .A(n5519), .B(n5518), .Z(n8954) );
  NANDN U9757 ( .A(n5521), .B(n5520), .Z(n5525) );
  NANDN U9758 ( .A(n5523), .B(n5522), .Z(n5524) );
  AND U9759 ( .A(n5525), .B(n5524), .Z(n6942) );
  NANDN U9760 ( .A(n5527), .B(n5526), .Z(n5531) );
  NANDN U9761 ( .A(n5529), .B(n5528), .Z(n5530) );
  AND U9762 ( .A(n5531), .B(n5530), .Z(n6940) );
  NANDN U9763 ( .A(n5533), .B(n5532), .Z(n5537) );
  NANDN U9764 ( .A(n5535), .B(n5534), .Z(n5536) );
  NAND U9765 ( .A(n5537), .B(n5536), .Z(n6941) );
  XOR U9766 ( .A(n6940), .B(n6941), .Z(n6943) );
  XOR U9767 ( .A(n6942), .B(n6943), .Z(n8955) );
  XNOR U9768 ( .A(n8954), .B(n8955), .Z(n8957) );
  NANDN U9769 ( .A(n5539), .B(n5538), .Z(n5543) );
  NAND U9770 ( .A(n5541), .B(n5540), .Z(n5542) );
  AND U9771 ( .A(n5543), .B(n5542), .Z(n8302) );
  NANDN U9772 ( .A(n5545), .B(n5544), .Z(n5549) );
  NAND U9773 ( .A(n5547), .B(n5546), .Z(n5548) );
  AND U9774 ( .A(n5549), .B(n5548), .Z(n8301) );
  XOR U9775 ( .A(n8302), .B(n8301), .Z(n8304) );
  NANDN U9776 ( .A(n5551), .B(n5550), .Z(n5555) );
  NAND U9777 ( .A(n5553), .B(n5552), .Z(n5554) );
  AND U9778 ( .A(n5555), .B(n5554), .Z(n8303) );
  XOR U9779 ( .A(n8304), .B(n8303), .Z(n6681) );
  NANDN U9780 ( .A(n5557), .B(n5556), .Z(n5561) );
  NAND U9781 ( .A(n5559), .B(n5558), .Z(n5560) );
  AND U9782 ( .A(n5561), .B(n5560), .Z(n8680) );
  NAND U9783 ( .A(n5563), .B(n5562), .Z(n5567) );
  NAND U9784 ( .A(n5565), .B(n5564), .Z(n5566) );
  AND U9785 ( .A(n5567), .B(n5566), .Z(n8679) );
  XOR U9786 ( .A(n8680), .B(n8679), .Z(n8682) );
  NAND U9787 ( .A(n5569), .B(n5568), .Z(n5573) );
  NAND U9788 ( .A(n5571), .B(n5570), .Z(n5572) );
  AND U9789 ( .A(n5573), .B(n5572), .Z(n8681) );
  XOR U9790 ( .A(n8682), .B(n8681), .Z(n6679) );
  NANDN U9791 ( .A(n5575), .B(n5574), .Z(n5579) );
  NANDN U9792 ( .A(n5577), .B(n5576), .Z(n5578) );
  AND U9793 ( .A(n5579), .B(n5578), .Z(n6678) );
  XNOR U9794 ( .A(n6679), .B(n6678), .Z(n6680) );
  XNOR U9795 ( .A(n6681), .B(n6680), .Z(n8956) );
  XNOR U9796 ( .A(n8957), .B(n8956), .Z(n8652) );
  NANDN U9797 ( .A(n5581), .B(n5580), .Z(n5585) );
  NANDN U9798 ( .A(n5583), .B(n5582), .Z(n5584) );
  AND U9799 ( .A(n5585), .B(n5584), .Z(n7997) );
  NANDN U9800 ( .A(n5587), .B(n5586), .Z(n5591) );
  NANDN U9801 ( .A(n5589), .B(n5588), .Z(n5590) );
  AND U9802 ( .A(n5591), .B(n5590), .Z(n7995) );
  NANDN U9803 ( .A(n5593), .B(n5592), .Z(n5597) );
  NANDN U9804 ( .A(n5595), .B(n5594), .Z(n5596) );
  NAND U9805 ( .A(n5597), .B(n5596), .Z(n7996) );
  XOR U9806 ( .A(n7995), .B(n7996), .Z(n7998) );
  XNOR U9807 ( .A(n7997), .B(n7998), .Z(n8589) );
  NAND U9808 ( .A(n5599), .B(n5598), .Z(n5603) );
  NAND U9809 ( .A(n5601), .B(n5600), .Z(n5602) );
  AND U9810 ( .A(n5603), .B(n5602), .Z(n6852) );
  NAND U9811 ( .A(n5605), .B(n5604), .Z(n5609) );
  NAND U9812 ( .A(n5607), .B(n5606), .Z(n5608) );
  NAND U9813 ( .A(n5609), .B(n5608), .Z(n6853) );
  XNOR U9814 ( .A(n6852), .B(n6853), .Z(n6855) );
  NANDN U9815 ( .A(n5611), .B(n5610), .Z(n5615) );
  NAND U9816 ( .A(n5613), .B(n5612), .Z(n5614) );
  AND U9817 ( .A(n5615), .B(n5614), .Z(n6854) );
  XOR U9818 ( .A(n6855), .B(n6854), .Z(n7357) );
  NANDN U9819 ( .A(n5617), .B(n5616), .Z(n5621) );
  NAND U9820 ( .A(n5619), .B(n5618), .Z(n5620) );
  AND U9821 ( .A(n5621), .B(n5620), .Z(n6858) );
  NANDN U9822 ( .A(n5623), .B(n5622), .Z(n5627) );
  NAND U9823 ( .A(n5625), .B(n5624), .Z(n5626) );
  NAND U9824 ( .A(n5627), .B(n5626), .Z(n6859) );
  XNOR U9825 ( .A(n6858), .B(n6859), .Z(n6861) );
  NAND U9826 ( .A(n5629), .B(n5628), .Z(n5633) );
  NAND U9827 ( .A(n5631), .B(n5630), .Z(n5632) );
  AND U9828 ( .A(n5633), .B(n5632), .Z(n6860) );
  XOR U9829 ( .A(n6861), .B(n6860), .Z(n7355) );
  NANDN U9830 ( .A(n5635), .B(n5634), .Z(n5639) );
  NANDN U9831 ( .A(n5637), .B(n5636), .Z(n5638) );
  AND U9832 ( .A(n5639), .B(n5638), .Z(n7354) );
  XNOR U9833 ( .A(n7355), .B(n7354), .Z(n7356) );
  XOR U9834 ( .A(n7357), .B(n7356), .Z(n8590) );
  XNOR U9835 ( .A(n8589), .B(n8590), .Z(n8592) );
  NANDN U9836 ( .A(n5641), .B(n5640), .Z(n5645) );
  NANDN U9837 ( .A(n5643), .B(n5642), .Z(n5644) );
  AND U9838 ( .A(n5645), .B(n5644), .Z(n8673) );
  NANDN U9839 ( .A(n5647), .B(n5646), .Z(n5651) );
  NAND U9840 ( .A(n5649), .B(n5648), .Z(n5650) );
  NAND U9841 ( .A(n5651), .B(n5650), .Z(n8674) );
  XNOR U9842 ( .A(n8673), .B(n8674), .Z(n8676) );
  NANDN U9843 ( .A(n5653), .B(n5652), .Z(n5657) );
  NAND U9844 ( .A(n5655), .B(n5654), .Z(n5656) );
  AND U9845 ( .A(n5657), .B(n5656), .Z(n8675) );
  XOR U9846 ( .A(n8676), .B(n8675), .Z(n7986) );
  NANDN U9847 ( .A(n5659), .B(n5658), .Z(n5663) );
  NANDN U9848 ( .A(n5661), .B(n5660), .Z(n5662) );
  AND U9849 ( .A(n5663), .B(n5662), .Z(n7983) );
  NANDN U9850 ( .A(n5665), .B(n5664), .Z(n5669) );
  NANDN U9851 ( .A(n5667), .B(n5666), .Z(n5668) );
  NAND U9852 ( .A(n5669), .B(n5668), .Z(n7984) );
  XNOR U9853 ( .A(n7983), .B(n7984), .Z(n7985) );
  XNOR U9854 ( .A(n7986), .B(n7985), .Z(n8591) );
  XNOR U9855 ( .A(n8592), .B(n8591), .Z(n8650) );
  NAND U9856 ( .A(n5671), .B(n5670), .Z(n5675) );
  NAND U9857 ( .A(n5673), .B(n5672), .Z(n5674) );
  AND U9858 ( .A(n5675), .B(n5674), .Z(n8649) );
  XOR U9859 ( .A(n8650), .B(n8649), .Z(n8651) );
  XOR U9860 ( .A(n8652), .B(n8651), .Z(n7123) );
  NANDN U9861 ( .A(n5677), .B(n5676), .Z(n5681) );
  NAND U9862 ( .A(n5679), .B(n5678), .Z(n5680) );
  AND U9863 ( .A(n5681), .B(n5680), .Z(n8463) );
  NAND U9864 ( .A(n5683), .B(n5682), .Z(n5687) );
  NAND U9865 ( .A(n5685), .B(n5684), .Z(n5686) );
  NAND U9866 ( .A(n5687), .B(n5686), .Z(n8464) );
  XNOR U9867 ( .A(n8463), .B(n8464), .Z(n8466) );
  NAND U9868 ( .A(n5689), .B(n5688), .Z(n5693) );
  NAND U9869 ( .A(n5691), .B(n5690), .Z(n5692) );
  AND U9870 ( .A(n5693), .B(n5692), .Z(n8465) );
  XOR U9871 ( .A(n8466), .B(n8465), .Z(n6996) );
  NANDN U9872 ( .A(n5695), .B(n5694), .Z(n5699) );
  NAND U9873 ( .A(n5697), .B(n5696), .Z(n5698) );
  AND U9874 ( .A(n5699), .B(n5698), .Z(n7800) );
  NANDN U9875 ( .A(n5701), .B(n5700), .Z(n5705) );
  NAND U9876 ( .A(n5703), .B(n5702), .Z(n5704) );
  NAND U9877 ( .A(n5705), .B(n5704), .Z(n7801) );
  XNOR U9878 ( .A(n7800), .B(n7801), .Z(n7803) );
  NANDN U9879 ( .A(n5707), .B(n5706), .Z(n5711) );
  NAND U9880 ( .A(n5709), .B(n5708), .Z(n5710) );
  AND U9881 ( .A(n5711), .B(n5710), .Z(n7802) );
  XOR U9882 ( .A(n7803), .B(n7802), .Z(n6995) );
  NANDN U9883 ( .A(n5713), .B(n5712), .Z(n5717) );
  NAND U9884 ( .A(n5715), .B(n5714), .Z(n5716) );
  AND U9885 ( .A(n5717), .B(n5716), .Z(n8247) );
  NANDN U9886 ( .A(n5719), .B(n5718), .Z(n5723) );
  NAND U9887 ( .A(n5721), .B(n5720), .Z(n5722) );
  NAND U9888 ( .A(n5723), .B(n5722), .Z(n8248) );
  XNOR U9889 ( .A(n8247), .B(n8248), .Z(n8250) );
  NANDN U9890 ( .A(n5725), .B(n5724), .Z(n5729) );
  NAND U9891 ( .A(n5727), .B(n5726), .Z(n5728) );
  AND U9892 ( .A(n5729), .B(n5728), .Z(n8249) );
  XNOR U9893 ( .A(n8250), .B(n8249), .Z(n6994) );
  XOR U9894 ( .A(n6995), .B(n6994), .Z(n6997) );
  XOR U9895 ( .A(n6996), .B(n6997), .Z(n6309) );
  NANDN U9896 ( .A(n5731), .B(n5730), .Z(n5735) );
  NAND U9897 ( .A(n5733), .B(n5732), .Z(n5734) );
  AND U9898 ( .A(n5735), .B(n5734), .Z(n8391) );
  NANDN U9899 ( .A(n5737), .B(n5736), .Z(n5741) );
  NAND U9900 ( .A(n5739), .B(n5738), .Z(n5740) );
  NAND U9901 ( .A(n5741), .B(n5740), .Z(n8392) );
  XNOR U9902 ( .A(n8391), .B(n8392), .Z(n8394) );
  NANDN U9903 ( .A(n5743), .B(n5742), .Z(n5747) );
  NAND U9904 ( .A(n5745), .B(n5744), .Z(n5746) );
  AND U9905 ( .A(n5747), .B(n5746), .Z(n8393) );
  XOR U9906 ( .A(n8394), .B(n8393), .Z(n7038) );
  NANDN U9907 ( .A(n5749), .B(n5748), .Z(n5753) );
  NANDN U9908 ( .A(n5751), .B(n5750), .Z(n5752) );
  AND U9909 ( .A(n5753), .B(n5752), .Z(n7036) );
  NANDN U9910 ( .A(n5755), .B(n5754), .Z(n5759) );
  NANDN U9911 ( .A(n5757), .B(n5756), .Z(n5758) );
  NAND U9912 ( .A(n5759), .B(n5758), .Z(n7037) );
  XOR U9913 ( .A(n7036), .B(n7037), .Z(n7039) );
  XOR U9914 ( .A(n7038), .B(n7039), .Z(n6307) );
  NANDN U9915 ( .A(n5761), .B(n5760), .Z(n5765) );
  NANDN U9916 ( .A(n5763), .B(n5762), .Z(n5764) );
  AND U9917 ( .A(n5765), .B(n5764), .Z(n7851) );
  NANDN U9918 ( .A(n5767), .B(n5766), .Z(n5771) );
  NAND U9919 ( .A(n5769), .B(n5768), .Z(n5770) );
  AND U9920 ( .A(n5771), .B(n5770), .Z(n8349) );
  NANDN U9921 ( .A(n5773), .B(n5772), .Z(n5777) );
  NAND U9922 ( .A(n5775), .B(n5774), .Z(n5776) );
  NAND U9923 ( .A(n5777), .B(n5776), .Z(n8350) );
  XNOR U9924 ( .A(n8349), .B(n8350), .Z(n8352) );
  NANDN U9925 ( .A(n5779), .B(n5778), .Z(n5783) );
  NAND U9926 ( .A(n5781), .B(n5780), .Z(n5782) );
  AND U9927 ( .A(n5783), .B(n5782), .Z(n8351) );
  XOR U9928 ( .A(n8352), .B(n8351), .Z(n7849) );
  NANDN U9929 ( .A(n5785), .B(n5784), .Z(n5789) );
  NAND U9930 ( .A(n5787), .B(n5786), .Z(n5788) );
  AND U9931 ( .A(n5789), .B(n5788), .Z(n8697) );
  NANDN U9932 ( .A(n5791), .B(n5790), .Z(n5795) );
  NANDN U9933 ( .A(n5793), .B(n5792), .Z(n5794) );
  NAND U9934 ( .A(n5795), .B(n5794), .Z(n8698) );
  XNOR U9935 ( .A(n8697), .B(n8698), .Z(n8700) );
  NANDN U9936 ( .A(n5797), .B(n5796), .Z(n5801) );
  NAND U9937 ( .A(n5799), .B(n5798), .Z(n5800) );
  AND U9938 ( .A(n5801), .B(n5800), .Z(n8699) );
  XNOR U9939 ( .A(n8700), .B(n8699), .Z(n7848) );
  XNOR U9940 ( .A(n7849), .B(n7848), .Z(n7850) );
  XNOR U9941 ( .A(n7851), .B(n7850), .Z(n6306) );
  XNOR U9942 ( .A(n6307), .B(n6306), .Z(n6308) );
  XOR U9943 ( .A(n6309), .B(n6308), .Z(n6560) );
  NANDN U9944 ( .A(n5803), .B(n5802), .Z(n5807) );
  NAND U9945 ( .A(n5805), .B(n5804), .Z(n5806) );
  AND U9946 ( .A(n5807), .B(n5806), .Z(n8853) );
  NANDN U9947 ( .A(n5809), .B(n5808), .Z(n5813) );
  NAND U9948 ( .A(n5811), .B(n5810), .Z(n5812) );
  NAND U9949 ( .A(n5813), .B(n5812), .Z(n8854) );
  XNOR U9950 ( .A(n8853), .B(n8854), .Z(n8856) );
  NANDN U9951 ( .A(n5815), .B(n5814), .Z(n5819) );
  NAND U9952 ( .A(n5817), .B(n5816), .Z(n5818) );
  AND U9953 ( .A(n5819), .B(n5818), .Z(n8855) );
  XOR U9954 ( .A(n8856), .B(n8855), .Z(n8051) );
  NANDN U9955 ( .A(n5821), .B(n5820), .Z(n5825) );
  NANDN U9956 ( .A(n5823), .B(n5822), .Z(n5824) );
  AND U9957 ( .A(n5825), .B(n5824), .Z(n8049) );
  NANDN U9958 ( .A(n5827), .B(n5826), .Z(n5831) );
  NANDN U9959 ( .A(n5829), .B(n5828), .Z(n5830) );
  NAND U9960 ( .A(n5831), .B(n5830), .Z(n8050) );
  XOR U9961 ( .A(n8049), .B(n8050), .Z(n8052) );
  XOR U9962 ( .A(n8051), .B(n8052), .Z(n6165) );
  NANDN U9963 ( .A(n5833), .B(n5832), .Z(n5837) );
  NAND U9964 ( .A(n5835), .B(n5834), .Z(n5836) );
  AND U9965 ( .A(n5837), .B(n5836), .Z(n8181) );
  NANDN U9966 ( .A(n5839), .B(n5838), .Z(n5843) );
  NAND U9967 ( .A(n5841), .B(n5840), .Z(n5842) );
  NAND U9968 ( .A(n5843), .B(n5842), .Z(n8182) );
  XNOR U9969 ( .A(n8181), .B(n8182), .Z(n8184) );
  NANDN U9970 ( .A(n5845), .B(n5844), .Z(n5849) );
  NAND U9971 ( .A(n5847), .B(n5846), .Z(n5848) );
  AND U9972 ( .A(n5849), .B(n5848), .Z(n8183) );
  XOR U9973 ( .A(n8184), .B(n8183), .Z(n7374) );
  NANDN U9974 ( .A(n5851), .B(n5850), .Z(n5855) );
  NANDN U9975 ( .A(n5853), .B(n5852), .Z(n5854) );
  AND U9976 ( .A(n5855), .B(n5854), .Z(n7372) );
  NANDN U9977 ( .A(n5857), .B(n5856), .Z(n5861) );
  NANDN U9978 ( .A(n5859), .B(n5858), .Z(n5860) );
  NAND U9979 ( .A(n5861), .B(n5860), .Z(n7373) );
  XOR U9980 ( .A(n7372), .B(n7373), .Z(n7375) );
  XOR U9981 ( .A(n7374), .B(n7375), .Z(n6163) );
  NANDN U9982 ( .A(n5863), .B(n5862), .Z(n5867) );
  NAND U9983 ( .A(n5865), .B(n5864), .Z(n5866) );
  NAND U9984 ( .A(n5867), .B(n5866), .Z(n6162) );
  XNOR U9985 ( .A(n6163), .B(n6162), .Z(n6164) );
  XOR U9986 ( .A(n6165), .B(n6164), .Z(n6558) );
  NAND U9987 ( .A(n5869), .B(n5868), .Z(n5873) );
  NAND U9988 ( .A(n5871), .B(n5870), .Z(n5872) );
  AND U9989 ( .A(n5873), .B(n5872), .Z(n6559) );
  XOR U9990 ( .A(n6558), .B(n6559), .Z(n6561) );
  XNOR U9991 ( .A(n6560), .B(n6561), .Z(n7120) );
  NANDN U9992 ( .A(n5875), .B(n5874), .Z(n5879) );
  NAND U9993 ( .A(n5877), .B(n5876), .Z(n5878) );
  AND U9994 ( .A(n5879), .B(n5878), .Z(n8091) );
  NANDN U9995 ( .A(n5881), .B(n5880), .Z(n5885) );
  NAND U9996 ( .A(n5883), .B(n5882), .Z(n5884) );
  NAND U9997 ( .A(n5885), .B(n5884), .Z(n8092) );
  XNOR U9998 ( .A(n8091), .B(n8092), .Z(n8094) );
  NANDN U9999 ( .A(n5887), .B(n5886), .Z(n5891) );
  NAND U10000 ( .A(n5889), .B(n5888), .Z(n5890) );
  AND U10001 ( .A(n5891), .B(n5890), .Z(n8093) );
  XOR U10002 ( .A(n8094), .B(n8093), .Z(n7206) );
  NANDN U10003 ( .A(n5893), .B(n5892), .Z(n5897) );
  NAND U10004 ( .A(n5895), .B(n5894), .Z(n5896) );
  AND U10005 ( .A(n5897), .B(n5896), .Z(n8109) );
  NANDN U10006 ( .A(n5899), .B(n5898), .Z(n5903) );
  NAND U10007 ( .A(n5901), .B(n5900), .Z(n5902) );
  NAND U10008 ( .A(n5903), .B(n5902), .Z(n8110) );
  XNOR U10009 ( .A(n8109), .B(n8110), .Z(n8112) );
  NANDN U10010 ( .A(n5905), .B(n5904), .Z(n5909) );
  NAND U10011 ( .A(n5907), .B(n5906), .Z(n5908) );
  AND U10012 ( .A(n5909), .B(n5908), .Z(n8111) );
  XOR U10013 ( .A(n8112), .B(n8111), .Z(n7205) );
  NANDN U10014 ( .A(n5911), .B(n5910), .Z(n5915) );
  NANDN U10015 ( .A(n5913), .B(n5912), .Z(n5914) );
  AND U10016 ( .A(n5915), .B(n5914), .Z(n7204) );
  XOR U10017 ( .A(n7205), .B(n7204), .Z(n7207) );
  XOR U10018 ( .A(n7206), .B(n7207), .Z(n7669) );
  NANDN U10019 ( .A(n5917), .B(n5916), .Z(n5921) );
  NAND U10020 ( .A(n5919), .B(n5918), .Z(n5920) );
  AND U10021 ( .A(n5921), .B(n5920), .Z(n8073) );
  NANDN U10022 ( .A(n5923), .B(n5922), .Z(n5927) );
  NAND U10023 ( .A(n5925), .B(n5924), .Z(n5926) );
  NAND U10024 ( .A(n5927), .B(n5926), .Z(n8074) );
  XNOR U10025 ( .A(n8073), .B(n8074), .Z(n8076) );
  NANDN U10026 ( .A(n5929), .B(n5928), .Z(n5933) );
  NAND U10027 ( .A(n5931), .B(n5930), .Z(n5932) );
  AND U10028 ( .A(n5933), .B(n5932), .Z(n8075) );
  XOR U10029 ( .A(n8076), .B(n8075), .Z(n7182) );
  NANDN U10030 ( .A(n5935), .B(n5934), .Z(n5939) );
  NANDN U10031 ( .A(n5937), .B(n5936), .Z(n5938) );
  AND U10032 ( .A(n5939), .B(n5938), .Z(n7180) );
  NANDN U10033 ( .A(n5941), .B(n5940), .Z(n5945) );
  NANDN U10034 ( .A(n5943), .B(n5942), .Z(n5944) );
  NAND U10035 ( .A(n5945), .B(n5944), .Z(n7181) );
  XOR U10036 ( .A(n7180), .B(n7181), .Z(n7183) );
  XOR U10037 ( .A(n7182), .B(n7183), .Z(n7667) );
  NANDN U10038 ( .A(n5947), .B(n5946), .Z(n5951) );
  NAND U10039 ( .A(n5949), .B(n5948), .Z(n5950) );
  NAND U10040 ( .A(n5951), .B(n5950), .Z(n7666) );
  XNOR U10041 ( .A(n7667), .B(n7666), .Z(n7668) );
  XNOR U10042 ( .A(n7669), .B(n7668), .Z(n8964) );
  NANDN U10043 ( .A(n5953), .B(n5952), .Z(n5957) );
  NAND U10044 ( .A(n5955), .B(n5954), .Z(n5956) );
  AND U10045 ( .A(n5957), .B(n5956), .Z(n6126) );
  NANDN U10046 ( .A(n5959), .B(n5958), .Z(n5963) );
  NANDN U10047 ( .A(n5961), .B(n5960), .Z(n5962) );
  AND U10048 ( .A(n5963), .B(n5962), .Z(n8045) );
  NANDN U10049 ( .A(n5965), .B(n5964), .Z(n5969) );
  NANDN U10050 ( .A(n5967), .B(n5966), .Z(n5968) );
  AND U10051 ( .A(n5969), .B(n5968), .Z(n8043) );
  NANDN U10052 ( .A(n5971), .B(n5970), .Z(n5975) );
  NANDN U10053 ( .A(n5973), .B(n5972), .Z(n5974) );
  NAND U10054 ( .A(n5975), .B(n5974), .Z(n8044) );
  XOR U10055 ( .A(n8043), .B(n8044), .Z(n8046) );
  XOR U10056 ( .A(n8045), .B(n8046), .Z(n6127) );
  XNOR U10057 ( .A(n6126), .B(n6127), .Z(n6129) );
  NANDN U10058 ( .A(n5977), .B(n5976), .Z(n5981) );
  NAND U10059 ( .A(n5979), .B(n5978), .Z(n5980) );
  AND U10060 ( .A(n5981), .B(n5980), .Z(n8619) );
  NANDN U10061 ( .A(n5983), .B(n5982), .Z(n5987) );
  NAND U10062 ( .A(n5985), .B(n5984), .Z(n5986) );
  NAND U10063 ( .A(n5987), .B(n5986), .Z(n8620) );
  XNOR U10064 ( .A(n8619), .B(n8620), .Z(n8622) );
  NANDN U10065 ( .A(n5989), .B(n5988), .Z(n5993) );
  NAND U10066 ( .A(n5991), .B(n5990), .Z(n5992) );
  AND U10067 ( .A(n5993), .B(n5992), .Z(n8621) );
  XOR U10068 ( .A(n8622), .B(n8621), .Z(n6393) );
  NAND U10069 ( .A(n5995), .B(n5994), .Z(n5999) );
  NAND U10070 ( .A(n5997), .B(n5996), .Z(n5998) );
  AND U10071 ( .A(n5999), .B(n5998), .Z(n7872) );
  NANDN U10072 ( .A(n6001), .B(n6000), .Z(n6005) );
  NAND U10073 ( .A(n6003), .B(n6002), .Z(n6004) );
  NAND U10074 ( .A(n6005), .B(n6004), .Z(n7873) );
  XNOR U10075 ( .A(n7872), .B(n7873), .Z(n7875) );
  NANDN U10076 ( .A(n6007), .B(n6006), .Z(n6011) );
  NAND U10077 ( .A(n6009), .B(n6008), .Z(n6010) );
  AND U10078 ( .A(n6011), .B(n6010), .Z(n7874) );
  XOR U10079 ( .A(n7875), .B(n7874), .Z(n6391) );
  NANDN U10080 ( .A(n6013), .B(n6012), .Z(n6017) );
  NANDN U10081 ( .A(n6015), .B(n6014), .Z(n6016) );
  AND U10082 ( .A(n6017), .B(n6016), .Z(n6390) );
  XNOR U10083 ( .A(n6391), .B(n6390), .Z(n6392) );
  XNOR U10084 ( .A(n6393), .B(n6392), .Z(n6128) );
  XNOR U10085 ( .A(n6129), .B(n6128), .Z(n8962) );
  NANDN U10086 ( .A(n6019), .B(n6018), .Z(n6023) );
  NAND U10087 ( .A(n6021), .B(n6020), .Z(n6022) );
  AND U10088 ( .A(n6023), .B(n6022), .Z(n7673) );
  NAND U10089 ( .A(n6025), .B(n6024), .Z(n6029) );
  NAND U10090 ( .A(n6027), .B(n6026), .Z(n6028) );
  NAND U10091 ( .A(n6029), .B(n6028), .Z(n6762) );
  NANDN U10092 ( .A(n6031), .B(n6030), .Z(n6035) );
  NANDN U10093 ( .A(n6033), .B(n6032), .Z(n6034) );
  AND U10094 ( .A(n6035), .B(n6034), .Z(n6763) );
  XOR U10095 ( .A(n6762), .B(n6763), .Z(n6765) );
  NANDN U10096 ( .A(n6037), .B(n6036), .Z(n6041) );
  NANDN U10097 ( .A(n6039), .B(n6038), .Z(n6040) );
  AND U10098 ( .A(n6041), .B(n6040), .Z(n6764) );
  XOR U10099 ( .A(n6765), .B(n6764), .Z(n7672) );
  XOR U10100 ( .A(n7673), .B(n7672), .Z(n7675) );
  NANDN U10101 ( .A(n6043), .B(n6042), .Z(n6047) );
  NAND U10102 ( .A(n6045), .B(n6044), .Z(n6046) );
  AND U10103 ( .A(n6047), .B(n6046), .Z(n8799) );
  NANDN U10104 ( .A(n6049), .B(n6048), .Z(n6053) );
  NAND U10105 ( .A(n6051), .B(n6050), .Z(n6052) );
  NAND U10106 ( .A(n6053), .B(n6052), .Z(n8800) );
  XNOR U10107 ( .A(n8799), .B(n8800), .Z(n8802) );
  NANDN U10108 ( .A(n6055), .B(n6054), .Z(n6059) );
  NAND U10109 ( .A(n6057), .B(n6056), .Z(n6058) );
  AND U10110 ( .A(n6059), .B(n6058), .Z(n8801) );
  XOR U10111 ( .A(n8802), .B(n8801), .Z(n6735) );
  NANDN U10112 ( .A(n6061), .B(n6060), .Z(n6065) );
  NANDN U10113 ( .A(n6063), .B(n6062), .Z(n6064) );
  AND U10114 ( .A(n6065), .B(n6064), .Z(n6732) );
  NANDN U10115 ( .A(n6067), .B(n6066), .Z(n6071) );
  NANDN U10116 ( .A(n6069), .B(n6068), .Z(n6070) );
  NAND U10117 ( .A(n6071), .B(n6070), .Z(n6733) );
  XNOR U10118 ( .A(n6732), .B(n6733), .Z(n6734) );
  XNOR U10119 ( .A(n6735), .B(n6734), .Z(n7674) );
  XNOR U10120 ( .A(n7675), .B(n7674), .Z(n8961) );
  XOR U10121 ( .A(n8962), .B(n8961), .Z(n8963) );
  XOR U10122 ( .A(n8964), .B(n8963), .Z(n7121) );
  XOR U10123 ( .A(n7120), .B(n7121), .Z(n7122) );
  XOR U10124 ( .A(n7123), .B(n7122), .Z(n7420) );
  XOR U10125 ( .A(n7421), .B(n7420), .Z(n7422) );
  XOR U10126 ( .A(n7423), .B(n7422), .Z(n7240) );
  XOR U10127 ( .A(n7241), .B(n7240), .Z(n7242) );
  XOR U10128 ( .A(n7243), .B(n7242), .Z(n7230) );
  XNOR U10129 ( .A(n7231), .B(n7230), .Z(o[1]) );
  NAND U10130 ( .A(n6073), .B(n6072), .Z(n6077) );
  NAND U10131 ( .A(n6075), .B(n6074), .Z(n6076) );
  NAND U10132 ( .A(n6077), .B(n6076), .Z(n9801) );
  NAND U10133 ( .A(n6079), .B(n6078), .Z(n6083) );
  NAND U10134 ( .A(n6081), .B(n6080), .Z(n6082) );
  AND U10135 ( .A(n6083), .B(n6082), .Z(n9800) );
  XOR U10136 ( .A(n9801), .B(n9800), .Z(n9803) );
  NANDN U10137 ( .A(n6085), .B(n6084), .Z(n6089) );
  OR U10138 ( .A(n6087), .B(n6086), .Z(n6088) );
  AND U10139 ( .A(n6089), .B(n6088), .Z(n9115) );
  NANDN U10140 ( .A(n6091), .B(n6090), .Z(n6095) );
  OR U10141 ( .A(n6093), .B(n6092), .Z(n6094) );
  AND U10142 ( .A(n6095), .B(n6094), .Z(n9112) );
  NANDN U10143 ( .A(n6097), .B(n6096), .Z(n6101) );
  NANDN U10144 ( .A(n6099), .B(n6098), .Z(n6100) );
  AND U10145 ( .A(n6101), .B(n6100), .Z(n9126) );
  NANDN U10146 ( .A(n6103), .B(n6102), .Z(n6107) );
  NANDN U10147 ( .A(n6105), .B(n6104), .Z(n6106) );
  AND U10148 ( .A(n6107), .B(n6106), .Z(n9124) );
  NANDN U10149 ( .A(n6109), .B(n6108), .Z(n6113) );
  OR U10150 ( .A(n6111), .B(n6110), .Z(n6112) );
  NAND U10151 ( .A(n6113), .B(n6112), .Z(n9125) );
  XOR U10152 ( .A(n9124), .B(n9125), .Z(n9127) );
  XOR U10153 ( .A(n9126), .B(n9127), .Z(n9113) );
  XNOR U10154 ( .A(n9112), .B(n9113), .Z(n9114) );
  XNOR U10155 ( .A(n9115), .B(n9114), .Z(n10505) );
  NAND U10156 ( .A(n6115), .B(n6114), .Z(n6119) );
  NAND U10157 ( .A(n6117), .B(n6116), .Z(n6118) );
  AND U10158 ( .A(n6119), .B(n6118), .Z(n10455) );
  NANDN U10159 ( .A(n6121), .B(n6120), .Z(n6125) );
  OR U10160 ( .A(n6123), .B(n6122), .Z(n6124) );
  AND U10161 ( .A(n6125), .B(n6124), .Z(n10517) );
  NANDN U10162 ( .A(n6127), .B(n6126), .Z(n6131) );
  NAND U10163 ( .A(n6129), .B(n6128), .Z(n6130) );
  AND U10164 ( .A(n6131), .B(n6130), .Z(n10515) );
  NANDN U10165 ( .A(n6133), .B(n6132), .Z(n6137) );
  OR U10166 ( .A(n6135), .B(n6134), .Z(n6136) );
  AND U10167 ( .A(n6137), .B(n6136), .Z(n10514) );
  XNOR U10168 ( .A(n10515), .B(n10514), .Z(n10516) );
  XOR U10169 ( .A(n10517), .B(n10516), .Z(n10454) );
  XOR U10170 ( .A(n10455), .B(n10454), .Z(n10457) );
  NAND U10171 ( .A(n6139), .B(n6138), .Z(n6143) );
  NAND U10172 ( .A(n6141), .B(n6140), .Z(n6142) );
  AND U10173 ( .A(n6143), .B(n6142), .Z(n10456) );
  XOR U10174 ( .A(n10457), .B(n10456), .Z(n10503) );
  NAND U10175 ( .A(n6145), .B(n6144), .Z(n6149) );
  NAND U10176 ( .A(n6147), .B(n6146), .Z(n6148) );
  AND U10177 ( .A(n6149), .B(n6148), .Z(n9247) );
  NANDN U10178 ( .A(n6151), .B(n6150), .Z(n6155) );
  NANDN U10179 ( .A(n6153), .B(n6152), .Z(n6154) );
  AND U10180 ( .A(n6155), .B(n6154), .Z(n9132) );
  NANDN U10181 ( .A(n6157), .B(n6156), .Z(n6161) );
  NANDN U10182 ( .A(n6159), .B(n6158), .Z(n6160) );
  AND U10183 ( .A(n6161), .B(n6160), .Z(n9130) );
  NANDN U10184 ( .A(n6163), .B(n6162), .Z(n6167) );
  NANDN U10185 ( .A(n6165), .B(n6164), .Z(n6166) );
  NAND U10186 ( .A(n6167), .B(n6166), .Z(n9131) );
  XOR U10187 ( .A(n9130), .B(n9131), .Z(n9133) );
  XOR U10188 ( .A(n9132), .B(n9133), .Z(n9245) );
  NAND U10189 ( .A(n6169), .B(n6168), .Z(n6173) );
  NAND U10190 ( .A(n6171), .B(n6170), .Z(n6172) );
  NAND U10191 ( .A(n6173), .B(n6172), .Z(n9244) );
  XOR U10192 ( .A(n9245), .B(n9244), .Z(n9246) );
  XNOR U10193 ( .A(n9247), .B(n9246), .Z(n10502) );
  XOR U10194 ( .A(n10503), .B(n10502), .Z(n10504) );
  XOR U10195 ( .A(n10505), .B(n10504), .Z(n9802) );
  XNOR U10196 ( .A(n9803), .B(n9802), .Z(n9235) );
  NAND U10197 ( .A(n6175), .B(n6174), .Z(n6179) );
  NAND U10198 ( .A(n6177), .B(n6176), .Z(n6178) );
  AND U10199 ( .A(n6179), .B(n6178), .Z(n9107) );
  NANDN U10200 ( .A(n6181), .B(n6180), .Z(n6185) );
  NANDN U10201 ( .A(n6183), .B(n6182), .Z(n6184) );
  AND U10202 ( .A(n6185), .B(n6184), .Z(n9096) );
  NANDN U10203 ( .A(n6187), .B(n6186), .Z(n6191) );
  NANDN U10204 ( .A(n6189), .B(n6188), .Z(n6190) );
  AND U10205 ( .A(n6191), .B(n6190), .Z(n9094) );
  NANDN U10206 ( .A(n6193), .B(n6192), .Z(n6197) );
  OR U10207 ( .A(n6195), .B(n6194), .Z(n6196) );
  AND U10208 ( .A(n6197), .B(n6196), .Z(n10534) );
  NANDN U10209 ( .A(n6199), .B(n6198), .Z(n6203) );
  NANDN U10210 ( .A(n6201), .B(n6200), .Z(n6202) );
  AND U10211 ( .A(n6203), .B(n6202), .Z(n10533) );
  NANDN U10212 ( .A(n6205), .B(n6204), .Z(n6209) );
  NANDN U10213 ( .A(n6207), .B(n6206), .Z(n6208) );
  AND U10214 ( .A(n6209), .B(n6208), .Z(n10532) );
  XOR U10215 ( .A(n10533), .B(n10532), .Z(n10535) );
  XOR U10216 ( .A(n10534), .B(n10535), .Z(n9095) );
  XOR U10217 ( .A(n9094), .B(n9095), .Z(n9097) );
  XNOR U10218 ( .A(n9096), .B(n9097), .Z(n9106) );
  NANDN U10219 ( .A(n6211), .B(n6210), .Z(n6215) );
  NANDN U10220 ( .A(n6213), .B(n6212), .Z(n6214) );
  AND U10221 ( .A(n6215), .B(n6214), .Z(n9120) );
  NANDN U10222 ( .A(n6217), .B(n6216), .Z(n6221) );
  NAND U10223 ( .A(n6219), .B(n6218), .Z(n6220) );
  AND U10224 ( .A(n6221), .B(n6220), .Z(n9118) );
  NANDN U10225 ( .A(n6223), .B(n6222), .Z(n6227) );
  OR U10226 ( .A(n6225), .B(n6224), .Z(n6226) );
  AND U10227 ( .A(n6227), .B(n6226), .Z(n10528) );
  NANDN U10228 ( .A(n6229), .B(n6228), .Z(n6233) );
  OR U10229 ( .A(n6231), .B(n6230), .Z(n6232) );
  AND U10230 ( .A(n6233), .B(n6232), .Z(n10526) );
  NANDN U10231 ( .A(n6235), .B(n6234), .Z(n6239) );
  NANDN U10232 ( .A(n6237), .B(n6236), .Z(n6238) );
  NAND U10233 ( .A(n6239), .B(n6238), .Z(n10527) );
  XOR U10234 ( .A(n10526), .B(n10527), .Z(n10529) );
  XOR U10235 ( .A(n10528), .B(n10529), .Z(n9119) );
  XOR U10236 ( .A(n9118), .B(n9119), .Z(n9121) );
  XNOR U10237 ( .A(n9120), .B(n9121), .Z(n9108) );
  XNOR U10238 ( .A(n9109), .B(n9108), .Z(n9233) );
  NANDN U10239 ( .A(n6241), .B(n6240), .Z(n6245) );
  OR U10240 ( .A(n6243), .B(n6242), .Z(n6244) );
  AND U10241 ( .A(n6245), .B(n6244), .Z(n9402) );
  NANDN U10242 ( .A(n6247), .B(n6246), .Z(n6251) );
  OR U10243 ( .A(n6249), .B(n6248), .Z(n6250) );
  AND U10244 ( .A(n6251), .B(n6250), .Z(n9399) );
  NANDN U10245 ( .A(n6253), .B(n6252), .Z(n6257) );
  OR U10246 ( .A(n6255), .B(n6254), .Z(n6256) );
  NAND U10247 ( .A(n6257), .B(n6256), .Z(n9400) );
  XNOR U10248 ( .A(n9399), .B(n9400), .Z(n9401) );
  XNOR U10249 ( .A(n9402), .B(n9401), .Z(n9223) );
  NANDN U10250 ( .A(n6259), .B(n6258), .Z(n6263) );
  OR U10251 ( .A(n6261), .B(n6260), .Z(n6262) );
  AND U10252 ( .A(n6263), .B(n6262), .Z(n9408) );
  NANDN U10253 ( .A(n6265), .B(n6264), .Z(n6269) );
  NANDN U10254 ( .A(n6267), .B(n6266), .Z(n6268) );
  AND U10255 ( .A(n6269), .B(n6268), .Z(n9405) );
  NANDN U10256 ( .A(n6271), .B(n6270), .Z(n6275) );
  OR U10257 ( .A(n6273), .B(n6272), .Z(n6274) );
  NAND U10258 ( .A(n6275), .B(n6274), .Z(n9406) );
  XNOR U10259 ( .A(n9405), .B(n9406), .Z(n9407) );
  XNOR U10260 ( .A(n9408), .B(n9407), .Z(n9221) );
  NAND U10261 ( .A(n6277), .B(n6276), .Z(n6281) );
  NAND U10262 ( .A(n6279), .B(n6278), .Z(n6280) );
  AND U10263 ( .A(n6281), .B(n6280), .Z(n9220) );
  XOR U10264 ( .A(n9221), .B(n9220), .Z(n9222) );
  XOR U10265 ( .A(n9223), .B(n9222), .Z(n10113) );
  NANDN U10266 ( .A(n6283), .B(n6282), .Z(n6287) );
  NAND U10267 ( .A(n6285), .B(n6284), .Z(n6286) );
  AND U10268 ( .A(n6287), .B(n6286), .Z(n9258) );
  NANDN U10269 ( .A(n6289), .B(n6288), .Z(n6293) );
  NAND U10270 ( .A(n6291), .B(n6290), .Z(n6292) );
  AND U10271 ( .A(n6293), .B(n6292), .Z(n9257) );
  NANDN U10272 ( .A(n6295), .B(n6294), .Z(n6299) );
  NANDN U10273 ( .A(n6297), .B(n6296), .Z(n6298) );
  AND U10274 ( .A(n6299), .B(n6298), .Z(n9256) );
  XOR U10275 ( .A(n9257), .B(n9256), .Z(n9259) );
  XOR U10276 ( .A(n9258), .B(n9259), .Z(n10545) );
  NANDN U10277 ( .A(n6301), .B(n6300), .Z(n6305) );
  NANDN U10278 ( .A(n6303), .B(n6302), .Z(n6304) );
  AND U10279 ( .A(n6305), .B(n6304), .Z(n10511) );
  NANDN U10280 ( .A(n6307), .B(n6306), .Z(n6311) );
  NANDN U10281 ( .A(n6309), .B(n6308), .Z(n6310) );
  AND U10282 ( .A(n6311), .B(n6310), .Z(n10508) );
  NANDN U10283 ( .A(n6313), .B(n6312), .Z(n6317) );
  NANDN U10284 ( .A(n6315), .B(n6314), .Z(n6316) );
  NAND U10285 ( .A(n6317), .B(n6316), .Z(n10509) );
  XNOR U10286 ( .A(n10508), .B(n10509), .Z(n10510) );
  XOR U10287 ( .A(n10511), .B(n10510), .Z(n10543) );
  NANDN U10288 ( .A(n6319), .B(n6318), .Z(n6323) );
  OR U10289 ( .A(n6321), .B(n6320), .Z(n6322) );
  AND U10290 ( .A(n6323), .B(n6322), .Z(n10349) );
  NANDN U10291 ( .A(n6325), .B(n6324), .Z(n6329) );
  NANDN U10292 ( .A(n6327), .B(n6326), .Z(n6328) );
  AND U10293 ( .A(n6329), .B(n6328), .Z(n10346) );
  NANDN U10294 ( .A(n6331), .B(n6330), .Z(n6335) );
  OR U10295 ( .A(n6333), .B(n6332), .Z(n6334) );
  NAND U10296 ( .A(n6335), .B(n6334), .Z(n10347) );
  XNOR U10297 ( .A(n10346), .B(n10347), .Z(n10348) );
  XNOR U10298 ( .A(n10349), .B(n10348), .Z(n10542) );
  XNOR U10299 ( .A(n10543), .B(n10542), .Z(n10544) );
  XNOR U10300 ( .A(n10545), .B(n10544), .Z(n10114) );
  XOR U10301 ( .A(n10113), .B(n10114), .Z(n10116) );
  NANDN U10302 ( .A(n6337), .B(n6336), .Z(n6341) );
  NAND U10303 ( .A(n6339), .B(n6338), .Z(n6340) );
  AND U10304 ( .A(n6341), .B(n6340), .Z(n9269) );
  NANDN U10305 ( .A(n6343), .B(n6342), .Z(n6347) );
  OR U10306 ( .A(n6345), .B(n6344), .Z(n6346) );
  AND U10307 ( .A(n6347), .B(n6346), .Z(n9443) );
  NAND U10308 ( .A(n6349), .B(n6348), .Z(n6353) );
  NAND U10309 ( .A(n6351), .B(n6350), .Z(n6352) );
  AND U10310 ( .A(n6353), .B(n6352), .Z(n9441) );
  NANDN U10311 ( .A(n6355), .B(n6354), .Z(n6359) );
  NAND U10312 ( .A(n6357), .B(n6356), .Z(n6358) );
  AND U10313 ( .A(n6359), .B(n6358), .Z(n9454) );
  NANDN U10314 ( .A(n6361), .B(n6360), .Z(n6365) );
  NAND U10315 ( .A(n6363), .B(n6362), .Z(n6364) );
  AND U10316 ( .A(n6365), .B(n6364), .Z(n9453) );
  NANDN U10317 ( .A(n6367), .B(n6366), .Z(n6371) );
  NAND U10318 ( .A(n6369), .B(n6368), .Z(n6370) );
  NAND U10319 ( .A(n6371), .B(n6370), .Z(n9452) );
  XOR U10320 ( .A(n9453), .B(n9452), .Z(n9455) );
  XNOR U10321 ( .A(n9454), .B(n9455), .Z(n9440) );
  XNOR U10322 ( .A(n9441), .B(n9440), .Z(n9442) );
  XNOR U10323 ( .A(n9443), .B(n9442), .Z(n9268) );
  XNOR U10324 ( .A(n9269), .B(n9268), .Z(n9271) );
  NANDN U10325 ( .A(n6373), .B(n6372), .Z(n6377) );
  NAND U10326 ( .A(n6375), .B(n6374), .Z(n6376) );
  AND U10327 ( .A(n6377), .B(n6376), .Z(n10229) );
  NANDN U10328 ( .A(n6379), .B(n6378), .Z(n6383) );
  NAND U10329 ( .A(n6381), .B(n6380), .Z(n6382) );
  AND U10330 ( .A(n6383), .B(n6382), .Z(n10228) );
  NANDN U10331 ( .A(n6385), .B(n6384), .Z(n6389) );
  NAND U10332 ( .A(n6387), .B(n6386), .Z(n6388) );
  NAND U10333 ( .A(n6389), .B(n6388), .Z(n10227) );
  XOR U10334 ( .A(n10228), .B(n10227), .Z(n10230) );
  XOR U10335 ( .A(n10229), .B(n10230), .Z(n10206) );
  NANDN U10336 ( .A(n6391), .B(n6390), .Z(n6395) );
  NANDN U10337 ( .A(n6393), .B(n6392), .Z(n6394) );
  AND U10338 ( .A(n6395), .B(n6394), .Z(n10204) );
  NANDN U10339 ( .A(n6397), .B(n6396), .Z(n6401) );
  NAND U10340 ( .A(n6399), .B(n6398), .Z(n6400) );
  AND U10341 ( .A(n6401), .B(n6400), .Z(n10199) );
  NANDN U10342 ( .A(n6403), .B(n6402), .Z(n6407) );
  NAND U10343 ( .A(n6405), .B(n6404), .Z(n6406) );
  AND U10344 ( .A(n6407), .B(n6406), .Z(n10198) );
  NANDN U10345 ( .A(n6409), .B(n6408), .Z(n6413) );
  NAND U10346 ( .A(n6411), .B(n6410), .Z(n6412) );
  NAND U10347 ( .A(n6413), .B(n6412), .Z(n10197) );
  XOR U10348 ( .A(n10198), .B(n10197), .Z(n10200) );
  XNOR U10349 ( .A(n10199), .B(n10200), .Z(n10203) );
  XNOR U10350 ( .A(n10204), .B(n10203), .Z(n10205) );
  XNOR U10351 ( .A(n10206), .B(n10205), .Z(n9270) );
  XNOR U10352 ( .A(n9271), .B(n9270), .Z(n10379) );
  NANDN U10353 ( .A(n6415), .B(n6414), .Z(n6419) );
  NANDN U10354 ( .A(n6417), .B(n6416), .Z(n6418) );
  AND U10355 ( .A(n6419), .B(n6418), .Z(n9274) );
  NANDN U10356 ( .A(n6421), .B(n6420), .Z(n6425) );
  NAND U10357 ( .A(n6423), .B(n6422), .Z(n6424) );
  AND U10358 ( .A(n6425), .B(n6424), .Z(n9473) );
  NANDN U10359 ( .A(n6427), .B(n6426), .Z(n6431) );
  OR U10360 ( .A(n6429), .B(n6428), .Z(n6430) );
  AND U10361 ( .A(n6431), .B(n6430), .Z(n9471) );
  NANDN U10362 ( .A(n6433), .B(n6432), .Z(n6437) );
  NAND U10363 ( .A(n6435), .B(n6434), .Z(n6436) );
  AND U10364 ( .A(n6437), .B(n6436), .Z(n10223) );
  NANDN U10365 ( .A(n6439), .B(n6438), .Z(n6443) );
  NAND U10366 ( .A(n6441), .B(n6440), .Z(n6442) );
  AND U10367 ( .A(n6443), .B(n6442), .Z(n10222) );
  NANDN U10368 ( .A(n6445), .B(n6444), .Z(n6449) );
  NAND U10369 ( .A(n6447), .B(n6446), .Z(n6448) );
  NAND U10370 ( .A(n6449), .B(n6448), .Z(n10221) );
  XOR U10371 ( .A(n10222), .B(n10221), .Z(n10224) );
  XNOR U10372 ( .A(n10223), .B(n10224), .Z(n9470) );
  XNOR U10373 ( .A(n9471), .B(n9470), .Z(n9472) );
  XOR U10374 ( .A(n9473), .B(n9472), .Z(n9275) );
  XNOR U10375 ( .A(n9274), .B(n9275), .Z(n9277) );
  NANDN U10376 ( .A(n6451), .B(n6450), .Z(n6455) );
  NANDN U10377 ( .A(n6453), .B(n6452), .Z(n6454) );
  AND U10378 ( .A(n6455), .B(n6454), .Z(n9833) );
  NANDN U10379 ( .A(n6457), .B(n6456), .Z(n6461) );
  NAND U10380 ( .A(n6459), .B(n6458), .Z(n6460) );
  AND U10381 ( .A(n6461), .B(n6460), .Z(n9831) );
  NANDN U10382 ( .A(n6463), .B(n6462), .Z(n6467) );
  NAND U10383 ( .A(n6465), .B(n6464), .Z(n6466) );
  NAND U10384 ( .A(n6467), .B(n6466), .Z(n9995) );
  NANDN U10385 ( .A(n6469), .B(n6468), .Z(n6473) );
  NAND U10386 ( .A(n6471), .B(n6470), .Z(n6472) );
  NAND U10387 ( .A(n6473), .B(n6472), .Z(n9994) );
  NANDN U10388 ( .A(n6475), .B(n6474), .Z(n6479) );
  NAND U10389 ( .A(n6477), .B(n6476), .Z(n6478) );
  NAND U10390 ( .A(n6479), .B(n6478), .Z(n9993) );
  XNOR U10391 ( .A(n9994), .B(n9993), .Z(n9996) );
  XOR U10392 ( .A(n9995), .B(n9996), .Z(n9830) );
  XNOR U10393 ( .A(n9831), .B(n9830), .Z(n9832) );
  XNOR U10394 ( .A(n9833), .B(n9832), .Z(n9276) );
  XNOR U10395 ( .A(n9277), .B(n9276), .Z(n10377) );
  NANDN U10396 ( .A(n6481), .B(n6480), .Z(n6485) );
  OR U10397 ( .A(n6483), .B(n6482), .Z(n6484) );
  AND U10398 ( .A(n6485), .B(n6484), .Z(n10248) );
  NANDN U10399 ( .A(n6487), .B(n6486), .Z(n6491) );
  OR U10400 ( .A(n6489), .B(n6488), .Z(n6490) );
  AND U10401 ( .A(n6491), .B(n6490), .Z(n10245) );
  NANDN U10402 ( .A(n6493), .B(n6492), .Z(n6497) );
  OR U10403 ( .A(n6495), .B(n6494), .Z(n6496) );
  NAND U10404 ( .A(n6497), .B(n6496), .Z(n10246) );
  XNOR U10405 ( .A(n10245), .B(n10246), .Z(n10247) );
  XOR U10406 ( .A(n10248), .B(n10247), .Z(n9251) );
  NANDN U10407 ( .A(n6499), .B(n6498), .Z(n6503) );
  NANDN U10408 ( .A(n6501), .B(n6500), .Z(n6502) );
  NAND U10409 ( .A(n6503), .B(n6502), .Z(n9250) );
  XNOR U10410 ( .A(n9251), .B(n9250), .Z(n9253) );
  NAND U10411 ( .A(n6505), .B(n6504), .Z(n6509) );
  NAND U10412 ( .A(n6507), .B(n6506), .Z(n6508) );
  AND U10413 ( .A(n6509), .B(n6508), .Z(n10188) );
  NANDN U10414 ( .A(n6511), .B(n6510), .Z(n6515) );
  NAND U10415 ( .A(n6513), .B(n6512), .Z(n6514) );
  AND U10416 ( .A(n6515), .B(n6514), .Z(n10186) );
  NANDN U10417 ( .A(n6517), .B(n6516), .Z(n6521) );
  NAND U10418 ( .A(n6519), .B(n6518), .Z(n6520) );
  NAND U10419 ( .A(n6521), .B(n6520), .Z(n10185) );
  XNOR U10420 ( .A(n10186), .B(n10185), .Z(n10187) );
  XOR U10421 ( .A(n10188), .B(n10187), .Z(n9436) );
  NANDN U10422 ( .A(n6523), .B(n6522), .Z(n6527) );
  NAND U10423 ( .A(n6525), .B(n6524), .Z(n6526) );
  NAND U10424 ( .A(n6527), .B(n6526), .Z(n9435) );
  NANDN U10425 ( .A(n6529), .B(n6528), .Z(n6533) );
  NAND U10426 ( .A(n6531), .B(n6530), .Z(n6532) );
  AND U10427 ( .A(n6533), .B(n6532), .Z(n9466) );
  NANDN U10428 ( .A(n6535), .B(n6534), .Z(n6539) );
  NAND U10429 ( .A(n6537), .B(n6536), .Z(n6538) );
  AND U10430 ( .A(n6539), .B(n6538), .Z(n9465) );
  NANDN U10431 ( .A(n6541), .B(n6540), .Z(n6545) );
  NAND U10432 ( .A(n6543), .B(n6542), .Z(n6544) );
  NAND U10433 ( .A(n6545), .B(n6544), .Z(n9464) );
  XOR U10434 ( .A(n9465), .B(n9464), .Z(n9467) );
  XNOR U10435 ( .A(n9466), .B(n9467), .Z(n9434) );
  XOR U10436 ( .A(n9435), .B(n9434), .Z(n9437) );
  XOR U10437 ( .A(n9436), .B(n9437), .Z(n9252) );
  XNOR U10438 ( .A(n9253), .B(n9252), .Z(n10376) );
  XOR U10439 ( .A(n10377), .B(n10376), .Z(n10378) );
  XOR U10440 ( .A(n10379), .B(n10378), .Z(n10115) );
  XOR U10441 ( .A(n10116), .B(n10115), .Z(n9232) );
  XOR U10442 ( .A(n9233), .B(n9232), .Z(n9234) );
  XNOR U10443 ( .A(n9235), .B(n9234), .Z(n9240) );
  NANDN U10444 ( .A(n6547), .B(n6546), .Z(n6551) );
  NANDN U10445 ( .A(n6549), .B(n6548), .Z(n6550) );
  AND U10446 ( .A(n6551), .B(n6550), .Z(n9372) );
  NANDN U10447 ( .A(n6553), .B(n6552), .Z(n6557) );
  NAND U10448 ( .A(n6555), .B(n6554), .Z(n6556) );
  AND U10449 ( .A(n6557), .B(n6556), .Z(n9370) );
  NAND U10450 ( .A(n6559), .B(n6558), .Z(n6563) );
  NAND U10451 ( .A(n6561), .B(n6560), .Z(n6562) );
  NAND U10452 ( .A(n6563), .B(n6562), .Z(n10451) );
  NAND U10453 ( .A(n6565), .B(n6564), .Z(n6569) );
  NAND U10454 ( .A(n6567), .B(n6566), .Z(n6568) );
  AND U10455 ( .A(n6569), .B(n6568), .Z(n10448) );
  NANDN U10456 ( .A(n6571), .B(n6570), .Z(n6575) );
  OR U10457 ( .A(n6573), .B(n6572), .Z(n6574) );
  AND U10458 ( .A(n6575), .B(n6574), .Z(n9749) );
  NANDN U10459 ( .A(n6577), .B(n6576), .Z(n6581) );
  NANDN U10460 ( .A(n6579), .B(n6578), .Z(n6580) );
  AND U10461 ( .A(n6581), .B(n6580), .Z(n9747) );
  NANDN U10462 ( .A(n6583), .B(n6582), .Z(n6587) );
  NAND U10463 ( .A(n6585), .B(n6584), .Z(n6586) );
  NAND U10464 ( .A(n6587), .B(n6586), .Z(n10121) );
  NAND U10465 ( .A(n6589), .B(n6588), .Z(n6593) );
  NAND U10466 ( .A(n6591), .B(n6590), .Z(n6592) );
  NAND U10467 ( .A(n6593), .B(n6592), .Z(n10120) );
  NANDN U10468 ( .A(n6595), .B(n6594), .Z(n6599) );
  NAND U10469 ( .A(n6597), .B(n6596), .Z(n6598) );
  NAND U10470 ( .A(n6599), .B(n6598), .Z(n10119) );
  XNOR U10471 ( .A(n10120), .B(n10119), .Z(n10122) );
  XOR U10472 ( .A(n10121), .B(n10122), .Z(n9746) );
  XNOR U10473 ( .A(n9747), .B(n9746), .Z(n9748) );
  XNOR U10474 ( .A(n9749), .B(n9748), .Z(n9082) );
  NANDN U10475 ( .A(n6601), .B(n6600), .Z(n6605) );
  OR U10476 ( .A(n6603), .B(n6602), .Z(n6604) );
  AND U10477 ( .A(n6605), .B(n6604), .Z(n9683) );
  NANDN U10478 ( .A(n6607), .B(n6606), .Z(n6611) );
  OR U10479 ( .A(n6609), .B(n6608), .Z(n6610) );
  AND U10480 ( .A(n6611), .B(n6610), .Z(n9681) );
  NANDN U10481 ( .A(n6613), .B(n6612), .Z(n6617) );
  NAND U10482 ( .A(n6615), .B(n6614), .Z(n6616) );
  AND U10483 ( .A(n6617), .B(n6616), .Z(n9168) );
  NAND U10484 ( .A(n6619), .B(n6618), .Z(n6623) );
  NAND U10485 ( .A(n6621), .B(n6620), .Z(n6622) );
  AND U10486 ( .A(n6623), .B(n6622), .Z(n9167) );
  NANDN U10487 ( .A(n6625), .B(n6624), .Z(n6629) );
  NAND U10488 ( .A(n6627), .B(n6626), .Z(n6628) );
  NAND U10489 ( .A(n6629), .B(n6628), .Z(n9166) );
  XOR U10490 ( .A(n9167), .B(n9166), .Z(n9169) );
  XNOR U10491 ( .A(n9168), .B(n9169), .Z(n9680) );
  XNOR U10492 ( .A(n9681), .B(n9680), .Z(n9682) );
  XOR U10493 ( .A(n9683), .B(n9682), .Z(n9083) );
  XNOR U10494 ( .A(n9082), .B(n9083), .Z(n9084) );
  NANDN U10495 ( .A(n6631), .B(n6630), .Z(n6635) );
  OR U10496 ( .A(n6633), .B(n6632), .Z(n6634) );
  AND U10497 ( .A(n6635), .B(n6634), .Z(n9497) );
  NANDN U10498 ( .A(n6637), .B(n6636), .Z(n6641) );
  NANDN U10499 ( .A(n6639), .B(n6638), .Z(n6640) );
  AND U10500 ( .A(n6641), .B(n6640), .Z(n9495) );
  NANDN U10501 ( .A(n6643), .B(n6642), .Z(n6647) );
  NAND U10502 ( .A(n6645), .B(n6644), .Z(n6646) );
  NAND U10503 ( .A(n6647), .B(n6646), .Z(n10133) );
  NANDN U10504 ( .A(n6649), .B(n6648), .Z(n6653) );
  NAND U10505 ( .A(n6651), .B(n6650), .Z(n6652) );
  NAND U10506 ( .A(n6653), .B(n6652), .Z(n10132) );
  NANDN U10507 ( .A(n6655), .B(n6654), .Z(n6659) );
  NAND U10508 ( .A(n6657), .B(n6656), .Z(n6658) );
  NAND U10509 ( .A(n6659), .B(n6658), .Z(n10131) );
  XNOR U10510 ( .A(n10132), .B(n10131), .Z(n10134) );
  XOR U10511 ( .A(n10133), .B(n10134), .Z(n9494) );
  XNOR U10512 ( .A(n9495), .B(n9494), .Z(n9496) );
  XOR U10513 ( .A(n9497), .B(n9496), .Z(n9085) );
  XNOR U10514 ( .A(n9084), .B(n9085), .Z(n10449) );
  XOR U10515 ( .A(n10448), .B(n10449), .Z(n10450) );
  XOR U10516 ( .A(n10451), .B(n10450), .Z(n9369) );
  NAND U10517 ( .A(n6661), .B(n6660), .Z(n6665) );
  NAND U10518 ( .A(n6663), .B(n6662), .Z(n6664) );
  AND U10519 ( .A(n6665), .B(n6664), .Z(n10443) );
  XOR U10520 ( .A(n10442), .B(n10443), .Z(n10445) );
  NANDN U10521 ( .A(n6667), .B(n6666), .Z(n6671) );
  NANDN U10522 ( .A(n6669), .B(n6668), .Z(n6670) );
  AND U10523 ( .A(n6671), .B(n6670), .Z(n9537) );
  NANDN U10524 ( .A(n6673), .B(n6672), .Z(n6677) );
  NANDN U10525 ( .A(n6675), .B(n6674), .Z(n6676) );
  AND U10526 ( .A(n6677), .B(n6676), .Z(n9858) );
  NANDN U10527 ( .A(n6679), .B(n6678), .Z(n6683) );
  NANDN U10528 ( .A(n6681), .B(n6680), .Z(n6682) );
  AND U10529 ( .A(n6683), .B(n6682), .Z(n9856) );
  NAND U10530 ( .A(n6685), .B(n6684), .Z(n6689) );
  NAND U10531 ( .A(n6687), .B(n6686), .Z(n6688) );
  NAND U10532 ( .A(n6689), .B(n6688), .Z(n9881) );
  NAND U10533 ( .A(n6691), .B(n6690), .Z(n6695) );
  NAND U10534 ( .A(n6693), .B(n6692), .Z(n6694) );
  NAND U10535 ( .A(n6695), .B(n6694), .Z(n9880) );
  NANDN U10536 ( .A(n6697), .B(n6696), .Z(n6701) );
  NAND U10537 ( .A(n6699), .B(n6698), .Z(n6700) );
  NAND U10538 ( .A(n6701), .B(n6700), .Z(n9879) );
  XNOR U10539 ( .A(n9880), .B(n9879), .Z(n9882) );
  XOR U10540 ( .A(n9881), .B(n9882), .Z(n9855) );
  XNOR U10541 ( .A(n9856), .B(n9855), .Z(n9857) );
  XNOR U10542 ( .A(n9858), .B(n9857), .Z(n9335) );
  NANDN U10543 ( .A(n6703), .B(n6702), .Z(n6707) );
  NAND U10544 ( .A(n6705), .B(n6704), .Z(n6706) );
  AND U10545 ( .A(n6707), .B(n6706), .Z(n9199) );
  NANDN U10546 ( .A(n6709), .B(n6708), .Z(n6713) );
  NANDN U10547 ( .A(n6711), .B(n6710), .Z(n6712) );
  AND U10548 ( .A(n6713), .B(n6712), .Z(n9197) );
  NANDN U10549 ( .A(n6715), .B(n6714), .Z(n6719) );
  NAND U10550 ( .A(n6717), .B(n6716), .Z(n6718) );
  AND U10551 ( .A(n6719), .B(n6718), .Z(n9162) );
  NANDN U10552 ( .A(n6721), .B(n6720), .Z(n6725) );
  NAND U10553 ( .A(n6723), .B(n6722), .Z(n6724) );
  AND U10554 ( .A(n6725), .B(n6724), .Z(n9161) );
  NANDN U10555 ( .A(n6727), .B(n6726), .Z(n6731) );
  NAND U10556 ( .A(n6729), .B(n6728), .Z(n6730) );
  NAND U10557 ( .A(n6731), .B(n6730), .Z(n9160) );
  XOR U10558 ( .A(n9161), .B(n9160), .Z(n9163) );
  XNOR U10559 ( .A(n9162), .B(n9163), .Z(n9196) );
  XNOR U10560 ( .A(n9197), .B(n9196), .Z(n9198) );
  XOR U10561 ( .A(n9199), .B(n9198), .Z(n9336) );
  XNOR U10562 ( .A(n9335), .B(n9336), .Z(n9337) );
  NANDN U10563 ( .A(n6733), .B(n6732), .Z(n6737) );
  NANDN U10564 ( .A(n6735), .B(n6734), .Z(n6736) );
  AND U10565 ( .A(n6737), .B(n6736), .Z(n9552) );
  NANDN U10566 ( .A(n6739), .B(n6738), .Z(n6743) );
  OR U10567 ( .A(n6741), .B(n6740), .Z(n6742) );
  AND U10568 ( .A(n6743), .B(n6742), .Z(n9550) );
  NANDN U10569 ( .A(n6745), .B(n6744), .Z(n6749) );
  NAND U10570 ( .A(n6747), .B(n6746), .Z(n6748) );
  AND U10571 ( .A(n6749), .B(n6748), .Z(n10103) );
  NANDN U10572 ( .A(n6751), .B(n6750), .Z(n6755) );
  NAND U10573 ( .A(n6753), .B(n6752), .Z(n6754) );
  AND U10574 ( .A(n6755), .B(n6754), .Z(n10102) );
  NAND U10575 ( .A(n6757), .B(n6756), .Z(n6761) );
  NAND U10576 ( .A(n6759), .B(n6758), .Z(n6760) );
  NAND U10577 ( .A(n6761), .B(n6760), .Z(n10101) );
  XOR U10578 ( .A(n10102), .B(n10101), .Z(n10104) );
  XNOR U10579 ( .A(n10103), .B(n10104), .Z(n9549) );
  XNOR U10580 ( .A(n9550), .B(n9549), .Z(n9551) );
  XOR U10581 ( .A(n9552), .B(n9551), .Z(n9338) );
  XOR U10582 ( .A(n9337), .B(n9338), .Z(n9538) );
  XNOR U10583 ( .A(n9537), .B(n9538), .Z(n9540) );
  NAND U10584 ( .A(n6763), .B(n6762), .Z(n6767) );
  NAND U10585 ( .A(n6765), .B(n6764), .Z(n6766) );
  NAND U10586 ( .A(n6767), .B(n6766), .Z(n9544) );
  NANDN U10587 ( .A(n6769), .B(n6768), .Z(n6773) );
  NAND U10588 ( .A(n6771), .B(n6770), .Z(n6772) );
  AND U10589 ( .A(n6773), .B(n6772), .Z(n9899) );
  NANDN U10590 ( .A(n6775), .B(n6774), .Z(n6779) );
  NAND U10591 ( .A(n6777), .B(n6776), .Z(n6778) );
  AND U10592 ( .A(n6779), .B(n6778), .Z(n9898) );
  NANDN U10593 ( .A(n6781), .B(n6780), .Z(n6785) );
  NAND U10594 ( .A(n6783), .B(n6782), .Z(n6784) );
  NAND U10595 ( .A(n6785), .B(n6784), .Z(n9897) );
  XOR U10596 ( .A(n9898), .B(n9897), .Z(n9900) );
  XNOR U10597 ( .A(n9899), .B(n9900), .Z(n9543) );
  XOR U10598 ( .A(n9544), .B(n9543), .Z(n9546) );
  NAND U10599 ( .A(n6787), .B(n6786), .Z(n6791) );
  NAND U10600 ( .A(n6789), .B(n6788), .Z(n6790) );
  NAND U10601 ( .A(n6791), .B(n6790), .Z(n9545) );
  XOR U10602 ( .A(n9546), .B(n9545), .Z(n9299) );
  NANDN U10603 ( .A(n6793), .B(n6792), .Z(n6797) );
  NAND U10604 ( .A(n6795), .B(n6794), .Z(n6796) );
  NAND U10605 ( .A(n6797), .B(n6796), .Z(n10109) );
  NANDN U10606 ( .A(n6799), .B(n6798), .Z(n6803) );
  NAND U10607 ( .A(n6801), .B(n6800), .Z(n6802) );
  NAND U10608 ( .A(n6803), .B(n6802), .Z(n10108) );
  NANDN U10609 ( .A(n6805), .B(n6804), .Z(n6809) );
  NAND U10610 ( .A(n6807), .B(n6806), .Z(n6808) );
  NAND U10611 ( .A(n6809), .B(n6808), .Z(n10107) );
  XOR U10612 ( .A(n10108), .B(n10107), .Z(n10110) );
  XNOR U10613 ( .A(n10109), .B(n10110), .Z(n10297) );
  NANDN U10614 ( .A(n6811), .B(n6810), .Z(n6815) );
  NANDN U10615 ( .A(n6813), .B(n6812), .Z(n6814) );
  AND U10616 ( .A(n6815), .B(n6814), .Z(n10295) );
  NANDN U10617 ( .A(n6817), .B(n6816), .Z(n6821) );
  NAND U10618 ( .A(n6819), .B(n6818), .Z(n6820) );
  NAND U10619 ( .A(n6821), .B(n6820), .Z(n10254) );
  NAND U10620 ( .A(n6823), .B(n6822), .Z(n6827) );
  NAND U10621 ( .A(n6825), .B(n6824), .Z(n6826) );
  NAND U10622 ( .A(n6827), .B(n6826), .Z(n10253) );
  NANDN U10623 ( .A(n6829), .B(n6828), .Z(n6833) );
  NAND U10624 ( .A(n6831), .B(n6830), .Z(n6832) );
  NAND U10625 ( .A(n6833), .B(n6832), .Z(n10252) );
  XNOR U10626 ( .A(n10253), .B(n10252), .Z(n10255) );
  XOR U10627 ( .A(n10254), .B(n10255), .Z(n10294) );
  XNOR U10628 ( .A(n10295), .B(n10294), .Z(n10296) );
  XOR U10629 ( .A(n10297), .B(n10296), .Z(n9298) );
  XOR U10630 ( .A(n9299), .B(n9298), .Z(n9300) );
  NANDN U10631 ( .A(n6835), .B(n6834), .Z(n6839) );
  NAND U10632 ( .A(n6837), .B(n6836), .Z(n6838) );
  AND U10633 ( .A(n6839), .B(n6838), .Z(n9935) );
  NANDN U10634 ( .A(n6841), .B(n6840), .Z(n6845) );
  NAND U10635 ( .A(n6843), .B(n6842), .Z(n6844) );
  AND U10636 ( .A(n6845), .B(n6844), .Z(n9934) );
  NANDN U10637 ( .A(n6847), .B(n6846), .Z(n6851) );
  NAND U10638 ( .A(n6849), .B(n6848), .Z(n6850) );
  NAND U10639 ( .A(n6851), .B(n6850), .Z(n9933) );
  XOR U10640 ( .A(n9934), .B(n9933), .Z(n9936) );
  XOR U10641 ( .A(n9935), .B(n9936), .Z(n9576) );
  NANDN U10642 ( .A(n6853), .B(n6852), .Z(n6857) );
  NAND U10643 ( .A(n6855), .B(n6854), .Z(n6856) );
  NAND U10644 ( .A(n6857), .B(n6856), .Z(n10272) );
  NANDN U10645 ( .A(n6859), .B(n6858), .Z(n6863) );
  NAND U10646 ( .A(n6861), .B(n6860), .Z(n6862) );
  NAND U10647 ( .A(n6863), .B(n6862), .Z(n10271) );
  NANDN U10648 ( .A(n6865), .B(n6864), .Z(n6869) );
  NAND U10649 ( .A(n6867), .B(n6866), .Z(n6868) );
  NAND U10650 ( .A(n6869), .B(n6868), .Z(n10270) );
  XOR U10651 ( .A(n10271), .B(n10270), .Z(n10273) );
  XNOR U10652 ( .A(n10272), .B(n10273), .Z(n9574) );
  NAND U10653 ( .A(n6871), .B(n6870), .Z(n6875) );
  NAND U10654 ( .A(n6873), .B(n6872), .Z(n6874) );
  AND U10655 ( .A(n6875), .B(n6874), .Z(n10085) );
  NANDN U10656 ( .A(n6877), .B(n6876), .Z(n6881) );
  NAND U10657 ( .A(n6879), .B(n6878), .Z(n6880) );
  AND U10658 ( .A(n6881), .B(n6880), .Z(n10084) );
  NANDN U10659 ( .A(n6883), .B(n6882), .Z(n6887) );
  NAND U10660 ( .A(n6885), .B(n6884), .Z(n6886) );
  NAND U10661 ( .A(n6887), .B(n6886), .Z(n10083) );
  XOR U10662 ( .A(n10084), .B(n10083), .Z(n10086) );
  XNOR U10663 ( .A(n10085), .B(n10086), .Z(n9573) );
  XOR U10664 ( .A(n9574), .B(n9573), .Z(n9575) );
  XOR U10665 ( .A(n9576), .B(n9575), .Z(n9301) );
  XNOR U10666 ( .A(n9300), .B(n9301), .Z(n9539) );
  XOR U10667 ( .A(n9540), .B(n9539), .Z(n9378) );
  NAND U10668 ( .A(n6889), .B(n6888), .Z(n6893) );
  NAND U10669 ( .A(n6891), .B(n6890), .Z(n6892) );
  NAND U10670 ( .A(n6893), .B(n6892), .Z(n10343) );
  NAND U10671 ( .A(n6895), .B(n6894), .Z(n6899) );
  NAND U10672 ( .A(n6897), .B(n6896), .Z(n6898) );
  NAND U10673 ( .A(n6899), .B(n6898), .Z(n10341) );
  NANDN U10674 ( .A(n6905), .B(n6904), .Z(n6909) );
  NANDN U10675 ( .A(n6907), .B(n6906), .Z(n6908) );
  AND U10676 ( .A(n6909), .B(n6908), .Z(n9719) );
  NANDN U10677 ( .A(n6911), .B(n6910), .Z(n6915) );
  NAND U10678 ( .A(n6913), .B(n6912), .Z(n6914) );
  AND U10679 ( .A(n6915), .B(n6914), .Z(n9717) );
  NANDN U10680 ( .A(n6917), .B(n6916), .Z(n6921) );
  NAND U10681 ( .A(n6919), .B(n6918), .Z(n6920) );
  AND U10682 ( .A(n6921), .B(n6920), .Z(n9953) );
  NANDN U10683 ( .A(n6923), .B(n6922), .Z(n6927) );
  NAND U10684 ( .A(n6925), .B(n6924), .Z(n6926) );
  AND U10685 ( .A(n6927), .B(n6926), .Z(n9952) );
  NANDN U10686 ( .A(n6929), .B(n6928), .Z(n6933) );
  NAND U10687 ( .A(n6931), .B(n6930), .Z(n6932) );
  NAND U10688 ( .A(n6933), .B(n6932), .Z(n9951) );
  XOR U10689 ( .A(n9952), .B(n9951), .Z(n9954) );
  XNOR U10690 ( .A(n9953), .B(n9954), .Z(n9716) );
  XNOR U10691 ( .A(n9717), .B(n9716), .Z(n9718) );
  XNOR U10692 ( .A(n9719), .B(n9718), .Z(n9320) );
  XNOR U10693 ( .A(n9321), .B(n9320), .Z(n9322) );
  NANDN U10694 ( .A(n6935), .B(n6934), .Z(n6939) );
  NANDN U10695 ( .A(n6937), .B(n6936), .Z(n6938) );
  AND U10696 ( .A(n6939), .B(n6938), .Z(n10481) );
  NANDN U10697 ( .A(n6941), .B(n6940), .Z(n6945) );
  NANDN U10698 ( .A(n6943), .B(n6942), .Z(n6944) );
  AND U10699 ( .A(n6945), .B(n6944), .Z(n10479) );
  NANDN U10700 ( .A(n6947), .B(n6946), .Z(n6951) );
  NANDN U10701 ( .A(n6949), .B(n6948), .Z(n6950) );
  NAND U10702 ( .A(n6951), .B(n6950), .Z(n10478) );
  XNOR U10703 ( .A(n10479), .B(n10478), .Z(n10480) );
  XOR U10704 ( .A(n10481), .B(n10480), .Z(n9323) );
  XNOR U10705 ( .A(n9322), .B(n9323), .Z(n10340) );
  XOR U10706 ( .A(n10341), .B(n10340), .Z(n10342) );
  XNOR U10707 ( .A(n10343), .B(n10342), .Z(n9376) );
  NAND U10708 ( .A(n6953), .B(n6952), .Z(n6957) );
  NANDN U10709 ( .A(n6955), .B(n6954), .Z(n6956) );
  NAND U10710 ( .A(n6957), .B(n6956), .Z(n9375) );
  XOR U10711 ( .A(n9376), .B(n9375), .Z(n9377) );
  XNOR U10712 ( .A(n10445), .B(n10444), .Z(n9239) );
  NAND U10713 ( .A(n6959), .B(n6958), .Z(n6963) );
  NAND U10714 ( .A(n6961), .B(n6960), .Z(n6962) );
  NAND U10715 ( .A(n6963), .B(n6962), .Z(n9143) );
  NAND U10716 ( .A(n6965), .B(n6964), .Z(n6969) );
  NAND U10717 ( .A(n6967), .B(n6966), .Z(n6968) );
  NAND U10718 ( .A(n6969), .B(n6968), .Z(n9771) );
  NANDN U10719 ( .A(n6971), .B(n6970), .Z(n6975) );
  NAND U10720 ( .A(n6973), .B(n6972), .Z(n6974) );
  AND U10721 ( .A(n6975), .B(n6974), .Z(n9737) );
  NANDN U10722 ( .A(n6977), .B(n6976), .Z(n6981) );
  NANDN U10723 ( .A(n6979), .B(n6978), .Z(n6980) );
  AND U10724 ( .A(n6981), .B(n6980), .Z(n9734) );
  NANDN U10725 ( .A(n6983), .B(n6982), .Z(n6987) );
  OR U10726 ( .A(n6985), .B(n6984), .Z(n6986) );
  AND U10727 ( .A(n6987), .B(n6986), .Z(n9912) );
  NANDN U10728 ( .A(n6989), .B(n6988), .Z(n6993) );
  OR U10729 ( .A(n6991), .B(n6990), .Z(n6992) );
  AND U10730 ( .A(n6993), .B(n6992), .Z(n9910) );
  NANDN U10731 ( .A(n6995), .B(n6994), .Z(n6999) );
  OR U10732 ( .A(n6997), .B(n6996), .Z(n6998) );
  NAND U10733 ( .A(n6999), .B(n6998), .Z(n9909) );
  XNOR U10734 ( .A(n9910), .B(n9909), .Z(n9911) );
  XOR U10735 ( .A(n9912), .B(n9911), .Z(n9735) );
  XNOR U10736 ( .A(n9734), .B(n9735), .Z(n9736) );
  XNOR U10737 ( .A(n9737), .B(n9736), .Z(n9770) );
  XOR U10738 ( .A(n9771), .B(n9770), .Z(n9772) );
  NANDN U10739 ( .A(n7001), .B(n7000), .Z(n7005) );
  NANDN U10740 ( .A(n7003), .B(n7002), .Z(n7004) );
  AND U10741 ( .A(n7005), .B(n7004), .Z(n9501) );
  NANDN U10742 ( .A(n7007), .B(n7006), .Z(n7011) );
  OR U10743 ( .A(n7009), .B(n7008), .Z(n7010) );
  AND U10744 ( .A(n7011), .B(n7010), .Z(n10158) );
  NANDN U10745 ( .A(n7013), .B(n7012), .Z(n7017) );
  OR U10746 ( .A(n7015), .B(n7014), .Z(n7016) );
  AND U10747 ( .A(n7017), .B(n7016), .Z(n10156) );
  NANDN U10748 ( .A(n7019), .B(n7018), .Z(n7023) );
  NANDN U10749 ( .A(n7021), .B(n7020), .Z(n7022) );
  NAND U10750 ( .A(n7023), .B(n7022), .Z(n10155) );
  XNOR U10751 ( .A(n10156), .B(n10155), .Z(n10157) );
  XOR U10752 ( .A(n10158), .B(n10157), .Z(n9502) );
  XNOR U10753 ( .A(n9501), .B(n9502), .Z(n9503) );
  NANDN U10754 ( .A(n7025), .B(n7024), .Z(n7029) );
  NANDN U10755 ( .A(n7027), .B(n7026), .Z(n7028) );
  AND U10756 ( .A(n7029), .B(n7028), .Z(n9978) );
  NANDN U10757 ( .A(n7031), .B(n7030), .Z(n7035) );
  NAND U10758 ( .A(n7033), .B(n7032), .Z(n7034) );
  AND U10759 ( .A(n7035), .B(n7034), .Z(n9976) );
  NANDN U10760 ( .A(n7037), .B(n7036), .Z(n7041) );
  OR U10761 ( .A(n7039), .B(n7038), .Z(n7040) );
  NAND U10762 ( .A(n7041), .B(n7040), .Z(n9975) );
  XNOR U10763 ( .A(n9976), .B(n9975), .Z(n9977) );
  XOR U10764 ( .A(n9978), .B(n9977), .Z(n9504) );
  XNOR U10765 ( .A(n9503), .B(n9504), .Z(n9773) );
  XOR U10766 ( .A(n9772), .B(n9773), .Z(n9142) );
  XOR U10767 ( .A(n9143), .B(n9142), .Z(n9145) );
  NAND U10768 ( .A(n7043), .B(n7042), .Z(n7047) );
  NAND U10769 ( .A(n7045), .B(n7044), .Z(n7046) );
  AND U10770 ( .A(n7047), .B(n7046), .Z(n9144) );
  XNOR U10771 ( .A(n9145), .B(n9144), .Z(n9388) );
  NAND U10772 ( .A(n7049), .B(n7048), .Z(n7053) );
  NAND U10773 ( .A(n7051), .B(n7050), .Z(n7052) );
  AND U10774 ( .A(n7053), .B(n7052), .Z(n9387) );
  XOR U10775 ( .A(n9388), .B(n9387), .Z(n9390) );
  NANDN U10776 ( .A(n7055), .B(n7054), .Z(n7059) );
  NANDN U10777 ( .A(n7057), .B(n7056), .Z(n7058) );
  AND U10778 ( .A(n7059), .B(n7058), .Z(n9101) );
  NANDN U10779 ( .A(n7061), .B(n7060), .Z(n7065) );
  NAND U10780 ( .A(n7063), .B(n7062), .Z(n7064) );
  AND U10781 ( .A(n7065), .B(n7064), .Z(n9100) );
  XNOR U10782 ( .A(n9101), .B(n9100), .Z(n9103) );
  NANDN U10783 ( .A(n7067), .B(n7066), .Z(n7071) );
  NANDN U10784 ( .A(n7069), .B(n7068), .Z(n7070) );
  AND U10785 ( .A(n7071), .B(n7070), .Z(n10325) );
  NAND U10786 ( .A(n7073), .B(n7072), .Z(n7077) );
  NAND U10787 ( .A(n7075), .B(n7074), .Z(n7076) );
  AND U10788 ( .A(n7077), .B(n7076), .Z(n9528) );
  NAND U10789 ( .A(n7079), .B(n7078), .Z(n7083) );
  NAND U10790 ( .A(n7081), .B(n7080), .Z(n7082) );
  AND U10791 ( .A(n7083), .B(n7082), .Z(n9526) );
  NANDN U10792 ( .A(n7085), .B(n7084), .Z(n7089) );
  NAND U10793 ( .A(n7087), .B(n7086), .Z(n7088) );
  NAND U10794 ( .A(n7089), .B(n7088), .Z(n9525) );
  XNOR U10795 ( .A(n9526), .B(n9525), .Z(n9527) );
  XOR U10796 ( .A(n9528), .B(n9527), .Z(n10326) );
  XNOR U10797 ( .A(n10325), .B(n10326), .Z(n10327) );
  NANDN U10798 ( .A(n7091), .B(n7090), .Z(n7095) );
  OR U10799 ( .A(n7093), .B(n7092), .Z(n7094) );
  AND U10800 ( .A(n7095), .B(n7094), .Z(n9677) );
  NANDN U10801 ( .A(n7097), .B(n7096), .Z(n7101) );
  NANDN U10802 ( .A(n7099), .B(n7098), .Z(n7100) );
  AND U10803 ( .A(n7101), .B(n7100), .Z(n9675) );
  NANDN U10804 ( .A(n7103), .B(n7102), .Z(n7107) );
  NANDN U10805 ( .A(n7105), .B(n7104), .Z(n7106) );
  NAND U10806 ( .A(n7107), .B(n7106), .Z(n9674) );
  XNOR U10807 ( .A(n9675), .B(n9674), .Z(n9676) );
  XOR U10808 ( .A(n9677), .B(n9676), .Z(n10328) );
  XNOR U10809 ( .A(n10327), .B(n10328), .Z(n9711) );
  NANDN U10810 ( .A(n7109), .B(n7108), .Z(n7113) );
  OR U10811 ( .A(n7111), .B(n7110), .Z(n7112) );
  AND U10812 ( .A(n7113), .B(n7112), .Z(n9710) );
  XOR U10813 ( .A(n9711), .B(n9710), .Z(n9713) );
  NANDN U10814 ( .A(n7115), .B(n7114), .Z(n7119) );
  OR U10815 ( .A(n7117), .B(n7116), .Z(n7118) );
  NAND U10816 ( .A(n7119), .B(n7118), .Z(n9712) );
  XOR U10817 ( .A(n9713), .B(n9712), .Z(n9102) );
  XNOR U10818 ( .A(n9103), .B(n9102), .Z(n10439) );
  NAND U10819 ( .A(n7121), .B(n7120), .Z(n7125) );
  NAND U10820 ( .A(n7123), .B(n7122), .Z(n7124) );
  NAND U10821 ( .A(n7125), .B(n7124), .Z(n10437) );
  NANDN U10822 ( .A(n7127), .B(n7126), .Z(n7131) );
  NAND U10823 ( .A(n7129), .B(n7128), .Z(n7130) );
  AND U10824 ( .A(n7131), .B(n7130), .Z(n9585) );
  NANDN U10825 ( .A(n7133), .B(n7132), .Z(n7137) );
  NANDN U10826 ( .A(n7135), .B(n7134), .Z(n7136) );
  AND U10827 ( .A(n7137), .B(n7136), .Z(n9583) );
  NANDN U10828 ( .A(n7139), .B(n7138), .Z(n7143) );
  NAND U10829 ( .A(n7141), .B(n7140), .Z(n7142) );
  AND U10830 ( .A(n7143), .B(n7142), .Z(n9701) );
  NANDN U10831 ( .A(n7145), .B(n7144), .Z(n7149) );
  NANDN U10832 ( .A(n7147), .B(n7146), .Z(n7148) );
  AND U10833 ( .A(n7149), .B(n7148), .Z(n9699) );
  NANDN U10834 ( .A(n7151), .B(n7150), .Z(n7155) );
  NANDN U10835 ( .A(n7153), .B(n7152), .Z(n7154) );
  NAND U10836 ( .A(n7155), .B(n7154), .Z(n9698) );
  XNOR U10837 ( .A(n9699), .B(n9698), .Z(n9700) );
  XOR U10838 ( .A(n9701), .B(n9700), .Z(n9584) );
  XOR U10839 ( .A(n9583), .B(n9584), .Z(n9586) );
  XNOR U10840 ( .A(n9585), .B(n9586), .Z(n9217) );
  NANDN U10841 ( .A(n7157), .B(n7156), .Z(n7161) );
  NAND U10842 ( .A(n7159), .B(n7158), .Z(n7160) );
  AND U10843 ( .A(n7161), .B(n7160), .Z(n10217) );
  NANDN U10844 ( .A(n7163), .B(n7162), .Z(n7167) );
  NAND U10845 ( .A(n7165), .B(n7164), .Z(n7166) );
  AND U10846 ( .A(n7167), .B(n7166), .Z(n10216) );
  NANDN U10847 ( .A(n7169), .B(n7168), .Z(n7173) );
  OR U10848 ( .A(n7171), .B(n7170), .Z(n7172) );
  AND U10849 ( .A(n7173), .B(n7172), .Z(n9193) );
  NANDN U10850 ( .A(n7175), .B(n7174), .Z(n7179) );
  NAND U10851 ( .A(n7177), .B(n7176), .Z(n7178) );
  AND U10852 ( .A(n7179), .B(n7178), .Z(n9191) );
  NANDN U10853 ( .A(n7181), .B(n7180), .Z(n7185) );
  OR U10854 ( .A(n7183), .B(n7182), .Z(n7184) );
  NAND U10855 ( .A(n7185), .B(n7184), .Z(n9190) );
  XNOR U10856 ( .A(n9191), .B(n9190), .Z(n9192) );
  XNOR U10857 ( .A(n9193), .B(n9192), .Z(n10215) );
  XOR U10858 ( .A(n10216), .B(n10215), .Z(n10218) );
  XNOR U10859 ( .A(n10217), .B(n10218), .Z(n9215) );
  NANDN U10860 ( .A(n7187), .B(n7186), .Z(n7191) );
  NANDN U10861 ( .A(n7189), .B(n7188), .Z(n7190) );
  AND U10862 ( .A(n7191), .B(n7190), .Z(n10065) );
  NANDN U10863 ( .A(n7193), .B(n7192), .Z(n7197) );
  NAND U10864 ( .A(n7195), .B(n7194), .Z(n7196) );
  AND U10865 ( .A(n7197), .B(n7196), .Z(n10056) );
  NANDN U10866 ( .A(n7199), .B(n7198), .Z(n7203) );
  NAND U10867 ( .A(n7201), .B(n7200), .Z(n7202) );
  AND U10868 ( .A(n7203), .B(n7202), .Z(n10054) );
  NANDN U10869 ( .A(n7205), .B(n7204), .Z(n7209) );
  OR U10870 ( .A(n7207), .B(n7206), .Z(n7208) );
  NAND U10871 ( .A(n7209), .B(n7208), .Z(n10053) );
  XNOR U10872 ( .A(n10054), .B(n10053), .Z(n10055) );
  XOR U10873 ( .A(n10056), .B(n10055), .Z(n10066) );
  XNOR U10874 ( .A(n10065), .B(n10066), .Z(n10068) );
  NANDN U10875 ( .A(n7211), .B(n7210), .Z(n7215) );
  NANDN U10876 ( .A(n7213), .B(n7212), .Z(n7214) );
  NAND U10877 ( .A(n7215), .B(n7214), .Z(n10426) );
  NANDN U10878 ( .A(n7217), .B(n7216), .Z(n7221) );
  NAND U10879 ( .A(n7219), .B(n7218), .Z(n7220) );
  NAND U10880 ( .A(n7221), .B(n7220), .Z(n10425) );
  NANDN U10881 ( .A(n7223), .B(n7222), .Z(n7227) );
  NANDN U10882 ( .A(n7225), .B(n7224), .Z(n7226) );
  NAND U10883 ( .A(n7227), .B(n7226), .Z(n10424) );
  XOR U10884 ( .A(n10425), .B(n10424), .Z(n10427) );
  XOR U10885 ( .A(n10426), .B(n10427), .Z(n10067) );
  XNOR U10886 ( .A(n10068), .B(n10067), .Z(n9214) );
  XOR U10887 ( .A(n9215), .B(n9214), .Z(n9216) );
  XOR U10888 ( .A(n9217), .B(n9216), .Z(n10436) );
  XOR U10889 ( .A(n10437), .B(n10436), .Z(n10438) );
  XOR U10890 ( .A(n10439), .B(n10438), .Z(n9389) );
  XNOR U10891 ( .A(n9390), .B(n9389), .Z(n9238) );
  XOR U10892 ( .A(n9239), .B(n9238), .Z(n9241) );
  XOR U10893 ( .A(n9240), .B(n9241), .Z(n10333) );
  NANDN U10894 ( .A(n7229), .B(n7228), .Z(n7233) );
  NAND U10895 ( .A(n7231), .B(n7230), .Z(n7232) );
  NAND U10896 ( .A(n7233), .B(n7232), .Z(n10331) );
  NAND U10897 ( .A(n7235), .B(n7234), .Z(n7239) );
  NAND U10898 ( .A(n7237), .B(n7236), .Z(n7238) );
  AND U10899 ( .A(n7239), .B(n7238), .Z(n10334) );
  NAND U10900 ( .A(n7241), .B(n7240), .Z(n7245) );
  NAND U10901 ( .A(n7243), .B(n7242), .Z(n7244) );
  AND U10902 ( .A(n7245), .B(n7244), .Z(n10335) );
  XOR U10903 ( .A(n10334), .B(n10335), .Z(n10337) );
  NAND U10904 ( .A(n7247), .B(n7246), .Z(n7251) );
  NAND U10905 ( .A(n7249), .B(n7248), .Z(n7250) );
  AND U10906 ( .A(n7251), .B(n7250), .Z(n9067) );
  NAND U10907 ( .A(n7253), .B(n7252), .Z(n7257) );
  NAND U10908 ( .A(n7255), .B(n7254), .Z(n7256) );
  AND U10909 ( .A(n7257), .B(n7256), .Z(n9065) );
  NAND U10910 ( .A(n7259), .B(n7258), .Z(n7263) );
  NAND U10911 ( .A(n7261), .B(n7260), .Z(n7262) );
  NAND U10912 ( .A(n7263), .B(n7262), .Z(n9229) );
  NAND U10913 ( .A(n7265), .B(n7264), .Z(n7269) );
  NAND U10914 ( .A(n7267), .B(n7266), .Z(n7268) );
  AND U10915 ( .A(n7269), .B(n7268), .Z(n9966) );
  NAND U10916 ( .A(n7271), .B(n7270), .Z(n7275) );
  NAND U10917 ( .A(n7273), .B(n7272), .Z(n7274) );
  AND U10918 ( .A(n7275), .B(n7274), .Z(n9963) );
  NAND U10919 ( .A(n7277), .B(n7276), .Z(n7281) );
  NANDN U10920 ( .A(n7279), .B(n7278), .Z(n7280) );
  AND U10921 ( .A(n7281), .B(n7280), .Z(n9964) );
  XOR U10922 ( .A(n9963), .B(n9964), .Z(n9965) );
  XNOR U10923 ( .A(n9966), .B(n9965), .Z(n9227) );
  NANDN U10924 ( .A(n7283), .B(n7282), .Z(n7287) );
  OR U10925 ( .A(n7285), .B(n7284), .Z(n7286) );
  AND U10926 ( .A(n7287), .B(n7286), .Z(n9695) );
  NANDN U10927 ( .A(n7289), .B(n7288), .Z(n7293) );
  NAND U10928 ( .A(n7291), .B(n7290), .Z(n7292) );
  AND U10929 ( .A(n7293), .B(n7292), .Z(n9693) );
  NANDN U10930 ( .A(n7295), .B(n7294), .Z(n7299) );
  OR U10931 ( .A(n7297), .B(n7296), .Z(n7298) );
  NAND U10932 ( .A(n7299), .B(n7298), .Z(n9692) );
  XNOR U10933 ( .A(n9693), .B(n9692), .Z(n9694) );
  XNOR U10934 ( .A(n9695), .B(n9694), .Z(n9446) );
  NANDN U10935 ( .A(n7301), .B(n7300), .Z(n7305) );
  NAND U10936 ( .A(n7303), .B(n7302), .Z(n7304) );
  AND U10937 ( .A(n7305), .B(n7304), .Z(n10367) );
  NANDN U10938 ( .A(n7307), .B(n7306), .Z(n7311) );
  NAND U10939 ( .A(n7309), .B(n7308), .Z(n7310) );
  AND U10940 ( .A(n7311), .B(n7310), .Z(n10365) );
  NANDN U10941 ( .A(n7313), .B(n7312), .Z(n7317) );
  OR U10942 ( .A(n7315), .B(n7314), .Z(n7316) );
  NAND U10943 ( .A(n7317), .B(n7316), .Z(n10364) );
  XNOR U10944 ( .A(n10365), .B(n10364), .Z(n10366) );
  XOR U10945 ( .A(n10367), .B(n10366), .Z(n9447) );
  XNOR U10946 ( .A(n9446), .B(n9447), .Z(n9449) );
  NANDN U10947 ( .A(n7319), .B(n7318), .Z(n7323) );
  NANDN U10948 ( .A(n7321), .B(n7320), .Z(n7322) );
  AND U10949 ( .A(n7323), .B(n7322), .Z(n10373) );
  NANDN U10950 ( .A(n7325), .B(n7324), .Z(n7329) );
  OR U10951 ( .A(n7327), .B(n7326), .Z(n7328) );
  AND U10952 ( .A(n7329), .B(n7328), .Z(n10371) );
  NANDN U10953 ( .A(n7331), .B(n7330), .Z(n7335) );
  NAND U10954 ( .A(n7333), .B(n7332), .Z(n7334) );
  NAND U10955 ( .A(n7335), .B(n7334), .Z(n10370) );
  XNOR U10956 ( .A(n10371), .B(n10370), .Z(n10372) );
  XNOR U10957 ( .A(n10373), .B(n10372), .Z(n9448) );
  XOR U10958 ( .A(n9449), .B(n9448), .Z(n9797) );
  NANDN U10959 ( .A(n7337), .B(n7336), .Z(n7341) );
  NAND U10960 ( .A(n7339), .B(n7338), .Z(n7340) );
  AND U10961 ( .A(n7341), .B(n7340), .Z(n10403) );
  NANDN U10962 ( .A(n7343), .B(n7342), .Z(n7347) );
  NANDN U10963 ( .A(n7345), .B(n7344), .Z(n7346) );
  AND U10964 ( .A(n7347), .B(n7346), .Z(n10401) );
  NANDN U10965 ( .A(n7349), .B(n7348), .Z(n7353) );
  NANDN U10966 ( .A(n7351), .B(n7350), .Z(n7352) );
  NAND U10967 ( .A(n7353), .B(n7352), .Z(n10400) );
  XNOR U10968 ( .A(n10401), .B(n10400), .Z(n10402) );
  XNOR U10969 ( .A(n10403), .B(n10402), .Z(n9915) );
  NANDN U10970 ( .A(n7355), .B(n7354), .Z(n7359) );
  NANDN U10971 ( .A(n7357), .B(n7356), .Z(n7358) );
  AND U10972 ( .A(n7359), .B(n7358), .Z(n10409) );
  NANDN U10973 ( .A(n7361), .B(n7360), .Z(n7365) );
  NAND U10974 ( .A(n7363), .B(n7362), .Z(n7364) );
  AND U10975 ( .A(n7365), .B(n7364), .Z(n10407) );
  NANDN U10976 ( .A(n7367), .B(n7366), .Z(n7371) );
  NANDN U10977 ( .A(n7369), .B(n7368), .Z(n7370) );
  NAND U10978 ( .A(n7371), .B(n7370), .Z(n10406) );
  XNOR U10979 ( .A(n10407), .B(n10406), .Z(n10408) );
  XOR U10980 ( .A(n10409), .B(n10408), .Z(n9916) );
  XNOR U10981 ( .A(n9915), .B(n9916), .Z(n9918) );
  NANDN U10982 ( .A(n7373), .B(n7372), .Z(n7377) );
  OR U10983 ( .A(n7375), .B(n7374), .Z(n7376) );
  AND U10984 ( .A(n7377), .B(n7376), .Z(n9689) );
  NANDN U10985 ( .A(n7379), .B(n7378), .Z(n7383) );
  NAND U10986 ( .A(n7381), .B(n7380), .Z(n7382) );
  AND U10987 ( .A(n7383), .B(n7382), .Z(n9687) );
  NANDN U10988 ( .A(n7385), .B(n7384), .Z(n7389) );
  NAND U10989 ( .A(n7387), .B(n7386), .Z(n7388) );
  NAND U10990 ( .A(n7389), .B(n7388), .Z(n9686) );
  XNOR U10991 ( .A(n9687), .B(n9686), .Z(n9688) );
  XNOR U10992 ( .A(n9689), .B(n9688), .Z(n9917) );
  XOR U10993 ( .A(n9918), .B(n9917), .Z(n9795) );
  NANDN U10994 ( .A(n7391), .B(n7390), .Z(n7395) );
  NANDN U10995 ( .A(n7393), .B(n7392), .Z(n7394) );
  AND U10996 ( .A(n7395), .B(n7394), .Z(n9972) );
  NANDN U10997 ( .A(n7397), .B(n7396), .Z(n7401) );
  OR U10998 ( .A(n7399), .B(n7398), .Z(n7400) );
  AND U10999 ( .A(n7401), .B(n7400), .Z(n9969) );
  NANDN U11000 ( .A(n7403), .B(n7402), .Z(n7407) );
  OR U11001 ( .A(n7405), .B(n7404), .Z(n7406) );
  AND U11002 ( .A(n7407), .B(n7406), .Z(n9151) );
  NANDN U11003 ( .A(n7409), .B(n7408), .Z(n7413) );
  OR U11004 ( .A(n7411), .B(n7410), .Z(n7412) );
  AND U11005 ( .A(n7413), .B(n7412), .Z(n9149) );
  NANDN U11006 ( .A(n7415), .B(n7414), .Z(n7419) );
  NANDN U11007 ( .A(n7417), .B(n7416), .Z(n7418) );
  NAND U11008 ( .A(n7419), .B(n7418), .Z(n9148) );
  XNOR U11009 ( .A(n9149), .B(n9148), .Z(n9150) );
  XOR U11010 ( .A(n9151), .B(n9150), .Z(n9970) );
  XNOR U11011 ( .A(n9969), .B(n9970), .Z(n9971) );
  XNOR U11012 ( .A(n9972), .B(n9971), .Z(n9794) );
  XNOR U11013 ( .A(n9795), .B(n9794), .Z(n9796) );
  XNOR U11014 ( .A(n9797), .B(n9796), .Z(n9226) );
  XOR U11015 ( .A(n9227), .B(n9226), .Z(n9228) );
  XOR U11016 ( .A(n9229), .B(n9228), .Z(n9064) );
  XOR U11017 ( .A(n9065), .B(n9064), .Z(n9066) );
  NAND U11018 ( .A(n7421), .B(n7420), .Z(n7425) );
  NAND U11019 ( .A(n7423), .B(n7422), .Z(n7424) );
  AND U11020 ( .A(n7425), .B(n7424), .Z(n9073) );
  NAND U11021 ( .A(n7427), .B(n7426), .Z(n7431) );
  NAND U11022 ( .A(n7429), .B(n7428), .Z(n7430) );
  NAND U11023 ( .A(n7431), .B(n7430), .Z(n9813) );
  NANDN U11024 ( .A(n7433), .B(n7432), .Z(n7437) );
  NANDN U11025 ( .A(n7435), .B(n7434), .Z(n7436) );
  AND U11026 ( .A(n7437), .B(n7436), .Z(n9138) );
  NANDN U11027 ( .A(n7439), .B(n7438), .Z(n7443) );
  NANDN U11028 ( .A(n7441), .B(n7440), .Z(n7442) );
  AND U11029 ( .A(n7443), .B(n7442), .Z(n9136) );
  NANDN U11030 ( .A(n7445), .B(n7444), .Z(n7449) );
  NAND U11031 ( .A(n7447), .B(n7446), .Z(n7448) );
  AND U11032 ( .A(n7449), .B(n7448), .Z(n10314) );
  NANDN U11033 ( .A(n7451), .B(n7450), .Z(n7455) );
  NAND U11034 ( .A(n7453), .B(n7452), .Z(n7454) );
  AND U11035 ( .A(n7455), .B(n7454), .Z(n10313) );
  NANDN U11036 ( .A(n7457), .B(n7456), .Z(n7461) );
  NAND U11037 ( .A(n7459), .B(n7458), .Z(n7460) );
  NAND U11038 ( .A(n7461), .B(n7460), .Z(n10312) );
  XOR U11039 ( .A(n10313), .B(n10312), .Z(n10315) );
  XOR U11040 ( .A(n10314), .B(n10315), .Z(n9743) );
  NANDN U11041 ( .A(n7463), .B(n7462), .Z(n7467) );
  NAND U11042 ( .A(n7465), .B(n7464), .Z(n7466) );
  NAND U11043 ( .A(n7467), .B(n7466), .Z(n10097) );
  NANDN U11044 ( .A(n7469), .B(n7468), .Z(n7473) );
  NAND U11045 ( .A(n7471), .B(n7470), .Z(n7472) );
  NAND U11046 ( .A(n7473), .B(n7472), .Z(n10096) );
  NAND U11047 ( .A(n7475), .B(n7474), .Z(n7479) );
  NAND U11048 ( .A(n7477), .B(n7476), .Z(n7478) );
  NAND U11049 ( .A(n7479), .B(n7478), .Z(n10095) );
  XOR U11050 ( .A(n10096), .B(n10095), .Z(n10098) );
  XNOR U11051 ( .A(n10097), .B(n10098), .Z(n9741) );
  NANDN U11052 ( .A(n7481), .B(n7480), .Z(n7485) );
  NAND U11053 ( .A(n7483), .B(n7482), .Z(n7484) );
  NAND U11054 ( .A(n7485), .B(n7484), .Z(n10175) );
  NANDN U11055 ( .A(n7487), .B(n7486), .Z(n7491) );
  NAND U11056 ( .A(n7489), .B(n7488), .Z(n7490) );
  NAND U11057 ( .A(n7491), .B(n7490), .Z(n10174) );
  NANDN U11058 ( .A(n7493), .B(n7492), .Z(n7497) );
  NAND U11059 ( .A(n7495), .B(n7494), .Z(n7496) );
  NAND U11060 ( .A(n7497), .B(n7496), .Z(n10173) );
  XNOR U11061 ( .A(n10174), .B(n10173), .Z(n10176) );
  XOR U11062 ( .A(n10175), .B(n10176), .Z(n9740) );
  XOR U11063 ( .A(n9741), .B(n9740), .Z(n9742) );
  XOR U11064 ( .A(n9743), .B(n9742), .Z(n9137) );
  XOR U11065 ( .A(n9136), .B(n9137), .Z(n9139) );
  XNOR U11066 ( .A(n9138), .B(n9139), .Z(n9812) );
  XOR U11067 ( .A(n9813), .B(n9812), .Z(n9815) );
  NANDN U11068 ( .A(n7499), .B(n7498), .Z(n7503) );
  NAND U11069 ( .A(n7501), .B(n7500), .Z(n7502) );
  AND U11070 ( .A(n7503), .B(n7502), .Z(n10523) );
  NANDN U11071 ( .A(n7505), .B(n7504), .Z(n7509) );
  NANDN U11072 ( .A(n7507), .B(n7506), .Z(n7508) );
  AND U11073 ( .A(n7509), .B(n7508), .Z(n10520) );
  NANDN U11074 ( .A(n7511), .B(n7510), .Z(n7515) );
  NANDN U11075 ( .A(n7513), .B(n7512), .Z(n7514) );
  AND U11076 ( .A(n7515), .B(n7514), .Z(n9755) );
  NANDN U11077 ( .A(n7517), .B(n7516), .Z(n7521) );
  NAND U11078 ( .A(n7519), .B(n7518), .Z(n7520) );
  NAND U11079 ( .A(n7521), .B(n7520), .Z(n9886) );
  NANDN U11080 ( .A(n7523), .B(n7522), .Z(n7527) );
  NAND U11081 ( .A(n7525), .B(n7524), .Z(n7526) );
  NAND U11082 ( .A(n7527), .B(n7526), .Z(n9885) );
  XOR U11083 ( .A(n9886), .B(n9885), .Z(n9888) );
  NANDN U11084 ( .A(n7529), .B(n7528), .Z(n7533) );
  NAND U11085 ( .A(n7531), .B(n7530), .Z(n7532) );
  NAND U11086 ( .A(n7533), .B(n7532), .Z(n9887) );
  XOR U11087 ( .A(n9888), .B(n9887), .Z(n9753) );
  NANDN U11088 ( .A(n7535), .B(n7534), .Z(n7539) );
  NAND U11089 ( .A(n7537), .B(n7536), .Z(n7538) );
  NAND U11090 ( .A(n7539), .B(n7538), .Z(n10181) );
  NANDN U11091 ( .A(n7541), .B(n7540), .Z(n7545) );
  NAND U11092 ( .A(n7543), .B(n7542), .Z(n7544) );
  NAND U11093 ( .A(n7545), .B(n7544), .Z(n10180) );
  NANDN U11094 ( .A(n7547), .B(n7546), .Z(n7551) );
  NAND U11095 ( .A(n7549), .B(n7548), .Z(n7550) );
  NAND U11096 ( .A(n7551), .B(n7550), .Z(n10179) );
  XNOR U11097 ( .A(n10180), .B(n10179), .Z(n10182) );
  XOR U11098 ( .A(n10181), .B(n10182), .Z(n9752) );
  XNOR U11099 ( .A(n9753), .B(n9752), .Z(n9754) );
  XOR U11100 ( .A(n9755), .B(n9754), .Z(n10521) );
  XNOR U11101 ( .A(n10520), .B(n10521), .Z(n10522) );
  XNOR U11102 ( .A(n10523), .B(n10522), .Z(n9814) );
  XOR U11103 ( .A(n9815), .B(n9814), .Z(n9382) );
  NANDN U11104 ( .A(n7553), .B(n7552), .Z(n7557) );
  NANDN U11105 ( .A(n7555), .B(n7554), .Z(n7556) );
  AND U11106 ( .A(n7557), .B(n7556), .Z(n10541) );
  NANDN U11107 ( .A(n7559), .B(n7558), .Z(n7563) );
  NANDN U11108 ( .A(n7561), .B(n7560), .Z(n7562) );
  AND U11109 ( .A(n7563), .B(n7562), .Z(n10539) );
  NANDN U11110 ( .A(n7565), .B(n7564), .Z(n7569) );
  NAND U11111 ( .A(n7567), .B(n7566), .Z(n7568) );
  NAND U11112 ( .A(n7569), .B(n7568), .Z(n10193) );
  NANDN U11113 ( .A(n7571), .B(n7570), .Z(n7575) );
  NAND U11114 ( .A(n7573), .B(n7572), .Z(n7574) );
  NAND U11115 ( .A(n7575), .B(n7574), .Z(n10192) );
  NANDN U11116 ( .A(n7577), .B(n7576), .Z(n7581) );
  NAND U11117 ( .A(n7579), .B(n7578), .Z(n7580) );
  NAND U11118 ( .A(n7581), .B(n7580), .Z(n10191) );
  XOR U11119 ( .A(n10192), .B(n10191), .Z(n10194) );
  XNOR U11120 ( .A(n10193), .B(n10194), .Z(n9827) );
  NANDN U11121 ( .A(n7583), .B(n7582), .Z(n7587) );
  NAND U11122 ( .A(n7585), .B(n7584), .Z(n7586) );
  NAND U11123 ( .A(n7587), .B(n7586), .Z(n10308) );
  NANDN U11124 ( .A(n7589), .B(n7588), .Z(n7593) );
  NAND U11125 ( .A(n7591), .B(n7590), .Z(n7592) );
  NAND U11126 ( .A(n7593), .B(n7592), .Z(n10307) );
  NANDN U11127 ( .A(n7595), .B(n7594), .Z(n7599) );
  NAND U11128 ( .A(n7597), .B(n7596), .Z(n7598) );
  NAND U11129 ( .A(n7599), .B(n7598), .Z(n10306) );
  XOR U11130 ( .A(n10307), .B(n10306), .Z(n10309) );
  XNOR U11131 ( .A(n10308), .B(n10309), .Z(n9825) );
  NANDN U11132 ( .A(n7601), .B(n7600), .Z(n7605) );
  NAND U11133 ( .A(n7603), .B(n7602), .Z(n7604) );
  NAND U11134 ( .A(n7605), .B(n7604), .Z(n10235) );
  NANDN U11135 ( .A(n7607), .B(n7606), .Z(n7611) );
  NAND U11136 ( .A(n7609), .B(n7608), .Z(n7610) );
  NAND U11137 ( .A(n7611), .B(n7610), .Z(n10234) );
  NANDN U11138 ( .A(n7613), .B(n7612), .Z(n7617) );
  NAND U11139 ( .A(n7615), .B(n7614), .Z(n7616) );
  NAND U11140 ( .A(n7617), .B(n7616), .Z(n10233) );
  XNOR U11141 ( .A(n10234), .B(n10233), .Z(n10236) );
  XOR U11142 ( .A(n10235), .B(n10236), .Z(n9824) );
  XOR U11143 ( .A(n9825), .B(n9824), .Z(n9826) );
  XOR U11144 ( .A(n9827), .B(n9826), .Z(n10538) );
  XOR U11145 ( .A(n10539), .B(n10538), .Z(n10540) );
  XNOR U11146 ( .A(n10541), .B(n10540), .Z(n9821) );
  NANDN U11147 ( .A(n7619), .B(n7618), .Z(n7623) );
  NANDN U11148 ( .A(n7621), .B(n7620), .Z(n7622) );
  AND U11149 ( .A(n7623), .B(n7622), .Z(n9414) );
  NANDN U11150 ( .A(n7625), .B(n7624), .Z(n7629) );
  NANDN U11151 ( .A(n7627), .B(n7626), .Z(n7628) );
  AND U11152 ( .A(n7629), .B(n7628), .Z(n9411) );
  NANDN U11153 ( .A(n7631), .B(n7630), .Z(n7635) );
  NAND U11154 ( .A(n7633), .B(n7632), .Z(n7634) );
  AND U11155 ( .A(n7635), .B(n7634), .Z(n9839) );
  NANDN U11156 ( .A(n7637), .B(n7636), .Z(n7641) );
  NANDN U11157 ( .A(n7639), .B(n7638), .Z(n7640) );
  AND U11158 ( .A(n7641), .B(n7640), .Z(n9837) );
  NANDN U11159 ( .A(n7643), .B(n7642), .Z(n7647) );
  NAND U11160 ( .A(n7645), .B(n7644), .Z(n7646) );
  NAND U11161 ( .A(n7647), .B(n7646), .Z(n9419) );
  NANDN U11162 ( .A(n7649), .B(n7648), .Z(n7653) );
  NAND U11163 ( .A(n7651), .B(n7650), .Z(n7652) );
  NAND U11164 ( .A(n7653), .B(n7652), .Z(n9418) );
  NANDN U11165 ( .A(n7655), .B(n7654), .Z(n7659) );
  NAND U11166 ( .A(n7657), .B(n7656), .Z(n7658) );
  NAND U11167 ( .A(n7659), .B(n7658), .Z(n9417) );
  XNOR U11168 ( .A(n9418), .B(n9417), .Z(n9420) );
  XOR U11169 ( .A(n9419), .B(n9420), .Z(n9836) );
  XNOR U11170 ( .A(n9837), .B(n9836), .Z(n9838) );
  XOR U11171 ( .A(n9839), .B(n9838), .Z(n9412) );
  XNOR U11172 ( .A(n9411), .B(n9412), .Z(n9413) );
  XNOR U11173 ( .A(n9414), .B(n9413), .Z(n9819) );
  NAND U11174 ( .A(n7661), .B(n7660), .Z(n7665) );
  NAND U11175 ( .A(n7663), .B(n7662), .Z(n7664) );
  AND U11176 ( .A(n7665), .B(n7664), .Z(n9818) );
  XOR U11177 ( .A(n9819), .B(n9818), .Z(n9820) );
  XOR U11178 ( .A(n9821), .B(n9820), .Z(n9381) );
  NANDN U11179 ( .A(n7667), .B(n7666), .Z(n7671) );
  NANDN U11180 ( .A(n7669), .B(n7668), .Z(n7670) );
  AND U11181 ( .A(n7671), .B(n7670), .Z(n9283) );
  NANDN U11182 ( .A(n7677), .B(n7676), .Z(n7681) );
  NAND U11183 ( .A(n7679), .B(n7678), .Z(n7680) );
  AND U11184 ( .A(n7681), .B(n7680), .Z(n9929) );
  NANDN U11185 ( .A(n7683), .B(n7682), .Z(n7687) );
  NAND U11186 ( .A(n7685), .B(n7684), .Z(n7686) );
  AND U11187 ( .A(n7687), .B(n7686), .Z(n9928) );
  NANDN U11188 ( .A(n7689), .B(n7688), .Z(n7693) );
  NAND U11189 ( .A(n7691), .B(n7690), .Z(n7692) );
  NAND U11190 ( .A(n7693), .B(n7692), .Z(n9927) );
  XOR U11191 ( .A(n9928), .B(n9927), .Z(n9930) );
  XOR U11192 ( .A(n9929), .B(n9930), .Z(n9479) );
  NANDN U11193 ( .A(n7695), .B(n7694), .Z(n7699) );
  NAND U11194 ( .A(n7697), .B(n7696), .Z(n7698) );
  AND U11195 ( .A(n7699), .B(n7698), .Z(n9477) );
  NANDN U11196 ( .A(n7701), .B(n7700), .Z(n7705) );
  NAND U11197 ( .A(n7703), .B(n7702), .Z(n7704) );
  AND U11198 ( .A(n7705), .B(n7704), .Z(n9941) );
  NANDN U11199 ( .A(n7707), .B(n7706), .Z(n7711) );
  NAND U11200 ( .A(n7709), .B(n7708), .Z(n7710) );
  AND U11201 ( .A(n7711), .B(n7710), .Z(n9940) );
  NANDN U11202 ( .A(n7713), .B(n7712), .Z(n7717) );
  NANDN U11203 ( .A(n7715), .B(n7714), .Z(n7716) );
  NAND U11204 ( .A(n7717), .B(n7716), .Z(n9939) );
  XOR U11205 ( .A(n9940), .B(n9939), .Z(n9942) );
  XNOR U11206 ( .A(n9941), .B(n9942), .Z(n9476) );
  XNOR U11207 ( .A(n9477), .B(n9476), .Z(n9478) );
  XNOR U11208 ( .A(n9479), .B(n9478), .Z(n9280) );
  XNOR U11209 ( .A(n9281), .B(n9280), .Z(n9282) );
  XNOR U11210 ( .A(n9283), .B(n9282), .Z(n9767) );
  NANDN U11211 ( .A(n7723), .B(n7722), .Z(n7727) );
  NAND U11212 ( .A(n7725), .B(n7724), .Z(n7726) );
  NAND U11213 ( .A(n7727), .B(n7726), .Z(n9875) );
  NAND U11214 ( .A(n7729), .B(n7728), .Z(n7733) );
  NAND U11215 ( .A(n7731), .B(n7730), .Z(n7732) );
  NAND U11216 ( .A(n7733), .B(n7732), .Z(n9874) );
  NANDN U11217 ( .A(n7735), .B(n7734), .Z(n7739) );
  NAND U11218 ( .A(n7737), .B(n7736), .Z(n7738) );
  NAND U11219 ( .A(n7739), .B(n7738), .Z(n9873) );
  XOR U11220 ( .A(n9874), .B(n9873), .Z(n9876) );
  XOR U11221 ( .A(n9875), .B(n9876), .Z(n9485) );
  NANDN U11222 ( .A(n7741), .B(n7740), .Z(n7745) );
  NANDN U11223 ( .A(n7743), .B(n7742), .Z(n7744) );
  AND U11224 ( .A(n7745), .B(n7744), .Z(n9482) );
  NANDN U11225 ( .A(n7747), .B(n7746), .Z(n7751) );
  NANDN U11226 ( .A(n7749), .B(n7748), .Z(n7750) );
  NAND U11227 ( .A(n7751), .B(n7750), .Z(n9483) );
  XNOR U11228 ( .A(n9482), .B(n9483), .Z(n9484) );
  XOR U11229 ( .A(n9485), .B(n9484), .Z(n9263) );
  NANDN U11230 ( .A(n7753), .B(n7752), .Z(n7757) );
  NANDN U11231 ( .A(n7755), .B(n7754), .Z(n7756) );
  AND U11232 ( .A(n7757), .B(n7756), .Z(n9262) );
  XOR U11233 ( .A(n9263), .B(n9262), .Z(n9265) );
  XNOR U11234 ( .A(n9264), .B(n9265), .Z(n9765) );
  NAND U11235 ( .A(n7759), .B(n7758), .Z(n7763) );
  NAND U11236 ( .A(n7761), .B(n7760), .Z(n7762) );
  NAND U11237 ( .A(n7763), .B(n7762), .Z(n9764) );
  XOR U11238 ( .A(n9765), .B(n9764), .Z(n9766) );
  XOR U11239 ( .A(n9767), .B(n9766), .Z(n9383) );
  XOR U11240 ( .A(n9384), .B(n9383), .Z(n9071) );
  NAND U11241 ( .A(n7765), .B(n7764), .Z(n7769) );
  NAND U11242 ( .A(n7767), .B(n7766), .Z(n7768) );
  AND U11243 ( .A(n7769), .B(n7768), .Z(n9806) );
  NANDN U11244 ( .A(n7771), .B(n7770), .Z(n7775) );
  NANDN U11245 ( .A(n7773), .B(n7772), .Z(n7774) );
  AND U11246 ( .A(n7775), .B(n7774), .Z(n10462) );
  NANDN U11247 ( .A(n7777), .B(n7776), .Z(n7781) );
  NANDN U11248 ( .A(n7779), .B(n7778), .Z(n7780) );
  AND U11249 ( .A(n7781), .B(n7780), .Z(n10460) );
  NANDN U11250 ( .A(n7783), .B(n7782), .Z(n7787) );
  NAND U11251 ( .A(n7785), .B(n7784), .Z(n7786) );
  AND U11252 ( .A(n7787), .B(n7786), .Z(n9597) );
  NAND U11253 ( .A(n7789), .B(n7788), .Z(n7793) );
  NAND U11254 ( .A(n7791), .B(n7790), .Z(n7792) );
  AND U11255 ( .A(n7793), .B(n7792), .Z(n9596) );
  NANDN U11256 ( .A(n7795), .B(n7794), .Z(n7799) );
  NAND U11257 ( .A(n7797), .B(n7796), .Z(n7798) );
  NAND U11258 ( .A(n7799), .B(n7798), .Z(n9595) );
  XOR U11259 ( .A(n9596), .B(n9595), .Z(n9598) );
  XOR U11260 ( .A(n9597), .B(n9598), .Z(n10493) );
  NANDN U11261 ( .A(n7801), .B(n7800), .Z(n7805) );
  NAND U11262 ( .A(n7803), .B(n7802), .Z(n7804) );
  AND U11263 ( .A(n7805), .B(n7804), .Z(n9591) );
  NAND U11264 ( .A(n7807), .B(n7806), .Z(n7811) );
  NAND U11265 ( .A(n7809), .B(n7808), .Z(n7810) );
  AND U11266 ( .A(n7811), .B(n7810), .Z(n9590) );
  NANDN U11267 ( .A(n7813), .B(n7812), .Z(n7817) );
  NAND U11268 ( .A(n7815), .B(n7814), .Z(n7816) );
  NAND U11269 ( .A(n7817), .B(n7816), .Z(n9589) );
  XOR U11270 ( .A(n9590), .B(n9589), .Z(n9592) );
  XOR U11271 ( .A(n9591), .B(n9592), .Z(n10491) );
  NANDN U11272 ( .A(n7819), .B(n7818), .Z(n7823) );
  NAND U11273 ( .A(n7821), .B(n7820), .Z(n7822) );
  AND U11274 ( .A(n7823), .B(n7822), .Z(n9460) );
  NANDN U11275 ( .A(n7825), .B(n7824), .Z(n7829) );
  NAND U11276 ( .A(n7827), .B(n7826), .Z(n7828) );
  AND U11277 ( .A(n7829), .B(n7828), .Z(n9459) );
  NANDN U11278 ( .A(n7831), .B(n7830), .Z(n7835) );
  NAND U11279 ( .A(n7833), .B(n7832), .Z(n7834) );
  NAND U11280 ( .A(n7835), .B(n7834), .Z(n9458) );
  XOR U11281 ( .A(n9459), .B(n9458), .Z(n9461) );
  XNOR U11282 ( .A(n9460), .B(n9461), .Z(n10490) );
  XNOR U11283 ( .A(n10491), .B(n10490), .Z(n10492) );
  XOR U11284 ( .A(n10493), .B(n10492), .Z(n10461) );
  XOR U11285 ( .A(n10460), .B(n10461), .Z(n10463) );
  XNOR U11286 ( .A(n10462), .B(n10463), .Z(n9807) );
  XOR U11287 ( .A(n9806), .B(n9807), .Z(n9809) );
  NANDN U11288 ( .A(n7837), .B(n7836), .Z(n7841) );
  NAND U11289 ( .A(n7839), .B(n7838), .Z(n7840) );
  AND U11290 ( .A(n7841), .B(n7840), .Z(n10355) );
  NANDN U11291 ( .A(n7843), .B(n7842), .Z(n7847) );
  NANDN U11292 ( .A(n7845), .B(n7844), .Z(n7846) );
  AND U11293 ( .A(n7847), .B(n7846), .Z(n10352) );
  NANDN U11294 ( .A(n7849), .B(n7848), .Z(n7853) );
  NAND U11295 ( .A(n7851), .B(n7850), .Z(n7852) );
  AND U11296 ( .A(n7853), .B(n7852), .Z(n10487) );
  NANDN U11297 ( .A(n7855), .B(n7854), .Z(n7859) );
  NAND U11298 ( .A(n7857), .B(n7856), .Z(n7858) );
  AND U11299 ( .A(n7859), .B(n7858), .Z(n10485) );
  NAND U11300 ( .A(n7861), .B(n7860), .Z(n7865) );
  NAND U11301 ( .A(n7863), .B(n7862), .Z(n7864) );
  AND U11302 ( .A(n7865), .B(n7864), .Z(n9651) );
  NAND U11303 ( .A(n7867), .B(n7866), .Z(n7871) );
  NAND U11304 ( .A(n7869), .B(n7868), .Z(n7870) );
  AND U11305 ( .A(n7871), .B(n7870), .Z(n9650) );
  NANDN U11306 ( .A(n7873), .B(n7872), .Z(n7877) );
  NAND U11307 ( .A(n7875), .B(n7874), .Z(n7876) );
  NAND U11308 ( .A(n7877), .B(n7876), .Z(n9649) );
  XOR U11309 ( .A(n9650), .B(n9649), .Z(n9652) );
  XNOR U11310 ( .A(n9651), .B(n9652), .Z(n10484) );
  XNOR U11311 ( .A(n10485), .B(n10484), .Z(n10486) );
  XOR U11312 ( .A(n10487), .B(n10486), .Z(n10353) );
  XNOR U11313 ( .A(n10352), .B(n10353), .Z(n10354) );
  XNOR U11314 ( .A(n10355), .B(n10354), .Z(n9808) );
  XNOR U11315 ( .A(n9809), .B(n9808), .Z(n9289) );
  NANDN U11316 ( .A(n7879), .B(n7878), .Z(n7883) );
  NANDN U11317 ( .A(n7881), .B(n7880), .Z(n7882) );
  AND U11318 ( .A(n7883), .B(n7882), .Z(n9210) );
  NANDN U11319 ( .A(n7885), .B(n7884), .Z(n7889) );
  NANDN U11320 ( .A(n7887), .B(n7886), .Z(n7888) );
  AND U11321 ( .A(n7889), .B(n7888), .Z(n9208) );
  NANDN U11322 ( .A(n7891), .B(n7890), .Z(n7895) );
  NAND U11323 ( .A(n7893), .B(n7892), .Z(n7894) );
  AND U11324 ( .A(n7895), .B(n7894), .Z(n10032) );
  NANDN U11325 ( .A(n7897), .B(n7896), .Z(n7901) );
  NAND U11326 ( .A(n7899), .B(n7898), .Z(n7900) );
  AND U11327 ( .A(n7901), .B(n7900), .Z(n10030) );
  NANDN U11328 ( .A(n7903), .B(n7902), .Z(n7907) );
  NANDN U11329 ( .A(n7905), .B(n7904), .Z(n7906) );
  NAND U11330 ( .A(n7907), .B(n7906), .Z(n10029) );
  XNOR U11331 ( .A(n10030), .B(n10029), .Z(n10031) );
  XOR U11332 ( .A(n10032), .B(n10031), .Z(n9209) );
  XOR U11333 ( .A(n9208), .B(n9209), .Z(n9211) );
  XNOR U11334 ( .A(n9210), .B(n9211), .Z(n9782) );
  NANDN U11335 ( .A(n7909), .B(n7908), .Z(n7913) );
  NANDN U11336 ( .A(n7911), .B(n7910), .Z(n7912) );
  AND U11337 ( .A(n7913), .B(n7912), .Z(n10152) );
  NANDN U11338 ( .A(n7918), .B(n7917), .Z(n7922) );
  NAND U11339 ( .A(n7920), .B(n7919), .Z(n7921) );
  AND U11340 ( .A(n7922), .B(n7921), .Z(n10140) );
  NANDN U11341 ( .A(n7924), .B(n7923), .Z(n7928) );
  NAND U11342 ( .A(n7926), .B(n7925), .Z(n7927) );
  AND U11343 ( .A(n7928), .B(n7927), .Z(n10138) );
  NANDN U11344 ( .A(n7930), .B(n7929), .Z(n7934) );
  NANDN U11345 ( .A(n7932), .B(n7931), .Z(n7933) );
  NAND U11346 ( .A(n7934), .B(n7933), .Z(n10137) );
  XNOR U11347 ( .A(n10138), .B(n10137), .Z(n10139) );
  XNOR U11348 ( .A(n10140), .B(n10139), .Z(n10149) );
  XNOR U11349 ( .A(n10150), .B(n10149), .Z(n10151) );
  XOR U11350 ( .A(n10152), .B(n10151), .Z(n9783) );
  XNOR U11351 ( .A(n9782), .B(n9783), .Z(n9785) );
  NANDN U11352 ( .A(n7936), .B(n7935), .Z(n7940) );
  NANDN U11353 ( .A(n7938), .B(n7937), .Z(n7939) );
  AND U11354 ( .A(n7940), .B(n7939), .Z(n9843) );
  NANDN U11355 ( .A(n7942), .B(n7941), .Z(n7946) );
  OR U11356 ( .A(n7944), .B(n7943), .Z(n7945) );
  AND U11357 ( .A(n7946), .B(n7945), .Z(n10074) );
  NANDN U11358 ( .A(n7948), .B(n7947), .Z(n7952) );
  OR U11359 ( .A(n7950), .B(n7949), .Z(n7951) );
  AND U11360 ( .A(n7952), .B(n7951), .Z(n10072) );
  NANDN U11361 ( .A(n7954), .B(n7953), .Z(n7958) );
  NANDN U11362 ( .A(n7956), .B(n7955), .Z(n7957) );
  NAND U11363 ( .A(n7958), .B(n7957), .Z(n10071) );
  XNOR U11364 ( .A(n10072), .B(n10071), .Z(n10073) );
  XOR U11365 ( .A(n10074), .B(n10073), .Z(n9844) );
  XNOR U11366 ( .A(n9843), .B(n9844), .Z(n9845) );
  NANDN U11367 ( .A(n7960), .B(n7959), .Z(n7964) );
  OR U11368 ( .A(n7962), .B(n7961), .Z(n7963) );
  AND U11369 ( .A(n7964), .B(n7963), .Z(n10291) );
  NANDN U11370 ( .A(n7966), .B(n7965), .Z(n7970) );
  OR U11371 ( .A(n7968), .B(n7967), .Z(n7969) );
  AND U11372 ( .A(n7970), .B(n7969), .Z(n10289) );
  NANDN U11373 ( .A(n7972), .B(n7971), .Z(n7976) );
  NANDN U11374 ( .A(n7974), .B(n7973), .Z(n7975) );
  NAND U11375 ( .A(n7976), .B(n7975), .Z(n10288) );
  XNOR U11376 ( .A(n10289), .B(n10288), .Z(n10290) );
  XOR U11377 ( .A(n10291), .B(n10290), .Z(n9846) );
  XNOR U11378 ( .A(n9845), .B(n9846), .Z(n9784) );
  XNOR U11379 ( .A(n9785), .B(n9784), .Z(n9287) );
  NANDN U11380 ( .A(n7978), .B(n7977), .Z(n7982) );
  NANDN U11381 ( .A(n7980), .B(n7979), .Z(n7981) );
  AND U11382 ( .A(n7982), .B(n7981), .Z(n10412) );
  NANDN U11383 ( .A(n7984), .B(n7983), .Z(n7988) );
  NANDN U11384 ( .A(n7986), .B(n7985), .Z(n7987) );
  AND U11385 ( .A(n7988), .B(n7987), .Z(n10475) );
  NANDN U11386 ( .A(n7990), .B(n7989), .Z(n7994) );
  NAND U11387 ( .A(n7992), .B(n7991), .Z(n7993) );
  AND U11388 ( .A(n7994), .B(n7993), .Z(n10473) );
  NANDN U11389 ( .A(n7996), .B(n7995), .Z(n8000) );
  NANDN U11390 ( .A(n7998), .B(n7997), .Z(n7999) );
  NAND U11391 ( .A(n8000), .B(n7999), .Z(n10472) );
  XNOR U11392 ( .A(n10473), .B(n10472), .Z(n10474) );
  XOR U11393 ( .A(n10475), .B(n10474), .Z(n10413) );
  XNOR U11394 ( .A(n10412), .B(n10413), .Z(n10414) );
  NANDN U11395 ( .A(n8002), .B(n8001), .Z(n8006) );
  OR U11396 ( .A(n8004), .B(n8003), .Z(n8005) );
  AND U11397 ( .A(n8006), .B(n8005), .Z(n10242) );
  NANDN U11398 ( .A(n8008), .B(n8007), .Z(n8012) );
  OR U11399 ( .A(n8010), .B(n8009), .Z(n8011) );
  AND U11400 ( .A(n8012), .B(n8011), .Z(n10240) );
  NANDN U11401 ( .A(n8014), .B(n8013), .Z(n8018) );
  OR U11402 ( .A(n8016), .B(n8015), .Z(n8017) );
  NAND U11403 ( .A(n8018), .B(n8017), .Z(n10239) );
  XNOR U11404 ( .A(n10240), .B(n10239), .Z(n10241) );
  XOR U11405 ( .A(n10242), .B(n10241), .Z(n10415) );
  XOR U11406 ( .A(n10414), .B(n10415), .Z(n9760) );
  NAND U11407 ( .A(n8020), .B(n8019), .Z(n8024) );
  NANDN U11408 ( .A(n8022), .B(n8021), .Z(n8023) );
  AND U11409 ( .A(n8024), .B(n8023), .Z(n9759) );
  NANDN U11410 ( .A(n8026), .B(n8025), .Z(n8030) );
  NANDN U11411 ( .A(n8028), .B(n8027), .Z(n8029) );
  AND U11412 ( .A(n8030), .B(n8029), .Z(n9706) );
  NANDN U11413 ( .A(n8032), .B(n8031), .Z(n8036) );
  NAND U11414 ( .A(n8034), .B(n8033), .Z(n8035) );
  AND U11415 ( .A(n8036), .B(n8035), .Z(n9705) );
  NANDN U11416 ( .A(n8038), .B(n8037), .Z(n8042) );
  OR U11417 ( .A(n8040), .B(n8039), .Z(n8041) );
  AND U11418 ( .A(n8042), .B(n8041), .Z(n10433) );
  NANDN U11419 ( .A(n8044), .B(n8043), .Z(n8048) );
  NANDN U11420 ( .A(n8046), .B(n8045), .Z(n8047) );
  AND U11421 ( .A(n8048), .B(n8047), .Z(n10431) );
  NANDN U11422 ( .A(n8050), .B(n8049), .Z(n8054) );
  OR U11423 ( .A(n8052), .B(n8051), .Z(n8053) );
  NAND U11424 ( .A(n8054), .B(n8053), .Z(n10430) );
  XNOR U11425 ( .A(n10431), .B(n10430), .Z(n10432) );
  XNOR U11426 ( .A(n10433), .B(n10432), .Z(n9704) );
  XOR U11427 ( .A(n9705), .B(n9704), .Z(n9707) );
  XOR U11428 ( .A(n9706), .B(n9707), .Z(n9758) );
  XOR U11429 ( .A(n9759), .B(n9758), .Z(n9761) );
  XOR U11430 ( .A(n9760), .B(n9761), .Z(n9286) );
  XOR U11431 ( .A(n9287), .B(n9286), .Z(n9288) );
  XOR U11432 ( .A(n9289), .B(n9288), .Z(n9070) );
  XOR U11433 ( .A(n9071), .B(n9070), .Z(n9072) );
  XOR U11434 ( .A(n9073), .B(n9072), .Z(n10548) );
  XOR U11435 ( .A(n10549), .B(n10548), .Z(n10551) );
  NANDN U11436 ( .A(n8056), .B(n8055), .Z(n8060) );
  NANDN U11437 ( .A(n8058), .B(n8057), .Z(n8059) );
  AND U11438 ( .A(n8060), .B(n8059), .Z(n9867) );
  NAND U11439 ( .A(n8062), .B(n8061), .Z(n8066) );
  NAND U11440 ( .A(n8064), .B(n8063), .Z(n8065) );
  AND U11441 ( .A(n8066), .B(n8065), .Z(n10079) );
  NANDN U11442 ( .A(n8068), .B(n8067), .Z(n8072) );
  NAND U11443 ( .A(n8070), .B(n8069), .Z(n8071) );
  AND U11444 ( .A(n8072), .B(n8071), .Z(n10078) );
  NANDN U11445 ( .A(n8074), .B(n8073), .Z(n8078) );
  NAND U11446 ( .A(n8076), .B(n8075), .Z(n8077) );
  NAND U11447 ( .A(n8078), .B(n8077), .Z(n10077) );
  XOR U11448 ( .A(n10078), .B(n10077), .Z(n10080) );
  XOR U11449 ( .A(n10079), .B(n10080), .Z(n9570) );
  NANDN U11450 ( .A(n8080), .B(n8079), .Z(n8084) );
  NAND U11451 ( .A(n8082), .B(n8081), .Z(n8083) );
  NAND U11452 ( .A(n8084), .B(n8083), .Z(n9670) );
  NANDN U11453 ( .A(n8086), .B(n8085), .Z(n8090) );
  NANDN U11454 ( .A(n8088), .B(n8087), .Z(n8089) );
  NAND U11455 ( .A(n8090), .B(n8089), .Z(n9669) );
  NANDN U11456 ( .A(n8092), .B(n8091), .Z(n8096) );
  NAND U11457 ( .A(n8094), .B(n8093), .Z(n8095) );
  NAND U11458 ( .A(n8096), .B(n8095), .Z(n9668) );
  XOR U11459 ( .A(n9669), .B(n9668), .Z(n9671) );
  XNOR U11460 ( .A(n9670), .B(n9671), .Z(n9568) );
  NAND U11461 ( .A(n8098), .B(n8097), .Z(n8102) );
  NAND U11462 ( .A(n8100), .B(n8099), .Z(n8101) );
  NAND U11463 ( .A(n8102), .B(n8101), .Z(n9658) );
  NAND U11464 ( .A(n8104), .B(n8103), .Z(n8108) );
  NAND U11465 ( .A(n8106), .B(n8105), .Z(n8107) );
  NAND U11466 ( .A(n8108), .B(n8107), .Z(n9657) );
  NANDN U11467 ( .A(n8110), .B(n8109), .Z(n8114) );
  NAND U11468 ( .A(n8112), .B(n8111), .Z(n8113) );
  NAND U11469 ( .A(n8114), .B(n8113), .Z(n9656) );
  XNOR U11470 ( .A(n9657), .B(n9656), .Z(n9659) );
  XOR U11471 ( .A(n9658), .B(n9659), .Z(n9567) );
  XOR U11472 ( .A(n9568), .B(n9567), .Z(n9569) );
  XNOR U11473 ( .A(n9570), .B(n9569), .Z(n9341) );
  NANDN U11474 ( .A(n8116), .B(n8115), .Z(n8120) );
  NANDN U11475 ( .A(n8118), .B(n8117), .Z(n8119) );
  AND U11476 ( .A(n8120), .B(n8119), .Z(n10146) );
  NANDN U11477 ( .A(n8122), .B(n8121), .Z(n8126) );
  NAND U11478 ( .A(n8124), .B(n8123), .Z(n8125) );
  AND U11479 ( .A(n8126), .B(n8125), .Z(n10144) );
  NANDN U11480 ( .A(n8128), .B(n8127), .Z(n8132) );
  NAND U11481 ( .A(n8130), .B(n8129), .Z(n8131) );
  AND U11482 ( .A(n8132), .B(n8131), .Z(n10007) );
  NANDN U11483 ( .A(n8134), .B(n8133), .Z(n8138) );
  NAND U11484 ( .A(n8136), .B(n8135), .Z(n8137) );
  AND U11485 ( .A(n8138), .B(n8137), .Z(n10006) );
  NANDN U11486 ( .A(n8140), .B(n8139), .Z(n8144) );
  NAND U11487 ( .A(n8142), .B(n8141), .Z(n8143) );
  NAND U11488 ( .A(n8144), .B(n8143), .Z(n10005) );
  XOR U11489 ( .A(n10006), .B(n10005), .Z(n10008) );
  XNOR U11490 ( .A(n10007), .B(n10008), .Z(n10143) );
  XNOR U11491 ( .A(n10144), .B(n10143), .Z(n10145) );
  XOR U11492 ( .A(n10146), .B(n10145), .Z(n9342) );
  XNOR U11493 ( .A(n9341), .B(n9342), .Z(n9343) );
  NANDN U11494 ( .A(n8146), .B(n8145), .Z(n8150) );
  NAND U11495 ( .A(n8148), .B(n8147), .Z(n8149) );
  AND U11496 ( .A(n8150), .B(n8149), .Z(n9558) );
  NANDN U11497 ( .A(n8152), .B(n8151), .Z(n8156) );
  NAND U11498 ( .A(n8154), .B(n8153), .Z(n8155) );
  AND U11499 ( .A(n8156), .B(n8155), .Z(n10266) );
  NAND U11500 ( .A(n8158), .B(n8157), .Z(n8162) );
  NAND U11501 ( .A(n8160), .B(n8159), .Z(n8161) );
  AND U11502 ( .A(n8162), .B(n8161), .Z(n10265) );
  NANDN U11503 ( .A(n8164), .B(n8163), .Z(n8168) );
  NAND U11504 ( .A(n8166), .B(n8165), .Z(n8167) );
  NAND U11505 ( .A(n8168), .B(n8167), .Z(n10264) );
  XOR U11506 ( .A(n10265), .B(n10264), .Z(n10267) );
  XOR U11507 ( .A(n10266), .B(n10267), .Z(n9556) );
  NANDN U11508 ( .A(n8170), .B(n8169), .Z(n8174) );
  NANDN U11509 ( .A(n8172), .B(n8171), .Z(n8173) );
  NAND U11510 ( .A(n8174), .B(n8173), .Z(n9555) );
  XNOR U11511 ( .A(n9556), .B(n9555), .Z(n9557) );
  XOR U11512 ( .A(n9558), .B(n9557), .Z(n9344) );
  XOR U11513 ( .A(n9343), .B(n9344), .Z(n9868) );
  XNOR U11514 ( .A(n9867), .B(n9868), .Z(n9870) );
  NANDN U11515 ( .A(n8176), .B(n8175), .Z(n8180) );
  OR U11516 ( .A(n8178), .B(n8177), .Z(n8179) );
  AND U11517 ( .A(n8180), .B(n8179), .Z(n9564) );
  NANDN U11518 ( .A(n8182), .B(n8181), .Z(n8186) );
  NAND U11519 ( .A(n8184), .B(n8183), .Z(n8185) );
  AND U11520 ( .A(n8186), .B(n8185), .Z(n10260) );
  NANDN U11521 ( .A(n8188), .B(n8187), .Z(n8192) );
  NAND U11522 ( .A(n8190), .B(n8189), .Z(n8191) );
  AND U11523 ( .A(n8192), .B(n8191), .Z(n10259) );
  NANDN U11524 ( .A(n8194), .B(n8193), .Z(n8198) );
  NAND U11525 ( .A(n8196), .B(n8195), .Z(n8197) );
  NAND U11526 ( .A(n8198), .B(n8197), .Z(n10258) );
  XOR U11527 ( .A(n10259), .B(n10258), .Z(n10261) );
  XOR U11528 ( .A(n10260), .B(n10261), .Z(n9562) );
  NANDN U11529 ( .A(n8200), .B(n8199), .Z(n8204) );
  NAND U11530 ( .A(n8202), .B(n8201), .Z(n8203) );
  NAND U11531 ( .A(n8204), .B(n8203), .Z(n9561) );
  XNOR U11532 ( .A(n9562), .B(n9561), .Z(n9563) );
  XNOR U11533 ( .A(n9564), .B(n9563), .Z(n9347) );
  NANDN U11534 ( .A(n8206), .B(n8205), .Z(n8210) );
  NANDN U11535 ( .A(n8208), .B(n8207), .Z(n8209) );
  AND U11536 ( .A(n8210), .B(n8209), .Z(n10062) );
  NANDN U11537 ( .A(n8212), .B(n8211), .Z(n8216) );
  OR U11538 ( .A(n8214), .B(n8213), .Z(n8215) );
  AND U11539 ( .A(n8216), .B(n8215), .Z(n10060) );
  NANDN U11540 ( .A(n8218), .B(n8217), .Z(n8222) );
  NAND U11541 ( .A(n8220), .B(n8219), .Z(n8221) );
  AND U11542 ( .A(n8222), .B(n8221), .Z(n9615) );
  NANDN U11543 ( .A(n8224), .B(n8223), .Z(n8228) );
  NAND U11544 ( .A(n8226), .B(n8225), .Z(n8227) );
  AND U11545 ( .A(n8228), .B(n8227), .Z(n9614) );
  NANDN U11546 ( .A(n8230), .B(n8229), .Z(n8234) );
  NAND U11547 ( .A(n8232), .B(n8231), .Z(n8233) );
  NAND U11548 ( .A(n8234), .B(n8233), .Z(n9613) );
  XOR U11549 ( .A(n9614), .B(n9613), .Z(n9616) );
  XNOR U11550 ( .A(n9615), .B(n9616), .Z(n10059) );
  XNOR U11551 ( .A(n10060), .B(n10059), .Z(n10061) );
  XOR U11552 ( .A(n10062), .B(n10061), .Z(n9348) );
  XNOR U11553 ( .A(n9347), .B(n9348), .Z(n9350) );
  NANDN U11554 ( .A(n8236), .B(n8235), .Z(n8240) );
  NAND U11555 ( .A(n8238), .B(n8237), .Z(n8239) );
  NAND U11556 ( .A(n8240), .B(n8239), .Z(n10127) );
  NANDN U11557 ( .A(n8242), .B(n8241), .Z(n8246) );
  NANDN U11558 ( .A(n8244), .B(n8243), .Z(n8245) );
  NAND U11559 ( .A(n8246), .B(n8245), .Z(n10126) );
  NANDN U11560 ( .A(n8248), .B(n8247), .Z(n8252) );
  NAND U11561 ( .A(n8250), .B(n8249), .Z(n8251) );
  NAND U11562 ( .A(n8252), .B(n8251), .Z(n10125) );
  XOR U11563 ( .A(n10126), .B(n10125), .Z(n10128) );
  XNOR U11564 ( .A(n10127), .B(n10128), .Z(n9864) );
  NANDN U11565 ( .A(n8254), .B(n8253), .Z(n8258) );
  NAND U11566 ( .A(n8256), .B(n8255), .Z(n8257) );
  AND U11567 ( .A(n8258), .B(n8257), .Z(n9862) );
  NAND U11568 ( .A(n8260), .B(n8259), .Z(n8264) );
  NAND U11569 ( .A(n8262), .B(n8261), .Z(n8263) );
  NAND U11570 ( .A(n8264), .B(n8263), .Z(n10037) );
  NANDN U11571 ( .A(n8266), .B(n8265), .Z(n8270) );
  NAND U11572 ( .A(n8268), .B(n8267), .Z(n8269) );
  NAND U11573 ( .A(n8270), .B(n8269), .Z(n10036) );
  NANDN U11574 ( .A(n8272), .B(n8271), .Z(n8276) );
  NAND U11575 ( .A(n8274), .B(n8273), .Z(n8275) );
  NAND U11576 ( .A(n8276), .B(n8275), .Z(n10035) );
  XNOR U11577 ( .A(n10036), .B(n10035), .Z(n10038) );
  XOR U11578 ( .A(n10037), .B(n10038), .Z(n9861) );
  XNOR U11579 ( .A(n9862), .B(n9861), .Z(n9863) );
  XOR U11580 ( .A(n9864), .B(n9863), .Z(n9349) );
  XOR U11581 ( .A(n9350), .B(n9349), .Z(n9869) );
  XNOR U11582 ( .A(n9870), .B(n9869), .Z(n9360) );
  NANDN U11583 ( .A(n8278), .B(n8277), .Z(n8282) );
  NAND U11584 ( .A(n8280), .B(n8279), .Z(n8281) );
  AND U11585 ( .A(n8282), .B(n8281), .Z(n9789) );
  NANDN U11586 ( .A(n8284), .B(n8283), .Z(n8288) );
  NANDN U11587 ( .A(n8286), .B(n8285), .Z(n8287) );
  AND U11588 ( .A(n8288), .B(n8287), .Z(n10468) );
  NANDN U11589 ( .A(n8290), .B(n8289), .Z(n8294) );
  NANDN U11590 ( .A(n8292), .B(n8291), .Z(n8293) );
  AND U11591 ( .A(n8294), .B(n8293), .Z(n10467) );
  NANDN U11592 ( .A(n8296), .B(n8295), .Z(n8300) );
  NAND U11593 ( .A(n8298), .B(n8297), .Z(n8299) );
  AND U11594 ( .A(n8300), .B(n8299), .Z(n10013) );
  NAND U11595 ( .A(n8302), .B(n8301), .Z(n8306) );
  NAND U11596 ( .A(n8304), .B(n8303), .Z(n8305) );
  AND U11597 ( .A(n8306), .B(n8305), .Z(n10012) );
  NAND U11598 ( .A(n8308), .B(n8307), .Z(n8312) );
  NAND U11599 ( .A(n8310), .B(n8309), .Z(n8311) );
  NAND U11600 ( .A(n8312), .B(n8311), .Z(n10011) );
  XOR U11601 ( .A(n10012), .B(n10011), .Z(n10014) );
  XNOR U11602 ( .A(n10013), .B(n10014), .Z(n10466) );
  XOR U11603 ( .A(n10467), .B(n10466), .Z(n10469) );
  XOR U11604 ( .A(n10468), .B(n10469), .Z(n9078) );
  NANDN U11605 ( .A(n8314), .B(n8313), .Z(n8318) );
  NAND U11606 ( .A(n8316), .B(n8315), .Z(n8317) );
  AND U11607 ( .A(n8318), .B(n8317), .Z(n9180) );
  NANDN U11608 ( .A(n8320), .B(n8319), .Z(n8324) );
  NAND U11609 ( .A(n8322), .B(n8321), .Z(n8323) );
  AND U11610 ( .A(n8324), .B(n8323), .Z(n9179) );
  NANDN U11611 ( .A(n8326), .B(n8325), .Z(n8330) );
  NAND U11612 ( .A(n8328), .B(n8327), .Z(n8329) );
  NAND U11613 ( .A(n8330), .B(n8329), .Z(n9178) );
  XOR U11614 ( .A(n9179), .B(n9178), .Z(n9181) );
  XOR U11615 ( .A(n9180), .B(n9181), .Z(n10025) );
  NANDN U11616 ( .A(n8332), .B(n8331), .Z(n8336) );
  NAND U11617 ( .A(n8334), .B(n8333), .Z(n8335) );
  AND U11618 ( .A(n8336), .B(n8335), .Z(n10024) );
  NANDN U11619 ( .A(n8338), .B(n8337), .Z(n8342) );
  NAND U11620 ( .A(n8340), .B(n8339), .Z(n8341) );
  AND U11621 ( .A(n8342), .B(n8341), .Z(n10043) );
  NAND U11622 ( .A(n8344), .B(n8343), .Z(n8348) );
  NAND U11623 ( .A(n8346), .B(n8345), .Z(n8347) );
  AND U11624 ( .A(n8348), .B(n8347), .Z(n10042) );
  NANDN U11625 ( .A(n8350), .B(n8349), .Z(n8354) );
  NAND U11626 ( .A(n8352), .B(n8351), .Z(n8353) );
  NAND U11627 ( .A(n8354), .B(n8353), .Z(n10041) );
  XOR U11628 ( .A(n10042), .B(n10041), .Z(n10044) );
  XNOR U11629 ( .A(n10043), .B(n10044), .Z(n10023) );
  XOR U11630 ( .A(n10024), .B(n10023), .Z(n10026) );
  XOR U11631 ( .A(n10025), .B(n10026), .Z(n9077) );
  NANDN U11632 ( .A(n8356), .B(n8355), .Z(n8360) );
  NAND U11633 ( .A(n8358), .B(n8357), .Z(n8359) );
  AND U11634 ( .A(n8360), .B(n8359), .Z(n10396) );
  NANDN U11635 ( .A(n8362), .B(n8361), .Z(n8366) );
  OR U11636 ( .A(n8364), .B(n8363), .Z(n8365) );
  AND U11637 ( .A(n8366), .B(n8365), .Z(n10395) );
  NAND U11638 ( .A(n8368), .B(n8367), .Z(n8372) );
  NAND U11639 ( .A(n8370), .B(n8369), .Z(n8371) );
  AND U11640 ( .A(n8372), .B(n8371), .Z(n9621) );
  NAND U11641 ( .A(n8374), .B(n8373), .Z(n8378) );
  NAND U11642 ( .A(n8376), .B(n8375), .Z(n8377) );
  AND U11643 ( .A(n8378), .B(n8377), .Z(n9620) );
  NANDN U11644 ( .A(n8380), .B(n8379), .Z(n8384) );
  NANDN U11645 ( .A(n8382), .B(n8381), .Z(n8383) );
  NAND U11646 ( .A(n8384), .B(n8383), .Z(n9619) );
  XOR U11647 ( .A(n9620), .B(n9619), .Z(n9622) );
  XNOR U11648 ( .A(n9621), .B(n9622), .Z(n10394) );
  XOR U11649 ( .A(n10395), .B(n10394), .Z(n10397) );
  XNOR U11650 ( .A(n10396), .B(n10397), .Z(n9076) );
  XOR U11651 ( .A(n9077), .B(n9076), .Z(n9079) );
  XNOR U11652 ( .A(n9078), .B(n9079), .Z(n9788) );
  XNOR U11653 ( .A(n9789), .B(n9788), .Z(n9791) );
  NAND U11654 ( .A(n8386), .B(n8385), .Z(n8390) );
  NAND U11655 ( .A(n8388), .B(n8387), .Z(n8389) );
  NAND U11656 ( .A(n8390), .B(n8389), .Z(n9515) );
  NANDN U11657 ( .A(n8392), .B(n8391), .Z(n8396) );
  NAND U11658 ( .A(n8394), .B(n8393), .Z(n8395) );
  NAND U11659 ( .A(n8396), .B(n8395), .Z(n9514) );
  NANDN U11660 ( .A(n8398), .B(n8397), .Z(n8402) );
  NAND U11661 ( .A(n8400), .B(n8399), .Z(n8401) );
  NAND U11662 ( .A(n8402), .B(n8401), .Z(n9513) );
  XOR U11663 ( .A(n9514), .B(n9513), .Z(n9516) );
  XOR U11664 ( .A(n9515), .B(n9516), .Z(n9582) );
  NANDN U11665 ( .A(n8404), .B(n8403), .Z(n8408) );
  NAND U11666 ( .A(n8406), .B(n8405), .Z(n8407) );
  NAND U11667 ( .A(n8408), .B(n8407), .Z(n9186) );
  NAND U11668 ( .A(n8410), .B(n8409), .Z(n8414) );
  NAND U11669 ( .A(n8412), .B(n8411), .Z(n8413) );
  NAND U11670 ( .A(n8414), .B(n8413), .Z(n9185) );
  NANDN U11671 ( .A(n8416), .B(n8415), .Z(n8420) );
  NAND U11672 ( .A(n8418), .B(n8417), .Z(n8419) );
  NAND U11673 ( .A(n8420), .B(n8419), .Z(n9184) );
  XOR U11674 ( .A(n9185), .B(n9184), .Z(n9187) );
  XOR U11675 ( .A(n9186), .B(n9187), .Z(n9580) );
  NANDN U11676 ( .A(n8422), .B(n8421), .Z(n8426) );
  NAND U11677 ( .A(n8424), .B(n8423), .Z(n8425) );
  NAND U11678 ( .A(n8426), .B(n8425), .Z(n9509) );
  NANDN U11679 ( .A(n8428), .B(n8427), .Z(n8432) );
  NAND U11680 ( .A(n8430), .B(n8429), .Z(n8431) );
  NAND U11681 ( .A(n8432), .B(n8431), .Z(n9508) );
  NAND U11682 ( .A(n8434), .B(n8433), .Z(n8438) );
  NAND U11683 ( .A(n8436), .B(n8435), .Z(n8437) );
  NAND U11684 ( .A(n8438), .B(n8437), .Z(n9507) );
  XOR U11685 ( .A(n9508), .B(n9507), .Z(n9510) );
  XOR U11686 ( .A(n9509), .B(n9510), .Z(n9579) );
  XOR U11687 ( .A(n9580), .B(n9579), .Z(n9581) );
  XOR U11688 ( .A(n9582), .B(n9581), .Z(n9309) );
  NANDN U11689 ( .A(n8440), .B(n8439), .Z(n8444) );
  NAND U11690 ( .A(n8442), .B(n8441), .Z(n8443) );
  AND U11691 ( .A(n8444), .B(n8443), .Z(n10020) );
  NANDN U11692 ( .A(n8446), .B(n8445), .Z(n8450) );
  NAND U11693 ( .A(n8448), .B(n8447), .Z(n8449) );
  AND U11694 ( .A(n8450), .B(n8449), .Z(n10018) );
  NANDN U11695 ( .A(n8452), .B(n8451), .Z(n8456) );
  NAND U11696 ( .A(n8454), .B(n8453), .Z(n8455) );
  AND U11697 ( .A(n8456), .B(n8455), .Z(n9989) );
  NANDN U11698 ( .A(n8458), .B(n8457), .Z(n8462) );
  NAND U11699 ( .A(n8460), .B(n8459), .Z(n8461) );
  AND U11700 ( .A(n8462), .B(n8461), .Z(n9988) );
  NANDN U11701 ( .A(n8464), .B(n8463), .Z(n8468) );
  NAND U11702 ( .A(n8466), .B(n8465), .Z(n8467) );
  NAND U11703 ( .A(n8468), .B(n8467), .Z(n9987) );
  XOR U11704 ( .A(n9988), .B(n9987), .Z(n9990) );
  XNOR U11705 ( .A(n9989), .B(n9990), .Z(n10017) );
  XNOR U11706 ( .A(n10018), .B(n10017), .Z(n10019) );
  XNOR U11707 ( .A(n10020), .B(n10019), .Z(n9308) );
  XNOR U11708 ( .A(n9309), .B(n9308), .Z(n9310) );
  NANDN U11709 ( .A(n8470), .B(n8469), .Z(n8474) );
  NANDN U11710 ( .A(n8472), .B(n8471), .Z(n8473) );
  AND U11711 ( .A(n8474), .B(n8473), .Z(n9852) );
  NANDN U11712 ( .A(n8476), .B(n8475), .Z(n8480) );
  NAND U11713 ( .A(n8478), .B(n8477), .Z(n8479) );
  NAND U11714 ( .A(n8480), .B(n8479), .Z(n9174) );
  NAND U11715 ( .A(n8482), .B(n8481), .Z(n8486) );
  NAND U11716 ( .A(n8484), .B(n8483), .Z(n8485) );
  NAND U11717 ( .A(n8486), .B(n8485), .Z(n9173) );
  NANDN U11718 ( .A(n8488), .B(n8487), .Z(n8492) );
  NAND U11719 ( .A(n8490), .B(n8489), .Z(n8491) );
  NAND U11720 ( .A(n8492), .B(n8491), .Z(n9172) );
  XOR U11721 ( .A(n9173), .B(n9172), .Z(n9175) );
  XNOR U11722 ( .A(n9174), .B(n9175), .Z(n9850) );
  NANDN U11723 ( .A(n8494), .B(n8493), .Z(n8498) );
  NAND U11724 ( .A(n8496), .B(n8495), .Z(n8497) );
  NAND U11725 ( .A(n8498), .B(n8497), .Z(n10049) );
  NANDN U11726 ( .A(n8500), .B(n8499), .Z(n8504) );
  NAND U11727 ( .A(n8502), .B(n8501), .Z(n8503) );
  NAND U11728 ( .A(n8504), .B(n8503), .Z(n10048) );
  NANDN U11729 ( .A(n8506), .B(n8505), .Z(n8510) );
  NAND U11730 ( .A(n8508), .B(n8507), .Z(n8509) );
  NAND U11731 ( .A(n8510), .B(n8509), .Z(n10047) );
  XNOR U11732 ( .A(n10048), .B(n10047), .Z(n10050) );
  XOR U11733 ( .A(n10049), .B(n10050), .Z(n9849) );
  XOR U11734 ( .A(n9850), .B(n9849), .Z(n9851) );
  XOR U11735 ( .A(n9852), .B(n9851), .Z(n9311) );
  XNOR U11736 ( .A(n9310), .B(n9311), .Z(n9790) );
  XNOR U11737 ( .A(n9791), .B(n9790), .Z(n9358) );
  NANDN U11738 ( .A(n8512), .B(n8511), .Z(n8516) );
  NANDN U11739 ( .A(n8514), .B(n8513), .Z(n8515) );
  AND U11740 ( .A(n8516), .B(n8515), .Z(n9088) );
  NANDN U11741 ( .A(n8518), .B(n8517), .Z(n8522) );
  NAND U11742 ( .A(n8520), .B(n8519), .Z(n8521) );
  AND U11743 ( .A(n8522), .B(n8521), .Z(n9924) );
  NANDN U11744 ( .A(n8524), .B(n8523), .Z(n8528) );
  NAND U11745 ( .A(n8526), .B(n8525), .Z(n8527) );
  NAND U11746 ( .A(n8528), .B(n8527), .Z(n10169) );
  NANDN U11747 ( .A(n8530), .B(n8529), .Z(n8534) );
  NAND U11748 ( .A(n8532), .B(n8531), .Z(n8533) );
  NAND U11749 ( .A(n8534), .B(n8533), .Z(n10168) );
  NANDN U11750 ( .A(n8536), .B(n8535), .Z(n8540) );
  NAND U11751 ( .A(n8538), .B(n8537), .Z(n8539) );
  NAND U11752 ( .A(n8540), .B(n8539), .Z(n10167) );
  XOR U11753 ( .A(n10168), .B(n10167), .Z(n10170) );
  XNOR U11754 ( .A(n10169), .B(n10170), .Z(n9922) );
  NANDN U11755 ( .A(n8542), .B(n8541), .Z(n8546) );
  NAND U11756 ( .A(n8544), .B(n8543), .Z(n8545) );
  NAND U11757 ( .A(n8546), .B(n8545), .Z(n9947) );
  NANDN U11758 ( .A(n8548), .B(n8547), .Z(n8552) );
  NAND U11759 ( .A(n8550), .B(n8549), .Z(n8551) );
  NAND U11760 ( .A(n8552), .B(n8551), .Z(n9946) );
  NANDN U11761 ( .A(n8554), .B(n8553), .Z(n8558) );
  NAND U11762 ( .A(n8556), .B(n8555), .Z(n8557) );
  NAND U11763 ( .A(n8558), .B(n8557), .Z(n9945) );
  XNOR U11764 ( .A(n9946), .B(n9945), .Z(n9948) );
  XOR U11765 ( .A(n9947), .B(n9948), .Z(n9921) );
  XOR U11766 ( .A(n9922), .B(n9921), .Z(n9923) );
  XOR U11767 ( .A(n9924), .B(n9923), .Z(n9089) );
  XNOR U11768 ( .A(n9088), .B(n9089), .Z(n9091) );
  NANDN U11769 ( .A(n8560), .B(n8559), .Z(n8564) );
  NAND U11770 ( .A(n8562), .B(n8561), .Z(n8563) );
  AND U11771 ( .A(n8564), .B(n8563), .Z(n10321) );
  NANDN U11772 ( .A(n8566), .B(n8565), .Z(n8570) );
  NAND U11773 ( .A(n8568), .B(n8567), .Z(n8569) );
  AND U11774 ( .A(n8570), .B(n8569), .Z(n10319) );
  NANDN U11775 ( .A(n8572), .B(n8571), .Z(n8576) );
  NAND U11776 ( .A(n8574), .B(n8573), .Z(n8575) );
  NAND U11777 ( .A(n8576), .B(n8575), .Z(n10278) );
  NANDN U11778 ( .A(n8578), .B(n8577), .Z(n8582) );
  NAND U11779 ( .A(n8580), .B(n8579), .Z(n8581) );
  NAND U11780 ( .A(n8582), .B(n8581), .Z(n10277) );
  NANDN U11781 ( .A(n8584), .B(n8583), .Z(n8588) );
  NAND U11782 ( .A(n8586), .B(n8585), .Z(n8587) );
  NAND U11783 ( .A(n8588), .B(n8587), .Z(n10276) );
  XNOR U11784 ( .A(n10277), .B(n10276), .Z(n10279) );
  XOR U11785 ( .A(n10278), .B(n10279), .Z(n10318) );
  XNOR U11786 ( .A(n10319), .B(n10318), .Z(n10320) );
  XNOR U11787 ( .A(n10321), .B(n10320), .Z(n9090) );
  XNOR U11788 ( .A(n9091), .B(n9090), .Z(n9779) );
  NANDN U11789 ( .A(n8590), .B(n8589), .Z(n8594) );
  NAND U11790 ( .A(n8592), .B(n8591), .Z(n8593) );
  AND U11791 ( .A(n8594), .B(n8593), .Z(n9328) );
  NANDN U11792 ( .A(n8596), .B(n8595), .Z(n8600) );
  NAND U11793 ( .A(n8598), .B(n8597), .Z(n8599) );
  AND U11794 ( .A(n8600), .B(n8599), .Z(n9327) );
  NANDN U11795 ( .A(n8602), .B(n8601), .Z(n8606) );
  NANDN U11796 ( .A(n8604), .B(n8603), .Z(n8605) );
  AND U11797 ( .A(n8606), .B(n8605), .Z(n10212) );
  NANDN U11798 ( .A(n8608), .B(n8607), .Z(n8612) );
  NANDN U11799 ( .A(n8610), .B(n8609), .Z(n8611) );
  AND U11800 ( .A(n8612), .B(n8611), .Z(n10210) );
  NANDN U11801 ( .A(n8614), .B(n8613), .Z(n8618) );
  NAND U11802 ( .A(n8616), .B(n8615), .Z(n8617) );
  AND U11803 ( .A(n8618), .B(n8617), .Z(n9959) );
  NANDN U11804 ( .A(n8620), .B(n8619), .Z(n8624) );
  NAND U11805 ( .A(n8622), .B(n8621), .Z(n8623) );
  AND U11806 ( .A(n8624), .B(n8623), .Z(n9958) );
  NANDN U11807 ( .A(n8626), .B(n8625), .Z(n8630) );
  NAND U11808 ( .A(n8628), .B(n8627), .Z(n8629) );
  NAND U11809 ( .A(n8630), .B(n8629), .Z(n9957) );
  XOR U11810 ( .A(n9958), .B(n9957), .Z(n9960) );
  XNOR U11811 ( .A(n9959), .B(n9960), .Z(n10209) );
  XNOR U11812 ( .A(n10210), .B(n10209), .Z(n10211) );
  XNOR U11813 ( .A(n10212), .B(n10211), .Z(n9326) );
  XOR U11814 ( .A(n9327), .B(n9326), .Z(n9329) );
  XNOR U11815 ( .A(n9328), .B(n9329), .Z(n9777) );
  NAND U11816 ( .A(n8632), .B(n8631), .Z(n8636) );
  NAND U11817 ( .A(n8634), .B(n8633), .Z(n8635) );
  AND U11818 ( .A(n8636), .B(n8635), .Z(n9776) );
  XOR U11819 ( .A(n9777), .B(n9776), .Z(n9778) );
  XOR U11820 ( .A(n9779), .B(n9778), .Z(n9357) );
  XOR U11821 ( .A(n9358), .B(n9357), .Z(n9359) );
  XNOR U11822 ( .A(n9360), .B(n9359), .Z(n9395) );
  NAND U11823 ( .A(n8638), .B(n8637), .Z(n8642) );
  NAND U11824 ( .A(n8640), .B(n8639), .Z(n8641) );
  AND U11825 ( .A(n8642), .B(n8641), .Z(n9354) );
  NAND U11826 ( .A(n8644), .B(n8643), .Z(n8648) );
  NAND U11827 ( .A(n8646), .B(n8645), .Z(n8647) );
  NAND U11828 ( .A(n8648), .B(n8647), .Z(n9352) );
  NAND U11829 ( .A(n8650), .B(n8649), .Z(n8654) );
  NAND U11830 ( .A(n8652), .B(n8651), .Z(n8653) );
  AND U11831 ( .A(n8654), .B(n8653), .Z(n10382) );
  NANDN U11832 ( .A(n8656), .B(n8655), .Z(n8660) );
  NAND U11833 ( .A(n8658), .B(n8657), .Z(n8659) );
  AND U11834 ( .A(n8660), .B(n8659), .Z(n10421) );
  NANDN U11835 ( .A(n8662), .B(n8661), .Z(n8666) );
  OR U11836 ( .A(n8664), .B(n8663), .Z(n8665) );
  AND U11837 ( .A(n8666), .B(n8665), .Z(n10419) );
  NAND U11838 ( .A(n8668), .B(n8667), .Z(n8672) );
  NAND U11839 ( .A(n8670), .B(n8669), .Z(n8671) );
  AND U11840 ( .A(n8672), .B(n8671), .Z(n10001) );
  NANDN U11841 ( .A(n8674), .B(n8673), .Z(n8678) );
  NAND U11842 ( .A(n8676), .B(n8675), .Z(n8677) );
  AND U11843 ( .A(n8678), .B(n8677), .Z(n10000) );
  NAND U11844 ( .A(n8680), .B(n8679), .Z(n8684) );
  NAND U11845 ( .A(n8682), .B(n8681), .Z(n8683) );
  NAND U11846 ( .A(n8684), .B(n8683), .Z(n9999) );
  XOR U11847 ( .A(n10000), .B(n9999), .Z(n10002) );
  XNOR U11848 ( .A(n10001), .B(n10002), .Z(n10418) );
  XNOR U11849 ( .A(n10419), .B(n10418), .Z(n10420) );
  XNOR U11850 ( .A(n10421), .B(n10420), .Z(n9292) );
  NANDN U11851 ( .A(n8686), .B(n8685), .Z(n8690) );
  NAND U11852 ( .A(n8688), .B(n8687), .Z(n8689) );
  AND U11853 ( .A(n8690), .B(n8689), .Z(n9521) );
  NANDN U11854 ( .A(n8692), .B(n8691), .Z(n8696) );
  NAND U11855 ( .A(n8694), .B(n8693), .Z(n8695) );
  AND U11856 ( .A(n8696), .B(n8695), .Z(n9520) );
  NANDN U11857 ( .A(n8698), .B(n8697), .Z(n8702) );
  NAND U11858 ( .A(n8700), .B(n8699), .Z(n8701) );
  NAND U11859 ( .A(n8702), .B(n8701), .Z(n9519) );
  XOR U11860 ( .A(n9520), .B(n9519), .Z(n9522) );
  XOR U11861 ( .A(n9521), .B(n9522), .Z(n10164) );
  NANDN U11862 ( .A(n8704), .B(n8703), .Z(n8708) );
  NAND U11863 ( .A(n8706), .B(n8705), .Z(n8707) );
  AND U11864 ( .A(n8708), .B(n8707), .Z(n9664) );
  NAND U11865 ( .A(n8710), .B(n8709), .Z(n8714) );
  NAND U11866 ( .A(n8712), .B(n8711), .Z(n8713) );
  AND U11867 ( .A(n8714), .B(n8713), .Z(n9663) );
  NANDN U11868 ( .A(n8716), .B(n8715), .Z(n8720) );
  NAND U11869 ( .A(n8718), .B(n8717), .Z(n8719) );
  NAND U11870 ( .A(n8720), .B(n8719), .Z(n9662) );
  XOR U11871 ( .A(n9663), .B(n9662), .Z(n9665) );
  XOR U11872 ( .A(n9664), .B(n9665), .Z(n10162) );
  NANDN U11873 ( .A(n8722), .B(n8721), .Z(n8726) );
  NAND U11874 ( .A(n8724), .B(n8723), .Z(n8725) );
  AND U11875 ( .A(n8726), .B(n8725), .Z(n10091) );
  NANDN U11876 ( .A(n8728), .B(n8727), .Z(n8732) );
  NAND U11877 ( .A(n8730), .B(n8729), .Z(n8731) );
  AND U11878 ( .A(n8732), .B(n8731), .Z(n10090) );
  NANDN U11879 ( .A(n8734), .B(n8733), .Z(n8738) );
  NAND U11880 ( .A(n8736), .B(n8735), .Z(n8737) );
  NAND U11881 ( .A(n8738), .B(n8737), .Z(n10089) );
  XOR U11882 ( .A(n10090), .B(n10089), .Z(n10092) );
  XNOR U11883 ( .A(n10091), .B(n10092), .Z(n10161) );
  XNOR U11884 ( .A(n10162), .B(n10161), .Z(n10163) );
  XOR U11885 ( .A(n10164), .B(n10163), .Z(n9293) );
  XNOR U11886 ( .A(n9292), .B(n9293), .Z(n9294) );
  NANDN U11887 ( .A(n8740), .B(n8739), .Z(n8744) );
  NAND U11888 ( .A(n8742), .B(n8741), .Z(n8743) );
  AND U11889 ( .A(n8744), .B(n8743), .Z(n9725) );
  NANDN U11890 ( .A(n8746), .B(n8745), .Z(n8750) );
  NAND U11891 ( .A(n8748), .B(n8747), .Z(n8749) );
  AND U11892 ( .A(n8750), .B(n8749), .Z(n10284) );
  NANDN U11893 ( .A(n8752), .B(n8751), .Z(n8756) );
  NAND U11894 ( .A(n8754), .B(n8753), .Z(n8755) );
  AND U11895 ( .A(n8756), .B(n8755), .Z(n10283) );
  NANDN U11896 ( .A(n8758), .B(n8757), .Z(n8762) );
  NAND U11897 ( .A(n8760), .B(n8759), .Z(n8761) );
  NAND U11898 ( .A(n8762), .B(n8761), .Z(n10282) );
  XOR U11899 ( .A(n10283), .B(n10282), .Z(n10285) );
  XOR U11900 ( .A(n10284), .B(n10285), .Z(n9723) );
  NANDN U11901 ( .A(n8764), .B(n8763), .Z(n8768) );
  NAND U11902 ( .A(n8766), .B(n8765), .Z(n8767) );
  AND U11903 ( .A(n8768), .B(n8767), .Z(n10302) );
  NANDN U11904 ( .A(n8770), .B(n8769), .Z(n8774) );
  NAND U11905 ( .A(n8772), .B(n8771), .Z(n8773) );
  AND U11906 ( .A(n8774), .B(n8773), .Z(n10301) );
  NANDN U11907 ( .A(n8776), .B(n8775), .Z(n8780) );
  NAND U11908 ( .A(n8778), .B(n8777), .Z(n8779) );
  NAND U11909 ( .A(n8780), .B(n8779), .Z(n10300) );
  XOR U11910 ( .A(n10301), .B(n10300), .Z(n10303) );
  XNOR U11911 ( .A(n10302), .B(n10303), .Z(n9722) );
  XNOR U11912 ( .A(n9723), .B(n9722), .Z(n9724) );
  XOR U11913 ( .A(n9725), .B(n9724), .Z(n9295) );
  XNOR U11914 ( .A(n9294), .B(n9295), .Z(n10383) );
  XOR U11915 ( .A(n10382), .B(n10383), .Z(n10385) );
  NANDN U11916 ( .A(n8782), .B(n8781), .Z(n8786) );
  OR U11917 ( .A(n8784), .B(n8783), .Z(n8785) );
  AND U11918 ( .A(n8786), .B(n8785), .Z(n10499) );
  NANDN U11919 ( .A(n8788), .B(n8787), .Z(n8792) );
  OR U11920 ( .A(n8790), .B(n8789), .Z(n8791) );
  AND U11921 ( .A(n8792), .B(n8791), .Z(n10497) );
  NANDN U11922 ( .A(n8794), .B(n8793), .Z(n8798) );
  NAND U11923 ( .A(n8796), .B(n8795), .Z(n8797) );
  AND U11924 ( .A(n8798), .B(n8797), .Z(n9983) );
  NANDN U11925 ( .A(n8800), .B(n8799), .Z(n8804) );
  NAND U11926 ( .A(n8802), .B(n8801), .Z(n8803) );
  AND U11927 ( .A(n8804), .B(n8803), .Z(n9982) );
  NANDN U11928 ( .A(n8806), .B(n8805), .Z(n8810) );
  NAND U11929 ( .A(n8808), .B(n8807), .Z(n8809) );
  NAND U11930 ( .A(n8810), .B(n8809), .Z(n9981) );
  XOR U11931 ( .A(n9982), .B(n9981), .Z(n9984) );
  XNOR U11932 ( .A(n9983), .B(n9984), .Z(n10496) );
  XNOR U11933 ( .A(n10497), .B(n10496), .Z(n10498) );
  XNOR U11934 ( .A(n10499), .B(n10498), .Z(n9314) );
  NANDN U11935 ( .A(n8812), .B(n8811), .Z(n8816) );
  OR U11936 ( .A(n8814), .B(n8813), .Z(n8815) );
  AND U11937 ( .A(n8816), .B(n8815), .Z(n9205) );
  NANDN U11938 ( .A(n8818), .B(n8817), .Z(n8822) );
  NANDN U11939 ( .A(n8820), .B(n8819), .Z(n8821) );
  AND U11940 ( .A(n8822), .B(n8821), .Z(n9203) );
  NANDN U11941 ( .A(n8824), .B(n8823), .Z(n8828) );
  NAND U11942 ( .A(n8826), .B(n8825), .Z(n8827) );
  NAND U11943 ( .A(n8828), .B(n8827), .Z(n9603) );
  NAND U11944 ( .A(n8830), .B(n8829), .Z(n8834) );
  NAND U11945 ( .A(n8832), .B(n8831), .Z(n8833) );
  NAND U11946 ( .A(n8834), .B(n8833), .Z(n9602) );
  NAND U11947 ( .A(n8836), .B(n8835), .Z(n8840) );
  NAND U11948 ( .A(n8838), .B(n8837), .Z(n8839) );
  NAND U11949 ( .A(n8840), .B(n8839), .Z(n9601) );
  XNOR U11950 ( .A(n9602), .B(n9601), .Z(n9604) );
  XOR U11951 ( .A(n9603), .B(n9604), .Z(n9202) );
  XNOR U11952 ( .A(n9203), .B(n9202), .Z(n9204) );
  XOR U11953 ( .A(n9205), .B(n9204), .Z(n9315) );
  XNOR U11954 ( .A(n9314), .B(n9315), .Z(n9316) );
  NANDN U11955 ( .A(n8842), .B(n8841), .Z(n8846) );
  OR U11956 ( .A(n8844), .B(n8843), .Z(n8845) );
  AND U11957 ( .A(n8846), .B(n8845), .Z(n10361) );
  NANDN U11958 ( .A(n8848), .B(n8847), .Z(n8852) );
  NAND U11959 ( .A(n8850), .B(n8849), .Z(n8851) );
  AND U11960 ( .A(n8852), .B(n8851), .Z(n10359) );
  NANDN U11961 ( .A(n8854), .B(n8853), .Z(n8858) );
  NAND U11962 ( .A(n8856), .B(n8855), .Z(n8857) );
  AND U11963 ( .A(n8858), .B(n8857), .Z(n9609) );
  NANDN U11964 ( .A(n8860), .B(n8859), .Z(n8864) );
  NAND U11965 ( .A(n8862), .B(n8861), .Z(n8863) );
  AND U11966 ( .A(n8864), .B(n8863), .Z(n9608) );
  NANDN U11967 ( .A(n8866), .B(n8865), .Z(n8870) );
  NAND U11968 ( .A(n8868), .B(n8867), .Z(n8869) );
  NAND U11969 ( .A(n8870), .B(n8869), .Z(n9607) );
  XOR U11970 ( .A(n9608), .B(n9607), .Z(n9610) );
  XNOR U11971 ( .A(n9609), .B(n9610), .Z(n10358) );
  XNOR U11972 ( .A(n10359), .B(n10358), .Z(n10360) );
  XOR U11973 ( .A(n10361), .B(n10360), .Z(n9317) );
  XNOR U11974 ( .A(n9316), .B(n9317), .Z(n10384) );
  XNOR U11975 ( .A(n10385), .B(n10384), .Z(n9351) );
  XOR U11976 ( .A(n9352), .B(n9351), .Z(n9353) );
  XNOR U11977 ( .A(n9354), .B(n9353), .Z(n9394) );
  NAND U11978 ( .A(n8872), .B(n8871), .Z(n8876) );
  NAND U11979 ( .A(n8874), .B(n8873), .Z(n8875) );
  AND U11980 ( .A(n8876), .B(n8875), .Z(n9366) );
  NANDN U11981 ( .A(n8878), .B(n8877), .Z(n8882) );
  NAND U11982 ( .A(n8880), .B(n8879), .Z(n8881) );
  AND U11983 ( .A(n8882), .B(n8881), .Z(n9425) );
  NAND U11984 ( .A(n8884), .B(n8883), .Z(n8888) );
  NAND U11985 ( .A(n8886), .B(n8885), .Z(n8887) );
  AND U11986 ( .A(n8888), .B(n8887), .Z(n9424) );
  NANDN U11987 ( .A(n8890), .B(n8889), .Z(n8894) );
  NAND U11988 ( .A(n8892), .B(n8891), .Z(n8893) );
  NAND U11989 ( .A(n8894), .B(n8893), .Z(n9423) );
  XOR U11990 ( .A(n9424), .B(n9423), .Z(n9426) );
  XOR U11991 ( .A(n9425), .B(n9426), .Z(n9627) );
  NANDN U11992 ( .A(n8896), .B(n8895), .Z(n8900) );
  OR U11993 ( .A(n8898), .B(n8897), .Z(n8899) );
  AND U11994 ( .A(n8900), .B(n8899), .Z(n9626) );
  NANDN U11995 ( .A(n8902), .B(n8901), .Z(n8906) );
  OR U11996 ( .A(n8904), .B(n8903), .Z(n8905) );
  AND U11997 ( .A(n8906), .B(n8905), .Z(n9646) );
  NANDN U11998 ( .A(n8907), .B(oglobal[1]), .Z(n8911) );
  NANDN U11999 ( .A(n8909), .B(n8908), .Z(n8910) );
  AND U12000 ( .A(n8911), .B(n8910), .Z(n9644) );
  NAND U12001 ( .A(n8913), .B(n8912), .Z(n8917) );
  NAND U12002 ( .A(n8915), .B(n8914), .Z(n8916) );
  AND U12003 ( .A(n8917), .B(n8916), .Z(n9643) );
  XNOR U12004 ( .A(n9644), .B(n9643), .Z(n9645) );
  XNOR U12005 ( .A(n9646), .B(n9645), .Z(n9625) );
  XOR U12006 ( .A(n9626), .B(n9625), .Z(n9628) );
  XNOR U12007 ( .A(n9627), .B(n9628), .Z(n9334) );
  NAND U12008 ( .A(n8919), .B(n8918), .Z(n8923) );
  NAND U12009 ( .A(n8921), .B(n8920), .Z(n8922) );
  AND U12010 ( .A(n8923), .B(n8922), .Z(n9430) );
  NANDN U12011 ( .A(n8925), .B(n8924), .Z(n8929) );
  NAND U12012 ( .A(n8927), .B(n8926), .Z(n8928) );
  NAND U12013 ( .A(n8929), .B(n8928), .Z(n9429) );
  XOR U12014 ( .A(oglobal[2]), .B(n9429), .Z(n9431) );
  XOR U12015 ( .A(n9430), .B(n9431), .Z(n9632) );
  NANDN U12016 ( .A(n8931), .B(n8930), .Z(n8935) );
  NANDN U12017 ( .A(n8933), .B(n8932), .Z(n8934) );
  AND U12018 ( .A(n8935), .B(n8934), .Z(n9631) );
  XNOR U12019 ( .A(n9632), .B(n9631), .Z(n9634) );
  NANDN U12020 ( .A(n8937), .B(n8936), .Z(n8941) );
  NAND U12021 ( .A(n8939), .B(n8938), .Z(n8940) );
  AND U12022 ( .A(n8941), .B(n8940), .Z(n9640) );
  NAND U12023 ( .A(n8943), .B(n8942), .Z(n8947) );
  NAND U12024 ( .A(n8945), .B(n8944), .Z(n8946) );
  AND U12025 ( .A(n8947), .B(n8946), .Z(n9637) );
  NAND U12026 ( .A(n8949), .B(n8948), .Z(n8953) );
  NAND U12027 ( .A(n8951), .B(n8950), .Z(n8952) );
  NAND U12028 ( .A(n8953), .B(n8952), .Z(n9638) );
  XNOR U12029 ( .A(n9637), .B(n9638), .Z(n9639) );
  XNOR U12030 ( .A(n9640), .B(n9639), .Z(n9633) );
  XOR U12031 ( .A(n9634), .B(n9633), .Z(n9333) );
  NANDN U12032 ( .A(n8955), .B(n8954), .Z(n8959) );
  NAND U12033 ( .A(n8957), .B(n8956), .Z(n8958) );
  NAND U12034 ( .A(n8959), .B(n8958), .Z(n9332) );
  XOR U12035 ( .A(n9333), .B(n9332), .Z(n8960) );
  XNOR U12036 ( .A(n9334), .B(n8960), .Z(n10391) );
  NAND U12037 ( .A(n8962), .B(n8961), .Z(n8966) );
  NAND U12038 ( .A(n8964), .B(n8963), .Z(n8965) );
  AND U12039 ( .A(n8966), .B(n8965), .Z(n10388) );
  NANDN U12040 ( .A(n8968), .B(n8967), .Z(n8972) );
  NAND U12041 ( .A(n8970), .B(n8969), .Z(n8971) );
  AND U12042 ( .A(n8972), .B(n8971), .Z(n9731) );
  NANDN U12043 ( .A(n8974), .B(n8973), .Z(n8978) );
  NAND U12044 ( .A(n8976), .B(n8975), .Z(n8977) );
  AND U12045 ( .A(n8978), .B(n8977), .Z(n9905) );
  NANDN U12046 ( .A(n8980), .B(n8979), .Z(n8984) );
  NAND U12047 ( .A(n8982), .B(n8981), .Z(n8983) );
  AND U12048 ( .A(n8984), .B(n8983), .Z(n9904) );
  NAND U12049 ( .A(n8986), .B(n8985), .Z(n8990) );
  NAND U12050 ( .A(n8988), .B(n8987), .Z(n8989) );
  NAND U12051 ( .A(n8990), .B(n8989), .Z(n9903) );
  XOR U12052 ( .A(n9904), .B(n9903), .Z(n9906) );
  XOR U12053 ( .A(n9905), .B(n9906), .Z(n9729) );
  NANDN U12054 ( .A(n8992), .B(n8991), .Z(n8996) );
  NAND U12055 ( .A(n8994), .B(n8993), .Z(n8995) );
  NAND U12056 ( .A(n8996), .B(n8995), .Z(n9728) );
  XNOR U12057 ( .A(n9729), .B(n9728), .Z(n9730) );
  XNOR U12058 ( .A(n9731), .B(n9730), .Z(n9302) );
  NANDN U12059 ( .A(n8998), .B(n8997), .Z(n9002) );
  OR U12060 ( .A(n9000), .B(n8999), .Z(n9001) );
  AND U12061 ( .A(n9002), .B(n9001), .Z(n9534) );
  NANDN U12062 ( .A(n9004), .B(n9003), .Z(n9008) );
  OR U12063 ( .A(n9006), .B(n9005), .Z(n9007) );
  AND U12064 ( .A(n9008), .B(n9007), .Z(n9532) );
  NANDN U12065 ( .A(n9010), .B(n9009), .Z(n9014) );
  NAND U12066 ( .A(n9012), .B(n9011), .Z(n9013) );
  AND U12067 ( .A(n9014), .B(n9013), .Z(n9156) );
  NANDN U12068 ( .A(n9016), .B(n9015), .Z(n9020) );
  NAND U12069 ( .A(n9018), .B(n9017), .Z(n9019) );
  AND U12070 ( .A(n9020), .B(n9019), .Z(n9155) );
  NANDN U12071 ( .A(n9022), .B(n9021), .Z(n9026) );
  NAND U12072 ( .A(n9024), .B(n9023), .Z(n9025) );
  NAND U12073 ( .A(n9026), .B(n9025), .Z(n9154) );
  XOR U12074 ( .A(n9155), .B(n9154), .Z(n9157) );
  XNOR U12075 ( .A(n9156), .B(n9157), .Z(n9531) );
  XNOR U12076 ( .A(n9532), .B(n9531), .Z(n9533) );
  XOR U12077 ( .A(n9534), .B(n9533), .Z(n9303) );
  XNOR U12078 ( .A(n9302), .B(n9303), .Z(n9304) );
  NANDN U12079 ( .A(n9028), .B(n9027), .Z(n9032) );
  OR U12080 ( .A(n9030), .B(n9029), .Z(n9031) );
  AND U12081 ( .A(n9032), .B(n9031), .Z(n9491) );
  NANDN U12082 ( .A(n9034), .B(n9033), .Z(n9038) );
  OR U12083 ( .A(n9036), .B(n9035), .Z(n9037) );
  AND U12084 ( .A(n9038), .B(n9037), .Z(n9489) );
  NANDN U12085 ( .A(n9040), .B(n9039), .Z(n9044) );
  NAND U12086 ( .A(n9042), .B(n9041), .Z(n9043) );
  NAND U12087 ( .A(n9044), .B(n9043), .Z(n9893) );
  NANDN U12088 ( .A(n9046), .B(n9045), .Z(n9050) );
  NAND U12089 ( .A(n9048), .B(n9047), .Z(n9049) );
  NAND U12090 ( .A(n9050), .B(n9049), .Z(n9892) );
  NANDN U12091 ( .A(n9052), .B(n9051), .Z(n9056) );
  NAND U12092 ( .A(n9054), .B(n9053), .Z(n9055) );
  NAND U12093 ( .A(n9056), .B(n9055), .Z(n9891) );
  XNOR U12094 ( .A(n9892), .B(n9891), .Z(n9894) );
  XOR U12095 ( .A(n9893), .B(n9894), .Z(n9488) );
  XNOR U12096 ( .A(n9489), .B(n9488), .Z(n9490) );
  XOR U12097 ( .A(n9491), .B(n9490), .Z(n9305) );
  XNOR U12098 ( .A(n9304), .B(n9305), .Z(n10389) );
  XOR U12099 ( .A(n10388), .B(n10389), .Z(n10390) );
  XNOR U12100 ( .A(n10391), .B(n10390), .Z(n9363) );
  NAND U12101 ( .A(n9058), .B(n9057), .Z(n9062) );
  NAND U12102 ( .A(n9060), .B(n9059), .Z(n9061) );
  AND U12103 ( .A(n9062), .B(n9061), .Z(n9364) );
  XOR U12104 ( .A(n9363), .B(n9364), .Z(n9365) );
  XOR U12105 ( .A(n9366), .B(n9365), .Z(n9393) );
  XOR U12106 ( .A(n9394), .B(n9393), .Z(n9396) );
  XOR U12107 ( .A(n9395), .B(n9396), .Z(n10550) );
  XOR U12108 ( .A(n10551), .B(n10550), .Z(n10336) );
  XOR U12109 ( .A(n10337), .B(n10336), .Z(n10332) );
  XOR U12110 ( .A(n10331), .B(n10332), .Z(n9063) );
  XNOR U12111 ( .A(n10333), .B(n9063), .Z(o[2]) );
  NAND U12112 ( .A(n9065), .B(n9064), .Z(n9069) );
  NANDN U12113 ( .A(n9067), .B(n9066), .Z(n9068) );
  NAND U12114 ( .A(n9069), .B(n9068), .Z(n10562) );
  NAND U12115 ( .A(n9071), .B(n9070), .Z(n9075) );
  NANDN U12116 ( .A(n9073), .B(n9072), .Z(n9074) );
  NAND U12117 ( .A(n9075), .B(n9074), .Z(n10561) );
  XOR U12118 ( .A(n10562), .B(n10561), .Z(n10564) );
  NANDN U12119 ( .A(n9077), .B(n9076), .Z(n9081) );
  OR U12120 ( .A(n9079), .B(n9078), .Z(n9080) );
  AND U12121 ( .A(n9081), .B(n9080), .Z(n10594) );
  NANDN U12122 ( .A(n9083), .B(n9082), .Z(n9087) );
  NANDN U12123 ( .A(n9085), .B(n9084), .Z(n9086) );
  AND U12124 ( .A(n9087), .B(n9086), .Z(n10592) );
  NANDN U12125 ( .A(n9089), .B(n9088), .Z(n9093) );
  NAND U12126 ( .A(n9091), .B(n9090), .Z(n9092) );
  NAND U12127 ( .A(n9093), .B(n9092), .Z(n10591) );
  XNOR U12128 ( .A(n10592), .B(n10591), .Z(n10593) );
  XOR U12129 ( .A(n10594), .B(n10593), .Z(n11232) );
  NANDN U12130 ( .A(n9095), .B(n9094), .Z(n9099) );
  NANDN U12131 ( .A(n9097), .B(n9096), .Z(n9098) );
  AND U12132 ( .A(n9099), .B(n9098), .Z(n11231) );
  XNOR U12133 ( .A(n11232), .B(n11231), .Z(n11234) );
  NANDN U12134 ( .A(n9101), .B(n9100), .Z(n9105) );
  NAND U12135 ( .A(n9103), .B(n9102), .Z(n9104) );
  AND U12136 ( .A(n9105), .B(n9104), .Z(n11233) );
  XOR U12137 ( .A(n11234), .B(n11233), .Z(n10831) );
  NANDN U12138 ( .A(n9107), .B(n9106), .Z(n9111) );
  NAND U12139 ( .A(n9109), .B(n9108), .Z(n9110) );
  AND U12140 ( .A(n9111), .B(n9110), .Z(n10829) );
  NANDN U12141 ( .A(n9113), .B(n9112), .Z(n9117) );
  NANDN U12142 ( .A(n9115), .B(n9114), .Z(n9116) );
  AND U12143 ( .A(n9117), .B(n9116), .Z(n10729) );
  NANDN U12144 ( .A(n9119), .B(n9118), .Z(n9123) );
  NANDN U12145 ( .A(n9121), .B(n9120), .Z(n9122) );
  AND U12146 ( .A(n9123), .B(n9122), .Z(n10727) );
  NANDN U12147 ( .A(n9125), .B(n9124), .Z(n9129) );
  NANDN U12148 ( .A(n9127), .B(n9126), .Z(n9128) );
  AND U12149 ( .A(n9129), .B(n9128), .Z(n10753) );
  NANDN U12150 ( .A(n9131), .B(n9130), .Z(n9135) );
  NANDN U12151 ( .A(n9133), .B(n9132), .Z(n9134) );
  AND U12152 ( .A(n9135), .B(n9134), .Z(n10751) );
  NANDN U12153 ( .A(n9137), .B(n9136), .Z(n9141) );
  NANDN U12154 ( .A(n9139), .B(n9138), .Z(n9140) );
  NAND U12155 ( .A(n9141), .B(n9140), .Z(n10750) );
  XNOR U12156 ( .A(n10751), .B(n10750), .Z(n10752) );
  XNOR U12157 ( .A(n10753), .B(n10752), .Z(n10726) );
  XNOR U12158 ( .A(n10727), .B(n10726), .Z(n10728) );
  XNOR U12159 ( .A(n10729), .B(n10728), .Z(n10828) );
  NAND U12160 ( .A(n9143), .B(n9142), .Z(n9147) );
  NAND U12161 ( .A(n9145), .B(n9144), .Z(n9146) );
  AND U12162 ( .A(n9147), .B(n9146), .Z(n10835) );
  NANDN U12163 ( .A(n9149), .B(n9148), .Z(n9153) );
  NANDN U12164 ( .A(n9151), .B(n9150), .Z(n9152) );
  AND U12165 ( .A(n9153), .B(n9152), .Z(n10793) );
  NANDN U12166 ( .A(n9155), .B(n9154), .Z(n9159) );
  OR U12167 ( .A(n9157), .B(n9156), .Z(n9158) );
  AND U12168 ( .A(n9159), .B(n9158), .Z(n11158) );
  NANDN U12169 ( .A(n9161), .B(n9160), .Z(n9165) );
  OR U12170 ( .A(n9163), .B(n9162), .Z(n9164) );
  AND U12171 ( .A(n9165), .B(n9164), .Z(n11156) );
  NANDN U12172 ( .A(n9167), .B(n9166), .Z(n9171) );
  OR U12173 ( .A(n9169), .B(n9168), .Z(n9170) );
  NAND U12174 ( .A(n9171), .B(n9170), .Z(n11157) );
  XOR U12175 ( .A(n11156), .B(n11157), .Z(n11159) );
  XNOR U12176 ( .A(n11158), .B(n11159), .Z(n10792) );
  XNOR U12177 ( .A(n10793), .B(n10792), .Z(n10795) );
  NAND U12178 ( .A(n9173), .B(n9172), .Z(n9177) );
  NAND U12179 ( .A(n9175), .B(n9174), .Z(n9176) );
  AND U12180 ( .A(n9177), .B(n9176), .Z(n11087) );
  NANDN U12181 ( .A(n9179), .B(n9178), .Z(n9183) );
  OR U12182 ( .A(n9181), .B(n9180), .Z(n9182) );
  AND U12183 ( .A(n9183), .B(n9182), .Z(n11085) );
  NAND U12184 ( .A(n9185), .B(n9184), .Z(n9189) );
  NAND U12185 ( .A(n9187), .B(n9186), .Z(n9188) );
  NAND U12186 ( .A(n9189), .B(n9188), .Z(n11086) );
  XOR U12187 ( .A(n11085), .B(n11086), .Z(n11088) );
  XNOR U12188 ( .A(n11087), .B(n11088), .Z(n10794) );
  XOR U12189 ( .A(n10795), .B(n10794), .Z(n10581) );
  NANDN U12190 ( .A(n9191), .B(n9190), .Z(n9195) );
  NANDN U12191 ( .A(n9193), .B(n9192), .Z(n9194) );
  AND U12192 ( .A(n9195), .B(n9194), .Z(n10798) );
  NANDN U12193 ( .A(n9197), .B(n9196), .Z(n9201) );
  NANDN U12194 ( .A(n9199), .B(n9198), .Z(n9200) );
  NAND U12195 ( .A(n9201), .B(n9200), .Z(n10799) );
  XNOR U12196 ( .A(n10798), .B(n10799), .Z(n10800) );
  NANDN U12197 ( .A(n9203), .B(n9202), .Z(n9207) );
  NANDN U12198 ( .A(n9205), .B(n9204), .Z(n9206) );
  NAND U12199 ( .A(n9207), .B(n9206), .Z(n10801) );
  XNOR U12200 ( .A(n10800), .B(n10801), .Z(n10579) );
  NANDN U12201 ( .A(n9209), .B(n9208), .Z(n9213) );
  NANDN U12202 ( .A(n9211), .B(n9210), .Z(n9212) );
  NAND U12203 ( .A(n9213), .B(n9212), .Z(n10580) );
  XOR U12204 ( .A(n10579), .B(n10580), .Z(n10582) );
  XNOR U12205 ( .A(n10581), .B(n10582), .Z(n10777) );
  NAND U12206 ( .A(n9215), .B(n9214), .Z(n9219) );
  NAND U12207 ( .A(n9217), .B(n9216), .Z(n9218) );
  AND U12208 ( .A(n9219), .B(n9218), .Z(n10774) );
  NAND U12209 ( .A(n9221), .B(n9220), .Z(n9225) );
  NAND U12210 ( .A(n9223), .B(n9222), .Z(n9224) );
  AND U12211 ( .A(n9225), .B(n9224), .Z(n10775) );
  XOR U12212 ( .A(n10774), .B(n10775), .Z(n10776) );
  XOR U12213 ( .A(n10777), .B(n10776), .Z(n10834) );
  NAND U12214 ( .A(n9227), .B(n9226), .Z(n9231) );
  NAND U12215 ( .A(n9229), .B(n9228), .Z(n9230) );
  AND U12216 ( .A(n9231), .B(n9230), .Z(n10836) );
  XNOR U12217 ( .A(n10837), .B(n10836), .Z(n11262) );
  NAND U12218 ( .A(n9233), .B(n9232), .Z(n9237) );
  NAND U12219 ( .A(n9235), .B(n9234), .Z(n9236) );
  NAND U12220 ( .A(n9237), .B(n9236), .Z(n11261) );
  XOR U12221 ( .A(n11262), .B(n11261), .Z(n11264) );
  XOR U12222 ( .A(n11263), .B(n11264), .Z(n10563) );
  XOR U12223 ( .A(n10564), .B(n10563), .Z(n10555) );
  NAND U12224 ( .A(n9239), .B(n9238), .Z(n9243) );
  NAND U12225 ( .A(n9241), .B(n9240), .Z(n9242) );
  AND U12226 ( .A(n9243), .B(n9242), .Z(n10556) );
  XOR U12227 ( .A(n10555), .B(n10556), .Z(n10558) );
  NAND U12228 ( .A(n9245), .B(n9244), .Z(n9249) );
  NAND U12229 ( .A(n9247), .B(n9246), .Z(n9248) );
  NAND U12230 ( .A(n9249), .B(n9248), .Z(n10575) );
  NANDN U12231 ( .A(n9251), .B(n9250), .Z(n9255) );
  NAND U12232 ( .A(n9253), .B(n9252), .Z(n9254) );
  AND U12233 ( .A(n9255), .B(n9254), .Z(n10873) );
  NANDN U12234 ( .A(n9257), .B(n9256), .Z(n9261) );
  OR U12235 ( .A(n9259), .B(n9258), .Z(n9260) );
  AND U12236 ( .A(n9261), .B(n9260), .Z(n10871) );
  NANDN U12237 ( .A(n9263), .B(n9262), .Z(n9267) );
  OR U12238 ( .A(n9265), .B(n9264), .Z(n9266) );
  NAND U12239 ( .A(n9267), .B(n9266), .Z(n10870) );
  XNOR U12240 ( .A(n10871), .B(n10870), .Z(n10872) );
  XOR U12241 ( .A(n10873), .B(n10872), .Z(n10574) );
  NANDN U12242 ( .A(n9269), .B(n9268), .Z(n9273) );
  NAND U12243 ( .A(n9271), .B(n9270), .Z(n9272) );
  AND U12244 ( .A(n9273), .B(n9272), .Z(n10644) );
  NANDN U12245 ( .A(n9275), .B(n9274), .Z(n9279) );
  NAND U12246 ( .A(n9277), .B(n9276), .Z(n9278) );
  AND U12247 ( .A(n9279), .B(n9278), .Z(n10643) );
  NANDN U12248 ( .A(n9281), .B(n9280), .Z(n9285) );
  NAND U12249 ( .A(n9283), .B(n9282), .Z(n9284) );
  NAND U12250 ( .A(n9285), .B(n9284), .Z(n10642) );
  XOR U12251 ( .A(n10643), .B(n10642), .Z(n10645) );
  XNOR U12252 ( .A(n10644), .B(n10645), .Z(n10573) );
  XOR U12253 ( .A(n10574), .B(n10573), .Z(n10576) );
  XOR U12254 ( .A(n10575), .B(n10576), .Z(n10612) );
  NAND U12255 ( .A(n9287), .B(n9286), .Z(n9291) );
  NAND U12256 ( .A(n9289), .B(n9288), .Z(n9290) );
  NAND U12257 ( .A(n9291), .B(n9290), .Z(n10610) );
  NANDN U12258 ( .A(n9293), .B(n9292), .Z(n9297) );
  NANDN U12259 ( .A(n9295), .B(n9294), .Z(n9296) );
  AND U12260 ( .A(n9297), .B(n9296), .Z(n10823) );
  XNOR U12261 ( .A(n10823), .B(n10822), .Z(n10825) );
  NANDN U12262 ( .A(n9303), .B(n9302), .Z(n9307) );
  NANDN U12263 ( .A(n9305), .B(n9304), .Z(n9306) );
  AND U12264 ( .A(n9307), .B(n9306), .Z(n10588) );
  NANDN U12265 ( .A(n9309), .B(n9308), .Z(n9313) );
  NANDN U12266 ( .A(n9311), .B(n9310), .Z(n9312) );
  AND U12267 ( .A(n9313), .B(n9312), .Z(n10586) );
  NANDN U12268 ( .A(n9315), .B(n9314), .Z(n9319) );
  NANDN U12269 ( .A(n9317), .B(n9316), .Z(n9318) );
  NAND U12270 ( .A(n9319), .B(n9318), .Z(n10585) );
  XNOR U12271 ( .A(n10586), .B(n10585), .Z(n10587) );
  XNOR U12272 ( .A(n10588), .B(n10587), .Z(n10824) );
  XOR U12273 ( .A(n10825), .B(n10824), .Z(n11246) );
  NANDN U12274 ( .A(n9321), .B(n9320), .Z(n9325) );
  NANDN U12275 ( .A(n9323), .B(n9322), .Z(n9324) );
  AND U12276 ( .A(n9325), .B(n9324), .Z(n10650) );
  NANDN U12277 ( .A(n9327), .B(n9326), .Z(n9331) );
  OR U12278 ( .A(n9329), .B(n9328), .Z(n9330) );
  AND U12279 ( .A(n9331), .B(n9330), .Z(n10649) );
  XOR U12280 ( .A(n10649), .B(n10648), .Z(n10651) );
  XOR U12281 ( .A(n10650), .B(n10651), .Z(n11244) );
  NANDN U12282 ( .A(n9336), .B(n9335), .Z(n9340) );
  NANDN U12283 ( .A(n9338), .B(n9337), .Z(n9339) );
  AND U12284 ( .A(n9340), .B(n9339), .Z(n10680) );
  NANDN U12285 ( .A(n9342), .B(n9341), .Z(n9346) );
  NANDN U12286 ( .A(n9344), .B(n9343), .Z(n9345) );
  AND U12287 ( .A(n9346), .B(n9345), .Z(n10679) );
  XOR U12288 ( .A(n10679), .B(n10678), .Z(n10681) );
  XNOR U12289 ( .A(n10680), .B(n10681), .Z(n11243) );
  XNOR U12290 ( .A(n11244), .B(n11243), .Z(n11245) );
  XNOR U12291 ( .A(n11246), .B(n11245), .Z(n10609) );
  XOR U12292 ( .A(n10610), .B(n10609), .Z(n10611) );
  XNOR U12293 ( .A(n10612), .B(n10611), .Z(n11106) );
  NAND U12294 ( .A(n9352), .B(n9351), .Z(n9356) );
  NAND U12295 ( .A(n9354), .B(n9353), .Z(n9355) );
  NAND U12296 ( .A(n9356), .B(n9355), .Z(n10771) );
  NAND U12297 ( .A(n9358), .B(n9357), .Z(n9362) );
  NAND U12298 ( .A(n9360), .B(n9359), .Z(n9361) );
  NAND U12299 ( .A(n9362), .B(n9361), .Z(n10769) );
  NAND U12300 ( .A(n9364), .B(n9363), .Z(n9368) );
  NANDN U12301 ( .A(n9366), .B(n9365), .Z(n9367) );
  NAND U12302 ( .A(n9368), .B(n9367), .Z(n10768) );
  XOR U12303 ( .A(n10769), .B(n10768), .Z(n10770) );
  XNOR U12304 ( .A(n10771), .B(n10770), .Z(n11104) );
  NANDN U12305 ( .A(n9370), .B(n9369), .Z(n9374) );
  NANDN U12306 ( .A(n9372), .B(n9371), .Z(n9373) );
  AND U12307 ( .A(n9374), .B(n9373), .Z(n10570) );
  NAND U12308 ( .A(n9376), .B(n9375), .Z(n9380) );
  NANDN U12309 ( .A(n9378), .B(n9377), .Z(n9379) );
  AND U12310 ( .A(n9380), .B(n9379), .Z(n10568) );
  NANDN U12311 ( .A(n9382), .B(n9381), .Z(n9386) );
  NAND U12312 ( .A(n9384), .B(n9383), .Z(n9385) );
  NAND U12313 ( .A(n9386), .B(n9385), .Z(n10567) );
  XNOR U12314 ( .A(n10570), .B(n10569), .Z(n11103) );
  XOR U12315 ( .A(n11104), .B(n11103), .Z(n11105) );
  XNOR U12316 ( .A(n11106), .B(n11105), .Z(n10629) );
  NAND U12317 ( .A(n9388), .B(n9387), .Z(n9392) );
  NAND U12318 ( .A(n9390), .B(n9389), .Z(n9391) );
  NAND U12319 ( .A(n9392), .B(n9391), .Z(n11270) );
  NAND U12320 ( .A(n9394), .B(n9393), .Z(n9398) );
  NAND U12321 ( .A(n9396), .B(n9395), .Z(n9397) );
  AND U12322 ( .A(n9398), .B(n9397), .Z(n11268) );
  NANDN U12323 ( .A(n9400), .B(n9399), .Z(n9404) );
  NAND U12324 ( .A(n9402), .B(n9401), .Z(n9403) );
  AND U12325 ( .A(n9404), .B(n9403), .Z(n10723) );
  NANDN U12326 ( .A(n9406), .B(n9405), .Z(n9410) );
  NAND U12327 ( .A(n9408), .B(n9407), .Z(n9409) );
  AND U12328 ( .A(n9410), .B(n9409), .Z(n10721) );
  NANDN U12329 ( .A(n9412), .B(n9411), .Z(n9416) );
  NAND U12330 ( .A(n9414), .B(n9413), .Z(n9415) );
  NAND U12331 ( .A(n9416), .B(n9415), .Z(n10720) );
  XNOR U12332 ( .A(n10721), .B(n10720), .Z(n10722) );
  XNOR U12333 ( .A(n10723), .B(n10722), .Z(n10672) );
  NAND U12334 ( .A(n9418), .B(n9417), .Z(n9422) );
  NANDN U12335 ( .A(n9420), .B(n9419), .Z(n9421) );
  AND U12336 ( .A(n9422), .B(n9421), .Z(n11198) );
  NANDN U12337 ( .A(n9424), .B(n9423), .Z(n9428) );
  OR U12338 ( .A(n9426), .B(n9425), .Z(n9427) );
  NAND U12339 ( .A(n9428), .B(n9427), .Z(n11199) );
  XNOR U12340 ( .A(n11198), .B(n11199), .Z(n11201) );
  NANDN U12341 ( .A(oglobal[2]), .B(n9429), .Z(n9433) );
  OR U12342 ( .A(n9431), .B(n9430), .Z(n9432) );
  AND U12343 ( .A(n9433), .B(n9432), .Z(n11200) );
  XOR U12344 ( .A(n11201), .B(n11200), .Z(n11151) );
  NAND U12345 ( .A(n9435), .B(n9434), .Z(n9439) );
  NAND U12346 ( .A(n9437), .B(n9436), .Z(n9438) );
  AND U12347 ( .A(n9439), .B(n9438), .Z(n11150) );
  XNOR U12348 ( .A(n11151), .B(n11150), .Z(n11153) );
  NANDN U12349 ( .A(n9441), .B(n9440), .Z(n9445) );
  NANDN U12350 ( .A(n9443), .B(n9442), .Z(n9444) );
  AND U12351 ( .A(n9445), .B(n9444), .Z(n11152) );
  XOR U12352 ( .A(n11153), .B(n11152), .Z(n11058) );
  NANDN U12353 ( .A(n9447), .B(n9446), .Z(n9451) );
  NAND U12354 ( .A(n9449), .B(n9448), .Z(n9450) );
  AND U12355 ( .A(n9451), .B(n9450), .Z(n11056) );
  NANDN U12356 ( .A(n9453), .B(n9452), .Z(n9457) );
  OR U12357 ( .A(n9455), .B(n9454), .Z(n9456) );
  AND U12358 ( .A(n9457), .B(n9456), .Z(n11189) );
  NANDN U12359 ( .A(n9459), .B(n9458), .Z(n9463) );
  OR U12360 ( .A(n9461), .B(n9460), .Z(n9462) );
  AND U12361 ( .A(n9463), .B(n9462), .Z(n11186) );
  NANDN U12362 ( .A(n9465), .B(n9464), .Z(n9469) );
  OR U12363 ( .A(n9467), .B(n9466), .Z(n9468) );
  NAND U12364 ( .A(n9469), .B(n9468), .Z(n11187) );
  XNOR U12365 ( .A(n11186), .B(n11187), .Z(n11188) );
  XOR U12366 ( .A(n11189), .B(n11188), .Z(n10889) );
  NANDN U12367 ( .A(n9471), .B(n9470), .Z(n9475) );
  NANDN U12368 ( .A(n9473), .B(n9472), .Z(n9474) );
  AND U12369 ( .A(n9475), .B(n9474), .Z(n10888) );
  XNOR U12370 ( .A(n10889), .B(n10888), .Z(n10891) );
  NANDN U12371 ( .A(n9477), .B(n9476), .Z(n9481) );
  NANDN U12372 ( .A(n9479), .B(n9478), .Z(n9480) );
  AND U12373 ( .A(n9481), .B(n9480), .Z(n10890) );
  XNOR U12374 ( .A(n10891), .B(n10890), .Z(n11055) );
  XNOR U12375 ( .A(n11056), .B(n11055), .Z(n11057) );
  XNOR U12376 ( .A(n11058), .B(n11057), .Z(n10673) );
  XOR U12377 ( .A(n10672), .B(n10673), .Z(n10675) );
  NANDN U12378 ( .A(n9483), .B(n9482), .Z(n9487) );
  NAND U12379 ( .A(n9485), .B(n9484), .Z(n9486) );
  AND U12380 ( .A(n9487), .B(n9486), .Z(n11126) );
  NANDN U12381 ( .A(n9489), .B(n9488), .Z(n9493) );
  NANDN U12382 ( .A(n9491), .B(n9490), .Z(n9492) );
  NAND U12383 ( .A(n9493), .B(n9492), .Z(n11125) );
  NANDN U12384 ( .A(n9495), .B(n9494), .Z(n9499) );
  NANDN U12385 ( .A(n9497), .B(n9496), .Z(n9498) );
  AND U12386 ( .A(n9499), .B(n9498), .Z(n11124) );
  XOR U12387 ( .A(n11125), .B(n11124), .Z(n9500) );
  XNOR U12388 ( .A(n11126), .B(n9500), .Z(n10656) );
  NANDN U12389 ( .A(n9502), .B(n9501), .Z(n9506) );
  NANDN U12390 ( .A(n9504), .B(n9503), .Z(n9505) );
  AND U12391 ( .A(n9506), .B(n9505), .Z(n10655) );
  NAND U12392 ( .A(n9508), .B(n9507), .Z(n9512) );
  NAND U12393 ( .A(n9510), .B(n9509), .Z(n9511) );
  AND U12394 ( .A(n9512), .B(n9511), .Z(n11195) );
  NAND U12395 ( .A(n9514), .B(n9513), .Z(n9518) );
  NAND U12396 ( .A(n9516), .B(n9515), .Z(n9517) );
  AND U12397 ( .A(n9518), .B(n9517), .Z(n11192) );
  NANDN U12398 ( .A(n9520), .B(n9519), .Z(n9524) );
  OR U12399 ( .A(n9522), .B(n9521), .Z(n9523) );
  NAND U12400 ( .A(n9524), .B(n9523), .Z(n11193) );
  XNOR U12401 ( .A(n11192), .B(n11193), .Z(n11194) );
  XOR U12402 ( .A(n11195), .B(n11194), .Z(n10956) );
  NANDN U12403 ( .A(n9526), .B(n9525), .Z(n9530) );
  NANDN U12404 ( .A(n9528), .B(n9527), .Z(n9529) );
  AND U12405 ( .A(n9530), .B(n9529), .Z(n10954) );
  NANDN U12406 ( .A(n9532), .B(n9531), .Z(n9536) );
  NANDN U12407 ( .A(n9534), .B(n9533), .Z(n9535) );
  NAND U12408 ( .A(n9536), .B(n9535), .Z(n10955) );
  XOR U12409 ( .A(n10954), .B(n10955), .Z(n10957) );
  XNOR U12410 ( .A(n10956), .B(n10957), .Z(n10654) );
  XOR U12411 ( .A(n10655), .B(n10654), .Z(n10657) );
  XNOR U12412 ( .A(n10656), .B(n10657), .Z(n10674) );
  XNOR U12413 ( .A(n10675), .B(n10674), .Z(n10921) );
  NANDN U12414 ( .A(n9538), .B(n9537), .Z(n9542) );
  NAND U12415 ( .A(n9540), .B(n9539), .Z(n9541) );
  AND U12416 ( .A(n9542), .B(n9541), .Z(n11238) );
  NAND U12417 ( .A(n9544), .B(n9543), .Z(n9548) );
  NAND U12418 ( .A(n9546), .B(n9545), .Z(n9547) );
  AND U12419 ( .A(n9548), .B(n9547), .Z(n10967) );
  NANDN U12420 ( .A(n9550), .B(n9549), .Z(n9554) );
  NANDN U12421 ( .A(n9552), .B(n9551), .Z(n9553) );
  AND U12422 ( .A(n9554), .B(n9553), .Z(n10936) );
  NANDN U12423 ( .A(n9556), .B(n9555), .Z(n9560) );
  NANDN U12424 ( .A(n9558), .B(n9557), .Z(n9559) );
  NAND U12425 ( .A(n9560), .B(n9559), .Z(n10937) );
  XNOR U12426 ( .A(n10936), .B(n10937), .Z(n10939) );
  NANDN U12427 ( .A(n9562), .B(n9561), .Z(n9566) );
  NANDN U12428 ( .A(n9564), .B(n9563), .Z(n9565) );
  AND U12429 ( .A(n9566), .B(n9565), .Z(n10938) );
  XNOR U12430 ( .A(n10939), .B(n10938), .Z(n10966) );
  XNOR U12431 ( .A(n10967), .B(n10966), .Z(n10968) );
  NAND U12432 ( .A(n9568), .B(n9567), .Z(n9572) );
  NANDN U12433 ( .A(n9570), .B(n9569), .Z(n9571) );
  AND U12434 ( .A(n9572), .B(n9571), .Z(n11137) );
  NAND U12435 ( .A(n9574), .B(n9573), .Z(n9578) );
  NANDN U12436 ( .A(n9576), .B(n9575), .Z(n9577) );
  AND U12437 ( .A(n9578), .B(n9577), .Z(n11135) );
  XNOR U12438 ( .A(n11135), .B(n11134), .Z(n11136) );
  XOR U12439 ( .A(n11137), .B(n11136), .Z(n10969) );
  XNOR U12440 ( .A(n10968), .B(n10969), .Z(n11237) );
  XNOR U12441 ( .A(n11238), .B(n11237), .Z(n11240) );
  NANDN U12442 ( .A(n9584), .B(n9583), .Z(n9588) );
  OR U12443 ( .A(n9586), .B(n9585), .Z(n9587) );
  AND U12444 ( .A(n9588), .B(n9587), .Z(n11181) );
  NANDN U12445 ( .A(n9590), .B(n9589), .Z(n9594) );
  OR U12446 ( .A(n9592), .B(n9591), .Z(n9593) );
  NAND U12447 ( .A(n9594), .B(n9593), .Z(n11216) );
  XNOR U12448 ( .A(oglobal[3]), .B(n11216), .Z(n11217) );
  NANDN U12449 ( .A(n9596), .B(n9595), .Z(n9600) );
  OR U12450 ( .A(n9598), .B(n9597), .Z(n9599) );
  NAND U12451 ( .A(n9600), .B(n9599), .Z(n11218) );
  XNOR U12452 ( .A(n11217), .B(n11218), .Z(n11022) );
  NAND U12453 ( .A(n9602), .B(n9601), .Z(n9606) );
  NANDN U12454 ( .A(n9604), .B(n9603), .Z(n9605) );
  AND U12455 ( .A(n9606), .B(n9605), .Z(n11020) );
  NANDN U12456 ( .A(n9608), .B(n9607), .Z(n9612) );
  OR U12457 ( .A(n9610), .B(n9609), .Z(n9611) );
  AND U12458 ( .A(n9612), .B(n9611), .Z(n11212) );
  NANDN U12459 ( .A(n9614), .B(n9613), .Z(n9618) );
  OR U12460 ( .A(n9616), .B(n9615), .Z(n9617) );
  AND U12461 ( .A(n9618), .B(n9617), .Z(n11210) );
  NANDN U12462 ( .A(n9620), .B(n9619), .Z(n9624) );
  OR U12463 ( .A(n9622), .B(n9621), .Z(n9623) );
  NAND U12464 ( .A(n9624), .B(n9623), .Z(n11211) );
  XOR U12465 ( .A(n11210), .B(n11211), .Z(n11213) );
  XOR U12466 ( .A(n11212), .B(n11213), .Z(n11021) );
  XOR U12467 ( .A(n11020), .B(n11021), .Z(n11023) );
  XNOR U12468 ( .A(n11022), .B(n11023), .Z(n11180) );
  XNOR U12469 ( .A(n11181), .B(n11180), .Z(n11182) );
  NANDN U12470 ( .A(n9626), .B(n9625), .Z(n9630) );
  OR U12471 ( .A(n9628), .B(n9627), .Z(n9629) );
  AND U12472 ( .A(n9630), .B(n9629), .Z(n11017) );
  NANDN U12473 ( .A(n9632), .B(n9631), .Z(n9636) );
  NAND U12474 ( .A(n9634), .B(n9633), .Z(n9635) );
  AND U12475 ( .A(n9636), .B(n9635), .Z(n11015) );
  NANDN U12476 ( .A(n9638), .B(n9637), .Z(n9642) );
  NANDN U12477 ( .A(n9640), .B(n9639), .Z(n9641) );
  AND U12478 ( .A(n9642), .B(n9641), .Z(n11223) );
  NANDN U12479 ( .A(n9644), .B(n9643), .Z(n9648) );
  NANDN U12480 ( .A(n9646), .B(n9645), .Z(n9647) );
  NAND U12481 ( .A(n9648), .B(n9647), .Z(n11221) );
  NANDN U12482 ( .A(n9650), .B(n9649), .Z(n9654) );
  OR U12483 ( .A(n9652), .B(n9651), .Z(n9653) );
  AND U12484 ( .A(n9654), .B(n9653), .Z(n11222) );
  XOR U12485 ( .A(n11221), .B(n11222), .Z(n9655) );
  XNOR U12486 ( .A(n11223), .B(n9655), .Z(n11014) );
  XNOR U12487 ( .A(n11015), .B(n11014), .Z(n11016) );
  XOR U12488 ( .A(n11017), .B(n11016), .Z(n11183) );
  XNOR U12489 ( .A(n11182), .B(n11183), .Z(n11239) );
  XNOR U12490 ( .A(n11240), .B(n11239), .Z(n10919) );
  NAND U12491 ( .A(n9657), .B(n9656), .Z(n9661) );
  NANDN U12492 ( .A(n9659), .B(n9658), .Z(n9660) );
  AND U12493 ( .A(n9661), .B(n9660), .Z(n11035) );
  NANDN U12494 ( .A(n9663), .B(n9662), .Z(n9667) );
  OR U12495 ( .A(n9665), .B(n9664), .Z(n9666) );
  AND U12496 ( .A(n9667), .B(n9666), .Z(n11032) );
  NAND U12497 ( .A(n9669), .B(n9668), .Z(n9673) );
  NAND U12498 ( .A(n9671), .B(n9670), .Z(n9672) );
  NAND U12499 ( .A(n9673), .B(n9672), .Z(n11033) );
  XNOR U12500 ( .A(n11032), .B(n11033), .Z(n11034) );
  XOR U12501 ( .A(n11035), .B(n11034), .Z(n10787) );
  NANDN U12502 ( .A(n9675), .B(n9674), .Z(n9679) );
  NANDN U12503 ( .A(n9677), .B(n9676), .Z(n9678) );
  AND U12504 ( .A(n9679), .B(n9678), .Z(n10786) );
  XNOR U12505 ( .A(n10787), .B(n10786), .Z(n10789) );
  NANDN U12506 ( .A(n9681), .B(n9680), .Z(n9685) );
  NANDN U12507 ( .A(n9683), .B(n9682), .Z(n9684) );
  AND U12508 ( .A(n9685), .B(n9684), .Z(n10788) );
  XOR U12509 ( .A(n10789), .B(n10788), .Z(n10710) );
  NANDN U12510 ( .A(n9687), .B(n9686), .Z(n9691) );
  NANDN U12511 ( .A(n9689), .B(n9688), .Z(n9690) );
  AND U12512 ( .A(n9691), .B(n9690), .Z(n10702) );
  NANDN U12513 ( .A(n9693), .B(n9692), .Z(n9697) );
  NANDN U12514 ( .A(n9695), .B(n9694), .Z(n9696) );
  NAND U12515 ( .A(n9697), .B(n9696), .Z(n10703) );
  XNOR U12516 ( .A(n10702), .B(n10703), .Z(n10705) );
  NANDN U12517 ( .A(n9699), .B(n9698), .Z(n9703) );
  NANDN U12518 ( .A(n9701), .B(n9700), .Z(n9702) );
  AND U12519 ( .A(n9703), .B(n9702), .Z(n10704) );
  XOR U12520 ( .A(n10705), .B(n10704), .Z(n10709) );
  NANDN U12521 ( .A(n9705), .B(n9704), .Z(n9709) );
  NANDN U12522 ( .A(n9707), .B(n9706), .Z(n9708) );
  NAND U12523 ( .A(n9709), .B(n9708), .Z(n10708) );
  XOR U12524 ( .A(n10709), .B(n10708), .Z(n10711) );
  XNOR U12525 ( .A(n10710), .B(n10711), .Z(n10669) );
  NAND U12526 ( .A(n9711), .B(n9710), .Z(n9715) );
  NAND U12527 ( .A(n9713), .B(n9712), .Z(n9714) );
  AND U12528 ( .A(n9715), .B(n9714), .Z(n10666) );
  NANDN U12529 ( .A(n9717), .B(n9716), .Z(n9721) );
  NANDN U12530 ( .A(n9719), .B(n9718), .Z(n9720) );
  AND U12531 ( .A(n9721), .B(n9720), .Z(n10894) );
  NANDN U12532 ( .A(n9723), .B(n9722), .Z(n9727) );
  NANDN U12533 ( .A(n9725), .B(n9724), .Z(n9726) );
  NAND U12534 ( .A(n9727), .B(n9726), .Z(n10895) );
  XNOR U12535 ( .A(n10894), .B(n10895), .Z(n10896) );
  NANDN U12536 ( .A(n9729), .B(n9728), .Z(n9733) );
  NANDN U12537 ( .A(n9731), .B(n9730), .Z(n9732) );
  NAND U12538 ( .A(n9733), .B(n9732), .Z(n10897) );
  XNOR U12539 ( .A(n10896), .B(n10897), .Z(n10756) );
  NANDN U12540 ( .A(n9735), .B(n9734), .Z(n9739) );
  NANDN U12541 ( .A(n9737), .B(n9736), .Z(n9738) );
  NAND U12542 ( .A(n9739), .B(n9738), .Z(n10757) );
  XNOR U12543 ( .A(n10756), .B(n10757), .Z(n10758) );
  NAND U12544 ( .A(n9741), .B(n9740), .Z(n9745) );
  NANDN U12545 ( .A(n9743), .B(n9742), .Z(n9744) );
  AND U12546 ( .A(n9745), .B(n9744), .Z(n11144) );
  NANDN U12547 ( .A(n9747), .B(n9746), .Z(n9751) );
  NANDN U12548 ( .A(n9749), .B(n9748), .Z(n9750) );
  NAND U12549 ( .A(n9751), .B(n9750), .Z(n11145) );
  XNOR U12550 ( .A(n11144), .B(n11145), .Z(n11146) );
  NANDN U12551 ( .A(n9753), .B(n9752), .Z(n9757) );
  NANDN U12552 ( .A(n9755), .B(n9754), .Z(n9756) );
  NAND U12553 ( .A(n9757), .B(n9756), .Z(n11147) );
  XOR U12554 ( .A(n11146), .B(n11147), .Z(n10759) );
  XNOR U12555 ( .A(n10758), .B(n10759), .Z(n10667) );
  XOR U12556 ( .A(n10666), .B(n10667), .Z(n10668) );
  XOR U12557 ( .A(n10669), .B(n10668), .Z(n10918) );
  XOR U12558 ( .A(n10919), .B(n10918), .Z(n10920) );
  XOR U12559 ( .A(n10921), .B(n10920), .Z(n11267) );
  XOR U12560 ( .A(n11268), .B(n11267), .Z(n11269) );
  XOR U12561 ( .A(n11270), .B(n11269), .Z(n10628) );
  NAND U12562 ( .A(n9759), .B(n9758), .Z(n9763) );
  NAND U12563 ( .A(n9761), .B(n9760), .Z(n9762) );
  AND U12564 ( .A(n9763), .B(n9762), .Z(n10604) );
  NAND U12565 ( .A(n9765), .B(n9764), .Z(n9769) );
  NAND U12566 ( .A(n9767), .B(n9766), .Z(n9768) );
  AND U12567 ( .A(n9769), .B(n9768), .Z(n10783) );
  NAND U12568 ( .A(n9771), .B(n9770), .Z(n9775) );
  NAND U12569 ( .A(n9773), .B(n9772), .Z(n9774) );
  NAND U12570 ( .A(n9775), .B(n9774), .Z(n10781) );
  NAND U12571 ( .A(n9777), .B(n9776), .Z(n9781) );
  NAND U12572 ( .A(n9779), .B(n9778), .Z(n9780) );
  AND U12573 ( .A(n9781), .B(n9780), .Z(n10780) );
  XOR U12574 ( .A(n10781), .B(n10780), .Z(n10782) );
  XOR U12575 ( .A(n10783), .B(n10782), .Z(n10603) );
  XOR U12576 ( .A(n10604), .B(n10603), .Z(n10606) );
  NANDN U12577 ( .A(n9783), .B(n9782), .Z(n9787) );
  NAND U12578 ( .A(n9785), .B(n9784), .Z(n9786) );
  AND U12579 ( .A(n9787), .B(n9786), .Z(n11258) );
  NANDN U12580 ( .A(n9789), .B(n9788), .Z(n9793) );
  NAND U12581 ( .A(n9791), .B(n9790), .Z(n9792) );
  AND U12582 ( .A(n9793), .B(n9792), .Z(n11256) );
  NANDN U12583 ( .A(n9795), .B(n9794), .Z(n9799) );
  NANDN U12584 ( .A(n9797), .B(n9796), .Z(n9798) );
  AND U12585 ( .A(n9799), .B(n9798), .Z(n11255) );
  XNOR U12586 ( .A(n11256), .B(n11255), .Z(n11257) );
  XNOR U12587 ( .A(n11258), .B(n11257), .Z(n10605) );
  XNOR U12588 ( .A(n10606), .B(n10605), .Z(n10909) );
  NAND U12589 ( .A(n9801), .B(n9800), .Z(n9805) );
  NAND U12590 ( .A(n9803), .B(n9802), .Z(n9804) );
  NAND U12591 ( .A(n9805), .B(n9804), .Z(n11228) );
  NAND U12592 ( .A(n9807), .B(n9806), .Z(n9811) );
  NAND U12593 ( .A(n9809), .B(n9808), .Z(n9810) );
  NAND U12594 ( .A(n9811), .B(n9810), .Z(n11111) );
  NAND U12595 ( .A(n9813), .B(n9812), .Z(n9817) );
  NAND U12596 ( .A(n9815), .B(n9814), .Z(n9816) );
  NAND U12597 ( .A(n9817), .B(n9816), .Z(n11109) );
  NAND U12598 ( .A(n9819), .B(n9818), .Z(n9823) );
  NAND U12599 ( .A(n9821), .B(n9820), .Z(n9822) );
  AND U12600 ( .A(n9823), .B(n9822), .Z(n11110) );
  XOR U12601 ( .A(n11109), .B(n11110), .Z(n11112) );
  XOR U12602 ( .A(n11111), .B(n11112), .Z(n11225) );
  NAND U12603 ( .A(n9825), .B(n9824), .Z(n9829) );
  NAND U12604 ( .A(n9827), .B(n9826), .Z(n9828) );
  NAND U12605 ( .A(n9829), .B(n9828), .Z(n11050) );
  NANDN U12606 ( .A(n9831), .B(n9830), .Z(n9835) );
  NANDN U12607 ( .A(n9833), .B(n9832), .Z(n9834) );
  NAND U12608 ( .A(n9835), .B(n9834), .Z(n11049) );
  NANDN U12609 ( .A(n9837), .B(n9836), .Z(n9841) );
  NANDN U12610 ( .A(n9839), .B(n9838), .Z(n9840) );
  AND U12611 ( .A(n9841), .B(n9840), .Z(n11048) );
  XOR U12612 ( .A(n11049), .B(n11048), .Z(n9842) );
  XOR U12613 ( .A(n11050), .B(n9842), .Z(n10747) );
  NANDN U12614 ( .A(n9844), .B(n9843), .Z(n9848) );
  NANDN U12615 ( .A(n9846), .B(n9845), .Z(n9847) );
  AND U12616 ( .A(n9848), .B(n9847), .Z(n10745) );
  NAND U12617 ( .A(n9850), .B(n9849), .Z(n9854) );
  NANDN U12618 ( .A(n9852), .B(n9851), .Z(n9853) );
  AND U12619 ( .A(n9854), .B(n9853), .Z(n11118) );
  NANDN U12620 ( .A(n9856), .B(n9855), .Z(n9860) );
  NANDN U12621 ( .A(n9858), .B(n9857), .Z(n9859) );
  AND U12622 ( .A(n9860), .B(n9859), .Z(n11116) );
  NANDN U12623 ( .A(n9862), .B(n9861), .Z(n9866) );
  NAND U12624 ( .A(n9864), .B(n9863), .Z(n9865) );
  NAND U12625 ( .A(n9866), .B(n9865), .Z(n11115) );
  XNOR U12626 ( .A(n11116), .B(n11115), .Z(n11117) );
  XNOR U12627 ( .A(n11118), .B(n11117), .Z(n10744) );
  XNOR U12628 ( .A(n10745), .B(n10744), .Z(n10746) );
  XNOR U12629 ( .A(n10747), .B(n10746), .Z(n11251) );
  NANDN U12630 ( .A(n9868), .B(n9867), .Z(n9872) );
  NAND U12631 ( .A(n9870), .B(n9869), .Z(n9871) );
  AND U12632 ( .A(n9872), .B(n9871), .Z(n11250) );
  NAND U12633 ( .A(n9874), .B(n9873), .Z(n9878) );
  NAND U12634 ( .A(n9876), .B(n9875), .Z(n9877) );
  AND U12635 ( .A(n9878), .B(n9877), .Z(n11011) );
  NAND U12636 ( .A(n9880), .B(n9879), .Z(n9884) );
  NANDN U12637 ( .A(n9882), .B(n9881), .Z(n9883) );
  AND U12638 ( .A(n9884), .B(n9883), .Z(n11008) );
  NAND U12639 ( .A(n9886), .B(n9885), .Z(n9890) );
  NAND U12640 ( .A(n9888), .B(n9887), .Z(n9889) );
  NAND U12641 ( .A(n9890), .B(n9889), .Z(n11009) );
  XNOR U12642 ( .A(n11008), .B(n11009), .Z(n11010) );
  XOR U12643 ( .A(n11011), .B(n11010), .Z(n10950) );
  NAND U12644 ( .A(n9892), .B(n9891), .Z(n9896) );
  NANDN U12645 ( .A(n9894), .B(n9893), .Z(n9895) );
  AND U12646 ( .A(n9896), .B(n9895), .Z(n10984) );
  NANDN U12647 ( .A(n9898), .B(n9897), .Z(n9902) );
  OR U12648 ( .A(n9900), .B(n9899), .Z(n9901) );
  NAND U12649 ( .A(n9902), .B(n9901), .Z(n10985) );
  XNOR U12650 ( .A(n10984), .B(n10985), .Z(n10987) );
  NANDN U12651 ( .A(n9904), .B(n9903), .Z(n9908) );
  OR U12652 ( .A(n9906), .B(n9905), .Z(n9907) );
  AND U12653 ( .A(n9908), .B(n9907), .Z(n10986) );
  XOR U12654 ( .A(n10987), .B(n10986), .Z(n10949) );
  NANDN U12655 ( .A(n9910), .B(n9909), .Z(n9914) );
  NANDN U12656 ( .A(n9912), .B(n9911), .Z(n9913) );
  AND U12657 ( .A(n9914), .B(n9913), .Z(n10948) );
  XOR U12658 ( .A(n10949), .B(n10948), .Z(n10951) );
  XOR U12659 ( .A(n10950), .B(n10951), .Z(n10963) );
  NANDN U12660 ( .A(n9916), .B(n9915), .Z(n9920) );
  NAND U12661 ( .A(n9918), .B(n9917), .Z(n9919) );
  AND U12662 ( .A(n9920), .B(n9919), .Z(n10961) );
  NAND U12663 ( .A(n9922), .B(n9921), .Z(n9926) );
  NANDN U12664 ( .A(n9924), .B(n9923), .Z(n9925) );
  AND U12665 ( .A(n9926), .B(n9925), .Z(n11045) );
  NANDN U12666 ( .A(n9928), .B(n9927), .Z(n9932) );
  OR U12667 ( .A(n9930), .B(n9929), .Z(n9931) );
  AND U12668 ( .A(n9932), .B(n9931), .Z(n10975) );
  NANDN U12669 ( .A(n9934), .B(n9933), .Z(n9938) );
  OR U12670 ( .A(n9936), .B(n9935), .Z(n9937) );
  AND U12671 ( .A(n9938), .B(n9937), .Z(n10973) );
  NANDN U12672 ( .A(n9940), .B(n9939), .Z(n9944) );
  OR U12673 ( .A(n9942), .B(n9941), .Z(n9943) );
  AND U12674 ( .A(n9944), .B(n9943), .Z(n10972) );
  XOR U12675 ( .A(n10973), .B(n10972), .Z(n10974) );
  XOR U12676 ( .A(n10975), .B(n10974), .Z(n11044) );
  XNOR U12677 ( .A(n11045), .B(n11044), .Z(n11047) );
  NAND U12678 ( .A(n9946), .B(n9945), .Z(n9950) );
  NANDN U12679 ( .A(n9948), .B(n9947), .Z(n9949) );
  AND U12680 ( .A(n9950), .B(n9949), .Z(n11005) );
  NANDN U12681 ( .A(n9952), .B(n9951), .Z(n9956) );
  OR U12682 ( .A(n9954), .B(n9953), .Z(n9955) );
  AND U12683 ( .A(n9956), .B(n9955), .Z(n11003) );
  NANDN U12684 ( .A(n9958), .B(n9957), .Z(n9962) );
  OR U12685 ( .A(n9960), .B(n9959), .Z(n9961) );
  AND U12686 ( .A(n9962), .B(n9961), .Z(n11002) );
  XOR U12687 ( .A(n11003), .B(n11002), .Z(n11004) );
  XOR U12688 ( .A(n11005), .B(n11004), .Z(n11046) );
  XOR U12689 ( .A(n11047), .B(n11046), .Z(n10960) );
  XNOR U12690 ( .A(n10961), .B(n10960), .Z(n10962) );
  XNOR U12691 ( .A(n10963), .B(n10962), .Z(n11249) );
  XOR U12692 ( .A(n11250), .B(n11249), .Z(n11252) );
  XNOR U12693 ( .A(n11251), .B(n11252), .Z(n11226) );
  XOR U12694 ( .A(n11225), .B(n11226), .Z(n11227) );
  XNOR U12695 ( .A(n11228), .B(n11227), .Z(n10906) );
  NAND U12696 ( .A(n9964), .B(n9963), .Z(n9968) );
  NAND U12697 ( .A(n9966), .B(n9965), .Z(n9967) );
  NAND U12698 ( .A(n9968), .B(n9967), .Z(n10597) );
  NANDN U12699 ( .A(n9970), .B(n9969), .Z(n9974) );
  NAND U12700 ( .A(n9972), .B(n9971), .Z(n9973) );
  AND U12701 ( .A(n9974), .B(n9973), .Z(n10685) );
  NANDN U12702 ( .A(n9976), .B(n9975), .Z(n9980) );
  NANDN U12703 ( .A(n9978), .B(n9977), .Z(n9979) );
  AND U12704 ( .A(n9980), .B(n9979), .Z(n10817) );
  NANDN U12705 ( .A(n9982), .B(n9981), .Z(n9986) );
  OR U12706 ( .A(n9984), .B(n9983), .Z(n9985) );
  AND U12707 ( .A(n9986), .B(n9985), .Z(n11063) );
  NANDN U12708 ( .A(n9988), .B(n9987), .Z(n9992) );
  OR U12709 ( .A(n9990), .B(n9989), .Z(n9991) );
  AND U12710 ( .A(n9992), .B(n9991), .Z(n11061) );
  NAND U12711 ( .A(n9994), .B(n9993), .Z(n9998) );
  NANDN U12712 ( .A(n9996), .B(n9995), .Z(n9997) );
  NAND U12713 ( .A(n9998), .B(n9997), .Z(n11062) );
  XOR U12714 ( .A(n11061), .B(n11062), .Z(n11064) );
  XNOR U12715 ( .A(n11063), .B(n11064), .Z(n10816) );
  XNOR U12716 ( .A(n10817), .B(n10816), .Z(n10818) );
  NANDN U12717 ( .A(n10000), .B(n9999), .Z(n10004) );
  OR U12718 ( .A(n10002), .B(n10001), .Z(n10003) );
  AND U12719 ( .A(n10004), .B(n10003), .Z(n11069) );
  NANDN U12720 ( .A(n10006), .B(n10005), .Z(n10010) );
  OR U12721 ( .A(n10008), .B(n10007), .Z(n10009) );
  AND U12722 ( .A(n10010), .B(n10009), .Z(n11067) );
  NANDN U12723 ( .A(n10012), .B(n10011), .Z(n10016) );
  OR U12724 ( .A(n10014), .B(n10013), .Z(n10015) );
  NAND U12725 ( .A(n10016), .B(n10015), .Z(n11068) );
  XOR U12726 ( .A(n11067), .B(n11068), .Z(n11070) );
  XOR U12727 ( .A(n11069), .B(n11070), .Z(n10819) );
  XNOR U12728 ( .A(n10818), .B(n10819), .Z(n10684) );
  XNOR U12729 ( .A(n10685), .B(n10684), .Z(n10686) );
  NANDN U12730 ( .A(n10018), .B(n10017), .Z(n10022) );
  NANDN U12731 ( .A(n10020), .B(n10019), .Z(n10021) );
  AND U12732 ( .A(n10022), .B(n10021), .Z(n10813) );
  NANDN U12733 ( .A(n10024), .B(n10023), .Z(n10028) );
  OR U12734 ( .A(n10026), .B(n10025), .Z(n10027) );
  AND U12735 ( .A(n10028), .B(n10027), .Z(n10811) );
  NANDN U12736 ( .A(n10030), .B(n10029), .Z(n10034) );
  NANDN U12737 ( .A(n10032), .B(n10031), .Z(n10033) );
  NAND U12738 ( .A(n10034), .B(n10033), .Z(n10810) );
  XNOR U12739 ( .A(n10811), .B(n10810), .Z(n10812) );
  XOR U12740 ( .A(n10813), .B(n10812), .Z(n10687) );
  XNOR U12741 ( .A(n10686), .B(n10687), .Z(n10598) );
  XOR U12742 ( .A(n10597), .B(n10598), .Z(n10600) );
  NAND U12743 ( .A(n10036), .B(n10035), .Z(n10040) );
  NANDN U12744 ( .A(n10038), .B(n10037), .Z(n10039) );
  AND U12745 ( .A(n10040), .B(n10039), .Z(n11076) );
  NANDN U12746 ( .A(n10042), .B(n10041), .Z(n10046) );
  OR U12747 ( .A(n10044), .B(n10043), .Z(n10045) );
  AND U12748 ( .A(n10046), .B(n10045), .Z(n11073) );
  NAND U12749 ( .A(n10048), .B(n10047), .Z(n10052) );
  NANDN U12750 ( .A(n10050), .B(n10049), .Z(n10051) );
  NAND U12751 ( .A(n10052), .B(n10051), .Z(n11074) );
  XNOR U12752 ( .A(n11073), .B(n11074), .Z(n11075) );
  XOR U12753 ( .A(n11076), .B(n11075), .Z(n10697) );
  NANDN U12754 ( .A(n10054), .B(n10053), .Z(n10058) );
  NANDN U12755 ( .A(n10056), .B(n10055), .Z(n10057) );
  AND U12756 ( .A(n10058), .B(n10057), .Z(n10696) );
  XNOR U12757 ( .A(n10697), .B(n10696), .Z(n10699) );
  NANDN U12758 ( .A(n10060), .B(n10059), .Z(n10064) );
  NANDN U12759 ( .A(n10062), .B(n10061), .Z(n10063) );
  AND U12760 ( .A(n10064), .B(n10063), .Z(n10698) );
  XOR U12761 ( .A(n10699), .B(n10698), .Z(n10867) );
  NANDN U12762 ( .A(n10066), .B(n10065), .Z(n10070) );
  NAND U12763 ( .A(n10068), .B(n10067), .Z(n10069) );
  AND U12764 ( .A(n10070), .B(n10069), .Z(n10865) );
  NANDN U12765 ( .A(n10072), .B(n10071), .Z(n10076) );
  NANDN U12766 ( .A(n10074), .B(n10073), .Z(n10075) );
  AND U12767 ( .A(n10076), .B(n10075), .Z(n11141) );
  NANDN U12768 ( .A(n10078), .B(n10077), .Z(n10082) );
  OR U12769 ( .A(n10080), .B(n10079), .Z(n10081) );
  AND U12770 ( .A(n10082), .B(n10081), .Z(n11165) );
  NANDN U12771 ( .A(n10084), .B(n10083), .Z(n10088) );
  OR U12772 ( .A(n10086), .B(n10085), .Z(n10087) );
  AND U12773 ( .A(n10088), .B(n10087), .Z(n11163) );
  NANDN U12774 ( .A(n10090), .B(n10089), .Z(n10094) );
  OR U12775 ( .A(n10092), .B(n10091), .Z(n10093) );
  AND U12776 ( .A(n10094), .B(n10093), .Z(n11162) );
  XOR U12777 ( .A(n11163), .B(n11162), .Z(n11164) );
  XOR U12778 ( .A(n11165), .B(n11164), .Z(n11140) );
  XNOR U12779 ( .A(n11141), .B(n11140), .Z(n11143) );
  NAND U12780 ( .A(n10096), .B(n10095), .Z(n10100) );
  NAND U12781 ( .A(n10098), .B(n10097), .Z(n10099) );
  AND U12782 ( .A(n10100), .B(n10099), .Z(n11041) );
  NANDN U12783 ( .A(n10102), .B(n10101), .Z(n10106) );
  OR U12784 ( .A(n10104), .B(n10103), .Z(n10105) );
  AND U12785 ( .A(n10106), .B(n10105), .Z(n11039) );
  NAND U12786 ( .A(n10108), .B(n10107), .Z(n10112) );
  NAND U12787 ( .A(n10110), .B(n10109), .Z(n10111) );
  AND U12788 ( .A(n10112), .B(n10111), .Z(n11038) );
  XOR U12789 ( .A(n11039), .B(n11038), .Z(n11040) );
  XOR U12790 ( .A(n11041), .B(n11040), .Z(n11142) );
  XOR U12791 ( .A(n11143), .B(n11142), .Z(n10864) );
  XNOR U12792 ( .A(n10865), .B(n10864), .Z(n10866) );
  XNOR U12793 ( .A(n10867), .B(n10866), .Z(n10599) );
  XNOR U12794 ( .A(n10600), .B(n10599), .Z(n10915) );
  NAND U12795 ( .A(n10114), .B(n10113), .Z(n10118) );
  NAND U12796 ( .A(n10116), .B(n10115), .Z(n10117) );
  NAND U12797 ( .A(n10118), .B(n10117), .Z(n10913) );
  NAND U12798 ( .A(n10120), .B(n10119), .Z(n10124) );
  NANDN U12799 ( .A(n10122), .B(n10121), .Z(n10123) );
  AND U12800 ( .A(n10124), .B(n10123), .Z(n11094) );
  NAND U12801 ( .A(n10126), .B(n10125), .Z(n10130) );
  NAND U12802 ( .A(n10128), .B(n10127), .Z(n10129) );
  AND U12803 ( .A(n10130), .B(n10129), .Z(n11091) );
  NAND U12804 ( .A(n10132), .B(n10131), .Z(n10136) );
  NANDN U12805 ( .A(n10134), .B(n10133), .Z(n10135) );
  NAND U12806 ( .A(n10136), .B(n10135), .Z(n11092) );
  XNOR U12807 ( .A(n11091), .B(n11092), .Z(n11093) );
  XOR U12808 ( .A(n11094), .B(n11093), .Z(n10805) );
  NANDN U12809 ( .A(n10138), .B(n10137), .Z(n10142) );
  NANDN U12810 ( .A(n10140), .B(n10139), .Z(n10141) );
  AND U12811 ( .A(n10142), .B(n10141), .Z(n10804) );
  XNOR U12812 ( .A(n10805), .B(n10804), .Z(n10807) );
  NANDN U12813 ( .A(n10144), .B(n10143), .Z(n10148) );
  NANDN U12814 ( .A(n10146), .B(n10145), .Z(n10147) );
  AND U12815 ( .A(n10148), .B(n10147), .Z(n10806) );
  XOR U12816 ( .A(n10807), .B(n10806), .Z(n10860) );
  NANDN U12817 ( .A(n10150), .B(n10149), .Z(n10154) );
  NANDN U12818 ( .A(n10152), .B(n10151), .Z(n10153) );
  AND U12819 ( .A(n10154), .B(n10153), .Z(n10859) );
  NANDN U12820 ( .A(n10156), .B(n10155), .Z(n10160) );
  NANDN U12821 ( .A(n10158), .B(n10157), .Z(n10159) );
  AND U12822 ( .A(n10160), .B(n10159), .Z(n10691) );
  NANDN U12823 ( .A(n10162), .B(n10161), .Z(n10166) );
  NANDN U12824 ( .A(n10164), .B(n10163), .Z(n10165) );
  NAND U12825 ( .A(n10166), .B(n10165), .Z(n10690) );
  XNOR U12826 ( .A(n10691), .B(n10690), .Z(n10692) );
  NAND U12827 ( .A(n10168), .B(n10167), .Z(n10172) );
  NAND U12828 ( .A(n10170), .B(n10169), .Z(n10171) );
  AND U12829 ( .A(n10172), .B(n10171), .Z(n10992) );
  NAND U12830 ( .A(n10174), .B(n10173), .Z(n10178) );
  NANDN U12831 ( .A(n10176), .B(n10175), .Z(n10177) );
  AND U12832 ( .A(n10178), .B(n10177), .Z(n10990) );
  NAND U12833 ( .A(n10180), .B(n10179), .Z(n10184) );
  NANDN U12834 ( .A(n10182), .B(n10181), .Z(n10183) );
  NAND U12835 ( .A(n10184), .B(n10183), .Z(n10991) );
  XOR U12836 ( .A(n10990), .B(n10991), .Z(n10993) );
  XOR U12837 ( .A(n10992), .B(n10993), .Z(n10693) );
  XNOR U12838 ( .A(n10692), .B(n10693), .Z(n10858) );
  XOR U12839 ( .A(n10859), .B(n10858), .Z(n10861) );
  XNOR U12840 ( .A(n10860), .B(n10861), .Z(n10639) );
  NANDN U12841 ( .A(n10186), .B(n10185), .Z(n10190) );
  NANDN U12842 ( .A(n10188), .B(n10187), .Z(n10189) );
  AND U12843 ( .A(n10190), .B(n10189), .Z(n11082) );
  NAND U12844 ( .A(n10192), .B(n10191), .Z(n10196) );
  NAND U12845 ( .A(n10194), .B(n10193), .Z(n10195) );
  AND U12846 ( .A(n10196), .B(n10195), .Z(n11079) );
  NANDN U12847 ( .A(n10198), .B(n10197), .Z(n10202) );
  OR U12848 ( .A(n10200), .B(n10199), .Z(n10201) );
  NAND U12849 ( .A(n10202), .B(n10201), .Z(n11080) );
  XNOR U12850 ( .A(n11079), .B(n11080), .Z(n11081) );
  XOR U12851 ( .A(n11082), .B(n11081), .Z(n10925) );
  NANDN U12852 ( .A(n10204), .B(n10203), .Z(n10208) );
  NANDN U12853 ( .A(n10206), .B(n10205), .Z(n10207) );
  AND U12854 ( .A(n10208), .B(n10207), .Z(n10924) );
  XNOR U12855 ( .A(n10925), .B(n10924), .Z(n10927) );
  NANDN U12856 ( .A(n10210), .B(n10209), .Z(n10214) );
  NANDN U12857 ( .A(n10212), .B(n10211), .Z(n10213) );
  AND U12858 ( .A(n10214), .B(n10213), .Z(n10926) );
  XOR U12859 ( .A(n10927), .B(n10926), .Z(n10878) );
  NANDN U12860 ( .A(n10216), .B(n10215), .Z(n10220) );
  OR U12861 ( .A(n10218), .B(n10217), .Z(n10219) );
  AND U12862 ( .A(n10220), .B(n10219), .Z(n10877) );
  NANDN U12863 ( .A(n10222), .B(n10221), .Z(n10226) );
  OR U12864 ( .A(n10224), .B(n10223), .Z(n10225) );
  NAND U12865 ( .A(n10226), .B(n10225), .Z(n11028) );
  NANDN U12866 ( .A(n10228), .B(n10227), .Z(n10232) );
  OR U12867 ( .A(n10230), .B(n10229), .Z(n10231) );
  NAND U12868 ( .A(n10232), .B(n10231), .Z(n11027) );
  NAND U12869 ( .A(n10234), .B(n10233), .Z(n10238) );
  NANDN U12870 ( .A(n10236), .B(n10235), .Z(n10237) );
  NAND U12871 ( .A(n10238), .B(n10237), .Z(n11026) );
  XOR U12872 ( .A(n11027), .B(n11026), .Z(n11029) );
  XOR U12873 ( .A(n11028), .B(n11029), .Z(n11123) );
  NANDN U12874 ( .A(n10240), .B(n10239), .Z(n10244) );
  NANDN U12875 ( .A(n10242), .B(n10241), .Z(n10243) );
  NAND U12876 ( .A(n10244), .B(n10243), .Z(n11121) );
  NANDN U12877 ( .A(n10246), .B(n10245), .Z(n10250) );
  NAND U12878 ( .A(n10248), .B(n10247), .Z(n10249) );
  AND U12879 ( .A(n10250), .B(n10249), .Z(n11122) );
  XOR U12880 ( .A(n11121), .B(n11122), .Z(n10251) );
  XNOR U12881 ( .A(n11123), .B(n10251), .Z(n10876) );
  XOR U12882 ( .A(n10877), .B(n10876), .Z(n10879) );
  XNOR U12883 ( .A(n10878), .B(n10879), .Z(n10637) );
  NAND U12884 ( .A(n10253), .B(n10252), .Z(n10257) );
  NANDN U12885 ( .A(n10255), .B(n10254), .Z(n10256) );
  AND U12886 ( .A(n10257), .B(n10256), .Z(n11168) );
  NANDN U12887 ( .A(n10259), .B(n10258), .Z(n10263) );
  OR U12888 ( .A(n10261), .B(n10260), .Z(n10262) );
  NAND U12889 ( .A(n10263), .B(n10262), .Z(n11169) );
  XNOR U12890 ( .A(n11168), .B(n11169), .Z(n11171) );
  NANDN U12891 ( .A(n10265), .B(n10264), .Z(n10269) );
  OR U12892 ( .A(n10267), .B(n10266), .Z(n10268) );
  AND U12893 ( .A(n10269), .B(n10268), .Z(n11170) );
  XOR U12894 ( .A(n11171), .B(n11170), .Z(n10945) );
  NAND U12895 ( .A(n10271), .B(n10270), .Z(n10275) );
  NAND U12896 ( .A(n10273), .B(n10272), .Z(n10274) );
  AND U12897 ( .A(n10275), .B(n10274), .Z(n10999) );
  NAND U12898 ( .A(n10277), .B(n10276), .Z(n10281) );
  NANDN U12899 ( .A(n10279), .B(n10278), .Z(n10280) );
  AND U12900 ( .A(n10281), .B(n10280), .Z(n10996) );
  NANDN U12901 ( .A(n10283), .B(n10282), .Z(n10287) );
  OR U12902 ( .A(n10285), .B(n10284), .Z(n10286) );
  NAND U12903 ( .A(n10287), .B(n10286), .Z(n10997) );
  XNOR U12904 ( .A(n10996), .B(n10997), .Z(n10998) );
  XOR U12905 ( .A(n10999), .B(n10998), .Z(n10943) );
  NANDN U12906 ( .A(n10289), .B(n10288), .Z(n10293) );
  NANDN U12907 ( .A(n10291), .B(n10290), .Z(n10292) );
  AND U12908 ( .A(n10293), .B(n10292), .Z(n10942) );
  XNOR U12909 ( .A(n10943), .B(n10942), .Z(n10944) );
  XNOR U12910 ( .A(n10945), .B(n10944), .Z(n11130) );
  NANDN U12911 ( .A(n10295), .B(n10294), .Z(n10299) );
  NAND U12912 ( .A(n10297), .B(n10296), .Z(n10298) );
  NAND U12913 ( .A(n10299), .B(n10298), .Z(n11053) );
  NANDN U12914 ( .A(n10301), .B(n10300), .Z(n10305) );
  OR U12915 ( .A(n10303), .B(n10302), .Z(n10304) );
  AND U12916 ( .A(n10305), .B(n10304), .Z(n10979) );
  NAND U12917 ( .A(n10307), .B(n10306), .Z(n10311) );
  NAND U12918 ( .A(n10309), .B(n10308), .Z(n10310) );
  AND U12919 ( .A(n10311), .B(n10310), .Z(n10978) );
  XOR U12920 ( .A(n10979), .B(n10978), .Z(n10981) );
  NANDN U12921 ( .A(n10313), .B(n10312), .Z(n10317) );
  OR U12922 ( .A(n10315), .B(n10314), .Z(n10316) );
  AND U12923 ( .A(n10317), .B(n10316), .Z(n10980) );
  XOR U12924 ( .A(n10981), .B(n10980), .Z(n11052) );
  NANDN U12925 ( .A(n10319), .B(n10318), .Z(n10323) );
  NANDN U12926 ( .A(n10321), .B(n10320), .Z(n10322) );
  AND U12927 ( .A(n10323), .B(n10322), .Z(n11051) );
  XNOR U12928 ( .A(n11052), .B(n11051), .Z(n10324) );
  XNOR U12929 ( .A(n11053), .B(n10324), .Z(n11128) );
  NANDN U12930 ( .A(n10326), .B(n10325), .Z(n10330) );
  NANDN U12931 ( .A(n10328), .B(n10327), .Z(n10329) );
  NAND U12932 ( .A(n10330), .B(n10329), .Z(n11129) );
  XOR U12933 ( .A(n11128), .B(n11129), .Z(n11131) );
  XNOR U12934 ( .A(n11130), .B(n11131), .Z(n10636) );
  XOR U12935 ( .A(n10637), .B(n10636), .Z(n10638) );
  XOR U12936 ( .A(n10639), .B(n10638), .Z(n10912) );
  XOR U12937 ( .A(n10913), .B(n10912), .Z(n10914) );
  XOR U12938 ( .A(n10915), .B(n10914), .Z(n10907) );
  XOR U12939 ( .A(n10906), .B(n10907), .Z(n10908) );
  XOR U12940 ( .A(n10909), .B(n10908), .Z(n10627) );
  XOR U12941 ( .A(n10628), .B(n10627), .Z(n10630) );
  XOR U12942 ( .A(n10629), .B(n10630), .Z(n10557) );
  XOR U12943 ( .A(n10558), .B(n10557), .Z(n10633) );
  NAND U12944 ( .A(n10335), .B(n10334), .Z(n10339) );
  NAND U12945 ( .A(n10337), .B(n10336), .Z(n10338) );
  NAND U12946 ( .A(n10339), .B(n10338), .Z(n11282) );
  NAND U12947 ( .A(n10341), .B(n10340), .Z(n10345) );
  NAND U12948 ( .A(n10343), .B(n10342), .Z(n10344) );
  AND U12949 ( .A(n10345), .B(n10344), .Z(n10765) );
  NANDN U12950 ( .A(n10347), .B(n10346), .Z(n10351) );
  NAND U12951 ( .A(n10349), .B(n10348), .Z(n10350) );
  AND U12952 ( .A(n10351), .B(n10350), .Z(n10843) );
  NANDN U12953 ( .A(n10353), .B(n10352), .Z(n10357) );
  NANDN U12954 ( .A(n10355), .B(n10354), .Z(n10356) );
  AND U12955 ( .A(n10357), .B(n10356), .Z(n10841) );
  NANDN U12956 ( .A(n10359), .B(n10358), .Z(n10363) );
  NANDN U12957 ( .A(n10361), .B(n10360), .Z(n10362) );
  AND U12958 ( .A(n10363), .B(n10362), .Z(n10930) );
  NANDN U12959 ( .A(n10365), .B(n10364), .Z(n10369) );
  NANDN U12960 ( .A(n10367), .B(n10366), .Z(n10368) );
  NAND U12961 ( .A(n10369), .B(n10368), .Z(n10931) );
  XNOR U12962 ( .A(n10930), .B(n10931), .Z(n10933) );
  NANDN U12963 ( .A(n10371), .B(n10370), .Z(n10375) );
  NANDN U12964 ( .A(n10373), .B(n10372), .Z(n10374) );
  AND U12965 ( .A(n10375), .B(n10374), .Z(n10932) );
  XNOR U12966 ( .A(n10933), .B(n10932), .Z(n10840) );
  XNOR U12967 ( .A(n10841), .B(n10840), .Z(n10842) );
  XOR U12968 ( .A(n10843), .B(n10842), .Z(n10763) );
  NAND U12969 ( .A(n10377), .B(n10376), .Z(n10381) );
  NAND U12970 ( .A(n10379), .B(n10378), .Z(n10380) );
  NAND U12971 ( .A(n10381), .B(n10380), .Z(n10762) );
  XOR U12972 ( .A(n10763), .B(n10762), .Z(n10764) );
  XNOR U12973 ( .A(n10765), .B(n10764), .Z(n10618) );
  NAND U12974 ( .A(n10383), .B(n10382), .Z(n10387) );
  NAND U12975 ( .A(n10385), .B(n10384), .Z(n10386) );
  NAND U12976 ( .A(n10387), .B(n10386), .Z(n10663) );
  NAND U12977 ( .A(n10389), .B(n10388), .Z(n10393) );
  NAND U12978 ( .A(n10391), .B(n10390), .Z(n10392) );
  NAND U12979 ( .A(n10393), .B(n10392), .Z(n10661) );
  NANDN U12980 ( .A(n10395), .B(n10394), .Z(n10399) );
  OR U12981 ( .A(n10397), .B(n10396), .Z(n10398) );
  AND U12982 ( .A(n10399), .B(n10398), .Z(n11097) );
  NANDN U12983 ( .A(n10401), .B(n10400), .Z(n10405) );
  NANDN U12984 ( .A(n10403), .B(n10402), .Z(n10404) );
  NAND U12985 ( .A(n10405), .B(n10404), .Z(n11098) );
  XNOR U12986 ( .A(n11097), .B(n11098), .Z(n11100) );
  NANDN U12987 ( .A(n10407), .B(n10406), .Z(n10411) );
  NANDN U12988 ( .A(n10409), .B(n10408), .Z(n10410) );
  AND U12989 ( .A(n10411), .B(n10410), .Z(n11099) );
  XOR U12990 ( .A(n11100), .B(n11099), .Z(n10849) );
  NANDN U12991 ( .A(n10413), .B(n10412), .Z(n10417) );
  NANDN U12992 ( .A(n10415), .B(n10414), .Z(n10416) );
  AND U12993 ( .A(n10417), .B(n10416), .Z(n10847) );
  NANDN U12994 ( .A(n10419), .B(n10418), .Z(n10423) );
  NANDN U12995 ( .A(n10421), .B(n10420), .Z(n10422) );
  AND U12996 ( .A(n10423), .B(n10422), .Z(n11174) );
  NAND U12997 ( .A(n10425), .B(n10424), .Z(n10429) );
  NAND U12998 ( .A(n10427), .B(n10426), .Z(n10428) );
  NAND U12999 ( .A(n10429), .B(n10428), .Z(n11175) );
  XNOR U13000 ( .A(n11174), .B(n11175), .Z(n11177) );
  NANDN U13001 ( .A(n10431), .B(n10430), .Z(n10435) );
  NANDN U13002 ( .A(n10433), .B(n10432), .Z(n10434) );
  AND U13003 ( .A(n10435), .B(n10434), .Z(n11176) );
  XNOR U13004 ( .A(n11177), .B(n11176), .Z(n10846) );
  XNOR U13005 ( .A(n10847), .B(n10846), .Z(n10848) );
  XNOR U13006 ( .A(n10849), .B(n10848), .Z(n10660) );
  XOR U13007 ( .A(n10661), .B(n10660), .Z(n10662) );
  XOR U13008 ( .A(n10663), .B(n10662), .Z(n10615) );
  NAND U13009 ( .A(n10437), .B(n10436), .Z(n10441) );
  NAND U13010 ( .A(n10439), .B(n10438), .Z(n10440) );
  AND U13011 ( .A(n10441), .B(n10440), .Z(n10616) );
  XOR U13012 ( .A(n10615), .B(n10616), .Z(n10617) );
  XNOR U13013 ( .A(n10618), .B(n10617), .Z(n11275) );
  NAND U13014 ( .A(n10443), .B(n10442), .Z(n10447) );
  NAND U13015 ( .A(n10445), .B(n10444), .Z(n10446) );
  NAND U13016 ( .A(n10447), .B(n10446), .Z(n11274) );
  NAND U13017 ( .A(n10449), .B(n10448), .Z(n10453) );
  NAND U13018 ( .A(n10451), .B(n10450), .Z(n10452) );
  NAND U13019 ( .A(n10453), .B(n10452), .Z(n10740) );
  NAND U13020 ( .A(n10455), .B(n10454), .Z(n10459) );
  NAND U13021 ( .A(n10457), .B(n10456), .Z(n10458) );
  NAND U13022 ( .A(n10459), .B(n10458), .Z(n10738) );
  NANDN U13023 ( .A(n10461), .B(n10460), .Z(n10465) );
  NANDN U13024 ( .A(n10463), .B(n10462), .Z(n10464) );
  AND U13025 ( .A(n10465), .B(n10464), .Z(n10853) );
  NANDN U13026 ( .A(n10467), .B(n10466), .Z(n10471) );
  OR U13027 ( .A(n10469), .B(n10468), .Z(n10470) );
  AND U13028 ( .A(n10471), .B(n10470), .Z(n11204) );
  NANDN U13029 ( .A(n10473), .B(n10472), .Z(n10477) );
  NANDN U13030 ( .A(n10475), .B(n10474), .Z(n10476) );
  NAND U13031 ( .A(n10477), .B(n10476), .Z(n11205) );
  XNOR U13032 ( .A(n11204), .B(n11205), .Z(n11207) );
  NANDN U13033 ( .A(n10479), .B(n10478), .Z(n10483) );
  NANDN U13034 ( .A(n10481), .B(n10480), .Z(n10482) );
  AND U13035 ( .A(n10483), .B(n10482), .Z(n11206) );
  XNOR U13036 ( .A(n11207), .B(n11206), .Z(n10852) );
  XNOR U13037 ( .A(n10853), .B(n10852), .Z(n10854) );
  NANDN U13038 ( .A(n10485), .B(n10484), .Z(n10489) );
  NANDN U13039 ( .A(n10487), .B(n10486), .Z(n10488) );
  AND U13040 ( .A(n10489), .B(n10488), .Z(n10903) );
  NANDN U13041 ( .A(n10491), .B(n10490), .Z(n10495) );
  NANDN U13042 ( .A(n10493), .B(n10492), .Z(n10494) );
  AND U13043 ( .A(n10495), .B(n10494), .Z(n10901) );
  NANDN U13044 ( .A(n10497), .B(n10496), .Z(n10501) );
  NANDN U13045 ( .A(n10499), .B(n10498), .Z(n10500) );
  NAND U13046 ( .A(n10501), .B(n10500), .Z(n10900) );
  XNOR U13047 ( .A(n10901), .B(n10900), .Z(n10902) );
  XOR U13048 ( .A(n10903), .B(n10902), .Z(n10855) );
  XNOR U13049 ( .A(n10854), .B(n10855), .Z(n10739) );
  XOR U13050 ( .A(n10738), .B(n10739), .Z(n10741) );
  XOR U13051 ( .A(n10740), .B(n10741), .Z(n10624) );
  NAND U13052 ( .A(n10503), .B(n10502), .Z(n10507) );
  NAND U13053 ( .A(n10505), .B(n10504), .Z(n10506) );
  NAND U13054 ( .A(n10507), .B(n10506), .Z(n10622) );
  NANDN U13055 ( .A(n10509), .B(n10508), .Z(n10513) );
  NAND U13056 ( .A(n10511), .B(n10510), .Z(n10512) );
  AND U13057 ( .A(n10513), .B(n10512), .Z(n10885) );
  NANDN U13058 ( .A(n10515), .B(n10514), .Z(n10519) );
  NAND U13059 ( .A(n10517), .B(n10516), .Z(n10518) );
  AND U13060 ( .A(n10519), .B(n10518), .Z(n10883) );
  NANDN U13061 ( .A(n10521), .B(n10520), .Z(n10525) );
  NANDN U13062 ( .A(n10523), .B(n10522), .Z(n10524) );
  NAND U13063 ( .A(n10525), .B(n10524), .Z(n10882) );
  XNOR U13064 ( .A(n10883), .B(n10882), .Z(n10884) );
  XNOR U13065 ( .A(n10885), .B(n10884), .Z(n10732) );
  NANDN U13066 ( .A(n10527), .B(n10526), .Z(n10531) );
  NANDN U13067 ( .A(n10529), .B(n10528), .Z(n10530) );
  AND U13068 ( .A(n10531), .B(n10530), .Z(n10717) );
  NANDN U13069 ( .A(n10533), .B(n10532), .Z(n10537) );
  NANDN U13070 ( .A(n10535), .B(n10534), .Z(n10536) );
  AND U13071 ( .A(n10537), .B(n10536), .Z(n10715) );
  XNOR U13072 ( .A(n10715), .B(n10714), .Z(n10716) );
  XOR U13073 ( .A(n10717), .B(n10716), .Z(n10733) );
  XNOR U13074 ( .A(n10732), .B(n10733), .Z(n10734) );
  NANDN U13075 ( .A(n10543), .B(n10542), .Z(n10547) );
  NANDN U13076 ( .A(n10545), .B(n10544), .Z(n10546) );
  NAND U13077 ( .A(n10547), .B(n10546), .Z(n10735) );
  XNOR U13078 ( .A(n10734), .B(n10735), .Z(n10621) );
  XOR U13079 ( .A(n10622), .B(n10621), .Z(n10623) );
  XNOR U13080 ( .A(n10624), .B(n10623), .Z(n11273) );
  XOR U13081 ( .A(n11274), .B(n11273), .Z(n11276) );
  XNOR U13082 ( .A(n11275), .B(n11276), .Z(n11280) );
  NAND U13083 ( .A(n10549), .B(n10548), .Z(n10553) );
  NAND U13084 ( .A(n10551), .B(n10550), .Z(n10552) );
  NAND U13085 ( .A(n10553), .B(n10552), .Z(n11279) );
  XOR U13086 ( .A(n11280), .B(n11279), .Z(n11281) );
  XOR U13087 ( .A(n11282), .B(n11281), .Z(n10635) );
  XNOR U13088 ( .A(n10634), .B(n10635), .Z(n10554) );
  XOR U13089 ( .A(n10633), .B(n10554), .Z(o[3]) );
  NAND U13090 ( .A(n10556), .B(n10555), .Z(n10560) );
  NAND U13091 ( .A(n10558), .B(n10557), .Z(n10559) );
  NAND U13092 ( .A(n10560), .B(n10559), .Z(n11385) );
  NAND U13093 ( .A(n10562), .B(n10561), .Z(n10566) );
  NAND U13094 ( .A(n10564), .B(n10563), .Z(n10565) );
  AND U13095 ( .A(n10566), .B(n10565), .Z(n11367) );
  NANDN U13096 ( .A(n10568), .B(n10567), .Z(n10572) );
  NAND U13097 ( .A(n10570), .B(n10569), .Z(n10571) );
  AND U13098 ( .A(n10572), .B(n10571), .Z(n11642) );
  NAND U13099 ( .A(n10574), .B(n10573), .Z(n10578) );
  NAND U13100 ( .A(n10576), .B(n10575), .Z(n10577) );
  AND U13101 ( .A(n10578), .B(n10577), .Z(n11307) );
  NANDN U13102 ( .A(n10580), .B(n10579), .Z(n10584) );
  OR U13103 ( .A(n10582), .B(n10581), .Z(n10583) );
  AND U13104 ( .A(n10584), .B(n10583), .Z(n11592) );
  NANDN U13105 ( .A(n10586), .B(n10585), .Z(n10590) );
  NANDN U13106 ( .A(n10588), .B(n10587), .Z(n10589) );
  AND U13107 ( .A(n10590), .B(n10589), .Z(n11591) );
  XNOR U13108 ( .A(n11592), .B(n11591), .Z(n11594) );
  NANDN U13109 ( .A(n10592), .B(n10591), .Z(n10596) );
  NAND U13110 ( .A(n10594), .B(n10593), .Z(n10595) );
  AND U13111 ( .A(n10596), .B(n10595), .Z(n11593) );
  XNOR U13112 ( .A(n11594), .B(n11593), .Z(n11305) );
  NAND U13113 ( .A(n10598), .B(n10597), .Z(n10602) );
  NAND U13114 ( .A(n10600), .B(n10599), .Z(n10601) );
  NAND U13115 ( .A(n10602), .B(n10601), .Z(n11304) );
  XOR U13116 ( .A(n11305), .B(n11304), .Z(n11306) );
  XOR U13117 ( .A(n11307), .B(n11306), .Z(n11640) );
  NAND U13118 ( .A(n10604), .B(n10603), .Z(n10608) );
  NAND U13119 ( .A(n10606), .B(n10605), .Z(n10607) );
  AND U13120 ( .A(n10608), .B(n10607), .Z(n11639) );
  NAND U13121 ( .A(n10610), .B(n10609), .Z(n10614) );
  NAND U13122 ( .A(n10612), .B(n10611), .Z(n10613) );
  AND U13123 ( .A(n10614), .B(n10613), .Z(n11319) );
  NAND U13124 ( .A(n10616), .B(n10615), .Z(n10620) );
  NAND U13125 ( .A(n10618), .B(n10617), .Z(n10619) );
  AND U13126 ( .A(n10620), .B(n10619), .Z(n11316) );
  NAND U13127 ( .A(n10622), .B(n10621), .Z(n10626) );
  NAND U13128 ( .A(n10624), .B(n10623), .Z(n10625) );
  AND U13129 ( .A(n10626), .B(n10625), .Z(n11317) );
  XOR U13130 ( .A(n11316), .B(n11317), .Z(n11318) );
  XOR U13131 ( .A(n11319), .B(n11318), .Z(n11364) );
  XOR U13132 ( .A(n11365), .B(n11364), .Z(n11366) );
  XNOR U13133 ( .A(n11367), .B(n11366), .Z(n11383) );
  NAND U13134 ( .A(n10628), .B(n10627), .Z(n10632) );
  NAND U13135 ( .A(n10630), .B(n10629), .Z(n10631) );
  NAND U13136 ( .A(n10632), .B(n10631), .Z(n11382) );
  XOR U13137 ( .A(n11383), .B(n11382), .Z(n11384) );
  XNOR U13138 ( .A(n11385), .B(n11384), .Z(n11645) );
  NAND U13139 ( .A(n10637), .B(n10636), .Z(n10641) );
  NAND U13140 ( .A(n10639), .B(n10638), .Z(n10640) );
  NAND U13141 ( .A(n10641), .B(n10640), .Z(n11409) );
  NANDN U13142 ( .A(n10643), .B(n10642), .Z(n10647) );
  OR U13143 ( .A(n10645), .B(n10644), .Z(n10646) );
  AND U13144 ( .A(n10647), .B(n10646), .Z(n11457) );
  NANDN U13145 ( .A(n10649), .B(n10648), .Z(n10653) );
  OR U13146 ( .A(n10651), .B(n10650), .Z(n10652) );
  AND U13147 ( .A(n10653), .B(n10652), .Z(n11456) );
  NANDN U13148 ( .A(n10655), .B(n10654), .Z(n10659) );
  NANDN U13149 ( .A(n10657), .B(n10656), .Z(n10658) );
  NAND U13150 ( .A(n10659), .B(n10658), .Z(n11455) );
  XOR U13151 ( .A(n11456), .B(n11455), .Z(n11458) );
  XNOR U13152 ( .A(n11457), .B(n11458), .Z(n11407) );
  NAND U13153 ( .A(n10661), .B(n10660), .Z(n10665) );
  NAND U13154 ( .A(n10663), .B(n10662), .Z(n10664) );
  AND U13155 ( .A(n10665), .B(n10664), .Z(n11406) );
  XOR U13156 ( .A(n11407), .B(n11406), .Z(n11408) );
  XOR U13157 ( .A(n11409), .B(n11408), .Z(n11289) );
  NAND U13158 ( .A(n10667), .B(n10666), .Z(n10671) );
  NAND U13159 ( .A(n10669), .B(n10668), .Z(n10670) );
  AND U13160 ( .A(n10671), .B(n10670), .Z(n11343) );
  NAND U13161 ( .A(n10673), .B(n10672), .Z(n10677) );
  NAND U13162 ( .A(n10675), .B(n10674), .Z(n10676) );
  NAND U13163 ( .A(n10677), .B(n10676), .Z(n11341) );
  NANDN U13164 ( .A(n10679), .B(n10678), .Z(n10683) );
  OR U13165 ( .A(n10681), .B(n10680), .Z(n10682) );
  AND U13166 ( .A(n10683), .B(n10682), .Z(n11549) );
  NANDN U13167 ( .A(n10685), .B(n10684), .Z(n10689) );
  NANDN U13168 ( .A(n10687), .B(n10686), .Z(n10688) );
  AND U13169 ( .A(n10689), .B(n10688), .Z(n11547) );
  NANDN U13170 ( .A(n10691), .B(n10690), .Z(n10695) );
  NANDN U13171 ( .A(n10693), .B(n10692), .Z(n10694) );
  AND U13172 ( .A(n10695), .B(n10694), .Z(n11598) );
  NANDN U13173 ( .A(n10697), .B(n10696), .Z(n10701) );
  NAND U13174 ( .A(n10699), .B(n10698), .Z(n10700) );
  AND U13175 ( .A(n10701), .B(n10700), .Z(n11597) );
  XNOR U13176 ( .A(n11598), .B(n11597), .Z(n11599) );
  NANDN U13177 ( .A(n10703), .B(n10702), .Z(n10707) );
  NAND U13178 ( .A(n10705), .B(n10704), .Z(n10706) );
  NAND U13179 ( .A(n10707), .B(n10706), .Z(n11600) );
  XNOR U13180 ( .A(n11599), .B(n11600), .Z(n11546) );
  XNOR U13181 ( .A(n11547), .B(n11546), .Z(n11548) );
  XNOR U13182 ( .A(n11549), .B(n11548), .Z(n11340) );
  XOR U13183 ( .A(n11341), .B(n11340), .Z(n11342) );
  XOR U13184 ( .A(n11343), .B(n11342), .Z(n11287) );
  NANDN U13185 ( .A(n10709), .B(n10708), .Z(n10713) );
  OR U13186 ( .A(n10711), .B(n10710), .Z(n10712) );
  AND U13187 ( .A(n10713), .B(n10712), .Z(n11635) );
  NANDN U13188 ( .A(n10715), .B(n10714), .Z(n10719) );
  NANDN U13189 ( .A(n10717), .B(n10716), .Z(n10718) );
  AND U13190 ( .A(n10719), .B(n10718), .Z(n11634) );
  NANDN U13191 ( .A(n10721), .B(n10720), .Z(n10725) );
  NANDN U13192 ( .A(n10723), .B(n10722), .Z(n10724) );
  NAND U13193 ( .A(n10725), .B(n10724), .Z(n11633) );
  XOR U13194 ( .A(n11634), .B(n11633), .Z(n11636) );
  XOR U13195 ( .A(n11635), .B(n11636), .Z(n11469) );
  NANDN U13196 ( .A(n10727), .B(n10726), .Z(n10731) );
  NANDN U13197 ( .A(n10729), .B(n10728), .Z(n10730) );
  AND U13198 ( .A(n10731), .B(n10730), .Z(n11468) );
  XNOR U13199 ( .A(n11469), .B(n11468), .Z(n11470) );
  NANDN U13200 ( .A(n10733), .B(n10732), .Z(n10737) );
  NANDN U13201 ( .A(n10735), .B(n10734), .Z(n10736) );
  NAND U13202 ( .A(n10737), .B(n10736), .Z(n11471) );
  XNOR U13203 ( .A(n11470), .B(n11471), .Z(n11286) );
  XOR U13204 ( .A(n11289), .B(n11288), .Z(n11353) );
  NAND U13205 ( .A(n10739), .B(n10738), .Z(n10743) );
  NAND U13206 ( .A(n10741), .B(n10740), .Z(n10742) );
  AND U13207 ( .A(n10743), .B(n10742), .Z(n11561) );
  NANDN U13208 ( .A(n10745), .B(n10744), .Z(n10749) );
  NANDN U13209 ( .A(n10747), .B(n10746), .Z(n10748) );
  AND U13210 ( .A(n10749), .B(n10748), .Z(n11630) );
  NANDN U13211 ( .A(n10751), .B(n10750), .Z(n10755) );
  NANDN U13212 ( .A(n10753), .B(n10752), .Z(n10754) );
  AND U13213 ( .A(n10755), .B(n10754), .Z(n11628) );
  NANDN U13214 ( .A(n10757), .B(n10756), .Z(n10761) );
  NANDN U13215 ( .A(n10759), .B(n10758), .Z(n10760) );
  AND U13216 ( .A(n10761), .B(n10760), .Z(n11627) );
  XNOR U13217 ( .A(n11628), .B(n11627), .Z(n11629) );
  XOR U13218 ( .A(n11630), .B(n11629), .Z(n11559) );
  NAND U13219 ( .A(n10763), .B(n10762), .Z(n10767) );
  NAND U13220 ( .A(n10765), .B(n10764), .Z(n10766) );
  NAND U13221 ( .A(n10767), .B(n10766), .Z(n11558) );
  XOR U13222 ( .A(n11559), .B(n11558), .Z(n11560) );
  XNOR U13223 ( .A(n11561), .B(n11560), .Z(n11395) );
  NAND U13224 ( .A(n10769), .B(n10768), .Z(n10773) );
  NAND U13225 ( .A(n10771), .B(n10770), .Z(n10772) );
  AND U13226 ( .A(n10773), .B(n10772), .Z(n11394) );
  XOR U13227 ( .A(n11395), .B(n11394), .Z(n11397) );
  NAND U13228 ( .A(n10775), .B(n10774), .Z(n10779) );
  NAND U13229 ( .A(n10777), .B(n10776), .Z(n10778) );
  NAND U13230 ( .A(n10779), .B(n10778), .Z(n11403) );
  NAND U13231 ( .A(n10781), .B(n10780), .Z(n10785) );
  NAND U13232 ( .A(n10783), .B(n10782), .Z(n10784) );
  NAND U13233 ( .A(n10785), .B(n10784), .Z(n11401) );
  NANDN U13234 ( .A(n10787), .B(n10786), .Z(n10791) );
  NAND U13235 ( .A(n10789), .B(n10788), .Z(n10790) );
  AND U13236 ( .A(n10791), .B(n10790), .Z(n11618) );
  NANDN U13237 ( .A(n10793), .B(n10792), .Z(n10797) );
  NAND U13238 ( .A(n10795), .B(n10794), .Z(n10796) );
  AND U13239 ( .A(n10797), .B(n10796), .Z(n11616) );
  NANDN U13240 ( .A(n10799), .B(n10798), .Z(n10803) );
  NANDN U13241 ( .A(n10801), .B(n10800), .Z(n10802) );
  AND U13242 ( .A(n10803), .B(n10802), .Z(n11615) );
  XNOR U13243 ( .A(n11616), .B(n11615), .Z(n11617) );
  XOR U13244 ( .A(n11618), .B(n11617), .Z(n11493) );
  NANDN U13245 ( .A(n10805), .B(n10804), .Z(n10809) );
  NAND U13246 ( .A(n10807), .B(n10806), .Z(n10808) );
  AND U13247 ( .A(n10809), .B(n10808), .Z(n11481) );
  NANDN U13248 ( .A(n10811), .B(n10810), .Z(n10815) );
  NANDN U13249 ( .A(n10813), .B(n10812), .Z(n10814) );
  AND U13250 ( .A(n10815), .B(n10814), .Z(n11480) );
  XNOR U13251 ( .A(n11481), .B(n11480), .Z(n11482) );
  NANDN U13252 ( .A(n10817), .B(n10816), .Z(n10821) );
  NANDN U13253 ( .A(n10819), .B(n10818), .Z(n10820) );
  NAND U13254 ( .A(n10821), .B(n10820), .Z(n11483) );
  XNOR U13255 ( .A(n11482), .B(n11483), .Z(n11492) );
  XNOR U13256 ( .A(n11493), .B(n11492), .Z(n11495) );
  NANDN U13257 ( .A(n10823), .B(n10822), .Z(n10827) );
  NAND U13258 ( .A(n10825), .B(n10824), .Z(n10826) );
  AND U13259 ( .A(n10827), .B(n10826), .Z(n11494) );
  XNOR U13260 ( .A(n11495), .B(n11494), .Z(n11400) );
  XOR U13261 ( .A(n11401), .B(n11400), .Z(n11402) );
  XOR U13262 ( .A(n11403), .B(n11402), .Z(n11396) );
  XOR U13263 ( .A(n11397), .B(n11396), .Z(n11352) );
  NANDN U13264 ( .A(n10829), .B(n10828), .Z(n10833) );
  NANDN U13265 ( .A(n10831), .B(n10830), .Z(n10832) );
  AND U13266 ( .A(n10833), .B(n10832), .Z(n11313) );
  NANDN U13267 ( .A(n10835), .B(n10834), .Z(n10839) );
  NAND U13268 ( .A(n10837), .B(n10836), .Z(n10838) );
  AND U13269 ( .A(n10839), .B(n10838), .Z(n11311) );
  NANDN U13270 ( .A(n10841), .B(n10840), .Z(n10845) );
  NANDN U13271 ( .A(n10843), .B(n10842), .Z(n10844) );
  AND U13272 ( .A(n10845), .B(n10844), .Z(n11531) );
  NANDN U13273 ( .A(n10847), .B(n10846), .Z(n10851) );
  NANDN U13274 ( .A(n10849), .B(n10848), .Z(n10850) );
  AND U13275 ( .A(n10851), .B(n10850), .Z(n11529) );
  NANDN U13276 ( .A(n10853), .B(n10852), .Z(n10857) );
  NANDN U13277 ( .A(n10855), .B(n10854), .Z(n10856) );
  NAND U13278 ( .A(n10857), .B(n10856), .Z(n11528) );
  XNOR U13279 ( .A(n11529), .B(n11528), .Z(n11530) );
  XNOR U13280 ( .A(n11531), .B(n11530), .Z(n11334) );
  NANDN U13281 ( .A(n10859), .B(n10858), .Z(n10863) );
  OR U13282 ( .A(n10861), .B(n10860), .Z(n10862) );
  AND U13283 ( .A(n10863), .B(n10862), .Z(n11525) );
  NANDN U13284 ( .A(n10865), .B(n10864), .Z(n10869) );
  NANDN U13285 ( .A(n10867), .B(n10866), .Z(n10868) );
  AND U13286 ( .A(n10869), .B(n10868), .Z(n11523) );
  NANDN U13287 ( .A(n10871), .B(n10870), .Z(n10875) );
  NANDN U13288 ( .A(n10873), .B(n10872), .Z(n10874) );
  NAND U13289 ( .A(n10875), .B(n10874), .Z(n11522) );
  XNOR U13290 ( .A(n11523), .B(n11522), .Z(n11524) );
  XNOR U13291 ( .A(n11525), .B(n11524), .Z(n11335) );
  XOR U13292 ( .A(n11334), .B(n11335), .Z(n11336) );
  NANDN U13293 ( .A(n10877), .B(n10876), .Z(n10881) );
  OR U13294 ( .A(n10879), .B(n10878), .Z(n10880) );
  AND U13295 ( .A(n10881), .B(n10880), .Z(n11624) );
  NANDN U13296 ( .A(n10883), .B(n10882), .Z(n10887) );
  NANDN U13297 ( .A(n10885), .B(n10884), .Z(n10886) );
  AND U13298 ( .A(n10887), .B(n10886), .Z(n11622) );
  NANDN U13299 ( .A(n10889), .B(n10888), .Z(n10893) );
  NAND U13300 ( .A(n10891), .B(n10890), .Z(n10892) );
  AND U13301 ( .A(n10893), .B(n10892), .Z(n11488) );
  NANDN U13302 ( .A(n10895), .B(n10894), .Z(n10899) );
  NANDN U13303 ( .A(n10897), .B(n10896), .Z(n10898) );
  AND U13304 ( .A(n10899), .B(n10898), .Z(n11487) );
  NANDN U13305 ( .A(n10901), .B(n10900), .Z(n10905) );
  NANDN U13306 ( .A(n10903), .B(n10902), .Z(n10904) );
  AND U13307 ( .A(n10905), .B(n10904), .Z(n11486) );
  XOR U13308 ( .A(n11487), .B(n11486), .Z(n11489) );
  XNOR U13309 ( .A(n11488), .B(n11489), .Z(n11621) );
  XNOR U13310 ( .A(n11622), .B(n11621), .Z(n11623) );
  XNOR U13311 ( .A(n11624), .B(n11623), .Z(n11337) );
  XOR U13312 ( .A(n11336), .B(n11337), .Z(n11310) );
  XNOR U13313 ( .A(n11355), .B(n11354), .Z(n11372) );
  NAND U13314 ( .A(n10907), .B(n10906), .Z(n10911) );
  NAND U13315 ( .A(n10909), .B(n10908), .Z(n10910) );
  NAND U13316 ( .A(n10911), .B(n10910), .Z(n11370) );
  NAND U13317 ( .A(n10913), .B(n10912), .Z(n10917) );
  NAND U13318 ( .A(n10915), .B(n10914), .Z(n10916) );
  AND U13319 ( .A(n10917), .B(n10916), .Z(n11391) );
  NAND U13320 ( .A(n10919), .B(n10918), .Z(n10923) );
  NAND U13321 ( .A(n10921), .B(n10920), .Z(n10922) );
  AND U13322 ( .A(n10923), .B(n10922), .Z(n11389) );
  NANDN U13323 ( .A(n10925), .B(n10924), .Z(n10929) );
  NAND U13324 ( .A(n10927), .B(n10926), .Z(n10928) );
  AND U13325 ( .A(n10929), .B(n10928), .Z(n11477) );
  NANDN U13326 ( .A(n10931), .B(n10930), .Z(n10935) );
  NAND U13327 ( .A(n10933), .B(n10932), .Z(n10934) );
  AND U13328 ( .A(n10935), .B(n10934), .Z(n11475) );
  NANDN U13329 ( .A(n10937), .B(n10936), .Z(n10941) );
  NAND U13330 ( .A(n10939), .B(n10938), .Z(n10940) );
  NAND U13331 ( .A(n10941), .B(n10940), .Z(n11474) );
  XNOR U13332 ( .A(n11475), .B(n11474), .Z(n11476) );
  XNOR U13333 ( .A(n11477), .B(n11476), .Z(n11537) );
  NANDN U13334 ( .A(n10943), .B(n10942), .Z(n10947) );
  NANDN U13335 ( .A(n10945), .B(n10944), .Z(n10946) );
  AND U13336 ( .A(n10947), .B(n10946), .Z(n11513) );
  NANDN U13337 ( .A(n10949), .B(n10948), .Z(n10953) );
  OR U13338 ( .A(n10951), .B(n10950), .Z(n10952) );
  AND U13339 ( .A(n10953), .B(n10952), .Z(n11510) );
  NANDN U13340 ( .A(n10955), .B(n10954), .Z(n10959) );
  OR U13341 ( .A(n10957), .B(n10956), .Z(n10958) );
  NAND U13342 ( .A(n10959), .B(n10958), .Z(n11511) );
  XNOR U13343 ( .A(n11510), .B(n11511), .Z(n11512) );
  XOR U13344 ( .A(n11513), .B(n11512), .Z(n11535) );
  NANDN U13345 ( .A(n10961), .B(n10960), .Z(n10965) );
  NANDN U13346 ( .A(n10963), .B(n10962), .Z(n10964) );
  AND U13347 ( .A(n10965), .B(n10964), .Z(n11534) );
  XNOR U13348 ( .A(n11535), .B(n11534), .Z(n11536) );
  XNOR U13349 ( .A(n11537), .B(n11536), .Z(n11329) );
  NANDN U13350 ( .A(n10967), .B(n10966), .Z(n10971) );
  NANDN U13351 ( .A(n10969), .B(n10968), .Z(n10970) );
  AND U13352 ( .A(n10971), .B(n10970), .Z(n11499) );
  NAND U13353 ( .A(n10973), .B(n10972), .Z(n10977) );
  NAND U13354 ( .A(n10975), .B(n10974), .Z(n10976) );
  AND U13355 ( .A(n10977), .B(n10976), .Z(n11427) );
  NAND U13356 ( .A(n10979), .B(n10978), .Z(n10983) );
  NAND U13357 ( .A(n10981), .B(n10980), .Z(n10982) );
  AND U13358 ( .A(n10983), .B(n10982), .Z(n11426) );
  NANDN U13359 ( .A(n10985), .B(n10984), .Z(n10989) );
  NAND U13360 ( .A(n10987), .B(n10986), .Z(n10988) );
  NAND U13361 ( .A(n10989), .B(n10988), .Z(n11425) );
  XOR U13362 ( .A(n11426), .B(n11425), .Z(n11428) );
  XOR U13363 ( .A(n11427), .B(n11428), .Z(n11572) );
  NANDN U13364 ( .A(n10991), .B(n10990), .Z(n10995) );
  NANDN U13365 ( .A(n10993), .B(n10992), .Z(n10994) );
  AND U13366 ( .A(n10995), .B(n10994), .Z(n11421) );
  NANDN U13367 ( .A(n10997), .B(n10996), .Z(n11001) );
  NAND U13368 ( .A(n10999), .B(n10998), .Z(n11000) );
  AND U13369 ( .A(n11001), .B(n11000), .Z(n11420) );
  NAND U13370 ( .A(n11003), .B(n11002), .Z(n11007) );
  NAND U13371 ( .A(n11005), .B(n11004), .Z(n11006) );
  NAND U13372 ( .A(n11007), .B(n11006), .Z(n11419) );
  XOR U13373 ( .A(n11420), .B(n11419), .Z(n11422) );
  XOR U13374 ( .A(n11421), .B(n11422), .Z(n11571) );
  NANDN U13375 ( .A(n11009), .B(n11008), .Z(n11013) );
  NAND U13376 ( .A(n11011), .B(n11010), .Z(n11012) );
  AND U13377 ( .A(n11013), .B(n11012), .Z(n11570) );
  XOR U13378 ( .A(n11571), .B(n11570), .Z(n11573) );
  XNOR U13379 ( .A(n11572), .B(n11573), .Z(n11498) );
  XNOR U13380 ( .A(n11499), .B(n11498), .Z(n11500) );
  NANDN U13381 ( .A(n11015), .B(n11014), .Z(n11019) );
  NANDN U13382 ( .A(n11017), .B(n11016), .Z(n11018) );
  AND U13383 ( .A(n11019), .B(n11018), .Z(n11567) );
  NANDN U13384 ( .A(n11021), .B(n11020), .Z(n11025) );
  NANDN U13385 ( .A(n11023), .B(n11022), .Z(n11024) );
  AND U13386 ( .A(n11025), .B(n11024), .Z(n11565) );
  NAND U13387 ( .A(n11027), .B(n11026), .Z(n11031) );
  NAND U13388 ( .A(n11029), .B(n11028), .Z(n11030) );
  AND U13389 ( .A(n11031), .B(n11030), .Z(n11415) );
  NANDN U13390 ( .A(n11033), .B(n11032), .Z(n11037) );
  NAND U13391 ( .A(n11035), .B(n11034), .Z(n11036) );
  AND U13392 ( .A(n11037), .B(n11036), .Z(n11414) );
  NAND U13393 ( .A(n11039), .B(n11038), .Z(n11043) );
  NAND U13394 ( .A(n11041), .B(n11040), .Z(n11042) );
  NAND U13395 ( .A(n11043), .B(n11042), .Z(n11413) );
  XOR U13396 ( .A(n11414), .B(n11413), .Z(n11416) );
  XNOR U13397 ( .A(n11415), .B(n11416), .Z(n11564) );
  XNOR U13398 ( .A(n11565), .B(n11564), .Z(n11566) );
  XOR U13399 ( .A(n11567), .B(n11566), .Z(n11501) );
  XNOR U13400 ( .A(n11500), .B(n11501), .Z(n11328) );
  XOR U13401 ( .A(n11329), .B(n11328), .Z(n11330) );
  XNOR U13402 ( .A(n11610), .B(n11609), .Z(n11054) );
  XOR U13403 ( .A(n11611), .B(n11054), .Z(n11543) );
  NANDN U13404 ( .A(n11056), .B(n11055), .Z(n11060) );
  NANDN U13405 ( .A(n11058), .B(n11057), .Z(n11059) );
  AND U13406 ( .A(n11060), .B(n11059), .Z(n11541) );
  NANDN U13407 ( .A(n11062), .B(n11061), .Z(n11066) );
  NANDN U13408 ( .A(n11064), .B(n11063), .Z(n11065) );
  AND U13409 ( .A(n11066), .B(n11065), .Z(n11439) );
  NANDN U13410 ( .A(n11068), .B(n11067), .Z(n11072) );
  NANDN U13411 ( .A(n11070), .B(n11069), .Z(n11071) );
  AND U13412 ( .A(n11072), .B(n11071), .Z(n11438) );
  NANDN U13413 ( .A(n11074), .B(n11073), .Z(n11078) );
  NAND U13414 ( .A(n11076), .B(n11075), .Z(n11077) );
  NAND U13415 ( .A(n11078), .B(n11077), .Z(n11437) );
  XOR U13416 ( .A(n11438), .B(n11437), .Z(n11440) );
  XOR U13417 ( .A(n11439), .B(n11440), .Z(n11445) );
  NANDN U13418 ( .A(n11080), .B(n11079), .Z(n11084) );
  NAND U13419 ( .A(n11082), .B(n11081), .Z(n11083) );
  AND U13420 ( .A(n11084), .B(n11083), .Z(n11433) );
  NANDN U13421 ( .A(n11086), .B(n11085), .Z(n11090) );
  NANDN U13422 ( .A(n11088), .B(n11087), .Z(n11089) );
  AND U13423 ( .A(n11090), .B(n11089), .Z(n11432) );
  NANDN U13424 ( .A(n11092), .B(n11091), .Z(n11096) );
  NAND U13425 ( .A(n11094), .B(n11093), .Z(n11095) );
  NAND U13426 ( .A(n11096), .B(n11095), .Z(n11431) );
  XOR U13427 ( .A(n11432), .B(n11431), .Z(n11434) );
  XOR U13428 ( .A(n11433), .B(n11434), .Z(n11444) );
  NANDN U13429 ( .A(n11098), .B(n11097), .Z(n11102) );
  NAND U13430 ( .A(n11100), .B(n11099), .Z(n11101) );
  NAND U13431 ( .A(n11102), .B(n11101), .Z(n11443) );
  XOR U13432 ( .A(n11444), .B(n11443), .Z(n11446) );
  XNOR U13433 ( .A(n11445), .B(n11446), .Z(n11540) );
  XNOR U13434 ( .A(n11541), .B(n11540), .Z(n11542) );
  XNOR U13435 ( .A(n11543), .B(n11542), .Z(n11331) );
  XOR U13436 ( .A(n11330), .B(n11331), .Z(n11388) );
  XOR U13437 ( .A(n11389), .B(n11388), .Z(n11390) );
  XOR U13438 ( .A(n11391), .B(n11390), .Z(n11361) );
  NAND U13439 ( .A(n11104), .B(n11103), .Z(n11108) );
  NAND U13440 ( .A(n11106), .B(n11105), .Z(n11107) );
  AND U13441 ( .A(n11108), .B(n11107), .Z(n11359) );
  NAND U13442 ( .A(n11110), .B(n11109), .Z(n11114) );
  NAND U13443 ( .A(n11112), .B(n11111), .Z(n11113) );
  NAND U13444 ( .A(n11114), .B(n11113), .Z(n11292) );
  NANDN U13445 ( .A(n11116), .B(n11115), .Z(n11120) );
  NANDN U13446 ( .A(n11118), .B(n11117), .Z(n11119) );
  AND U13447 ( .A(n11120), .B(n11119), .Z(n11614) );
  XNOR U13448 ( .A(n11613), .B(n11612), .Z(n11127) );
  XOR U13449 ( .A(n11614), .B(n11127), .Z(n11553) );
  NANDN U13450 ( .A(n11129), .B(n11128), .Z(n11133) );
  NANDN U13451 ( .A(n11131), .B(n11130), .Z(n11132) );
  AND U13452 ( .A(n11133), .B(n11132), .Z(n11552) );
  XNOR U13453 ( .A(n11553), .B(n11552), .Z(n11554) );
  NANDN U13454 ( .A(n11135), .B(n11134), .Z(n11139) );
  NANDN U13455 ( .A(n11137), .B(n11136), .Z(n11138) );
  AND U13456 ( .A(n11139), .B(n11138), .Z(n11606) );
  NANDN U13457 ( .A(n11145), .B(n11144), .Z(n11149) );
  NANDN U13458 ( .A(n11147), .B(n11146), .Z(n11148) );
  AND U13459 ( .A(n11149), .B(n11148), .Z(n11603) );
  XNOR U13460 ( .A(n11604), .B(n11603), .Z(n11605) );
  XOR U13461 ( .A(n11606), .B(n11605), .Z(n11555) );
  XNOR U13462 ( .A(n11554), .B(n11555), .Z(n11293) );
  XOR U13463 ( .A(n11292), .B(n11293), .Z(n11295) );
  NANDN U13464 ( .A(n11151), .B(n11150), .Z(n11155) );
  NAND U13465 ( .A(n11153), .B(n11152), .Z(n11154) );
  AND U13466 ( .A(n11155), .B(n11154), .Z(n11506) );
  NANDN U13467 ( .A(n11157), .B(n11156), .Z(n11161) );
  NANDN U13468 ( .A(n11159), .B(n11158), .Z(n11160) );
  AND U13469 ( .A(n11161), .B(n11160), .Z(n11577) );
  NAND U13470 ( .A(n11163), .B(n11162), .Z(n11167) );
  NAND U13471 ( .A(n11165), .B(n11164), .Z(n11166) );
  NAND U13472 ( .A(n11167), .B(n11166), .Z(n11576) );
  XNOR U13473 ( .A(n11577), .B(n11576), .Z(n11579) );
  NANDN U13474 ( .A(n11169), .B(n11168), .Z(n11173) );
  NAND U13475 ( .A(n11171), .B(n11170), .Z(n11172) );
  NAND U13476 ( .A(n11173), .B(n11172), .Z(n11412) );
  XOR U13477 ( .A(n11412), .B(oglobal[4]), .Z(n11578) );
  XOR U13478 ( .A(n11579), .B(n11578), .Z(n11505) );
  NANDN U13479 ( .A(n11175), .B(n11174), .Z(n11179) );
  NAND U13480 ( .A(n11177), .B(n11176), .Z(n11178) );
  NAND U13481 ( .A(n11179), .B(n11178), .Z(n11504) );
  XOR U13482 ( .A(n11505), .B(n11504), .Z(n11507) );
  XOR U13483 ( .A(n11506), .B(n11507), .Z(n11452) );
  NANDN U13484 ( .A(n11181), .B(n11180), .Z(n11185) );
  NANDN U13485 ( .A(n11183), .B(n11182), .Z(n11184) );
  AND U13486 ( .A(n11185), .B(n11184), .Z(n11450) );
  NANDN U13487 ( .A(n11187), .B(n11186), .Z(n11191) );
  NAND U13488 ( .A(n11189), .B(n11188), .Z(n11190) );
  AND U13489 ( .A(n11191), .B(n11190), .Z(n11587) );
  NANDN U13490 ( .A(n11193), .B(n11192), .Z(n11197) );
  NAND U13491 ( .A(n11195), .B(n11194), .Z(n11196) );
  AND U13492 ( .A(n11197), .B(n11196), .Z(n11586) );
  NANDN U13493 ( .A(n11199), .B(n11198), .Z(n11203) );
  NAND U13494 ( .A(n11201), .B(n11200), .Z(n11202) );
  NAND U13495 ( .A(n11203), .B(n11202), .Z(n11585) );
  XOR U13496 ( .A(n11586), .B(n11585), .Z(n11588) );
  XOR U13497 ( .A(n11587), .B(n11588), .Z(n11518) );
  NANDN U13498 ( .A(n11205), .B(n11204), .Z(n11209) );
  NAND U13499 ( .A(n11207), .B(n11206), .Z(n11208) );
  AND U13500 ( .A(n11209), .B(n11208), .Z(n11517) );
  NANDN U13501 ( .A(n11211), .B(n11210), .Z(n11215) );
  NANDN U13502 ( .A(n11213), .B(n11212), .Z(n11214) );
  AND U13503 ( .A(n11215), .B(n11214), .Z(n11584) );
  NANDN U13504 ( .A(n11216), .B(oglobal[3]), .Z(n11220) );
  NANDN U13505 ( .A(n11218), .B(n11217), .Z(n11219) );
  NAND U13506 ( .A(n11220), .B(n11219), .Z(n11582) );
  XOR U13507 ( .A(n11582), .B(n11583), .Z(n11224) );
  XNOR U13508 ( .A(n11584), .B(n11224), .Z(n11516) );
  XOR U13509 ( .A(n11517), .B(n11516), .Z(n11519) );
  XNOR U13510 ( .A(n11518), .B(n11519), .Z(n11449) );
  XNOR U13511 ( .A(n11450), .B(n11449), .Z(n11451) );
  XNOR U13512 ( .A(n11452), .B(n11451), .Z(n11294) );
  XNOR U13513 ( .A(n11295), .B(n11294), .Z(n11323) );
  NAND U13514 ( .A(n11226), .B(n11225), .Z(n11230) );
  NAND U13515 ( .A(n11228), .B(n11227), .Z(n11229) );
  AND U13516 ( .A(n11230), .B(n11229), .Z(n11322) );
  XOR U13517 ( .A(n11323), .B(n11322), .Z(n11324) );
  NANDN U13518 ( .A(n11232), .B(n11231), .Z(n11236) );
  NAND U13519 ( .A(n11234), .B(n11233), .Z(n11235) );
  AND U13520 ( .A(n11236), .B(n11235), .Z(n11299) );
  NANDN U13521 ( .A(n11238), .B(n11237), .Z(n11242) );
  NAND U13522 ( .A(n11240), .B(n11239), .Z(n11241) );
  NAND U13523 ( .A(n11242), .B(n11241), .Z(n11298) );
  XOR U13524 ( .A(n11299), .B(n11298), .Z(n11301) );
  NANDN U13525 ( .A(n11244), .B(n11243), .Z(n11248) );
  NANDN U13526 ( .A(n11246), .B(n11245), .Z(n11247) );
  AND U13527 ( .A(n11248), .B(n11247), .Z(n11300) );
  XOR U13528 ( .A(n11301), .B(n11300), .Z(n11465) );
  NANDN U13529 ( .A(n11250), .B(n11249), .Z(n11254) );
  NANDN U13530 ( .A(n11252), .B(n11251), .Z(n11253) );
  AND U13531 ( .A(n11254), .B(n11253), .Z(n11462) );
  NANDN U13532 ( .A(n11256), .B(n11255), .Z(n11260) );
  NANDN U13533 ( .A(n11258), .B(n11257), .Z(n11259) );
  NAND U13534 ( .A(n11260), .B(n11259), .Z(n11463) );
  XNOR U13535 ( .A(n11462), .B(n11463), .Z(n11464) );
  XNOR U13536 ( .A(n11465), .B(n11464), .Z(n11325) );
  XOR U13537 ( .A(n11324), .B(n11325), .Z(n11358) );
  XOR U13538 ( .A(n11359), .B(n11358), .Z(n11360) );
  XOR U13539 ( .A(n11370), .B(n11371), .Z(n11373) );
  XOR U13540 ( .A(n11372), .B(n11373), .Z(n11378) );
  NAND U13541 ( .A(n11262), .B(n11261), .Z(n11266) );
  NAND U13542 ( .A(n11264), .B(n11263), .Z(n11265) );
  AND U13543 ( .A(n11266), .B(n11265), .Z(n11349) );
  NAND U13544 ( .A(n11268), .B(n11267), .Z(n11272) );
  NAND U13545 ( .A(n11270), .B(n11269), .Z(n11271) );
  AND U13546 ( .A(n11272), .B(n11271), .Z(n11347) );
  NAND U13547 ( .A(n11274), .B(n11273), .Z(n11278) );
  NAND U13548 ( .A(n11276), .B(n11275), .Z(n11277) );
  NAND U13549 ( .A(n11278), .B(n11277), .Z(n11346) );
  NAND U13550 ( .A(n11280), .B(n11279), .Z(n11284) );
  NAND U13551 ( .A(n11282), .B(n11281), .Z(n11283) );
  NAND U13552 ( .A(n11284), .B(n11283), .Z(n11376) );
  XOR U13553 ( .A(n11377), .B(n11376), .Z(n11379) );
  XOR U13554 ( .A(n11378), .B(n11379), .Z(n11647) );
  XNOR U13555 ( .A(n11646), .B(n11647), .Z(n11285) );
  XNOR U13556 ( .A(n11645), .B(n11285), .Z(o[4]) );
  NANDN U13557 ( .A(n11287), .B(n11286), .Z(n11291) );
  NAND U13558 ( .A(n11289), .B(n11288), .Z(n11290) );
  NAND U13559 ( .A(n11291), .B(n11290), .Z(n11663) );
  NAND U13560 ( .A(n11293), .B(n11292), .Z(n11297) );
  NAND U13561 ( .A(n11295), .B(n11294), .Z(n11296) );
  NAND U13562 ( .A(n11297), .B(n11296), .Z(n11695) );
  NAND U13563 ( .A(n11299), .B(n11298), .Z(n11303) );
  NAND U13564 ( .A(n11301), .B(n11300), .Z(n11302) );
  NAND U13565 ( .A(n11303), .B(n11302), .Z(n11693) );
  NAND U13566 ( .A(n11305), .B(n11304), .Z(n11309) );
  NAND U13567 ( .A(n11307), .B(n11306), .Z(n11308) );
  NAND U13568 ( .A(n11309), .B(n11308), .Z(n11692) );
  XOR U13569 ( .A(n11693), .B(n11692), .Z(n11694) );
  XOR U13570 ( .A(n11695), .B(n11694), .Z(n11662) );
  NANDN U13571 ( .A(n11311), .B(n11310), .Z(n11315) );
  NANDN U13572 ( .A(n11313), .B(n11312), .Z(n11314) );
  AND U13573 ( .A(n11315), .B(n11314), .Z(n11661) );
  XOR U13574 ( .A(n11663), .B(n11664), .Z(n11708) );
  NAND U13575 ( .A(n11317), .B(n11316), .Z(n11321) );
  NANDN U13576 ( .A(n11319), .B(n11318), .Z(n11320) );
  AND U13577 ( .A(n11321), .B(n11320), .Z(n11716) );
  NAND U13578 ( .A(n11323), .B(n11322), .Z(n11327) );
  NAND U13579 ( .A(n11325), .B(n11324), .Z(n11326) );
  NAND U13580 ( .A(n11327), .B(n11326), .Z(n11714) );
  NAND U13581 ( .A(n11329), .B(n11328), .Z(n11333) );
  NAND U13582 ( .A(n11331), .B(n11330), .Z(n11332) );
  NAND U13583 ( .A(n11333), .B(n11332), .Z(n11682) );
  NAND U13584 ( .A(n11335), .B(n11334), .Z(n11339) );
  NAND U13585 ( .A(n11337), .B(n11336), .Z(n11338) );
  NAND U13586 ( .A(n11339), .B(n11338), .Z(n11681) );
  NAND U13587 ( .A(n11341), .B(n11340), .Z(n11345) );
  NAND U13588 ( .A(n11343), .B(n11342), .Z(n11344) );
  NAND U13589 ( .A(n11345), .B(n11344), .Z(n11680) );
  XNOR U13590 ( .A(n11681), .B(n11680), .Z(n11683) );
  XOR U13591 ( .A(n11682), .B(n11683), .Z(n11713) );
  XOR U13592 ( .A(n11714), .B(n11713), .Z(n11715) );
  XOR U13593 ( .A(n11716), .B(n11715), .Z(n11707) );
  XOR U13594 ( .A(n11708), .B(n11707), .Z(n11709) );
  NANDN U13595 ( .A(n11347), .B(n11346), .Z(n11351) );
  NANDN U13596 ( .A(n11349), .B(n11348), .Z(n11350) );
  NAND U13597 ( .A(n11351), .B(n11350), .Z(n11710) );
  NANDN U13598 ( .A(n11353), .B(n11352), .Z(n11357) );
  NAND U13599 ( .A(n11355), .B(n11354), .Z(n11356) );
  AND U13600 ( .A(n11357), .B(n11356), .Z(n11658) );
  NAND U13601 ( .A(n11359), .B(n11358), .Z(n11363) );
  NANDN U13602 ( .A(n11361), .B(n11360), .Z(n11362) );
  AND U13603 ( .A(n11363), .B(n11362), .Z(n11656) );
  NAND U13604 ( .A(n11365), .B(n11364), .Z(n11369) );
  NAND U13605 ( .A(n11367), .B(n11366), .Z(n11368) );
  AND U13606 ( .A(n11369), .B(n11368), .Z(n11655) );
  XOR U13607 ( .A(n11658), .B(n11657), .Z(n11650) );
  NANDN U13608 ( .A(n11371), .B(n11370), .Z(n11375) );
  NANDN U13609 ( .A(n11373), .B(n11372), .Z(n11374) );
  AND U13610 ( .A(n11375), .B(n11374), .Z(n11651) );
  XNOR U13611 ( .A(n11652), .B(n11651), .Z(n11706) );
  NAND U13612 ( .A(n11377), .B(n11376), .Z(n11381) );
  NAND U13613 ( .A(n11379), .B(n11378), .Z(n11380) );
  AND U13614 ( .A(n11381), .B(n11380), .Z(n11700) );
  NAND U13615 ( .A(n11383), .B(n11382), .Z(n11387) );
  NAND U13616 ( .A(n11385), .B(n11384), .Z(n11386) );
  NAND U13617 ( .A(n11387), .B(n11386), .Z(n11698) );
  NAND U13618 ( .A(n11389), .B(n11388), .Z(n11393) );
  NAND U13619 ( .A(n11391), .B(n11390), .Z(n11392) );
  NAND U13620 ( .A(n11393), .B(n11392), .Z(n11675) );
  IV U13621 ( .A(n11675), .Z(n11673) );
  NAND U13622 ( .A(n11395), .B(n11394), .Z(n11399) );
  NAND U13623 ( .A(n11397), .B(n11396), .Z(n11398) );
  AND U13624 ( .A(n11399), .B(n11398), .Z(n11677) );
  NAND U13625 ( .A(n11401), .B(n11400), .Z(n11405) );
  NAND U13626 ( .A(n11403), .B(n11402), .Z(n11404) );
  AND U13627 ( .A(n11405), .B(n11404), .Z(n11722) );
  NAND U13628 ( .A(n11407), .B(n11406), .Z(n11411) );
  NAND U13629 ( .A(n11409), .B(n11408), .Z(n11410) );
  NAND U13630 ( .A(n11411), .B(n11410), .Z(n11720) );
  AND U13631 ( .A(oglobal[4]), .B(n11412), .Z(n11773) );
  XOR U13632 ( .A(n11773), .B(oglobal[5]), .Z(n11762) );
  NANDN U13633 ( .A(n11414), .B(n11413), .Z(n11418) );
  NANDN U13634 ( .A(n11416), .B(n11415), .Z(n11417) );
  AND U13635 ( .A(n11418), .B(n11417), .Z(n11761) );
  XNOR U13636 ( .A(n11762), .B(n11761), .Z(n11764) );
  NANDN U13637 ( .A(n11420), .B(n11419), .Z(n11424) );
  OR U13638 ( .A(n11422), .B(n11421), .Z(n11423) );
  AND U13639 ( .A(n11424), .B(n11423), .Z(n11763) );
  XOR U13640 ( .A(n11764), .B(n11763), .Z(n11782) );
  NANDN U13641 ( .A(n11426), .B(n11425), .Z(n11430) );
  OR U13642 ( .A(n11428), .B(n11427), .Z(n11429) );
  AND U13643 ( .A(n11430), .B(n11429), .Z(n11767) );
  NANDN U13644 ( .A(n11432), .B(n11431), .Z(n11436) );
  OR U13645 ( .A(n11434), .B(n11433), .Z(n11435) );
  NAND U13646 ( .A(n11436), .B(n11435), .Z(n11768) );
  XNOR U13647 ( .A(n11767), .B(n11768), .Z(n11770) );
  NANDN U13648 ( .A(n11438), .B(n11437), .Z(n11442) );
  OR U13649 ( .A(n11440), .B(n11439), .Z(n11441) );
  AND U13650 ( .A(n11442), .B(n11441), .Z(n11769) );
  XOR U13651 ( .A(n11770), .B(n11769), .Z(n11781) );
  NANDN U13652 ( .A(n11444), .B(n11443), .Z(n11448) );
  OR U13653 ( .A(n11446), .B(n11445), .Z(n11447) );
  AND U13654 ( .A(n11448), .B(n11447), .Z(n11780) );
  XOR U13655 ( .A(n11781), .B(n11780), .Z(n11783) );
  XOR U13656 ( .A(n11782), .B(n11783), .Z(n11740) );
  NANDN U13657 ( .A(n11450), .B(n11449), .Z(n11454) );
  NANDN U13658 ( .A(n11452), .B(n11451), .Z(n11453) );
  AND U13659 ( .A(n11454), .B(n11453), .Z(n11737) );
  NANDN U13660 ( .A(n11456), .B(n11455), .Z(n11460) );
  OR U13661 ( .A(n11458), .B(n11457), .Z(n11459) );
  NAND U13662 ( .A(n11460), .B(n11459), .Z(n11738) );
  XNOR U13663 ( .A(n11737), .B(n11738), .Z(n11739) );
  XNOR U13664 ( .A(n11740), .B(n11739), .Z(n11719) );
  XOR U13665 ( .A(n11720), .B(n11719), .Z(n11721) );
  XNOR U13666 ( .A(n11722), .B(n11721), .Z(n11674) );
  XOR U13667 ( .A(n11677), .B(n11674), .Z(n11461) );
  XOR U13668 ( .A(n11673), .B(n11461), .Z(n11830) );
  NANDN U13669 ( .A(n11463), .B(n11462), .Z(n11467) );
  NANDN U13670 ( .A(n11465), .B(n11464), .Z(n11466) );
  AND U13671 ( .A(n11467), .B(n11466), .Z(n11824) );
  NANDN U13672 ( .A(n11469), .B(n11468), .Z(n11473) );
  NANDN U13673 ( .A(n11471), .B(n11470), .Z(n11472) );
  AND U13674 ( .A(n11473), .B(n11472), .Z(n11823) );
  NANDN U13675 ( .A(n11475), .B(n11474), .Z(n11479) );
  NANDN U13676 ( .A(n11477), .B(n11476), .Z(n11478) );
  AND U13677 ( .A(n11479), .B(n11478), .Z(n11777) );
  NANDN U13678 ( .A(n11481), .B(n11480), .Z(n11485) );
  NANDN U13679 ( .A(n11483), .B(n11482), .Z(n11484) );
  AND U13680 ( .A(n11485), .B(n11484), .Z(n11774) );
  NANDN U13681 ( .A(n11487), .B(n11486), .Z(n11491) );
  OR U13682 ( .A(n11489), .B(n11488), .Z(n11490) );
  NAND U13683 ( .A(n11491), .B(n11490), .Z(n11775) );
  XNOR U13684 ( .A(n11774), .B(n11775), .Z(n11776) );
  XOR U13685 ( .A(n11777), .B(n11776), .Z(n11799) );
  NANDN U13686 ( .A(n11493), .B(n11492), .Z(n11497) );
  NAND U13687 ( .A(n11495), .B(n11494), .Z(n11496) );
  NAND U13688 ( .A(n11497), .B(n11496), .Z(n11798) );
  XNOR U13689 ( .A(n11799), .B(n11798), .Z(n11800) );
  NANDN U13690 ( .A(n11499), .B(n11498), .Z(n11503) );
  NANDN U13691 ( .A(n11501), .B(n11500), .Z(n11502) );
  NAND U13692 ( .A(n11503), .B(n11502), .Z(n11801) );
  XNOR U13693 ( .A(n11800), .B(n11801), .Z(n11822) );
  XOR U13694 ( .A(n11823), .B(n11822), .Z(n11825) );
  XNOR U13695 ( .A(n11824), .B(n11825), .Z(n11670) );
  NANDN U13696 ( .A(n11505), .B(n11504), .Z(n11509) );
  OR U13697 ( .A(n11507), .B(n11506), .Z(n11508) );
  AND U13698 ( .A(n11509), .B(n11508), .Z(n11793) );
  NANDN U13699 ( .A(n11511), .B(n11510), .Z(n11515) );
  NAND U13700 ( .A(n11513), .B(n11512), .Z(n11514) );
  NAND U13701 ( .A(n11515), .B(n11514), .Z(n11792) );
  XOR U13702 ( .A(n11793), .B(n11792), .Z(n11795) );
  NANDN U13703 ( .A(n11517), .B(n11516), .Z(n11521) );
  OR U13704 ( .A(n11519), .B(n11518), .Z(n11520) );
  AND U13705 ( .A(n11521), .B(n11520), .Z(n11794) );
  XOR U13706 ( .A(n11795), .B(n11794), .Z(n11732) );
  NANDN U13707 ( .A(n11523), .B(n11522), .Z(n11527) );
  NANDN U13708 ( .A(n11525), .B(n11524), .Z(n11526) );
  AND U13709 ( .A(n11527), .B(n11526), .Z(n11731) );
  XNOR U13710 ( .A(n11732), .B(n11731), .Z(n11733) );
  NANDN U13711 ( .A(n11529), .B(n11528), .Z(n11533) );
  NANDN U13712 ( .A(n11531), .B(n11530), .Z(n11532) );
  NAND U13713 ( .A(n11533), .B(n11532), .Z(n11734) );
  XNOR U13714 ( .A(n11733), .B(n11734), .Z(n11819) );
  NANDN U13715 ( .A(n11535), .B(n11534), .Z(n11539) );
  NAND U13716 ( .A(n11537), .B(n11536), .Z(n11538) );
  AND U13717 ( .A(n11539), .B(n11538), .Z(n11728) );
  NANDN U13718 ( .A(n11541), .B(n11540), .Z(n11545) );
  NANDN U13719 ( .A(n11543), .B(n11542), .Z(n11544) );
  AND U13720 ( .A(n11545), .B(n11544), .Z(n11726) );
  NANDN U13721 ( .A(n11547), .B(n11546), .Z(n11551) );
  NANDN U13722 ( .A(n11549), .B(n11548), .Z(n11550) );
  NAND U13723 ( .A(n11551), .B(n11550), .Z(n11725) );
  XNOR U13724 ( .A(n11726), .B(n11725), .Z(n11727) );
  XOR U13725 ( .A(n11728), .B(n11727), .Z(n11817) );
  NANDN U13726 ( .A(n11553), .B(n11552), .Z(n11557) );
  NANDN U13727 ( .A(n11555), .B(n11554), .Z(n11556) );
  AND U13728 ( .A(n11557), .B(n11556), .Z(n11816) );
  XNOR U13729 ( .A(n11817), .B(n11816), .Z(n11818) );
  XNOR U13730 ( .A(n11819), .B(n11818), .Z(n11668) );
  NAND U13731 ( .A(n11559), .B(n11558), .Z(n11563) );
  NAND U13732 ( .A(n11561), .B(n11560), .Z(n11562) );
  NAND U13733 ( .A(n11563), .B(n11562), .Z(n11687) );
  NANDN U13734 ( .A(n11565), .B(n11564), .Z(n11569) );
  NANDN U13735 ( .A(n11567), .B(n11566), .Z(n11568) );
  AND U13736 ( .A(n11569), .B(n11568), .Z(n11788) );
  NANDN U13737 ( .A(n11571), .B(n11570), .Z(n11575) );
  OR U13738 ( .A(n11573), .B(n11572), .Z(n11574) );
  AND U13739 ( .A(n11575), .B(n11574), .Z(n11786) );
  NANDN U13740 ( .A(n11577), .B(n11576), .Z(n11581) );
  NAND U13741 ( .A(n11579), .B(n11578), .Z(n11580) );
  AND U13742 ( .A(n11581), .B(n11580), .Z(n11758) );
  NANDN U13743 ( .A(n11586), .B(n11585), .Z(n11590) );
  OR U13744 ( .A(n11588), .B(n11587), .Z(n11589) );
  NAND U13745 ( .A(n11590), .B(n11589), .Z(n11755) );
  XNOR U13746 ( .A(n11756), .B(n11755), .Z(n11757) );
  XOR U13747 ( .A(n11758), .B(n11757), .Z(n11787) );
  XOR U13748 ( .A(n11786), .B(n11787), .Z(n11789) );
  XOR U13749 ( .A(n11788), .B(n11789), .Z(n11811) );
  NANDN U13750 ( .A(n11592), .B(n11591), .Z(n11596) );
  NAND U13751 ( .A(n11594), .B(n11593), .Z(n11595) );
  NAND U13752 ( .A(n11596), .B(n11595), .Z(n11810) );
  XNOR U13753 ( .A(n11811), .B(n11810), .Z(n11812) );
  NANDN U13754 ( .A(n11598), .B(n11597), .Z(n11602) );
  NANDN U13755 ( .A(n11600), .B(n11599), .Z(n11601) );
  AND U13756 ( .A(n11602), .B(n11601), .Z(n11743) );
  NANDN U13757 ( .A(n11604), .B(n11603), .Z(n11608) );
  NANDN U13758 ( .A(n11606), .B(n11605), .Z(n11607) );
  AND U13759 ( .A(n11608), .B(n11607), .Z(n11751) );
  XNOR U13760 ( .A(n11750), .B(n11749), .Z(n11752) );
  XOR U13761 ( .A(n11751), .B(n11752), .Z(n11744) );
  XNOR U13762 ( .A(n11743), .B(n11744), .Z(n11745) );
  NANDN U13763 ( .A(n11616), .B(n11615), .Z(n11620) );
  NAND U13764 ( .A(n11618), .B(n11617), .Z(n11619) );
  NAND U13765 ( .A(n11620), .B(n11619), .Z(n11746) );
  XOR U13766 ( .A(n11745), .B(n11746), .Z(n11813) );
  XNOR U13767 ( .A(n11812), .B(n11813), .Z(n11686) );
  XOR U13768 ( .A(n11687), .B(n11686), .Z(n11689) );
  NANDN U13769 ( .A(n11622), .B(n11621), .Z(n11626) );
  NANDN U13770 ( .A(n11624), .B(n11623), .Z(n11625) );
  AND U13771 ( .A(n11626), .B(n11625), .Z(n11806) );
  NANDN U13772 ( .A(n11628), .B(n11627), .Z(n11632) );
  NANDN U13773 ( .A(n11630), .B(n11629), .Z(n11631) );
  AND U13774 ( .A(n11632), .B(n11631), .Z(n11804) );
  NANDN U13775 ( .A(n11634), .B(n11633), .Z(n11638) );
  OR U13776 ( .A(n11636), .B(n11635), .Z(n11637) );
  NAND U13777 ( .A(n11638), .B(n11637), .Z(n11805) );
  XOR U13778 ( .A(n11804), .B(n11805), .Z(n11807) );
  XNOR U13779 ( .A(n11806), .B(n11807), .Z(n11688) );
  XNOR U13780 ( .A(n11689), .B(n11688), .Z(n11667) );
  XOR U13781 ( .A(n11668), .B(n11667), .Z(n11669) );
  XOR U13782 ( .A(n11670), .B(n11669), .Z(n11828) );
  NANDN U13783 ( .A(n11640), .B(n11639), .Z(n11644) );
  NANDN U13784 ( .A(n11642), .B(n11641), .Z(n11643) );
  NAND U13785 ( .A(n11644), .B(n11643), .Z(n11829) );
  XOR U13786 ( .A(n11830), .B(n11831), .Z(n11699) );
  XNOR U13787 ( .A(n11700), .B(n11701), .Z(n11705) );
  XNOR U13788 ( .A(n11705), .B(n11704), .Z(n11648) );
  XNOR U13789 ( .A(n11706), .B(n11648), .Z(o[5]) );
  NANDN U13790 ( .A(n11650), .B(n11649), .Z(n11654) );
  NAND U13791 ( .A(n11652), .B(n11651), .Z(n11653) );
  NAND U13792 ( .A(n11654), .B(n11653), .Z(n11922) );
  NANDN U13793 ( .A(n11656), .B(n11655), .Z(n11660) );
  NAND U13794 ( .A(n11658), .B(n11657), .Z(n11659) );
  AND U13795 ( .A(n11660), .B(n11659), .Z(n11844) );
  NANDN U13796 ( .A(n11662), .B(n11661), .Z(n11666) );
  NANDN U13797 ( .A(n11664), .B(n11663), .Z(n11665) );
  AND U13798 ( .A(n11666), .B(n11665), .Z(n11842) );
  NAND U13799 ( .A(n11668), .B(n11667), .Z(n11672) );
  NAND U13800 ( .A(n11670), .B(n11669), .Z(n11671) );
  AND U13801 ( .A(n11672), .B(n11671), .Z(n11903) );
  NANDN U13802 ( .A(n11673), .B(n11674), .Z(n11679) );
  NOR U13803 ( .A(n11675), .B(n11674), .Z(n11676) );
  OR U13804 ( .A(n11677), .B(n11676), .Z(n11678) );
  AND U13805 ( .A(n11679), .B(n11678), .Z(n11901) );
  NAND U13806 ( .A(n11681), .B(n11680), .Z(n11685) );
  NANDN U13807 ( .A(n11683), .B(n11682), .Z(n11684) );
  AND U13808 ( .A(n11685), .B(n11684), .Z(n11908) );
  NAND U13809 ( .A(n11687), .B(n11686), .Z(n11691) );
  NAND U13810 ( .A(n11689), .B(n11688), .Z(n11690) );
  NAND U13811 ( .A(n11691), .B(n11690), .Z(n11906) );
  NAND U13812 ( .A(n11693), .B(n11692), .Z(n11697) );
  NAND U13813 ( .A(n11695), .B(n11694), .Z(n11696) );
  AND U13814 ( .A(n11697), .B(n11696), .Z(n11907) );
  XNOR U13815 ( .A(n11906), .B(n11907), .Z(n11909) );
  XOR U13816 ( .A(n11901), .B(n11900), .Z(n11902) );
  XOR U13817 ( .A(n11903), .B(n11902), .Z(n11841) );
  XOR U13818 ( .A(n11844), .B(n11843), .Z(n11921) );
  XOR U13819 ( .A(n11922), .B(n11921), .Z(n11924) );
  NANDN U13820 ( .A(n11699), .B(n11698), .Z(n11703) );
  NANDN U13821 ( .A(n11701), .B(n11700), .Z(n11702) );
  AND U13822 ( .A(n11703), .B(n11702), .Z(n11923) );
  XNOR U13823 ( .A(n11924), .B(n11923), .Z(n11920) );
  NAND U13824 ( .A(n11708), .B(n11707), .Z(n11712) );
  NANDN U13825 ( .A(n11710), .B(n11709), .Z(n11711) );
  AND U13826 ( .A(n11712), .B(n11711), .Z(n11838) );
  NAND U13827 ( .A(n11714), .B(n11713), .Z(n11718) );
  NANDN U13828 ( .A(n11716), .B(n11715), .Z(n11717) );
  AND U13829 ( .A(n11718), .B(n11717), .Z(n11897) );
  NAND U13830 ( .A(n11720), .B(n11719), .Z(n11724) );
  NAND U13831 ( .A(n11722), .B(n11721), .Z(n11723) );
  NAND U13832 ( .A(n11724), .B(n11723), .Z(n11913) );
  NANDN U13833 ( .A(n11726), .B(n11725), .Z(n11730) );
  NAND U13834 ( .A(n11728), .B(n11727), .Z(n11729) );
  AND U13835 ( .A(n11730), .B(n11729), .Z(n11867) );
  NANDN U13836 ( .A(n11732), .B(n11731), .Z(n11736) );
  NANDN U13837 ( .A(n11734), .B(n11733), .Z(n11735) );
  AND U13838 ( .A(n11736), .B(n11735), .Z(n11865) );
  NANDN U13839 ( .A(n11738), .B(n11737), .Z(n11742) );
  NANDN U13840 ( .A(n11740), .B(n11739), .Z(n11741) );
  NAND U13841 ( .A(n11742), .B(n11741), .Z(n11866) );
  XOR U13842 ( .A(n11865), .B(n11866), .Z(n11868) );
  XNOR U13843 ( .A(n11867), .B(n11868), .Z(n11912) );
  XOR U13844 ( .A(n11913), .B(n11912), .Z(n11915) );
  NANDN U13845 ( .A(n11744), .B(n11743), .Z(n11748) );
  NANDN U13846 ( .A(n11746), .B(n11745), .Z(n11747) );
  AND U13847 ( .A(n11748), .B(n11747), .Z(n11880) );
  NAND U13848 ( .A(n11750), .B(n11749), .Z(n11754) );
  NANDN U13849 ( .A(n11752), .B(n11751), .Z(n11753) );
  AND U13850 ( .A(n11754), .B(n11753), .Z(n11878) );
  NANDN U13851 ( .A(n11756), .B(n11755), .Z(n11760) );
  NANDN U13852 ( .A(n11758), .B(n11757), .Z(n11759) );
  NAND U13853 ( .A(n11760), .B(n11759), .Z(n11888) );
  NANDN U13854 ( .A(n11762), .B(n11761), .Z(n11766) );
  NAND U13855 ( .A(n11764), .B(n11763), .Z(n11765) );
  AND U13856 ( .A(n11766), .B(n11765), .Z(n11889) );
  XOR U13857 ( .A(n11888), .B(n11889), .Z(n11891) );
  NANDN U13858 ( .A(n11768), .B(n11767), .Z(n11772) );
  NAND U13859 ( .A(n11770), .B(n11769), .Z(n11771) );
  AND U13860 ( .A(n11772), .B(n11771), .Z(n11885) );
  AND U13861 ( .A(n11773), .B(oglobal[5]), .Z(n11883) );
  XOR U13862 ( .A(n11883), .B(oglobal[6]), .Z(n11884) );
  XOR U13863 ( .A(n11885), .B(n11884), .Z(n11890) );
  XNOR U13864 ( .A(n11891), .B(n11890), .Z(n11877) );
  XNOR U13865 ( .A(n11878), .B(n11877), .Z(n11879) );
  XNOR U13866 ( .A(n11880), .B(n11879), .Z(n11855) );
  NANDN U13867 ( .A(n11775), .B(n11774), .Z(n11779) );
  NAND U13868 ( .A(n11777), .B(n11776), .Z(n11778) );
  AND U13869 ( .A(n11779), .B(n11778), .Z(n11873) );
  NANDN U13870 ( .A(n11781), .B(n11780), .Z(n11785) );
  OR U13871 ( .A(n11783), .B(n11782), .Z(n11784) );
  AND U13872 ( .A(n11785), .B(n11784), .Z(n11871) );
  NANDN U13873 ( .A(n11787), .B(n11786), .Z(n11791) );
  OR U13874 ( .A(n11789), .B(n11788), .Z(n11790) );
  NAND U13875 ( .A(n11791), .B(n11790), .Z(n11872) );
  XOR U13876 ( .A(n11871), .B(n11872), .Z(n11874) );
  XNOR U13877 ( .A(n11873), .B(n11874), .Z(n11853) );
  NAND U13878 ( .A(n11793), .B(n11792), .Z(n11797) );
  NAND U13879 ( .A(n11795), .B(n11794), .Z(n11796) );
  NAND U13880 ( .A(n11797), .B(n11796), .Z(n11854) );
  XOR U13881 ( .A(n11853), .B(n11854), .Z(n11856) );
  XNOR U13882 ( .A(n11855), .B(n11856), .Z(n11914) );
  XNOR U13883 ( .A(n11915), .B(n11914), .Z(n11895) );
  NANDN U13884 ( .A(n11799), .B(n11798), .Z(n11803) );
  NANDN U13885 ( .A(n11801), .B(n11800), .Z(n11802) );
  AND U13886 ( .A(n11803), .B(n11802), .Z(n11861) );
  NANDN U13887 ( .A(n11805), .B(n11804), .Z(n11809) );
  NANDN U13888 ( .A(n11807), .B(n11806), .Z(n11808) );
  AND U13889 ( .A(n11809), .B(n11808), .Z(n11860) );
  NANDN U13890 ( .A(n11811), .B(n11810), .Z(n11815) );
  NANDN U13891 ( .A(n11813), .B(n11812), .Z(n11814) );
  NAND U13892 ( .A(n11815), .B(n11814), .Z(n11859) );
  XOR U13893 ( .A(n11860), .B(n11859), .Z(n11862) );
  XOR U13894 ( .A(n11861), .B(n11862), .Z(n11848) );
  NANDN U13895 ( .A(n11817), .B(n11816), .Z(n11821) );
  NAND U13896 ( .A(n11819), .B(n11818), .Z(n11820) );
  AND U13897 ( .A(n11821), .B(n11820), .Z(n11847) );
  XNOR U13898 ( .A(n11848), .B(n11847), .Z(n11849) );
  NANDN U13899 ( .A(n11823), .B(n11822), .Z(n11827) );
  OR U13900 ( .A(n11825), .B(n11824), .Z(n11826) );
  NAND U13901 ( .A(n11827), .B(n11826), .Z(n11850) );
  XNOR U13902 ( .A(n11849), .B(n11850), .Z(n11894) );
  XOR U13903 ( .A(n11895), .B(n11894), .Z(n11896) );
  XOR U13904 ( .A(n11897), .B(n11896), .Z(n11836) );
  NANDN U13905 ( .A(n11829), .B(n11828), .Z(n11833) );
  NAND U13906 ( .A(n11831), .B(n11830), .Z(n11832) );
  AND U13907 ( .A(n11833), .B(n11832), .Z(n11835) );
  XOR U13908 ( .A(n11838), .B(n11837), .Z(n11918) );
  XOR U13909 ( .A(n11919), .B(n11918), .Z(n11834) );
  XNOR U13910 ( .A(n11920), .B(n11834), .Z(o[6]) );
  NANDN U13911 ( .A(n11836), .B(n11835), .Z(n11840) );
  NAND U13912 ( .A(n11838), .B(n11837), .Z(n11839) );
  NAND U13913 ( .A(n11840), .B(n11839), .Z(n11930) );
  NANDN U13914 ( .A(n11842), .B(n11841), .Z(n11846) );
  NANDN U13915 ( .A(n11844), .B(n11843), .Z(n11845) );
  NAND U13916 ( .A(n11846), .B(n11845), .Z(n11928) );
  NANDN U13917 ( .A(n11848), .B(n11847), .Z(n11852) );
  NANDN U13918 ( .A(n11850), .B(n11849), .Z(n11851) );
  AND U13919 ( .A(n11852), .B(n11851), .Z(n11945) );
  NANDN U13920 ( .A(n11854), .B(n11853), .Z(n11858) );
  NANDN U13921 ( .A(n11856), .B(n11855), .Z(n11857) );
  AND U13922 ( .A(n11858), .B(n11857), .Z(n11943) );
  NANDN U13923 ( .A(n11860), .B(n11859), .Z(n11864) );
  OR U13924 ( .A(n11862), .B(n11861), .Z(n11863) );
  AND U13925 ( .A(n11864), .B(n11863), .Z(n11951) );
  NANDN U13926 ( .A(n11866), .B(n11865), .Z(n11870) );
  OR U13927 ( .A(n11868), .B(n11867), .Z(n11869) );
  AND U13928 ( .A(n11870), .B(n11869), .Z(n11950) );
  NANDN U13929 ( .A(n11872), .B(n11871), .Z(n11876) );
  NANDN U13930 ( .A(n11874), .B(n11873), .Z(n11875) );
  AND U13931 ( .A(n11876), .B(n11875), .Z(n11963) );
  NANDN U13932 ( .A(n11878), .B(n11877), .Z(n11882) );
  NANDN U13933 ( .A(n11880), .B(n11879), .Z(n11881) );
  AND U13934 ( .A(n11882), .B(n11881), .Z(n11961) );
  NAND U13935 ( .A(n11883), .B(oglobal[6]), .Z(n11887) );
  NAND U13936 ( .A(n11885), .B(n11884), .Z(n11886) );
  NAND U13937 ( .A(n11887), .B(n11886), .Z(n11955) );
  XOR U13938 ( .A(n11955), .B(oglobal[7]), .Z(n11957) );
  NAND U13939 ( .A(n11889), .B(n11888), .Z(n11893) );
  NAND U13940 ( .A(n11891), .B(n11890), .Z(n11892) );
  NAND U13941 ( .A(n11893), .B(n11892), .Z(n11956) );
  XOR U13942 ( .A(n11957), .B(n11956), .Z(n11960) );
  XOR U13943 ( .A(n11961), .B(n11960), .Z(n11962) );
  XOR U13944 ( .A(n11963), .B(n11962), .Z(n11949) );
  XOR U13945 ( .A(n11950), .B(n11949), .Z(n11952) );
  XOR U13946 ( .A(n11951), .B(n11952), .Z(n11944) );
  XOR U13947 ( .A(n11943), .B(n11944), .Z(n11946) );
  XNOR U13948 ( .A(n11945), .B(n11946), .Z(n11938) );
  NAND U13949 ( .A(n11895), .B(n11894), .Z(n11899) );
  NAND U13950 ( .A(n11897), .B(n11896), .Z(n11898) );
  AND U13951 ( .A(n11899), .B(n11898), .Z(n11937) );
  XOR U13952 ( .A(n11938), .B(n11937), .Z(n11940) );
  NAND U13953 ( .A(n11901), .B(n11900), .Z(n11905) );
  NAND U13954 ( .A(n11903), .B(n11902), .Z(n11904) );
  NAND U13955 ( .A(n11905), .B(n11904), .Z(n11966) );
  NAND U13956 ( .A(n11907), .B(n11906), .Z(n11911) );
  NANDN U13957 ( .A(n11909), .B(n11908), .Z(n11910) );
  NAND U13958 ( .A(n11911), .B(n11910), .Z(n11965) );
  NAND U13959 ( .A(n11913), .B(n11912), .Z(n11917) );
  NAND U13960 ( .A(n11915), .B(n11914), .Z(n11916) );
  NAND U13961 ( .A(n11917), .B(n11916), .Z(n11964) );
  XOR U13962 ( .A(n11965), .B(n11964), .Z(n11967) );
  XOR U13963 ( .A(n11966), .B(n11967), .Z(n11939) );
  XOR U13964 ( .A(n11940), .B(n11939), .Z(n11929) );
  XOR U13965 ( .A(n11928), .B(n11929), .Z(n11931) );
  XOR U13966 ( .A(n11930), .B(n11931), .Z(n11934) );
  NAND U13967 ( .A(n11922), .B(n11921), .Z(n11926) );
  NAND U13968 ( .A(n11924), .B(n11923), .Z(n11925) );
  AND U13969 ( .A(n11926), .B(n11925), .Z(n11936) );
  XNOR U13970 ( .A(n11935), .B(n11936), .Z(n11927) );
  XOR U13971 ( .A(n11934), .B(n11927), .Z(o[7]) );
  NAND U13972 ( .A(n11929), .B(n11928), .Z(n11933) );
  NAND U13973 ( .A(n11931), .B(n11930), .Z(n11932) );
  AND U13974 ( .A(n11933), .B(n11932), .Z(n11991) );
  NAND U13975 ( .A(n11938), .B(n11937), .Z(n11942) );
  NAND U13976 ( .A(n11940), .B(n11939), .Z(n11941) );
  NAND U13977 ( .A(n11942), .B(n11941), .Z(n11973) );
  NANDN U13978 ( .A(n11944), .B(n11943), .Z(n11948) );
  OR U13979 ( .A(n11946), .B(n11945), .Z(n11947) );
  AND U13980 ( .A(n11948), .B(n11947), .Z(n11980) );
  NANDN U13981 ( .A(n11950), .B(n11949), .Z(n11954) );
  NANDN U13982 ( .A(n11952), .B(n11951), .Z(n11953) );
  AND U13983 ( .A(n11954), .B(n11953), .Z(n11978) );
  NAND U13984 ( .A(oglobal[7]), .B(n11955), .Z(n11959) );
  NAND U13985 ( .A(n11957), .B(n11956), .Z(n11958) );
  AND U13986 ( .A(n11959), .B(n11958), .Z(n11985) );
  XNOR U13987 ( .A(n11983), .B(oglobal[8]), .Z(n11984) );
  XNOR U13988 ( .A(n11985), .B(n11984), .Z(n11977) );
  XNOR U13989 ( .A(n11978), .B(n11977), .Z(n11979) );
  XOR U13990 ( .A(n11980), .B(n11979), .Z(n11972) );
  NAND U13991 ( .A(n11965), .B(n11964), .Z(n11969) );
  NAND U13992 ( .A(n11967), .B(n11966), .Z(n11968) );
  NAND U13993 ( .A(n11969), .B(n11968), .Z(n11971) );
  XNOR U13994 ( .A(n11972), .B(n11971), .Z(n11974) );
  IV U13995 ( .A(n11990), .Z(n11988) );
  XOR U13996 ( .A(n11989), .B(n11988), .Z(n11970) );
  XNOR U13997 ( .A(n11991), .B(n11970), .Z(o[8]) );
  NAND U13998 ( .A(n11972), .B(n11971), .Z(n11976) );
  NANDN U13999 ( .A(n11974), .B(n11973), .Z(n11975) );
  AND U14000 ( .A(n11976), .B(n11975), .Z(n11998) );
  NANDN U14001 ( .A(n11978), .B(n11977), .Z(n11982) );
  NANDN U14002 ( .A(n11980), .B(n11979), .Z(n11981) );
  AND U14003 ( .A(n11982), .B(n11981), .Z(n12001) );
  NANDN U14004 ( .A(n11983), .B(oglobal[8]), .Z(n11987) );
  NANDN U14005 ( .A(n11985), .B(n11984), .Z(n11986) );
  AND U14006 ( .A(n11987), .B(n11986), .Z(n11999) );
  XNOR U14007 ( .A(n11999), .B(oglobal[9]), .Z(n12000) );
  XOR U14008 ( .A(n12001), .B(n12000), .Z(n11996) );
  NANDN U14009 ( .A(n11988), .B(n11989), .Z(n11994) );
  NOR U14010 ( .A(n11990), .B(n11989), .Z(n11992) );
  OR U14011 ( .A(n11992), .B(n11991), .Z(n11993) );
  AND U14012 ( .A(n11994), .B(n11993), .Z(n11997) );
  XOR U14013 ( .A(n11996), .B(n11997), .Z(n11995) );
  XNOR U14014 ( .A(n11998), .B(n11995), .Z(o[9]) );
  NANDN U14015 ( .A(n11999), .B(oglobal[9]), .Z(n12003) );
  NANDN U14016 ( .A(n12001), .B(n12000), .Z(n12002) );
  AND U14017 ( .A(n12003), .B(n12002), .Z(n12004) );
  XNOR U14018 ( .A(n12004), .B(oglobal[10]), .Z(n12005) );
  XOR U14019 ( .A(n12006), .B(n12005), .Z(o[10]) );
  NANDN U14020 ( .A(n12004), .B(oglobal[10]), .Z(n12008) );
  NAND U14021 ( .A(n12006), .B(n12005), .Z(n12007) );
  NAND U14022 ( .A(n12008), .B(n12007), .Z(n12009) );
  XOR U14023 ( .A(oglobal[11]), .B(n12009), .Z(o[11]) );
  NAND U14024 ( .A(oglobal[11]), .B(n12009), .Z(n12010) );
  XNOR U14025 ( .A(oglobal[12]), .B(n12010), .Z(o[12]) );
  NANDN U14026 ( .A(n12010), .B(oglobal[12]), .Z(n12011) );
  XNOR U14027 ( .A(oglobal[13]), .B(n12011), .Z(o[13]) );
endmodule

