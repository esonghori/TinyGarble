
module mult_N128_CC8 ( clk, rst, a, b, c );
  input [127:0] a;
  input [15:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032;
  wire   [255:0] sreg;

  DFF \sreg_reg[239]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[238]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[237]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[236]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[235]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[234]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[233]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[232]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[231]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[230]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[229]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[228]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[227]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[226]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[225]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[224]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[223]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[222]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[221]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[220]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[219]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[218]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[217]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[216]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[215]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[214]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[213]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[212]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[211]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[210]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[209]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[208]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[207]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[206]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[205]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[204]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[203]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[202]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[201]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[200]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[199]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[198]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[197]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[196]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[195]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[194]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[193]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[192]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[191]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U19 ( .A(n9600), .B(n9599), .Z(n1) );
  NANDN U20 ( .A(n9598), .B(n9597), .Z(n2) );
  NAND U21 ( .A(n1), .B(n2), .Z(n9618) );
  NAND U22 ( .A(n9985), .B(n9986), .Z(n3) );
  NAND U23 ( .A(n9984), .B(n10000), .Z(n4) );
  NAND U24 ( .A(n3), .B(n4), .Z(n10013) );
  NAND U25 ( .A(sreg[126]), .B(n637), .Z(n5) );
  XOR U26 ( .A(sreg[126]), .B(n637), .Z(n6) );
  NANDN U27 ( .A(n636), .B(n6), .Z(n7) );
  NAND U28 ( .A(n5), .B(n7), .Z(n708) );
  NAND U29 ( .A(n9575), .B(n9574), .Z(n8) );
  NANDN U30 ( .A(n9573), .B(n9572), .Z(n9) );
  NAND U31 ( .A(n8), .B(n9), .Z(n9622) );
  NAND U32 ( .A(n9616), .B(n9615), .Z(n10) );
  NAND U33 ( .A(n9614), .B(n9613), .Z(n11) );
  AND U34 ( .A(n10), .B(n11), .Z(n9664) );
  NAND U35 ( .A(n93), .B(n94), .Z(n12) );
  XOR U36 ( .A(n93), .B(n94), .Z(n13) );
  NANDN U37 ( .A(n92), .B(n13), .Z(n14) );
  NAND U38 ( .A(n12), .B(n14), .Z(n106) );
  NAND U39 ( .A(sreg[127]), .B(n708), .Z(n15) );
  XOR U40 ( .A(sreg[127]), .B(n708), .Z(n16) );
  NANDN U41 ( .A(n707), .B(n16), .Z(n17) );
  NAND U42 ( .A(n15), .B(n17), .Z(n710) );
  NAND U43 ( .A(n10017), .B(n10018), .Z(n18) );
  NANDN U44 ( .A(n10020), .B(n10019), .Z(n19) );
  NAND U45 ( .A(n18), .B(n19), .Z(n10032) );
  NANDN U46 ( .A(b[0]), .B(a[127]), .Z(n20) );
  NAND U47 ( .A(b[1]), .B(n20), .Z(n9362) );
  NAND U48 ( .A(n629), .B(n628), .Z(n21) );
  NANDN U49 ( .A(n627), .B(n626), .Z(n22) );
  NAND U50 ( .A(n21), .B(n22), .Z(n645) );
  NAND U51 ( .A(n9618), .B(n9617), .Z(n23) );
  NANDN U52 ( .A(n9620), .B(n9619), .Z(n24) );
  AND U53 ( .A(n23), .B(n24), .Z(n9671) );
  XOR U54 ( .A(n9739), .B(n9740), .Z(n25) );
  NAND U55 ( .A(n25), .B(n9738), .Z(n26) );
  NAND U56 ( .A(n9739), .B(n9740), .Z(n27) );
  AND U57 ( .A(n26), .B(n27), .Z(n9784) );
  NAND U58 ( .A(n9966), .B(n9967), .Z(n28) );
  NANDN U59 ( .A(n9965), .B(n9964), .Z(n29) );
  AND U60 ( .A(n28), .B(n29), .Z(n9993) );
  NAND U61 ( .A(sreg[115]), .B(n91), .Z(n30) );
  XOR U62 ( .A(sreg[115]), .B(n91), .Z(n31) );
  NANDN U63 ( .A(n90), .B(n31), .Z(n32) );
  NAND U64 ( .A(n30), .B(n32), .Z(n127) );
  NAND U65 ( .A(n9610), .B(n9609), .Z(n33) );
  NANDN U66 ( .A(n9612), .B(n9611), .Z(n34) );
  AND U67 ( .A(n33), .B(n34), .Z(n9665) );
  XOR U68 ( .A(n443), .B(sreg[124]), .Z(n35) );
  NANDN U69 ( .A(n444), .B(n35), .Z(n36) );
  NAND U70 ( .A(n443), .B(sreg[124]), .Z(n37) );
  AND U71 ( .A(n36), .B(n37), .Z(n566) );
  XOR U72 ( .A(sreg[128]), .B(n710), .Z(n38) );
  NANDN U73 ( .A(n711), .B(n38), .Z(n39) );
  NAND U74 ( .A(sreg[128]), .B(n710), .Z(n40) );
  AND U75 ( .A(n39), .B(n40), .Z(n858) );
  NAND U76 ( .A(sreg[131]), .B(n940), .Z(n41) );
  XOR U77 ( .A(sreg[131]), .B(n940), .Z(n42) );
  NANDN U78 ( .A(n939), .B(n42), .Z(n43) );
  NAND U79 ( .A(n41), .B(n43), .Z(n1087) );
  XNOR U80 ( .A(a[127]), .B(a[126]), .Z(n44) );
  XNOR U81 ( .A(n10023), .B(n44), .Z(n45) );
  AND U82 ( .A(n45), .B(b[15]), .Z(n46) );
  NANDN U83 ( .A(n10026), .B(n10027), .Z(n47) );
  NANDN U84 ( .A(n10024), .B(n10025), .Z(n48) );
  AND U85 ( .A(n47), .B(n48), .Z(n49) );
  NOR U86 ( .A(n10032), .B(n10031), .Z(n50) );
  NANDN U87 ( .A(n10028), .B(n10031), .Z(n51) );
  OR U88 ( .A(n50), .B(n10029), .Z(n52) );
  NAND U89 ( .A(n51), .B(n52), .Z(n53) );
  OR U90 ( .A(n10029), .B(n51), .Z(n54) );
  NANDN U91 ( .A(n10030), .B(n54), .Z(n55) );
  NAND U92 ( .A(n53), .B(n55), .Z(n56) );
  XNOR U93 ( .A(n46), .B(n49), .Z(n57) );
  XNOR U94 ( .A(n56), .B(n57), .Z(c[255]) );
  AND U95 ( .A(b[0]), .B(a[0]), .Z(n59) );
  XOR U96 ( .A(n59), .B(sreg[112]), .Z(c[112]) );
  AND U97 ( .A(b[0]), .B(a[1]), .Z(n66) );
  NAND U98 ( .A(a[0]), .B(b[1]), .Z(n58) );
  XOR U99 ( .A(n66), .B(n58), .Z(n60) );
  XNOR U100 ( .A(sreg[113]), .B(n60), .Z(n62) );
  AND U101 ( .A(n59), .B(sreg[112]), .Z(n61) );
  XOR U102 ( .A(n62), .B(n61), .Z(c[113]) );
  NANDN U103 ( .A(n60), .B(sreg[113]), .Z(n64) );
  NAND U104 ( .A(n62), .B(n61), .Z(n63) );
  AND U105 ( .A(n64), .B(n63), .Z(n72) );
  XNOR U106 ( .A(n72), .B(sreg[114]), .Z(n74) );
  NAND U107 ( .A(a[0]), .B(b[2]), .Z(n65) );
  XNOR U108 ( .A(b[1]), .B(n65), .Z(n68) );
  NANDN U109 ( .A(a[0]), .B(n66), .Z(n67) );
  NAND U110 ( .A(n68), .B(n67), .Z(n78) );
  NAND U111 ( .A(b[0]), .B(a[2]), .Z(n69) );
  XNOR U112 ( .A(b[1]), .B(n69), .Z(n71) );
  NANDN U113 ( .A(b[0]), .B(a[1]), .Z(n70) );
  NAND U114 ( .A(n71), .B(n70), .Z(n77) );
  XOR U115 ( .A(n78), .B(n77), .Z(n73) );
  XOR U116 ( .A(n74), .B(n73), .Z(c[114]) );
  NANDN U117 ( .A(n72), .B(sreg[114]), .Z(n76) );
  NAND U118 ( .A(n74), .B(n73), .Z(n75) );
  NAND U119 ( .A(n76), .B(n75), .Z(n91) );
  NOR U120 ( .A(n78), .B(n77), .Z(n94) );
  NAND U121 ( .A(b[1]), .B(b[2]), .Z(n79) );
  AND U122 ( .A(b[3]), .B(n79), .Z(n9567) );
  XOR U123 ( .A(b[1]), .B(b[2]), .Z(n9421) );
  IV U124 ( .A(n9421), .Z(n9375) );
  NANDN U125 ( .A(n9375), .B(a[0]), .Z(n80) );
  AND U126 ( .A(n9567), .B(n80), .Z(n93) );
  NAND U127 ( .A(b[0]), .B(a[3]), .Z(n81) );
  XNOR U128 ( .A(b[1]), .B(n81), .Z(n83) );
  NANDN U129 ( .A(b[0]), .B(a[2]), .Z(n82) );
  NAND U130 ( .A(n83), .B(n82), .Z(n103) );
  XOR U131 ( .A(b[3]), .B(b[2]), .Z(n95) );
  XOR U132 ( .A(b[3]), .B(a[0]), .Z(n84) );
  NAND U133 ( .A(n95), .B(n84), .Z(n85) );
  OR U134 ( .A(n85), .B(n9421), .Z(n87) );
  XOR U135 ( .A(b[3]), .B(a[1]), .Z(n96) );
  NAND U136 ( .A(n9421), .B(n96), .Z(n86) );
  NAND U137 ( .A(n87), .B(n86), .Z(n102) );
  XOR U138 ( .A(n103), .B(n102), .Z(n92) );
  XOR U139 ( .A(n93), .B(n92), .Z(n88) );
  XOR U140 ( .A(n94), .B(n88), .Z(n90) );
  XOR U141 ( .A(sreg[115]), .B(n90), .Z(n89) );
  XNOR U142 ( .A(n91), .B(n89), .Z(c[115]) );
  XOR U143 ( .A(n127), .B(sreg[116]), .Z(n129) );
  ANDN U144 ( .B(n95), .A(n9421), .Z(n9420) );
  IV U145 ( .A(n9420), .Z(n9374) );
  NANDN U146 ( .A(n9374), .B(n96), .Z(n98) );
  XOR U147 ( .A(b[3]), .B(a[2]), .Z(n110) );
  NANDN U148 ( .A(n9375), .B(n110), .Z(n97) );
  AND U149 ( .A(n98), .B(n97), .Z(n124) );
  XOR U150 ( .A(b[4]), .B(b[3]), .Z(n9581) );
  IV U151 ( .A(n9581), .Z(n9503) );
  ANDN U152 ( .B(a[0]), .A(n9503), .Z(n121) );
  NAND U153 ( .A(b[0]), .B(a[4]), .Z(n99) );
  XNOR U154 ( .A(b[1]), .B(n99), .Z(n101) );
  NANDN U155 ( .A(b[0]), .B(a[3]), .Z(n100) );
  NAND U156 ( .A(n101), .B(n100), .Z(n122) );
  XNOR U157 ( .A(n121), .B(n122), .Z(n123) );
  XNOR U158 ( .A(n124), .B(n123), .Z(n104) );
  NANDN U159 ( .A(n103), .B(n102), .Z(n105) );
  XOR U160 ( .A(n104), .B(n105), .Z(n107) );
  XNOR U161 ( .A(n106), .B(n107), .Z(n128) );
  XOR U162 ( .A(n129), .B(n128), .Z(c[116]) );
  NANDN U163 ( .A(n105), .B(n104), .Z(n109) );
  NANDN U164 ( .A(n107), .B(n106), .Z(n108) );
  AND U165 ( .A(n109), .B(n108), .Z(n140) );
  NANDN U166 ( .A(n9374), .B(n110), .Z(n112) );
  XOR U167 ( .A(b[3]), .B(a[3]), .Z(n149) );
  NANDN U168 ( .A(n9375), .B(n149), .Z(n111) );
  AND U169 ( .A(n112), .B(n111), .Z(n156) );
  NAND U170 ( .A(b[3]), .B(b[4]), .Z(n113) );
  AND U171 ( .A(b[5]), .B(n113), .Z(n9706) );
  ANDN U172 ( .B(n9706), .A(n121), .Z(n155) );
  XNOR U173 ( .A(n156), .B(n155), .Z(n158) );
  NAND U174 ( .A(b[0]), .B(a[5]), .Z(n114) );
  XNOR U175 ( .A(b[1]), .B(n114), .Z(n116) );
  NANDN U176 ( .A(b[0]), .B(a[4]), .Z(n115) );
  NAND U177 ( .A(n116), .B(n115), .Z(n147) );
  XOR U178 ( .A(b[5]), .B(b[4]), .Z(n143) );
  XOR U179 ( .A(b[5]), .B(a[0]), .Z(n117) );
  NAND U180 ( .A(n143), .B(n117), .Z(n118) );
  OR U181 ( .A(n118), .B(n9581), .Z(n120) );
  XOR U182 ( .A(b[5]), .B(a[1]), .Z(n144) );
  NAND U183 ( .A(n9581), .B(n144), .Z(n119) );
  NAND U184 ( .A(n120), .B(n119), .Z(n148) );
  XNOR U185 ( .A(n147), .B(n148), .Z(n157) );
  XOR U186 ( .A(n158), .B(n157), .Z(n138) );
  NANDN U187 ( .A(n122), .B(n121), .Z(n126) );
  NANDN U188 ( .A(n124), .B(n123), .Z(n125) );
  AND U189 ( .A(n126), .B(n125), .Z(n137) );
  XNOR U190 ( .A(n138), .B(n137), .Z(n139) );
  XOR U191 ( .A(n140), .B(n139), .Z(n132) );
  XNOR U192 ( .A(n132), .B(sreg[117]), .Z(n134) );
  NAND U193 ( .A(n127), .B(sreg[116]), .Z(n131) );
  NAND U194 ( .A(n129), .B(n128), .Z(n130) );
  NAND U195 ( .A(n131), .B(n130), .Z(n133) );
  XOR U196 ( .A(n134), .B(n133), .Z(c[117]) );
  NANDN U197 ( .A(n132), .B(sreg[117]), .Z(n136) );
  NAND U198 ( .A(n134), .B(n133), .Z(n135) );
  AND U199 ( .A(n136), .B(n135), .Z(n195) );
  XNOR U200 ( .A(n195), .B(sreg[118]), .Z(n197) );
  NANDN U201 ( .A(n138), .B(n137), .Z(n142) );
  NAND U202 ( .A(n140), .B(n139), .Z(n141) );
  AND U203 ( .A(n142), .B(n141), .Z(n163) );
  ANDN U204 ( .B(n143), .A(n9581), .Z(n9580) );
  IV U205 ( .A(n9580), .Z(n9437) );
  NANDN U206 ( .A(n9437), .B(n144), .Z(n146) );
  XOR U207 ( .A(b[5]), .B(a[2]), .Z(n167) );
  NANDN U208 ( .A(n9503), .B(n167), .Z(n145) );
  AND U209 ( .A(n146), .B(n145), .Z(n190) );
  ANDN U210 ( .B(n148), .A(n147), .Z(n189) );
  XNOR U211 ( .A(n190), .B(n189), .Z(n192) );
  NANDN U212 ( .A(n9374), .B(n149), .Z(n151) );
  XOR U213 ( .A(b[3]), .B(a[4]), .Z(n180) );
  NANDN U214 ( .A(n9375), .B(n180), .Z(n150) );
  AND U215 ( .A(n151), .B(n150), .Z(n186) );
  XOR U216 ( .A(b[6]), .B(b[5]), .Z(n9696) );
  IV U217 ( .A(n9696), .Z(n9639) );
  ANDN U218 ( .B(a[0]), .A(n9639), .Z(n183) );
  NAND U219 ( .A(b[0]), .B(a[6]), .Z(n152) );
  XNOR U220 ( .A(b[1]), .B(n152), .Z(n154) );
  NANDN U221 ( .A(b[0]), .B(a[5]), .Z(n153) );
  NAND U222 ( .A(n154), .B(n153), .Z(n184) );
  XNOR U223 ( .A(n183), .B(n184), .Z(n185) );
  XNOR U224 ( .A(n186), .B(n185), .Z(n191) );
  XOR U225 ( .A(n192), .B(n191), .Z(n162) );
  NANDN U226 ( .A(n156), .B(n155), .Z(n160) );
  NAND U227 ( .A(n158), .B(n157), .Z(n159) );
  AND U228 ( .A(n160), .B(n159), .Z(n161) );
  XOR U229 ( .A(n162), .B(n161), .Z(n164) );
  XNOR U230 ( .A(n163), .B(n164), .Z(n196) );
  XOR U231 ( .A(n197), .B(n196), .Z(c[118]) );
  NANDN U232 ( .A(n162), .B(n161), .Z(n166) );
  OR U233 ( .A(n164), .B(n163), .Z(n165) );
  AND U234 ( .A(n166), .B(n165), .Z(n207) );
  NANDN U235 ( .A(n9437), .B(n167), .Z(n169) );
  XOR U236 ( .A(b[5]), .B(a[3]), .Z(n235) );
  NANDN U237 ( .A(n9503), .B(n235), .Z(n168) );
  AND U238 ( .A(n169), .B(n168), .Z(n230) );
  XOR U239 ( .A(b[7]), .B(a[1]), .Z(n224) );
  NANDN U240 ( .A(n9639), .B(n224), .Z(n176) );
  ANDN U241 ( .B(b[6]), .A(b[7]), .Z(n170) );
  NAND U242 ( .A(n170), .B(a[0]), .Z(n173) );
  NAND U243 ( .A(b[5]), .B(b[6]), .Z(n171) );
  NAND U244 ( .A(b[7]), .B(n171), .Z(n9765) );
  OR U245 ( .A(a[0]), .B(n9765), .Z(n172) );
  NAND U246 ( .A(n173), .B(n172), .Z(n174) );
  NAND U247 ( .A(n9639), .B(n174), .Z(n175) );
  AND U248 ( .A(n176), .B(n175), .Z(n231) );
  XOR U249 ( .A(n230), .B(n231), .Z(n220) );
  NOR U250 ( .A(n9765), .B(n183), .Z(n218) );
  NAND U251 ( .A(b[0]), .B(a[7]), .Z(n177) );
  XNOR U252 ( .A(b[1]), .B(n177), .Z(n179) );
  NANDN U253 ( .A(b[0]), .B(a[6]), .Z(n178) );
  NAND U254 ( .A(n179), .B(n178), .Z(n217) );
  XNOR U255 ( .A(n218), .B(n217), .Z(n219) );
  XNOR U256 ( .A(n220), .B(n219), .Z(n211) );
  NAND U257 ( .A(n9420), .B(n180), .Z(n182) );
  XNOR U258 ( .A(b[3]), .B(a[5]), .Z(n227) );
  NANDN U259 ( .A(n227), .B(n9421), .Z(n181) );
  NAND U260 ( .A(n182), .B(n181), .Z(n212) );
  XNOR U261 ( .A(n211), .B(n212), .Z(n213) );
  NANDN U262 ( .A(n184), .B(n183), .Z(n188) );
  NANDN U263 ( .A(n186), .B(n185), .Z(n187) );
  NAND U264 ( .A(n188), .B(n187), .Z(n214) );
  XNOR U265 ( .A(n213), .B(n214), .Z(n205) );
  NANDN U266 ( .A(n190), .B(n189), .Z(n194) );
  NAND U267 ( .A(n192), .B(n191), .Z(n193) );
  NAND U268 ( .A(n194), .B(n193), .Z(n206) );
  XOR U269 ( .A(n205), .B(n206), .Z(n208) );
  XOR U270 ( .A(n207), .B(n208), .Z(n200) );
  XNOR U271 ( .A(n200), .B(sreg[119]), .Z(n202) );
  NANDN U272 ( .A(n195), .B(sreg[118]), .Z(n199) );
  NAND U273 ( .A(n197), .B(n196), .Z(n198) );
  NAND U274 ( .A(n199), .B(n198), .Z(n201) );
  XOR U275 ( .A(n202), .B(n201), .Z(c[119]) );
  NANDN U276 ( .A(n200), .B(sreg[119]), .Z(n204) );
  NAND U277 ( .A(n202), .B(n201), .Z(n203) );
  AND U278 ( .A(n204), .B(n203), .Z(n279) );
  XNOR U279 ( .A(n279), .B(sreg[120]), .Z(n281) );
  NANDN U280 ( .A(n206), .B(n205), .Z(n210) );
  OR U281 ( .A(n208), .B(n207), .Z(n209) );
  AND U282 ( .A(n210), .B(n209), .Z(n275) );
  NANDN U283 ( .A(n212), .B(n211), .Z(n216) );
  NANDN U284 ( .A(n214), .B(n213), .Z(n215) );
  AND U285 ( .A(n216), .B(n215), .Z(n274) );
  NANDN U286 ( .A(n218), .B(n217), .Z(n222) );
  NANDN U287 ( .A(n220), .B(n219), .Z(n221) );
  AND U288 ( .A(n222), .B(n221), .Z(n241) );
  XOR U289 ( .A(b[6]), .B(b[7]), .Z(n223) );
  ANDN U290 ( .B(n223), .A(n9696), .Z(n9695) );
  IV U291 ( .A(n9695), .Z(n9588) );
  NANDN U292 ( .A(n9588), .B(n224), .Z(n226) );
  XOR U293 ( .A(b[7]), .B(a[2]), .Z(n259) );
  NANDN U294 ( .A(n9639), .B(n259), .Z(n225) );
  AND U295 ( .A(n226), .B(n225), .Z(n245) );
  NANDN U296 ( .A(n227), .B(n9420), .Z(n229) );
  XOR U297 ( .A(b[3]), .B(a[6]), .Z(n270) );
  NANDN U298 ( .A(n9375), .B(n270), .Z(n228) );
  NAND U299 ( .A(n229), .B(n228), .Z(n244) );
  XNOR U300 ( .A(n245), .B(n244), .Z(n247) );
  NOR U301 ( .A(n231), .B(n230), .Z(n246) );
  XOR U302 ( .A(n247), .B(n246), .Z(n239) );
  NAND U303 ( .A(b[0]), .B(a[8]), .Z(n232) );
  XNOR U304 ( .A(b[1]), .B(n232), .Z(n234) );
  NANDN U305 ( .A(b[0]), .B(a[7]), .Z(n233) );
  NAND U306 ( .A(n234), .B(n233), .Z(n252) );
  XOR U307 ( .A(b[8]), .B(b[7]), .Z(n9804) );
  IV U308 ( .A(n9804), .Z(n9758) );
  ANDN U309 ( .B(a[0]), .A(n9758), .Z(n263) );
  NANDN U310 ( .A(n9437), .B(n235), .Z(n237) );
  XOR U311 ( .A(b[5]), .B(a[4]), .Z(n264) );
  NANDN U312 ( .A(n9503), .B(n264), .Z(n236) );
  AND U313 ( .A(n237), .B(n236), .Z(n250) );
  XOR U314 ( .A(n263), .B(n250), .Z(n251) );
  XNOR U315 ( .A(n252), .B(n251), .Z(n238) );
  XNOR U316 ( .A(n239), .B(n238), .Z(n240) );
  XNOR U317 ( .A(n241), .B(n240), .Z(n273) );
  XOR U318 ( .A(n274), .B(n273), .Z(n276) );
  XNOR U319 ( .A(n275), .B(n276), .Z(n280) );
  XOR U320 ( .A(n281), .B(n280), .Z(c[120]) );
  NANDN U321 ( .A(n239), .B(n238), .Z(n243) );
  NANDN U322 ( .A(n241), .B(n240), .Z(n242) );
  AND U323 ( .A(n243), .B(n242), .Z(n289) );
  NANDN U324 ( .A(n245), .B(n244), .Z(n249) );
  NAND U325 ( .A(n247), .B(n246), .Z(n248) );
  AND U326 ( .A(n249), .B(n248), .Z(n328) );
  NANDN U327 ( .A(n250), .B(n263), .Z(n254) );
  OR U328 ( .A(n252), .B(n251), .Z(n253) );
  AND U329 ( .A(n254), .B(n253), .Z(n326) );
  XOR U330 ( .A(b[9]), .B(b[8]), .Z(n316) );
  XOR U331 ( .A(b[9]), .B(a[0]), .Z(n255) );
  NAND U332 ( .A(n316), .B(n255), .Z(n256) );
  OR U333 ( .A(n256), .B(n9804), .Z(n258) );
  XOR U334 ( .A(b[9]), .B(a[1]), .Z(n317) );
  NAND U335 ( .A(n9804), .B(n317), .Z(n257) );
  AND U336 ( .A(n258), .B(n257), .Z(n320) );
  NANDN U337 ( .A(n9588), .B(n259), .Z(n261) );
  XOR U338 ( .A(b[7]), .B(a[3]), .Z(n310) );
  NANDN U339 ( .A(n9639), .B(n310), .Z(n260) );
  NAND U340 ( .A(n261), .B(n260), .Z(n321) );
  XOR U341 ( .A(n320), .B(n321), .Z(n297) );
  NAND U342 ( .A(b[7]), .B(b[8]), .Z(n262) );
  NAND U343 ( .A(b[9]), .B(n262), .Z(n9866) );
  NOR U344 ( .A(n9866), .B(n263), .Z(n296) );
  NANDN U345 ( .A(n9437), .B(n264), .Z(n266) );
  XOR U346 ( .A(b[5]), .B(a[5]), .Z(n313) );
  NANDN U347 ( .A(n9503), .B(n313), .Z(n265) );
  AND U348 ( .A(n266), .B(n265), .Z(n295) );
  XOR U349 ( .A(n296), .B(n295), .Z(n298) );
  XOR U350 ( .A(n297), .B(n298), .Z(n304) );
  NAND U351 ( .A(b[0]), .B(a[9]), .Z(n267) );
  XNOR U352 ( .A(b[1]), .B(n267), .Z(n269) );
  NANDN U353 ( .A(b[0]), .B(a[8]), .Z(n268) );
  NAND U354 ( .A(n269), .B(n268), .Z(n302) );
  NANDN U355 ( .A(n9374), .B(n270), .Z(n272) );
  XOR U356 ( .A(b[3]), .B(a[7]), .Z(n322) );
  NANDN U357 ( .A(n9375), .B(n322), .Z(n271) );
  NAND U358 ( .A(n272), .B(n271), .Z(n301) );
  XNOR U359 ( .A(n302), .B(n301), .Z(n303) );
  XOR U360 ( .A(n304), .B(n303), .Z(n325) );
  XNOR U361 ( .A(n326), .B(n325), .Z(n327) );
  XOR U362 ( .A(n328), .B(n327), .Z(n290) );
  XNOR U363 ( .A(n289), .B(n290), .Z(n291) );
  NANDN U364 ( .A(n274), .B(n273), .Z(n278) );
  OR U365 ( .A(n276), .B(n275), .Z(n277) );
  NAND U366 ( .A(n278), .B(n277), .Z(n292) );
  XOR U367 ( .A(n291), .B(n292), .Z(n284) );
  XNOR U368 ( .A(sreg[121]), .B(n284), .Z(n286) );
  NANDN U369 ( .A(n279), .B(sreg[120]), .Z(n283) );
  NAND U370 ( .A(n281), .B(n280), .Z(n282) );
  NAND U371 ( .A(n283), .B(n282), .Z(n285) );
  XOR U372 ( .A(n286), .B(n285), .Z(c[121]) );
  NANDN U373 ( .A(n284), .B(sreg[121]), .Z(n288) );
  NAND U374 ( .A(n286), .B(n285), .Z(n287) );
  AND U375 ( .A(n288), .B(n287), .Z(n381) );
  XNOR U376 ( .A(sreg[122]), .B(n381), .Z(n383) );
  NANDN U377 ( .A(n290), .B(n289), .Z(n294) );
  NANDN U378 ( .A(n292), .B(n291), .Z(n293) );
  AND U379 ( .A(n294), .B(n293), .Z(n333) );
  NANDN U380 ( .A(n296), .B(n295), .Z(n300) );
  NANDN U381 ( .A(n298), .B(n297), .Z(n299) );
  AND U382 ( .A(n300), .B(n299), .Z(n376) );
  NANDN U383 ( .A(n302), .B(n301), .Z(n306) );
  NAND U384 ( .A(n304), .B(n303), .Z(n305) );
  AND U385 ( .A(n306), .B(n305), .Z(n375) );
  XNOR U386 ( .A(n376), .B(n375), .Z(n377) );
  NAND U387 ( .A(b[0]), .B(a[10]), .Z(n307) );
  XNOR U388 ( .A(b[1]), .B(n307), .Z(n309) );
  NANDN U389 ( .A(b[0]), .B(a[9]), .Z(n308) );
  NAND U390 ( .A(n309), .B(n308), .Z(n345) );
  XNOR U391 ( .A(b[9]), .B(b[10]), .Z(n9856) );
  ANDN U392 ( .B(a[0]), .A(n9856), .Z(n374) );
  NANDN U393 ( .A(n9588), .B(n310), .Z(n312) );
  XOR U394 ( .A(b[7]), .B(a[4]), .Z(n370) );
  NANDN U395 ( .A(n9639), .B(n370), .Z(n311) );
  AND U396 ( .A(n312), .B(n311), .Z(n343) );
  XOR U397 ( .A(n374), .B(n343), .Z(n344) );
  XOR U398 ( .A(n345), .B(n344), .Z(n340) );
  NANDN U399 ( .A(n9437), .B(n313), .Z(n315) );
  XOR U400 ( .A(b[5]), .B(a[6]), .Z(n364) );
  NANDN U401 ( .A(n9503), .B(n364), .Z(n314) );
  AND U402 ( .A(n315), .B(n314), .Z(n349) );
  ANDN U403 ( .B(n316), .A(n9804), .Z(n9803) );
  IV U404 ( .A(n9803), .Z(n9685) );
  NANDN U405 ( .A(n9685), .B(n317), .Z(n319) );
  XOR U406 ( .A(b[9]), .B(a[2]), .Z(n358) );
  NANDN U407 ( .A(n9758), .B(n358), .Z(n318) );
  NAND U408 ( .A(n319), .B(n318), .Z(n348) );
  XNOR U409 ( .A(n349), .B(n348), .Z(n351) );
  ANDN U410 ( .B(n321), .A(n320), .Z(n350) );
  XOR U411 ( .A(n351), .B(n350), .Z(n338) );
  NAND U412 ( .A(n9420), .B(n322), .Z(n324) );
  XNOR U413 ( .A(b[3]), .B(a[8]), .Z(n367) );
  NANDN U414 ( .A(n367), .B(n9421), .Z(n323) );
  AND U415 ( .A(n324), .B(n323), .Z(n337) );
  XNOR U416 ( .A(n338), .B(n337), .Z(n339) );
  XOR U417 ( .A(n340), .B(n339), .Z(n378) );
  XNOR U418 ( .A(n377), .B(n378), .Z(n331) );
  NANDN U419 ( .A(n326), .B(n325), .Z(n330) );
  NANDN U420 ( .A(n328), .B(n327), .Z(n329) );
  NAND U421 ( .A(n330), .B(n329), .Z(n332) );
  XOR U422 ( .A(n331), .B(n332), .Z(n334) );
  XNOR U423 ( .A(n333), .B(n334), .Z(n382) );
  XNOR U424 ( .A(n383), .B(n382), .Z(c[122]) );
  NANDN U425 ( .A(n332), .B(n331), .Z(n336) );
  NANDN U426 ( .A(n334), .B(n333), .Z(n335) );
  AND U427 ( .A(n336), .B(n335), .Z(n388) );
  NANDN U428 ( .A(n338), .B(n337), .Z(n342) );
  NANDN U429 ( .A(n340), .B(n339), .Z(n341) );
  AND U430 ( .A(n342), .B(n341), .Z(n434) );
  NANDN U431 ( .A(n343), .B(n374), .Z(n347) );
  OR U432 ( .A(n345), .B(n344), .Z(n346) );
  AND U433 ( .A(n347), .B(n346), .Z(n432) );
  NANDN U434 ( .A(n349), .B(n348), .Z(n353) );
  NAND U435 ( .A(n351), .B(n350), .Z(n352) );
  AND U436 ( .A(n353), .B(n352), .Z(n428) );
  XOR U437 ( .A(b[11]), .B(b[10]), .Z(n403) );
  XOR U438 ( .A(b[11]), .B(a[0]), .Z(n354) );
  NAND U439 ( .A(n403), .B(n354), .Z(n355) );
  OR U440 ( .A(n355), .B(n9882), .Z(n357) );
  XOR U441 ( .A(b[11]), .B(a[1]), .Z(n404) );
  NAND U442 ( .A(n9882), .B(n404), .Z(n356) );
  AND U443 ( .A(n357), .B(n356), .Z(n393) );
  NANDN U444 ( .A(n9685), .B(n358), .Z(n360) );
  XOR U445 ( .A(b[9]), .B(a[3]), .Z(n410) );
  NANDN U446 ( .A(n9758), .B(n410), .Z(n359) );
  AND U447 ( .A(n360), .B(n359), .Z(n392) );
  XOR U448 ( .A(n393), .B(n392), .Z(n415) );
  NAND U449 ( .A(b[0]), .B(a[11]), .Z(n361) );
  XNOR U450 ( .A(b[1]), .B(n361), .Z(n363) );
  NANDN U451 ( .A(b[0]), .B(a[10]), .Z(n362) );
  NAND U452 ( .A(n363), .B(n362), .Z(n413) );
  NAND U453 ( .A(n9580), .B(n364), .Z(n366) );
  XNOR U454 ( .A(b[5]), .B(a[7]), .Z(n400) );
  NANDN U455 ( .A(n400), .B(n9581), .Z(n365) );
  NAND U456 ( .A(n366), .B(n365), .Z(n414) );
  XOR U457 ( .A(n413), .B(n414), .Z(n416) );
  XOR U458 ( .A(n415), .B(n416), .Z(n426) );
  NANDN U459 ( .A(n367), .B(n9420), .Z(n369) );
  XOR U460 ( .A(b[3]), .B(a[9]), .Z(n394) );
  NANDN U461 ( .A(n9375), .B(n394), .Z(n368) );
  AND U462 ( .A(n369), .B(n368), .Z(n422) );
  NANDN U463 ( .A(n9588), .B(n370), .Z(n372) );
  XOR U464 ( .A(b[7]), .B(a[5]), .Z(n397) );
  NANDN U465 ( .A(n9639), .B(n397), .Z(n371) );
  AND U466 ( .A(n372), .B(n371), .Z(n420) );
  NAND U467 ( .A(b[9]), .B(b[10]), .Z(n373) );
  AND U468 ( .A(b[11]), .B(n373), .Z(n9965) );
  ANDN U469 ( .B(n9965), .A(n374), .Z(n419) );
  XNOR U470 ( .A(n420), .B(n419), .Z(n421) );
  XNOR U471 ( .A(n422), .B(n421), .Z(n425) );
  XNOR U472 ( .A(n426), .B(n425), .Z(n427) );
  XNOR U473 ( .A(n428), .B(n427), .Z(n431) );
  XNOR U474 ( .A(n432), .B(n431), .Z(n433) );
  XOR U475 ( .A(n434), .B(n433), .Z(n387) );
  NANDN U476 ( .A(n376), .B(n375), .Z(n380) );
  NANDN U477 ( .A(n378), .B(n377), .Z(n379) );
  NAND U478 ( .A(n380), .B(n379), .Z(n386) );
  XOR U479 ( .A(n387), .B(n386), .Z(n389) );
  XOR U480 ( .A(n388), .B(n389), .Z(n437) );
  XNOR U481 ( .A(n437), .B(sreg[123]), .Z(n439) );
  NANDN U482 ( .A(sreg[122]), .B(n381), .Z(n385) );
  NAND U483 ( .A(n383), .B(n382), .Z(n384) );
  AND U484 ( .A(n385), .B(n384), .Z(n438) );
  XOR U485 ( .A(n439), .B(n438), .Z(c[123]) );
  NANDN U486 ( .A(n387), .B(n386), .Z(n391) );
  OR U487 ( .A(n389), .B(n388), .Z(n390) );
  AND U488 ( .A(n391), .B(n390), .Z(n448) );
  NOR U489 ( .A(n393), .B(n392), .Z(n494) );
  NAND U490 ( .A(n9420), .B(n394), .Z(n396) );
  XNOR U491 ( .A(b[3]), .B(a[10]), .Z(n476) );
  NANDN U492 ( .A(n476), .B(n9421), .Z(n395) );
  AND U493 ( .A(n396), .B(n395), .Z(n492) );
  NAND U494 ( .A(n9695), .B(n397), .Z(n399) );
  XNOR U495 ( .A(b[7]), .B(a[6]), .Z(n466) );
  NANDN U496 ( .A(n466), .B(n9696), .Z(n398) );
  NAND U497 ( .A(n399), .B(n398), .Z(n493) );
  XOR U498 ( .A(n492), .B(n493), .Z(n495) );
  XOR U499 ( .A(n494), .B(n495), .Z(n460) );
  NANDN U500 ( .A(n400), .B(n9580), .Z(n402) );
  XOR U501 ( .A(b[5]), .B(a[8]), .Z(n483) );
  NANDN U502 ( .A(n9503), .B(n483), .Z(n401) );
  AND U503 ( .A(n402), .B(n401), .Z(n458) );
  ANDN U504 ( .B(n403), .A(n9882), .Z(n9883) );
  NAND U505 ( .A(n404), .B(n9883), .Z(n406) );
  XOR U506 ( .A(b[11]), .B(a[2]), .Z(n469) );
  NANDN U507 ( .A(n9856), .B(n469), .Z(n405) );
  NAND U508 ( .A(n406), .B(n405), .Z(n457) );
  XNOR U509 ( .A(n458), .B(n457), .Z(n459) );
  XNOR U510 ( .A(n460), .B(n459), .Z(n454) );
  NAND U511 ( .A(b[0]), .B(a[12]), .Z(n407) );
  XNOR U512 ( .A(b[1]), .B(n407), .Z(n409) );
  NANDN U513 ( .A(b[0]), .B(a[11]), .Z(n408) );
  NAND U514 ( .A(n409), .B(n408), .Z(n489) );
  XOR U515 ( .A(b[12]), .B(b[11]), .Z(n9973) );
  IV U516 ( .A(n9973), .Z(n9935) );
  ANDN U517 ( .B(a[0]), .A(n9935), .Z(n486) );
  NANDN U518 ( .A(n9685), .B(n410), .Z(n412) );
  XOR U519 ( .A(b[9]), .B(a[4]), .Z(n479) );
  NANDN U520 ( .A(n9758), .B(n479), .Z(n411) );
  AND U521 ( .A(n412), .B(n411), .Z(n487) );
  XNOR U522 ( .A(n486), .B(n487), .Z(n488) );
  XNOR U523 ( .A(n489), .B(n488), .Z(n451) );
  NANDN U524 ( .A(n414), .B(n413), .Z(n418) );
  OR U525 ( .A(n416), .B(n415), .Z(n417) );
  NAND U526 ( .A(n418), .B(n417), .Z(n452) );
  XNOR U527 ( .A(n451), .B(n452), .Z(n453) );
  XOR U528 ( .A(n454), .B(n453), .Z(n501) );
  NANDN U529 ( .A(n420), .B(n419), .Z(n424) );
  NANDN U530 ( .A(n422), .B(n421), .Z(n423) );
  AND U531 ( .A(n424), .B(n423), .Z(n498) );
  NANDN U532 ( .A(n426), .B(n425), .Z(n430) );
  NANDN U533 ( .A(n428), .B(n427), .Z(n429) );
  NAND U534 ( .A(n430), .B(n429), .Z(n499) );
  XNOR U535 ( .A(n498), .B(n499), .Z(n500) );
  XNOR U536 ( .A(n501), .B(n500), .Z(n445) );
  NANDN U537 ( .A(n432), .B(n431), .Z(n436) );
  NAND U538 ( .A(n434), .B(n433), .Z(n435) );
  NAND U539 ( .A(n436), .B(n435), .Z(n446) );
  XNOR U540 ( .A(n445), .B(n446), .Z(n447) );
  XNOR U541 ( .A(n448), .B(n447), .Z(n444) );
  NANDN U542 ( .A(n437), .B(sreg[123]), .Z(n441) );
  NAND U543 ( .A(n439), .B(n438), .Z(n440) );
  NAND U544 ( .A(n441), .B(n440), .Z(n443) );
  XOR U545 ( .A(n443), .B(sreg[124]), .Z(n442) );
  XNOR U546 ( .A(n444), .B(n442), .Z(c[124]) );
  NANDN U547 ( .A(n446), .B(n445), .Z(n450) );
  NANDN U548 ( .A(n448), .B(n447), .Z(n449) );
  AND U549 ( .A(n450), .B(n449), .Z(n507) );
  NANDN U550 ( .A(n452), .B(n451), .Z(n456) );
  NAND U551 ( .A(n454), .B(n453), .Z(n455) );
  AND U552 ( .A(n456), .B(n455), .Z(n560) );
  NANDN U553 ( .A(n458), .B(n457), .Z(n462) );
  NANDN U554 ( .A(n460), .B(n459), .Z(n461) );
  AND U555 ( .A(n462), .B(n461), .Z(n559) );
  NAND U556 ( .A(b[0]), .B(a[13]), .Z(n463) );
  XNOR U557 ( .A(b[1]), .B(n463), .Z(n465) );
  NANDN U558 ( .A(b[0]), .B(a[12]), .Z(n464) );
  NAND U559 ( .A(n465), .B(n464), .Z(n544) );
  NANDN U560 ( .A(n466), .B(n9695), .Z(n468) );
  XOR U561 ( .A(b[7]), .B(a[7]), .Z(n537) );
  NANDN U562 ( .A(n9639), .B(n537), .Z(n467) );
  NAND U563 ( .A(n468), .B(n467), .Z(n543) );
  XNOR U564 ( .A(n544), .B(n543), .Z(n546) );
  NAND U565 ( .A(n469), .B(n9883), .Z(n471) );
  XOR U566 ( .A(b[11]), .B(a[3]), .Z(n531) );
  NANDN U567 ( .A(n9856), .B(n531), .Z(n470) );
  AND U568 ( .A(n471), .B(n470), .Z(n556) );
  XOR U569 ( .A(b[13]), .B(b[12]), .Z(n549) );
  XOR U570 ( .A(b[13]), .B(a[0]), .Z(n472) );
  NAND U571 ( .A(n549), .B(n472), .Z(n473) );
  OR U572 ( .A(n473), .B(n9973), .Z(n475) );
  XOR U573 ( .A(b[13]), .B(a[1]), .Z(n550) );
  NAND U574 ( .A(n9973), .B(n550), .Z(n474) );
  NAND U575 ( .A(n475), .B(n474), .Z(n557) );
  XNOR U576 ( .A(n556), .B(n557), .Z(n545) );
  XOR U577 ( .A(n546), .B(n545), .Z(n518) );
  NANDN U578 ( .A(n476), .B(n9420), .Z(n478) );
  XOR U579 ( .A(b[3]), .B(a[11]), .Z(n540) );
  NANDN U580 ( .A(n9375), .B(n540), .Z(n477) );
  AND U581 ( .A(n478), .B(n477), .Z(n523) );
  NANDN U582 ( .A(n9685), .B(n479), .Z(n481) );
  XOR U583 ( .A(b[9]), .B(a[5]), .Z(n553) );
  NANDN U584 ( .A(n9758), .B(n553), .Z(n480) );
  NAND U585 ( .A(n481), .B(n480), .Z(n522) );
  XNOR U586 ( .A(n523), .B(n522), .Z(n525) );
  NAND U587 ( .A(b[11]), .B(b[12]), .Z(n482) );
  AND U588 ( .A(b[13]), .B(n482), .Z(n9999) );
  ANDN U589 ( .B(n9999), .A(n486), .Z(n524) );
  XOR U590 ( .A(n525), .B(n524), .Z(n517) );
  NAND U591 ( .A(n9580), .B(n483), .Z(n485) );
  XNOR U592 ( .A(b[5]), .B(a[9]), .Z(n534) );
  NANDN U593 ( .A(n534), .B(n9581), .Z(n484) );
  AND U594 ( .A(n485), .B(n484), .Z(n516) );
  XOR U595 ( .A(n517), .B(n516), .Z(n519) );
  XOR U596 ( .A(n518), .B(n519), .Z(n513) );
  NANDN U597 ( .A(n487), .B(n486), .Z(n491) );
  NANDN U598 ( .A(n489), .B(n488), .Z(n490) );
  AND U599 ( .A(n491), .B(n490), .Z(n511) );
  NANDN U600 ( .A(n493), .B(n492), .Z(n497) );
  OR U601 ( .A(n495), .B(n494), .Z(n496) );
  AND U602 ( .A(n497), .B(n496), .Z(n510) );
  XNOR U603 ( .A(n511), .B(n510), .Z(n512) );
  XNOR U604 ( .A(n513), .B(n512), .Z(n558) );
  XOR U605 ( .A(n559), .B(n558), .Z(n561) );
  XOR U606 ( .A(n560), .B(n561), .Z(n505) );
  NANDN U607 ( .A(n499), .B(n498), .Z(n503) );
  NANDN U608 ( .A(n501), .B(n500), .Z(n502) );
  NAND U609 ( .A(n503), .B(n502), .Z(n504) );
  XNOR U610 ( .A(n505), .B(n504), .Z(n506) );
  XNOR U611 ( .A(n507), .B(n506), .Z(n564) );
  XNOR U612 ( .A(sreg[125]), .B(n564), .Z(n565) );
  XNOR U613 ( .A(n566), .B(n565), .Z(c[125]) );
  NANDN U614 ( .A(n505), .B(n504), .Z(n509) );
  NANDN U615 ( .A(n507), .B(n506), .Z(n508) );
  AND U616 ( .A(n509), .B(n508), .Z(n572) );
  NANDN U617 ( .A(n511), .B(n510), .Z(n515) );
  NANDN U618 ( .A(n513), .B(n512), .Z(n514) );
  AND U619 ( .A(n515), .B(n514), .Z(n632) );
  NANDN U620 ( .A(n517), .B(n516), .Z(n521) );
  OR U621 ( .A(n519), .B(n518), .Z(n520) );
  AND U622 ( .A(n521), .B(n520), .Z(n630) );
  NANDN U623 ( .A(n523), .B(n522), .Z(n527) );
  NAND U624 ( .A(n525), .B(n524), .Z(n526) );
  AND U625 ( .A(n527), .B(n526), .Z(n617) );
  NAND U626 ( .A(b[0]), .B(a[14]), .Z(n528) );
  XNOR U627 ( .A(b[1]), .B(n528), .Z(n530) );
  NANDN U628 ( .A(b[0]), .B(a[13]), .Z(n529) );
  NAND U629 ( .A(n530), .B(n529), .Z(n623) );
  XOR U630 ( .A(b[13]), .B(b[14]), .Z(n9989) );
  IV U631 ( .A(n9989), .Z(n10006) );
  ANDN U632 ( .B(a[0]), .A(n10006), .Z(n620) );
  NAND U633 ( .A(n531), .B(n9883), .Z(n533) );
  XOR U634 ( .A(b[11]), .B(a[4]), .Z(n592) );
  NANDN U635 ( .A(n9856), .B(n592), .Z(n532) );
  AND U636 ( .A(n533), .B(n532), .Z(n621) );
  XNOR U637 ( .A(n620), .B(n621), .Z(n622) );
  XNOR U638 ( .A(n623), .B(n622), .Z(n614) );
  NANDN U639 ( .A(n534), .B(n9580), .Z(n536) );
  XOR U640 ( .A(b[5]), .B(a[10]), .Z(n586) );
  NANDN U641 ( .A(n9503), .B(n586), .Z(n535) );
  AND U642 ( .A(n536), .B(n535), .Z(n598) );
  NANDN U643 ( .A(n9588), .B(n537), .Z(n539) );
  XOR U644 ( .A(b[7]), .B(a[8]), .Z(n582) );
  NANDN U645 ( .A(n9639), .B(n582), .Z(n538) );
  AND U646 ( .A(n539), .B(n538), .Z(n596) );
  NANDN U647 ( .A(n9374), .B(n540), .Z(n542) );
  XOR U648 ( .A(b[3]), .B(a[12]), .Z(n589) );
  NANDN U649 ( .A(n9375), .B(n589), .Z(n541) );
  NAND U650 ( .A(n542), .B(n541), .Z(n595) );
  XNOR U651 ( .A(n596), .B(n595), .Z(n597) );
  XOR U652 ( .A(n598), .B(n597), .Z(n615) );
  XNOR U653 ( .A(n614), .B(n615), .Z(n616) );
  XNOR U654 ( .A(n617), .B(n616), .Z(n578) );
  NANDN U655 ( .A(n544), .B(n543), .Z(n548) );
  NAND U656 ( .A(n546), .B(n545), .Z(n547) );
  AND U657 ( .A(n548), .B(n547), .Z(n577) );
  ANDN U658 ( .B(n549), .A(n9973), .Z(n9972) );
  IV U659 ( .A(n9972), .Z(n9891) );
  NANDN U660 ( .A(n9891), .B(n550), .Z(n552) );
  XOR U661 ( .A(b[13]), .B(a[2]), .Z(n601) );
  NANDN U662 ( .A(n9935), .B(n601), .Z(n551) );
  AND U663 ( .A(n552), .B(n551), .Z(n627) );
  NANDN U664 ( .A(n9685), .B(n553), .Z(n555) );
  XOR U665 ( .A(b[9]), .B(a[6]), .Z(n611) );
  NANDN U666 ( .A(n9758), .B(n611), .Z(n554) );
  NAND U667 ( .A(n555), .B(n554), .Z(n626) );
  XNOR U668 ( .A(n627), .B(n626), .Z(n629) );
  ANDN U669 ( .B(n557), .A(n556), .Z(n628) );
  XOR U670 ( .A(n629), .B(n628), .Z(n576) );
  XOR U671 ( .A(n577), .B(n576), .Z(n579) );
  XOR U672 ( .A(n578), .B(n579), .Z(n631) );
  XOR U673 ( .A(n630), .B(n631), .Z(n633) );
  XOR U674 ( .A(n632), .B(n633), .Z(n571) );
  NANDN U675 ( .A(n559), .B(n558), .Z(n563) );
  OR U676 ( .A(n561), .B(n560), .Z(n562) );
  AND U677 ( .A(n563), .B(n562), .Z(n570) );
  XOR U678 ( .A(n571), .B(n570), .Z(n573) );
  XNOR U679 ( .A(n572), .B(n573), .Z(n637) );
  NANDN U680 ( .A(sreg[125]), .B(n564), .Z(n568) );
  NAND U681 ( .A(n566), .B(n565), .Z(n567) );
  NAND U682 ( .A(n568), .B(n567), .Z(n636) );
  XOR U683 ( .A(sreg[126]), .B(n636), .Z(n569) );
  XNOR U684 ( .A(n637), .B(n569), .Z(c[126]) );
  NANDN U685 ( .A(n571), .B(n570), .Z(n575) );
  OR U686 ( .A(n573), .B(n572), .Z(n574) );
  AND U687 ( .A(n575), .B(n574), .Z(n641) );
  NANDN U688 ( .A(n577), .B(n576), .Z(n581) );
  NANDN U689 ( .A(n579), .B(n578), .Z(n580) );
  AND U690 ( .A(n581), .B(n580), .Z(n702) );
  NANDN U691 ( .A(n9588), .B(n582), .Z(n584) );
  XOR U692 ( .A(b[7]), .B(a[9]), .Z(n689) );
  NANDN U693 ( .A(n9639), .B(n689), .Z(n583) );
  AND U694 ( .A(n584), .B(n583), .Z(n676) );
  NAND U695 ( .A(b[13]), .B(b[14]), .Z(n10023) );
  ANDN U696 ( .B(n10023), .A(n620), .Z(n585) );
  AND U697 ( .A(b[15]), .B(n585), .Z(n675) );
  XNOR U698 ( .A(n676), .B(n675), .Z(n678) );
  NANDN U699 ( .A(n9437), .B(n586), .Z(n588) );
  XOR U700 ( .A(b[5]), .B(a[11]), .Z(n698) );
  NANDN U701 ( .A(n9503), .B(n698), .Z(n587) );
  AND U702 ( .A(n588), .B(n587), .Z(n672) );
  NANDN U703 ( .A(n9374), .B(n589), .Z(n591) );
  XOR U704 ( .A(b[3]), .B(a[13]), .Z(n683) );
  NANDN U705 ( .A(n9375), .B(n683), .Z(n590) );
  AND U706 ( .A(n591), .B(n590), .Z(n670) );
  NAND U707 ( .A(n592), .B(n9883), .Z(n594) );
  XOR U708 ( .A(b[11]), .B(a[5]), .Z(n692) );
  NANDN U709 ( .A(n9856), .B(n692), .Z(n593) );
  NAND U710 ( .A(n594), .B(n593), .Z(n669) );
  XNOR U711 ( .A(n670), .B(n669), .Z(n671) );
  XNOR U712 ( .A(n672), .B(n671), .Z(n677) );
  XOR U713 ( .A(n678), .B(n677), .Z(n653) );
  NANDN U714 ( .A(n596), .B(n595), .Z(n600) );
  NANDN U715 ( .A(n598), .B(n597), .Z(n599) );
  AND U716 ( .A(n600), .B(n599), .Z(n651) );
  NANDN U717 ( .A(n9891), .B(n601), .Z(n603) );
  XOR U718 ( .A(b[13]), .B(a[3]), .Z(n666) );
  NANDN U719 ( .A(n9935), .B(n666), .Z(n602) );
  AND U720 ( .A(n603), .B(n602), .Z(n682) );
  XOR U721 ( .A(b[14]), .B(b[15]), .Z(n604) );
  ANDN U722 ( .B(n604), .A(n9989), .Z(n9987) );
  IV U723 ( .A(n9987), .Z(n10005) );
  XOR U724 ( .A(a[0]), .B(b[15]), .Z(n605) );
  NANDN U725 ( .A(n10005), .B(n605), .Z(n607) );
  XOR U726 ( .A(b[15]), .B(a[1]), .Z(n695) );
  ANDN U727 ( .B(n695), .A(n10006), .Z(n606) );
  ANDN U728 ( .B(n607), .A(n606), .Z(n681) );
  XOR U729 ( .A(n682), .B(n681), .Z(n660) );
  NAND U730 ( .A(b[0]), .B(a[15]), .Z(n608) );
  XNOR U731 ( .A(b[1]), .B(n608), .Z(n610) );
  NANDN U732 ( .A(b[0]), .B(a[14]), .Z(n609) );
  NAND U733 ( .A(n610), .B(n609), .Z(n657) );
  NAND U734 ( .A(n9803), .B(n611), .Z(n613) );
  XNOR U735 ( .A(b[9]), .B(a[7]), .Z(n686) );
  NANDN U736 ( .A(n686), .B(n9804), .Z(n612) );
  NAND U737 ( .A(n613), .B(n612), .Z(n658) );
  XNOR U738 ( .A(n657), .B(n658), .Z(n659) );
  XOR U739 ( .A(n660), .B(n659), .Z(n652) );
  XOR U740 ( .A(n651), .B(n652), .Z(n654) );
  XNOR U741 ( .A(n653), .B(n654), .Z(n701) );
  XNOR U742 ( .A(n702), .B(n701), .Z(n704) );
  NANDN U743 ( .A(n615), .B(n614), .Z(n619) );
  NANDN U744 ( .A(n617), .B(n616), .Z(n618) );
  AND U745 ( .A(n619), .B(n618), .Z(n648) );
  NANDN U746 ( .A(n621), .B(n620), .Z(n625) );
  NANDN U747 ( .A(n623), .B(n622), .Z(n624) );
  AND U748 ( .A(n625), .B(n624), .Z(n646) );
  XNOR U749 ( .A(n646), .B(n645), .Z(n647) );
  XNOR U750 ( .A(n648), .B(n647), .Z(n703) );
  XOR U751 ( .A(n704), .B(n703), .Z(n640) );
  NANDN U752 ( .A(n631), .B(n630), .Z(n635) );
  OR U753 ( .A(n633), .B(n632), .Z(n634) );
  AND U754 ( .A(n635), .B(n634), .Z(n639) );
  XOR U755 ( .A(n640), .B(n639), .Z(n642) );
  XOR U756 ( .A(n641), .B(n642), .Z(n707) );
  XNOR U757 ( .A(sreg[127]), .B(n708), .Z(n638) );
  XOR U758 ( .A(n707), .B(n638), .Z(c[127]) );
  NANDN U759 ( .A(n640), .B(n639), .Z(n644) );
  OR U760 ( .A(n642), .B(n641), .Z(n643) );
  AND U761 ( .A(n644), .B(n643), .Z(n715) );
  NANDN U762 ( .A(n646), .B(n645), .Z(n650) );
  NANDN U763 ( .A(n648), .B(n647), .Z(n649) );
  AND U764 ( .A(n650), .B(n649), .Z(n780) );
  NANDN U765 ( .A(n652), .B(n651), .Z(n656) );
  OR U766 ( .A(n654), .B(n653), .Z(n655) );
  AND U767 ( .A(n656), .B(n655), .Z(n778) );
  NANDN U768 ( .A(n658), .B(n657), .Z(n662) );
  NANDN U769 ( .A(n660), .B(n659), .Z(n661) );
  AND U770 ( .A(n662), .B(n661), .Z(n773) );
  NAND U771 ( .A(b[0]), .B(a[16]), .Z(n663) );
  XNOR U772 ( .A(b[1]), .B(n663), .Z(n665) );
  NANDN U773 ( .A(b[0]), .B(a[15]), .Z(n664) );
  NAND U774 ( .A(n665), .B(n664), .Z(n721) );
  NANDN U775 ( .A(n9891), .B(n666), .Z(n668) );
  XOR U776 ( .A(b[13]), .B(a[4]), .Z(n727) );
  NANDN U777 ( .A(n9935), .B(n727), .Z(n667) );
  AND U778 ( .A(n668), .B(n667), .Z(n719) );
  AND U779 ( .A(b[15]), .B(a[0]), .Z(n718) );
  XOR U780 ( .A(n719), .B(n718), .Z(n720) );
  XNOR U781 ( .A(n721), .B(n720), .Z(n772) );
  XNOR U782 ( .A(n773), .B(n772), .Z(n775) );
  NANDN U783 ( .A(n670), .B(n669), .Z(n674) );
  NANDN U784 ( .A(n672), .B(n671), .Z(n673) );
  AND U785 ( .A(n674), .B(n673), .Z(n774) );
  XOR U786 ( .A(n775), .B(n774), .Z(n769) );
  NANDN U787 ( .A(n676), .B(n675), .Z(n680) );
  NAND U788 ( .A(n678), .B(n677), .Z(n679) );
  AND U789 ( .A(n680), .B(n679), .Z(n767) );
  NOR U790 ( .A(n682), .B(n681), .Z(n747) );
  NAND U791 ( .A(n9420), .B(n683), .Z(n685) );
  XNOR U792 ( .A(b[3]), .B(a[14]), .Z(n736) );
  NANDN U793 ( .A(n736), .B(n9421), .Z(n684) );
  AND U794 ( .A(n685), .B(n684), .Z(n745) );
  NANDN U795 ( .A(n686), .B(n9803), .Z(n688) );
  XNOR U796 ( .A(b[9]), .B(a[8]), .Z(n757) );
  NANDN U797 ( .A(n757), .B(n9804), .Z(n687) );
  NAND U798 ( .A(n688), .B(n687), .Z(n746) );
  XOR U799 ( .A(n745), .B(n746), .Z(n748) );
  XOR U800 ( .A(n747), .B(n748), .Z(n742) );
  NANDN U801 ( .A(n9588), .B(n689), .Z(n691) );
  XOR U802 ( .A(b[7]), .B(a[10]), .Z(n733) );
  NANDN U803 ( .A(n9639), .B(n733), .Z(n690) );
  AND U804 ( .A(n691), .B(n690), .Z(n740) );
  NAND U805 ( .A(n692), .B(n9883), .Z(n694) );
  XOR U806 ( .A(b[11]), .B(a[6]), .Z(n751) );
  NANDN U807 ( .A(n9856), .B(n751), .Z(n693) );
  AND U808 ( .A(n694), .B(n693), .Z(n763) );
  NANDN U809 ( .A(n10005), .B(n695), .Z(n697) );
  XOR U810 ( .A(b[15]), .B(a[2]), .Z(n754) );
  NANDN U811 ( .A(n10006), .B(n754), .Z(n696) );
  AND U812 ( .A(n697), .B(n696), .Z(n761) );
  NANDN U813 ( .A(n9437), .B(n698), .Z(n700) );
  XOR U814 ( .A(b[5]), .B(a[12]), .Z(n730) );
  NANDN U815 ( .A(n9503), .B(n730), .Z(n699) );
  NAND U816 ( .A(n700), .B(n699), .Z(n760) );
  XNOR U817 ( .A(n761), .B(n760), .Z(n762) );
  XNOR U818 ( .A(n763), .B(n762), .Z(n739) );
  XNOR U819 ( .A(n740), .B(n739), .Z(n741) );
  XNOR U820 ( .A(n742), .B(n741), .Z(n766) );
  XNOR U821 ( .A(n767), .B(n766), .Z(n768) );
  XOR U822 ( .A(n769), .B(n768), .Z(n779) );
  XOR U823 ( .A(n778), .B(n779), .Z(n781) );
  XOR U824 ( .A(n780), .B(n781), .Z(n713) );
  NANDN U825 ( .A(n702), .B(n701), .Z(n706) );
  NAND U826 ( .A(n704), .B(n703), .Z(n705) );
  AND U827 ( .A(n706), .B(n705), .Z(n712) );
  XNOR U828 ( .A(n713), .B(n712), .Z(n714) );
  XNOR U829 ( .A(n715), .B(n714), .Z(n711) );
  XOR U830 ( .A(n710), .B(sreg[128]), .Z(n709) );
  XNOR U831 ( .A(n711), .B(n709), .Z(c[128]) );
  NANDN U832 ( .A(n713), .B(n712), .Z(n717) );
  NANDN U833 ( .A(n715), .B(n714), .Z(n716) );
  AND U834 ( .A(n717), .B(n716), .Z(n787) );
  NANDN U835 ( .A(n719), .B(n718), .Z(n723) );
  OR U836 ( .A(n721), .B(n720), .Z(n722) );
  AND U837 ( .A(n723), .B(n722), .Z(n819) );
  NAND U838 ( .A(b[0]), .B(a[17]), .Z(n724) );
  XNOR U839 ( .A(b[1]), .B(n724), .Z(n726) );
  NANDN U840 ( .A(b[0]), .B(a[16]), .Z(n725) );
  NAND U841 ( .A(n726), .B(n725), .Z(n799) );
  NANDN U842 ( .A(n9891), .B(n727), .Z(n729) );
  XOR U843 ( .A(b[13]), .B(a[5]), .Z(n805) );
  NANDN U844 ( .A(n9935), .B(n805), .Z(n728) );
  AND U845 ( .A(n729), .B(n728), .Z(n797) );
  AND U846 ( .A(b[15]), .B(a[1]), .Z(n796) );
  XNOR U847 ( .A(n797), .B(n796), .Z(n798) );
  XNOR U848 ( .A(n799), .B(n798), .Z(n817) );
  NANDN U849 ( .A(n9437), .B(n730), .Z(n732) );
  XOR U850 ( .A(b[5]), .B(a[13]), .Z(n808) );
  NANDN U851 ( .A(n9503), .B(n808), .Z(n731) );
  AND U852 ( .A(n732), .B(n731), .Z(n841) );
  NANDN U853 ( .A(n9588), .B(n733), .Z(n735) );
  XOR U854 ( .A(b[7]), .B(a[11]), .Z(n811) );
  NANDN U855 ( .A(n9639), .B(n811), .Z(n734) );
  AND U856 ( .A(n735), .B(n734), .Z(n839) );
  NANDN U857 ( .A(n736), .B(n9420), .Z(n738) );
  XOR U858 ( .A(b[3]), .B(a[15]), .Z(n814) );
  NANDN U859 ( .A(n9375), .B(n814), .Z(n737) );
  NAND U860 ( .A(n738), .B(n737), .Z(n838) );
  XNOR U861 ( .A(n839), .B(n838), .Z(n840) );
  XOR U862 ( .A(n841), .B(n840), .Z(n818) );
  XOR U863 ( .A(n817), .B(n818), .Z(n820) );
  XOR U864 ( .A(n819), .B(n820), .Z(n791) );
  NANDN U865 ( .A(n740), .B(n739), .Z(n744) );
  NANDN U866 ( .A(n742), .B(n741), .Z(n743) );
  AND U867 ( .A(n744), .B(n743), .Z(n790) );
  XNOR U868 ( .A(n791), .B(n790), .Z(n793) );
  NANDN U869 ( .A(n746), .B(n745), .Z(n750) );
  OR U870 ( .A(n748), .B(n747), .Z(n749) );
  AND U871 ( .A(n750), .B(n749), .Z(n845) );
  NAND U872 ( .A(n751), .B(n9883), .Z(n753) );
  XOR U873 ( .A(b[11]), .B(a[7]), .Z(n823) );
  NANDN U874 ( .A(n9856), .B(n823), .Z(n752) );
  AND U875 ( .A(n753), .B(n752), .Z(n834) );
  NANDN U876 ( .A(n10005), .B(n754), .Z(n756) );
  XOR U877 ( .A(b[15]), .B(a[3]), .Z(n826) );
  NANDN U878 ( .A(n10006), .B(n826), .Z(n755) );
  AND U879 ( .A(n756), .B(n755), .Z(n833) );
  NANDN U880 ( .A(n757), .B(n9803), .Z(n759) );
  XOR U881 ( .A(b[9]), .B(a[9]), .Z(n829) );
  NANDN U882 ( .A(n9758), .B(n829), .Z(n758) );
  NAND U883 ( .A(n759), .B(n758), .Z(n832) );
  XOR U884 ( .A(n833), .B(n832), .Z(n835) );
  XNOR U885 ( .A(n834), .B(n835), .Z(n844) );
  XNOR U886 ( .A(n845), .B(n844), .Z(n846) );
  NANDN U887 ( .A(n761), .B(n760), .Z(n765) );
  NANDN U888 ( .A(n763), .B(n762), .Z(n764) );
  NAND U889 ( .A(n765), .B(n764), .Z(n847) );
  XNOR U890 ( .A(n846), .B(n847), .Z(n792) );
  XOR U891 ( .A(n793), .B(n792), .Z(n852) );
  NANDN U892 ( .A(n767), .B(n766), .Z(n771) );
  NANDN U893 ( .A(n769), .B(n768), .Z(n770) );
  AND U894 ( .A(n771), .B(n770), .Z(n851) );
  NANDN U895 ( .A(n773), .B(n772), .Z(n777) );
  NAND U896 ( .A(n775), .B(n774), .Z(n776) );
  AND U897 ( .A(n777), .B(n776), .Z(n850) );
  XOR U898 ( .A(n851), .B(n850), .Z(n853) );
  XOR U899 ( .A(n852), .B(n853), .Z(n785) );
  NANDN U900 ( .A(n779), .B(n778), .Z(n783) );
  OR U901 ( .A(n781), .B(n780), .Z(n782) );
  AND U902 ( .A(n783), .B(n782), .Z(n784) );
  XNOR U903 ( .A(n785), .B(n784), .Z(n786) );
  XNOR U904 ( .A(n787), .B(n786), .Z(n856) );
  XNOR U905 ( .A(sreg[129]), .B(n856), .Z(n857) );
  XNOR U906 ( .A(n858), .B(n857), .Z(c[129]) );
  NANDN U907 ( .A(n785), .B(n784), .Z(n789) );
  NANDN U908 ( .A(n787), .B(n786), .Z(n788) );
  AND U909 ( .A(n789), .B(n788), .Z(n864) );
  NANDN U910 ( .A(n791), .B(n790), .Z(n795) );
  NAND U911 ( .A(n793), .B(n792), .Z(n794) );
  AND U912 ( .A(n795), .B(n794), .Z(n930) );
  NANDN U913 ( .A(n797), .B(n796), .Z(n801) );
  NANDN U914 ( .A(n799), .B(n798), .Z(n800) );
  AND U915 ( .A(n801), .B(n800), .Z(n896) );
  NAND U916 ( .A(b[0]), .B(a[18]), .Z(n802) );
  XNOR U917 ( .A(b[1]), .B(n802), .Z(n804) );
  NANDN U918 ( .A(b[0]), .B(a[17]), .Z(n803) );
  NAND U919 ( .A(n804), .B(n803), .Z(n876) );
  NANDN U920 ( .A(n9891), .B(n805), .Z(n807) );
  XOR U921 ( .A(b[13]), .B(a[6]), .Z(n882) );
  NANDN U922 ( .A(n9935), .B(n882), .Z(n806) );
  AND U923 ( .A(n807), .B(n806), .Z(n874) );
  AND U924 ( .A(b[15]), .B(a[2]), .Z(n873) );
  XNOR U925 ( .A(n874), .B(n873), .Z(n875) );
  XNOR U926 ( .A(n876), .B(n875), .Z(n894) );
  NANDN U927 ( .A(n9437), .B(n808), .Z(n810) );
  XOR U928 ( .A(b[5]), .B(a[14]), .Z(n885) );
  NANDN U929 ( .A(n9503), .B(n885), .Z(n809) );
  AND U930 ( .A(n810), .B(n809), .Z(n918) );
  NANDN U931 ( .A(n9588), .B(n811), .Z(n813) );
  XOR U932 ( .A(b[7]), .B(a[12]), .Z(n888) );
  NANDN U933 ( .A(n9639), .B(n888), .Z(n812) );
  AND U934 ( .A(n813), .B(n812), .Z(n916) );
  NANDN U935 ( .A(n9374), .B(n814), .Z(n816) );
  XOR U936 ( .A(b[3]), .B(a[16]), .Z(n891) );
  NANDN U937 ( .A(n9375), .B(n891), .Z(n815) );
  NAND U938 ( .A(n816), .B(n815), .Z(n915) );
  XNOR U939 ( .A(n916), .B(n915), .Z(n917) );
  XOR U940 ( .A(n918), .B(n917), .Z(n895) );
  XOR U941 ( .A(n894), .B(n895), .Z(n897) );
  XOR U942 ( .A(n896), .B(n897), .Z(n868) );
  NANDN U943 ( .A(n818), .B(n817), .Z(n822) );
  OR U944 ( .A(n820), .B(n819), .Z(n821) );
  AND U945 ( .A(n822), .B(n821), .Z(n867) );
  XNOR U946 ( .A(n868), .B(n867), .Z(n870) );
  NAND U947 ( .A(n823), .B(n9883), .Z(n825) );
  XOR U948 ( .A(b[11]), .B(a[8]), .Z(n900) );
  NANDN U949 ( .A(n9856), .B(n900), .Z(n824) );
  AND U950 ( .A(n825), .B(n824), .Z(n911) );
  NANDN U951 ( .A(n10005), .B(n826), .Z(n828) );
  XOR U952 ( .A(b[15]), .B(a[4]), .Z(n903) );
  NANDN U953 ( .A(n10006), .B(n903), .Z(n827) );
  AND U954 ( .A(n828), .B(n827), .Z(n910) );
  NANDN U955 ( .A(n9685), .B(n829), .Z(n831) );
  XOR U956 ( .A(b[9]), .B(a[10]), .Z(n906) );
  NANDN U957 ( .A(n9758), .B(n906), .Z(n830) );
  NAND U958 ( .A(n831), .B(n830), .Z(n909) );
  XOR U959 ( .A(n910), .B(n909), .Z(n912) );
  XOR U960 ( .A(n911), .B(n912), .Z(n922) );
  NANDN U961 ( .A(n833), .B(n832), .Z(n837) );
  OR U962 ( .A(n835), .B(n834), .Z(n836) );
  AND U963 ( .A(n837), .B(n836), .Z(n921) );
  XNOR U964 ( .A(n922), .B(n921), .Z(n923) );
  NANDN U965 ( .A(n839), .B(n838), .Z(n843) );
  NANDN U966 ( .A(n841), .B(n840), .Z(n842) );
  NAND U967 ( .A(n843), .B(n842), .Z(n924) );
  XNOR U968 ( .A(n923), .B(n924), .Z(n869) );
  XOR U969 ( .A(n870), .B(n869), .Z(n928) );
  NANDN U970 ( .A(n845), .B(n844), .Z(n849) );
  NANDN U971 ( .A(n847), .B(n846), .Z(n848) );
  AND U972 ( .A(n849), .B(n848), .Z(n927) );
  XNOR U973 ( .A(n928), .B(n927), .Z(n929) );
  XOR U974 ( .A(n930), .B(n929), .Z(n862) );
  NANDN U975 ( .A(n851), .B(n850), .Z(n855) );
  OR U976 ( .A(n853), .B(n852), .Z(n854) );
  AND U977 ( .A(n855), .B(n854), .Z(n861) );
  XNOR U978 ( .A(n862), .B(n861), .Z(n863) );
  XNOR U979 ( .A(n864), .B(n863), .Z(n933) );
  XNOR U980 ( .A(sreg[130]), .B(n933), .Z(n935) );
  NANDN U981 ( .A(sreg[129]), .B(n856), .Z(n860) );
  NAND U982 ( .A(n858), .B(n857), .Z(n859) );
  NAND U983 ( .A(n860), .B(n859), .Z(n934) );
  XNOR U984 ( .A(n935), .B(n934), .Z(c[130]) );
  NANDN U985 ( .A(n862), .B(n861), .Z(n866) );
  NANDN U986 ( .A(n864), .B(n863), .Z(n865) );
  AND U987 ( .A(n866), .B(n865), .Z(n943) );
  NANDN U988 ( .A(n868), .B(n867), .Z(n872) );
  NAND U989 ( .A(n870), .B(n869), .Z(n871) );
  AND U990 ( .A(n872), .B(n871), .Z(n1010) );
  NANDN U991 ( .A(n874), .B(n873), .Z(n878) );
  NANDN U992 ( .A(n876), .B(n875), .Z(n877) );
  AND U993 ( .A(n878), .B(n877), .Z(n976) );
  NAND U994 ( .A(b[0]), .B(a[19]), .Z(n879) );
  XNOR U995 ( .A(b[1]), .B(n879), .Z(n881) );
  NANDN U996 ( .A(b[0]), .B(a[18]), .Z(n880) );
  NAND U997 ( .A(n881), .B(n880), .Z(n956) );
  NANDN U998 ( .A(n9891), .B(n882), .Z(n884) );
  XOR U999 ( .A(b[13]), .B(a[7]), .Z(n962) );
  NANDN U1000 ( .A(n9935), .B(n962), .Z(n883) );
  AND U1001 ( .A(n884), .B(n883), .Z(n954) );
  AND U1002 ( .A(b[15]), .B(a[3]), .Z(n953) );
  XNOR U1003 ( .A(n954), .B(n953), .Z(n955) );
  XNOR U1004 ( .A(n956), .B(n955), .Z(n974) );
  NANDN U1005 ( .A(n9437), .B(n885), .Z(n887) );
  XOR U1006 ( .A(b[5]), .B(a[15]), .Z(n965) );
  NANDN U1007 ( .A(n9503), .B(n965), .Z(n886) );
  AND U1008 ( .A(n887), .B(n886), .Z(n998) );
  NANDN U1009 ( .A(n9588), .B(n888), .Z(n890) );
  XOR U1010 ( .A(b[7]), .B(a[13]), .Z(n968) );
  NANDN U1011 ( .A(n9639), .B(n968), .Z(n889) );
  AND U1012 ( .A(n890), .B(n889), .Z(n996) );
  NANDN U1013 ( .A(n9374), .B(n891), .Z(n893) );
  XOR U1014 ( .A(b[3]), .B(a[17]), .Z(n971) );
  NANDN U1015 ( .A(n9375), .B(n971), .Z(n892) );
  NAND U1016 ( .A(n893), .B(n892), .Z(n995) );
  XNOR U1017 ( .A(n996), .B(n995), .Z(n997) );
  XOR U1018 ( .A(n998), .B(n997), .Z(n975) );
  XOR U1019 ( .A(n974), .B(n975), .Z(n977) );
  XOR U1020 ( .A(n976), .B(n977), .Z(n948) );
  NANDN U1021 ( .A(n895), .B(n894), .Z(n899) );
  OR U1022 ( .A(n897), .B(n896), .Z(n898) );
  AND U1023 ( .A(n899), .B(n898), .Z(n947) );
  XNOR U1024 ( .A(n948), .B(n947), .Z(n950) );
  NAND U1025 ( .A(n900), .B(n9883), .Z(n902) );
  XOR U1026 ( .A(b[11]), .B(a[9]), .Z(n980) );
  NANDN U1027 ( .A(n9856), .B(n980), .Z(n901) );
  AND U1028 ( .A(n902), .B(n901), .Z(n991) );
  NANDN U1029 ( .A(n10005), .B(n903), .Z(n905) );
  XOR U1030 ( .A(b[15]), .B(a[5]), .Z(n983) );
  NANDN U1031 ( .A(n10006), .B(n983), .Z(n904) );
  AND U1032 ( .A(n905), .B(n904), .Z(n990) );
  NANDN U1033 ( .A(n9685), .B(n906), .Z(n908) );
  XOR U1034 ( .A(b[9]), .B(a[11]), .Z(n986) );
  NANDN U1035 ( .A(n9758), .B(n986), .Z(n907) );
  NAND U1036 ( .A(n908), .B(n907), .Z(n989) );
  XOR U1037 ( .A(n990), .B(n989), .Z(n992) );
  XOR U1038 ( .A(n991), .B(n992), .Z(n1002) );
  NANDN U1039 ( .A(n910), .B(n909), .Z(n914) );
  OR U1040 ( .A(n912), .B(n911), .Z(n913) );
  AND U1041 ( .A(n914), .B(n913), .Z(n1001) );
  XNOR U1042 ( .A(n1002), .B(n1001), .Z(n1003) );
  NANDN U1043 ( .A(n916), .B(n915), .Z(n920) );
  NANDN U1044 ( .A(n918), .B(n917), .Z(n919) );
  NAND U1045 ( .A(n920), .B(n919), .Z(n1004) );
  XNOR U1046 ( .A(n1003), .B(n1004), .Z(n949) );
  XOR U1047 ( .A(n950), .B(n949), .Z(n1008) );
  NANDN U1048 ( .A(n922), .B(n921), .Z(n926) );
  NANDN U1049 ( .A(n924), .B(n923), .Z(n925) );
  AND U1050 ( .A(n926), .B(n925), .Z(n1007) );
  XNOR U1051 ( .A(n1008), .B(n1007), .Z(n1009) );
  XOR U1052 ( .A(n1010), .B(n1009), .Z(n942) );
  NANDN U1053 ( .A(n928), .B(n927), .Z(n932) );
  NAND U1054 ( .A(n930), .B(n929), .Z(n931) );
  AND U1055 ( .A(n932), .B(n931), .Z(n941) );
  XOR U1056 ( .A(n942), .B(n941), .Z(n944) );
  XOR U1057 ( .A(n943), .B(n944), .Z(n939) );
  NANDN U1058 ( .A(sreg[130]), .B(n933), .Z(n937) );
  NAND U1059 ( .A(n935), .B(n934), .Z(n936) );
  AND U1060 ( .A(n937), .B(n936), .Z(n940) );
  XNOR U1061 ( .A(sreg[131]), .B(n940), .Z(n938) );
  XOR U1062 ( .A(n939), .B(n938), .Z(c[131]) );
  NANDN U1063 ( .A(n942), .B(n941), .Z(n946) );
  OR U1064 ( .A(n944), .B(n943), .Z(n945) );
  AND U1065 ( .A(n946), .B(n945), .Z(n1016) );
  NANDN U1066 ( .A(n948), .B(n947), .Z(n952) );
  NAND U1067 ( .A(n950), .B(n949), .Z(n951) );
  AND U1068 ( .A(n952), .B(n951), .Z(n1082) );
  NANDN U1069 ( .A(n954), .B(n953), .Z(n958) );
  NANDN U1070 ( .A(n956), .B(n955), .Z(n957) );
  AND U1071 ( .A(n958), .B(n957), .Z(n1048) );
  NAND U1072 ( .A(b[0]), .B(a[20]), .Z(n959) );
  XNOR U1073 ( .A(b[1]), .B(n959), .Z(n961) );
  NANDN U1074 ( .A(b[0]), .B(a[19]), .Z(n960) );
  NAND U1075 ( .A(n961), .B(n960), .Z(n1028) );
  NANDN U1076 ( .A(n9891), .B(n962), .Z(n964) );
  XOR U1077 ( .A(b[13]), .B(a[8]), .Z(n1031) );
  NANDN U1078 ( .A(n9935), .B(n1031), .Z(n963) );
  AND U1079 ( .A(n964), .B(n963), .Z(n1026) );
  AND U1080 ( .A(b[15]), .B(a[4]), .Z(n1025) );
  XNOR U1081 ( .A(n1026), .B(n1025), .Z(n1027) );
  XNOR U1082 ( .A(n1028), .B(n1027), .Z(n1046) );
  NANDN U1083 ( .A(n9437), .B(n965), .Z(n967) );
  XOR U1084 ( .A(b[5]), .B(a[16]), .Z(n1037) );
  NANDN U1085 ( .A(n9503), .B(n1037), .Z(n966) );
  AND U1086 ( .A(n967), .B(n966), .Z(n1070) );
  NANDN U1087 ( .A(n9588), .B(n968), .Z(n970) );
  XOR U1088 ( .A(b[7]), .B(a[14]), .Z(n1040) );
  NANDN U1089 ( .A(n9639), .B(n1040), .Z(n969) );
  AND U1090 ( .A(n970), .B(n969), .Z(n1068) );
  NANDN U1091 ( .A(n9374), .B(n971), .Z(n973) );
  XOR U1092 ( .A(b[3]), .B(a[18]), .Z(n1043) );
  NANDN U1093 ( .A(n9375), .B(n1043), .Z(n972) );
  NAND U1094 ( .A(n973), .B(n972), .Z(n1067) );
  XNOR U1095 ( .A(n1068), .B(n1067), .Z(n1069) );
  XOR U1096 ( .A(n1070), .B(n1069), .Z(n1047) );
  XOR U1097 ( .A(n1046), .B(n1047), .Z(n1049) );
  XOR U1098 ( .A(n1048), .B(n1049), .Z(n1020) );
  NANDN U1099 ( .A(n975), .B(n974), .Z(n979) );
  OR U1100 ( .A(n977), .B(n976), .Z(n978) );
  AND U1101 ( .A(n979), .B(n978), .Z(n1019) );
  XNOR U1102 ( .A(n1020), .B(n1019), .Z(n1022) );
  NAND U1103 ( .A(n980), .B(n9883), .Z(n982) );
  XOR U1104 ( .A(b[11]), .B(a[10]), .Z(n1052) );
  NANDN U1105 ( .A(n9856), .B(n1052), .Z(n981) );
  AND U1106 ( .A(n982), .B(n981), .Z(n1063) );
  NANDN U1107 ( .A(n10005), .B(n983), .Z(n985) );
  XOR U1108 ( .A(b[15]), .B(a[6]), .Z(n1055) );
  NANDN U1109 ( .A(n10006), .B(n1055), .Z(n984) );
  AND U1110 ( .A(n985), .B(n984), .Z(n1062) );
  NANDN U1111 ( .A(n9685), .B(n986), .Z(n988) );
  XOR U1112 ( .A(b[9]), .B(a[12]), .Z(n1058) );
  NANDN U1113 ( .A(n9758), .B(n1058), .Z(n987) );
  NAND U1114 ( .A(n988), .B(n987), .Z(n1061) );
  XOR U1115 ( .A(n1062), .B(n1061), .Z(n1064) );
  XOR U1116 ( .A(n1063), .B(n1064), .Z(n1074) );
  NANDN U1117 ( .A(n990), .B(n989), .Z(n994) );
  OR U1118 ( .A(n992), .B(n991), .Z(n993) );
  AND U1119 ( .A(n994), .B(n993), .Z(n1073) );
  XNOR U1120 ( .A(n1074), .B(n1073), .Z(n1075) );
  NANDN U1121 ( .A(n996), .B(n995), .Z(n1000) );
  NANDN U1122 ( .A(n998), .B(n997), .Z(n999) );
  NAND U1123 ( .A(n1000), .B(n999), .Z(n1076) );
  XNOR U1124 ( .A(n1075), .B(n1076), .Z(n1021) );
  XOR U1125 ( .A(n1022), .B(n1021), .Z(n1080) );
  NANDN U1126 ( .A(n1002), .B(n1001), .Z(n1006) );
  NANDN U1127 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U1128 ( .A(n1006), .B(n1005), .Z(n1079) );
  XNOR U1129 ( .A(n1080), .B(n1079), .Z(n1081) );
  XOR U1130 ( .A(n1082), .B(n1081), .Z(n1014) );
  NANDN U1131 ( .A(n1008), .B(n1007), .Z(n1012) );
  NAND U1132 ( .A(n1010), .B(n1009), .Z(n1011) );
  AND U1133 ( .A(n1012), .B(n1011), .Z(n1013) );
  XNOR U1134 ( .A(n1014), .B(n1013), .Z(n1015) );
  XNOR U1135 ( .A(n1016), .B(n1015), .Z(n1085) );
  XNOR U1136 ( .A(sreg[132]), .B(n1085), .Z(n1086) );
  XOR U1137 ( .A(n1087), .B(n1086), .Z(c[132]) );
  NANDN U1138 ( .A(n1014), .B(n1013), .Z(n1018) );
  NANDN U1139 ( .A(n1016), .B(n1015), .Z(n1017) );
  AND U1140 ( .A(n1018), .B(n1017), .Z(n1093) );
  NANDN U1141 ( .A(n1020), .B(n1019), .Z(n1024) );
  NAND U1142 ( .A(n1022), .B(n1021), .Z(n1023) );
  AND U1143 ( .A(n1024), .B(n1023), .Z(n1159) );
  NANDN U1144 ( .A(n1026), .B(n1025), .Z(n1030) );
  NANDN U1145 ( .A(n1028), .B(n1027), .Z(n1029) );
  AND U1146 ( .A(n1030), .B(n1029), .Z(n1125) );
  NANDN U1147 ( .A(n9891), .B(n1031), .Z(n1033) );
  XOR U1148 ( .A(b[13]), .B(a[9]), .Z(n1111) );
  NANDN U1149 ( .A(n9935), .B(n1111), .Z(n1032) );
  AND U1150 ( .A(n1033), .B(n1032), .Z(n1103) );
  AND U1151 ( .A(b[15]), .B(a[5]), .Z(n1102) );
  XNOR U1152 ( .A(n1103), .B(n1102), .Z(n1104) );
  NAND U1153 ( .A(b[0]), .B(a[21]), .Z(n1034) );
  XNOR U1154 ( .A(b[1]), .B(n1034), .Z(n1036) );
  NANDN U1155 ( .A(b[0]), .B(a[20]), .Z(n1035) );
  NAND U1156 ( .A(n1036), .B(n1035), .Z(n1105) );
  XNOR U1157 ( .A(n1104), .B(n1105), .Z(n1123) );
  NANDN U1158 ( .A(n9437), .B(n1037), .Z(n1039) );
  XOR U1159 ( .A(b[5]), .B(a[17]), .Z(n1114) );
  NANDN U1160 ( .A(n9503), .B(n1114), .Z(n1038) );
  AND U1161 ( .A(n1039), .B(n1038), .Z(n1147) );
  NANDN U1162 ( .A(n9588), .B(n1040), .Z(n1042) );
  XOR U1163 ( .A(b[7]), .B(a[15]), .Z(n1117) );
  NANDN U1164 ( .A(n9639), .B(n1117), .Z(n1041) );
  AND U1165 ( .A(n1042), .B(n1041), .Z(n1145) );
  NANDN U1166 ( .A(n9374), .B(n1043), .Z(n1045) );
  XOR U1167 ( .A(b[3]), .B(a[19]), .Z(n1120) );
  NANDN U1168 ( .A(n9375), .B(n1120), .Z(n1044) );
  NAND U1169 ( .A(n1045), .B(n1044), .Z(n1144) );
  XNOR U1170 ( .A(n1145), .B(n1144), .Z(n1146) );
  XOR U1171 ( .A(n1147), .B(n1146), .Z(n1124) );
  XOR U1172 ( .A(n1123), .B(n1124), .Z(n1126) );
  XOR U1173 ( .A(n1125), .B(n1126), .Z(n1097) );
  NANDN U1174 ( .A(n1047), .B(n1046), .Z(n1051) );
  OR U1175 ( .A(n1049), .B(n1048), .Z(n1050) );
  AND U1176 ( .A(n1051), .B(n1050), .Z(n1096) );
  XNOR U1177 ( .A(n1097), .B(n1096), .Z(n1099) );
  NAND U1178 ( .A(n1052), .B(n9883), .Z(n1054) );
  XOR U1179 ( .A(b[11]), .B(a[11]), .Z(n1129) );
  NANDN U1180 ( .A(n9856), .B(n1129), .Z(n1053) );
  AND U1181 ( .A(n1054), .B(n1053), .Z(n1140) );
  NANDN U1182 ( .A(n10005), .B(n1055), .Z(n1057) );
  XOR U1183 ( .A(b[15]), .B(a[7]), .Z(n1132) );
  NANDN U1184 ( .A(n10006), .B(n1132), .Z(n1056) );
  AND U1185 ( .A(n1057), .B(n1056), .Z(n1139) );
  NANDN U1186 ( .A(n9685), .B(n1058), .Z(n1060) );
  XOR U1187 ( .A(b[9]), .B(a[13]), .Z(n1135) );
  NANDN U1188 ( .A(n9758), .B(n1135), .Z(n1059) );
  NAND U1189 ( .A(n1060), .B(n1059), .Z(n1138) );
  XOR U1190 ( .A(n1139), .B(n1138), .Z(n1141) );
  XOR U1191 ( .A(n1140), .B(n1141), .Z(n1151) );
  NANDN U1192 ( .A(n1062), .B(n1061), .Z(n1066) );
  OR U1193 ( .A(n1064), .B(n1063), .Z(n1065) );
  AND U1194 ( .A(n1066), .B(n1065), .Z(n1150) );
  XNOR U1195 ( .A(n1151), .B(n1150), .Z(n1152) );
  NANDN U1196 ( .A(n1068), .B(n1067), .Z(n1072) );
  NANDN U1197 ( .A(n1070), .B(n1069), .Z(n1071) );
  NAND U1198 ( .A(n1072), .B(n1071), .Z(n1153) );
  XNOR U1199 ( .A(n1152), .B(n1153), .Z(n1098) );
  XOR U1200 ( .A(n1099), .B(n1098), .Z(n1157) );
  NANDN U1201 ( .A(n1074), .B(n1073), .Z(n1078) );
  NANDN U1202 ( .A(n1076), .B(n1075), .Z(n1077) );
  AND U1203 ( .A(n1078), .B(n1077), .Z(n1156) );
  XNOR U1204 ( .A(n1157), .B(n1156), .Z(n1158) );
  XOR U1205 ( .A(n1159), .B(n1158), .Z(n1091) );
  NANDN U1206 ( .A(n1080), .B(n1079), .Z(n1084) );
  NAND U1207 ( .A(n1082), .B(n1081), .Z(n1083) );
  AND U1208 ( .A(n1084), .B(n1083), .Z(n1090) );
  XNOR U1209 ( .A(n1091), .B(n1090), .Z(n1092) );
  XNOR U1210 ( .A(n1093), .B(n1092), .Z(n1162) );
  XNOR U1211 ( .A(sreg[133]), .B(n1162), .Z(n1164) );
  NANDN U1212 ( .A(sreg[132]), .B(n1085), .Z(n1089) );
  NANDN U1213 ( .A(n1087), .B(n1086), .Z(n1088) );
  NAND U1214 ( .A(n1089), .B(n1088), .Z(n1163) );
  XNOR U1215 ( .A(n1164), .B(n1163), .Z(c[133]) );
  NANDN U1216 ( .A(n1091), .B(n1090), .Z(n1095) );
  NANDN U1217 ( .A(n1093), .B(n1092), .Z(n1094) );
  AND U1218 ( .A(n1095), .B(n1094), .Z(n1170) );
  NANDN U1219 ( .A(n1097), .B(n1096), .Z(n1101) );
  NAND U1220 ( .A(n1099), .B(n1098), .Z(n1100) );
  AND U1221 ( .A(n1101), .B(n1100), .Z(n1236) );
  NANDN U1222 ( .A(n1103), .B(n1102), .Z(n1107) );
  NANDN U1223 ( .A(n1105), .B(n1104), .Z(n1106) );
  AND U1224 ( .A(n1107), .B(n1106), .Z(n1202) );
  NAND U1225 ( .A(b[0]), .B(a[22]), .Z(n1108) );
  XNOR U1226 ( .A(b[1]), .B(n1108), .Z(n1110) );
  NANDN U1227 ( .A(b[0]), .B(a[21]), .Z(n1109) );
  NAND U1228 ( .A(n1110), .B(n1109), .Z(n1182) );
  NANDN U1229 ( .A(n9891), .B(n1111), .Z(n1113) );
  XOR U1230 ( .A(b[13]), .B(a[10]), .Z(n1188) );
  NANDN U1231 ( .A(n9935), .B(n1188), .Z(n1112) );
  AND U1232 ( .A(n1113), .B(n1112), .Z(n1180) );
  AND U1233 ( .A(b[15]), .B(a[6]), .Z(n1179) );
  XNOR U1234 ( .A(n1180), .B(n1179), .Z(n1181) );
  XNOR U1235 ( .A(n1182), .B(n1181), .Z(n1200) );
  NANDN U1236 ( .A(n9437), .B(n1114), .Z(n1116) );
  XOR U1237 ( .A(b[5]), .B(a[18]), .Z(n1191) );
  NANDN U1238 ( .A(n9503), .B(n1191), .Z(n1115) );
  AND U1239 ( .A(n1116), .B(n1115), .Z(n1224) );
  NANDN U1240 ( .A(n9588), .B(n1117), .Z(n1119) );
  XOR U1241 ( .A(b[7]), .B(a[16]), .Z(n1194) );
  NANDN U1242 ( .A(n9639), .B(n1194), .Z(n1118) );
  AND U1243 ( .A(n1119), .B(n1118), .Z(n1222) );
  NANDN U1244 ( .A(n9374), .B(n1120), .Z(n1122) );
  XOR U1245 ( .A(b[3]), .B(a[20]), .Z(n1197) );
  NANDN U1246 ( .A(n9375), .B(n1197), .Z(n1121) );
  NAND U1247 ( .A(n1122), .B(n1121), .Z(n1221) );
  XNOR U1248 ( .A(n1222), .B(n1221), .Z(n1223) );
  XOR U1249 ( .A(n1224), .B(n1223), .Z(n1201) );
  XOR U1250 ( .A(n1200), .B(n1201), .Z(n1203) );
  XOR U1251 ( .A(n1202), .B(n1203), .Z(n1174) );
  NANDN U1252 ( .A(n1124), .B(n1123), .Z(n1128) );
  OR U1253 ( .A(n1126), .B(n1125), .Z(n1127) );
  AND U1254 ( .A(n1128), .B(n1127), .Z(n1173) );
  XNOR U1255 ( .A(n1174), .B(n1173), .Z(n1176) );
  NAND U1256 ( .A(n1129), .B(n9883), .Z(n1131) );
  XOR U1257 ( .A(b[11]), .B(a[12]), .Z(n1206) );
  NANDN U1258 ( .A(n9856), .B(n1206), .Z(n1130) );
  AND U1259 ( .A(n1131), .B(n1130), .Z(n1217) );
  NANDN U1260 ( .A(n10005), .B(n1132), .Z(n1134) );
  XOR U1261 ( .A(b[15]), .B(a[8]), .Z(n1209) );
  NANDN U1262 ( .A(n10006), .B(n1209), .Z(n1133) );
  AND U1263 ( .A(n1134), .B(n1133), .Z(n1216) );
  NANDN U1264 ( .A(n9685), .B(n1135), .Z(n1137) );
  XOR U1265 ( .A(b[9]), .B(a[14]), .Z(n1212) );
  NANDN U1266 ( .A(n9758), .B(n1212), .Z(n1136) );
  NAND U1267 ( .A(n1137), .B(n1136), .Z(n1215) );
  XOR U1268 ( .A(n1216), .B(n1215), .Z(n1218) );
  XOR U1269 ( .A(n1217), .B(n1218), .Z(n1228) );
  NANDN U1270 ( .A(n1139), .B(n1138), .Z(n1143) );
  OR U1271 ( .A(n1141), .B(n1140), .Z(n1142) );
  AND U1272 ( .A(n1143), .B(n1142), .Z(n1227) );
  XNOR U1273 ( .A(n1228), .B(n1227), .Z(n1229) );
  NANDN U1274 ( .A(n1145), .B(n1144), .Z(n1149) );
  NANDN U1275 ( .A(n1147), .B(n1146), .Z(n1148) );
  NAND U1276 ( .A(n1149), .B(n1148), .Z(n1230) );
  XNOR U1277 ( .A(n1229), .B(n1230), .Z(n1175) );
  XOR U1278 ( .A(n1176), .B(n1175), .Z(n1234) );
  NANDN U1279 ( .A(n1151), .B(n1150), .Z(n1155) );
  NANDN U1280 ( .A(n1153), .B(n1152), .Z(n1154) );
  AND U1281 ( .A(n1155), .B(n1154), .Z(n1233) );
  XNOR U1282 ( .A(n1234), .B(n1233), .Z(n1235) );
  XOR U1283 ( .A(n1236), .B(n1235), .Z(n1168) );
  NANDN U1284 ( .A(n1157), .B(n1156), .Z(n1161) );
  NAND U1285 ( .A(n1159), .B(n1158), .Z(n1160) );
  AND U1286 ( .A(n1161), .B(n1160), .Z(n1167) );
  XNOR U1287 ( .A(n1168), .B(n1167), .Z(n1169) );
  XNOR U1288 ( .A(n1170), .B(n1169), .Z(n1239) );
  XNOR U1289 ( .A(sreg[134]), .B(n1239), .Z(n1241) );
  NANDN U1290 ( .A(sreg[133]), .B(n1162), .Z(n1166) );
  NAND U1291 ( .A(n1164), .B(n1163), .Z(n1165) );
  NAND U1292 ( .A(n1166), .B(n1165), .Z(n1240) );
  XNOR U1293 ( .A(n1241), .B(n1240), .Z(c[134]) );
  NANDN U1294 ( .A(n1168), .B(n1167), .Z(n1172) );
  NANDN U1295 ( .A(n1170), .B(n1169), .Z(n1171) );
  AND U1296 ( .A(n1172), .B(n1171), .Z(n1247) );
  NANDN U1297 ( .A(n1174), .B(n1173), .Z(n1178) );
  NAND U1298 ( .A(n1176), .B(n1175), .Z(n1177) );
  AND U1299 ( .A(n1178), .B(n1177), .Z(n1313) );
  NANDN U1300 ( .A(n1180), .B(n1179), .Z(n1184) );
  NANDN U1301 ( .A(n1182), .B(n1181), .Z(n1183) );
  AND U1302 ( .A(n1184), .B(n1183), .Z(n1279) );
  NAND U1303 ( .A(b[0]), .B(a[23]), .Z(n1185) );
  XNOR U1304 ( .A(b[1]), .B(n1185), .Z(n1187) );
  NANDN U1305 ( .A(b[0]), .B(a[22]), .Z(n1186) );
  NAND U1306 ( .A(n1187), .B(n1186), .Z(n1259) );
  NANDN U1307 ( .A(n9891), .B(n1188), .Z(n1190) );
  XOR U1308 ( .A(b[13]), .B(a[11]), .Z(n1265) );
  NANDN U1309 ( .A(n9935), .B(n1265), .Z(n1189) );
  AND U1310 ( .A(n1190), .B(n1189), .Z(n1257) );
  AND U1311 ( .A(b[15]), .B(a[7]), .Z(n1256) );
  XNOR U1312 ( .A(n1257), .B(n1256), .Z(n1258) );
  XNOR U1313 ( .A(n1259), .B(n1258), .Z(n1277) );
  NANDN U1314 ( .A(n9437), .B(n1191), .Z(n1193) );
  XOR U1315 ( .A(b[5]), .B(a[19]), .Z(n1268) );
  NANDN U1316 ( .A(n9503), .B(n1268), .Z(n1192) );
  AND U1317 ( .A(n1193), .B(n1192), .Z(n1301) );
  NANDN U1318 ( .A(n9588), .B(n1194), .Z(n1196) );
  XOR U1319 ( .A(b[7]), .B(a[17]), .Z(n1271) );
  NANDN U1320 ( .A(n9639), .B(n1271), .Z(n1195) );
  AND U1321 ( .A(n1196), .B(n1195), .Z(n1299) );
  NANDN U1322 ( .A(n9374), .B(n1197), .Z(n1199) );
  XOR U1323 ( .A(b[3]), .B(a[21]), .Z(n1274) );
  NANDN U1324 ( .A(n9375), .B(n1274), .Z(n1198) );
  NAND U1325 ( .A(n1199), .B(n1198), .Z(n1298) );
  XNOR U1326 ( .A(n1299), .B(n1298), .Z(n1300) );
  XOR U1327 ( .A(n1301), .B(n1300), .Z(n1278) );
  XOR U1328 ( .A(n1277), .B(n1278), .Z(n1280) );
  XOR U1329 ( .A(n1279), .B(n1280), .Z(n1251) );
  NANDN U1330 ( .A(n1201), .B(n1200), .Z(n1205) );
  OR U1331 ( .A(n1203), .B(n1202), .Z(n1204) );
  AND U1332 ( .A(n1205), .B(n1204), .Z(n1250) );
  XNOR U1333 ( .A(n1251), .B(n1250), .Z(n1253) );
  NAND U1334 ( .A(n1206), .B(n9883), .Z(n1208) );
  XOR U1335 ( .A(b[11]), .B(a[13]), .Z(n1283) );
  NANDN U1336 ( .A(n9856), .B(n1283), .Z(n1207) );
  AND U1337 ( .A(n1208), .B(n1207), .Z(n1294) );
  NANDN U1338 ( .A(n10005), .B(n1209), .Z(n1211) );
  XOR U1339 ( .A(b[15]), .B(a[9]), .Z(n1286) );
  NANDN U1340 ( .A(n10006), .B(n1286), .Z(n1210) );
  AND U1341 ( .A(n1211), .B(n1210), .Z(n1293) );
  NANDN U1342 ( .A(n9685), .B(n1212), .Z(n1214) );
  XOR U1343 ( .A(b[9]), .B(a[15]), .Z(n1289) );
  NANDN U1344 ( .A(n9758), .B(n1289), .Z(n1213) );
  NAND U1345 ( .A(n1214), .B(n1213), .Z(n1292) );
  XOR U1346 ( .A(n1293), .B(n1292), .Z(n1295) );
  XOR U1347 ( .A(n1294), .B(n1295), .Z(n1305) );
  NANDN U1348 ( .A(n1216), .B(n1215), .Z(n1220) );
  OR U1349 ( .A(n1218), .B(n1217), .Z(n1219) );
  AND U1350 ( .A(n1220), .B(n1219), .Z(n1304) );
  XNOR U1351 ( .A(n1305), .B(n1304), .Z(n1306) );
  NANDN U1352 ( .A(n1222), .B(n1221), .Z(n1226) );
  NANDN U1353 ( .A(n1224), .B(n1223), .Z(n1225) );
  NAND U1354 ( .A(n1226), .B(n1225), .Z(n1307) );
  XNOR U1355 ( .A(n1306), .B(n1307), .Z(n1252) );
  XOR U1356 ( .A(n1253), .B(n1252), .Z(n1311) );
  NANDN U1357 ( .A(n1228), .B(n1227), .Z(n1232) );
  NANDN U1358 ( .A(n1230), .B(n1229), .Z(n1231) );
  AND U1359 ( .A(n1232), .B(n1231), .Z(n1310) );
  XNOR U1360 ( .A(n1311), .B(n1310), .Z(n1312) );
  XOR U1361 ( .A(n1313), .B(n1312), .Z(n1245) );
  NANDN U1362 ( .A(n1234), .B(n1233), .Z(n1238) );
  NAND U1363 ( .A(n1236), .B(n1235), .Z(n1237) );
  AND U1364 ( .A(n1238), .B(n1237), .Z(n1244) );
  XNOR U1365 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U1366 ( .A(n1247), .B(n1246), .Z(n1316) );
  XNOR U1367 ( .A(sreg[135]), .B(n1316), .Z(n1318) );
  NANDN U1368 ( .A(sreg[134]), .B(n1239), .Z(n1243) );
  NAND U1369 ( .A(n1241), .B(n1240), .Z(n1242) );
  NAND U1370 ( .A(n1243), .B(n1242), .Z(n1317) );
  XNOR U1371 ( .A(n1318), .B(n1317), .Z(c[135]) );
  NANDN U1372 ( .A(n1245), .B(n1244), .Z(n1249) );
  NANDN U1373 ( .A(n1247), .B(n1246), .Z(n1248) );
  AND U1374 ( .A(n1249), .B(n1248), .Z(n1324) );
  NANDN U1375 ( .A(n1251), .B(n1250), .Z(n1255) );
  NAND U1376 ( .A(n1253), .B(n1252), .Z(n1254) );
  AND U1377 ( .A(n1255), .B(n1254), .Z(n1390) );
  NANDN U1378 ( .A(n1257), .B(n1256), .Z(n1261) );
  NANDN U1379 ( .A(n1259), .B(n1258), .Z(n1260) );
  AND U1380 ( .A(n1261), .B(n1260), .Z(n1356) );
  NAND U1381 ( .A(b[0]), .B(a[24]), .Z(n1262) );
  XNOR U1382 ( .A(b[1]), .B(n1262), .Z(n1264) );
  NANDN U1383 ( .A(b[0]), .B(a[23]), .Z(n1263) );
  NAND U1384 ( .A(n1264), .B(n1263), .Z(n1336) );
  NANDN U1385 ( .A(n9891), .B(n1265), .Z(n1267) );
  XOR U1386 ( .A(b[13]), .B(a[12]), .Z(n1342) );
  NANDN U1387 ( .A(n9935), .B(n1342), .Z(n1266) );
  AND U1388 ( .A(n1267), .B(n1266), .Z(n1334) );
  AND U1389 ( .A(b[15]), .B(a[8]), .Z(n1333) );
  XNOR U1390 ( .A(n1334), .B(n1333), .Z(n1335) );
  XNOR U1391 ( .A(n1336), .B(n1335), .Z(n1354) );
  NANDN U1392 ( .A(n9437), .B(n1268), .Z(n1270) );
  XOR U1393 ( .A(b[5]), .B(a[20]), .Z(n1345) );
  NANDN U1394 ( .A(n9503), .B(n1345), .Z(n1269) );
  AND U1395 ( .A(n1270), .B(n1269), .Z(n1378) );
  NANDN U1396 ( .A(n9588), .B(n1271), .Z(n1273) );
  XOR U1397 ( .A(b[7]), .B(a[18]), .Z(n1348) );
  NANDN U1398 ( .A(n9639), .B(n1348), .Z(n1272) );
  AND U1399 ( .A(n1273), .B(n1272), .Z(n1376) );
  NANDN U1400 ( .A(n9374), .B(n1274), .Z(n1276) );
  XOR U1401 ( .A(b[3]), .B(a[22]), .Z(n1351) );
  NANDN U1402 ( .A(n9375), .B(n1351), .Z(n1275) );
  NAND U1403 ( .A(n1276), .B(n1275), .Z(n1375) );
  XNOR U1404 ( .A(n1376), .B(n1375), .Z(n1377) );
  XOR U1405 ( .A(n1378), .B(n1377), .Z(n1355) );
  XOR U1406 ( .A(n1354), .B(n1355), .Z(n1357) );
  XOR U1407 ( .A(n1356), .B(n1357), .Z(n1328) );
  NANDN U1408 ( .A(n1278), .B(n1277), .Z(n1282) );
  OR U1409 ( .A(n1280), .B(n1279), .Z(n1281) );
  AND U1410 ( .A(n1282), .B(n1281), .Z(n1327) );
  XNOR U1411 ( .A(n1328), .B(n1327), .Z(n1330) );
  NAND U1412 ( .A(n1283), .B(n9883), .Z(n1285) );
  XOR U1413 ( .A(b[11]), .B(a[14]), .Z(n1360) );
  NANDN U1414 ( .A(n9856), .B(n1360), .Z(n1284) );
  AND U1415 ( .A(n1285), .B(n1284), .Z(n1371) );
  NANDN U1416 ( .A(n10005), .B(n1286), .Z(n1288) );
  XOR U1417 ( .A(b[15]), .B(a[10]), .Z(n1363) );
  NANDN U1418 ( .A(n10006), .B(n1363), .Z(n1287) );
  AND U1419 ( .A(n1288), .B(n1287), .Z(n1370) );
  NANDN U1420 ( .A(n9685), .B(n1289), .Z(n1291) );
  XOR U1421 ( .A(b[9]), .B(a[16]), .Z(n1366) );
  NANDN U1422 ( .A(n9758), .B(n1366), .Z(n1290) );
  NAND U1423 ( .A(n1291), .B(n1290), .Z(n1369) );
  XOR U1424 ( .A(n1370), .B(n1369), .Z(n1372) );
  XOR U1425 ( .A(n1371), .B(n1372), .Z(n1382) );
  NANDN U1426 ( .A(n1293), .B(n1292), .Z(n1297) );
  OR U1427 ( .A(n1295), .B(n1294), .Z(n1296) );
  AND U1428 ( .A(n1297), .B(n1296), .Z(n1381) );
  XNOR U1429 ( .A(n1382), .B(n1381), .Z(n1383) );
  NANDN U1430 ( .A(n1299), .B(n1298), .Z(n1303) );
  NANDN U1431 ( .A(n1301), .B(n1300), .Z(n1302) );
  NAND U1432 ( .A(n1303), .B(n1302), .Z(n1384) );
  XNOR U1433 ( .A(n1383), .B(n1384), .Z(n1329) );
  XOR U1434 ( .A(n1330), .B(n1329), .Z(n1388) );
  NANDN U1435 ( .A(n1305), .B(n1304), .Z(n1309) );
  NANDN U1436 ( .A(n1307), .B(n1306), .Z(n1308) );
  AND U1437 ( .A(n1309), .B(n1308), .Z(n1387) );
  XNOR U1438 ( .A(n1388), .B(n1387), .Z(n1389) );
  XOR U1439 ( .A(n1390), .B(n1389), .Z(n1322) );
  NANDN U1440 ( .A(n1311), .B(n1310), .Z(n1315) );
  NAND U1441 ( .A(n1313), .B(n1312), .Z(n1314) );
  AND U1442 ( .A(n1315), .B(n1314), .Z(n1321) );
  XNOR U1443 ( .A(n1322), .B(n1321), .Z(n1323) );
  XNOR U1444 ( .A(n1324), .B(n1323), .Z(n1393) );
  XNOR U1445 ( .A(sreg[136]), .B(n1393), .Z(n1395) );
  NANDN U1446 ( .A(sreg[135]), .B(n1316), .Z(n1320) );
  NAND U1447 ( .A(n1318), .B(n1317), .Z(n1319) );
  NAND U1448 ( .A(n1320), .B(n1319), .Z(n1394) );
  XNOR U1449 ( .A(n1395), .B(n1394), .Z(c[136]) );
  NANDN U1450 ( .A(n1322), .B(n1321), .Z(n1326) );
  NANDN U1451 ( .A(n1324), .B(n1323), .Z(n1325) );
  AND U1452 ( .A(n1326), .B(n1325), .Z(n1401) );
  NANDN U1453 ( .A(n1328), .B(n1327), .Z(n1332) );
  NAND U1454 ( .A(n1330), .B(n1329), .Z(n1331) );
  AND U1455 ( .A(n1332), .B(n1331), .Z(n1467) );
  NANDN U1456 ( .A(n1334), .B(n1333), .Z(n1338) );
  NANDN U1457 ( .A(n1336), .B(n1335), .Z(n1337) );
  AND U1458 ( .A(n1338), .B(n1337), .Z(n1433) );
  NAND U1459 ( .A(b[0]), .B(a[25]), .Z(n1339) );
  XNOR U1460 ( .A(b[1]), .B(n1339), .Z(n1341) );
  NANDN U1461 ( .A(b[0]), .B(a[24]), .Z(n1340) );
  NAND U1462 ( .A(n1341), .B(n1340), .Z(n1413) );
  NANDN U1463 ( .A(n9891), .B(n1342), .Z(n1344) );
  XOR U1464 ( .A(b[13]), .B(a[13]), .Z(n1416) );
  NANDN U1465 ( .A(n9935), .B(n1416), .Z(n1343) );
  AND U1466 ( .A(n1344), .B(n1343), .Z(n1411) );
  AND U1467 ( .A(b[15]), .B(a[9]), .Z(n1410) );
  XNOR U1468 ( .A(n1411), .B(n1410), .Z(n1412) );
  XNOR U1469 ( .A(n1413), .B(n1412), .Z(n1431) );
  NANDN U1470 ( .A(n9437), .B(n1345), .Z(n1347) );
  XOR U1471 ( .A(b[5]), .B(a[21]), .Z(n1422) );
  NANDN U1472 ( .A(n9503), .B(n1422), .Z(n1346) );
  AND U1473 ( .A(n1347), .B(n1346), .Z(n1455) );
  NANDN U1474 ( .A(n9588), .B(n1348), .Z(n1350) );
  XOR U1475 ( .A(b[7]), .B(a[19]), .Z(n1425) );
  NANDN U1476 ( .A(n9639), .B(n1425), .Z(n1349) );
  AND U1477 ( .A(n1350), .B(n1349), .Z(n1453) );
  NANDN U1478 ( .A(n9374), .B(n1351), .Z(n1353) );
  XOR U1479 ( .A(b[3]), .B(a[23]), .Z(n1428) );
  NANDN U1480 ( .A(n9375), .B(n1428), .Z(n1352) );
  NAND U1481 ( .A(n1353), .B(n1352), .Z(n1452) );
  XNOR U1482 ( .A(n1453), .B(n1452), .Z(n1454) );
  XOR U1483 ( .A(n1455), .B(n1454), .Z(n1432) );
  XOR U1484 ( .A(n1431), .B(n1432), .Z(n1434) );
  XOR U1485 ( .A(n1433), .B(n1434), .Z(n1405) );
  NANDN U1486 ( .A(n1355), .B(n1354), .Z(n1359) );
  OR U1487 ( .A(n1357), .B(n1356), .Z(n1358) );
  AND U1488 ( .A(n1359), .B(n1358), .Z(n1404) );
  XNOR U1489 ( .A(n1405), .B(n1404), .Z(n1407) );
  NAND U1490 ( .A(n1360), .B(n9883), .Z(n1362) );
  XOR U1491 ( .A(b[11]), .B(a[15]), .Z(n1437) );
  NANDN U1492 ( .A(n9856), .B(n1437), .Z(n1361) );
  AND U1493 ( .A(n1362), .B(n1361), .Z(n1448) );
  NANDN U1494 ( .A(n10005), .B(n1363), .Z(n1365) );
  XOR U1495 ( .A(b[15]), .B(a[11]), .Z(n1440) );
  NANDN U1496 ( .A(n10006), .B(n1440), .Z(n1364) );
  AND U1497 ( .A(n1365), .B(n1364), .Z(n1447) );
  NANDN U1498 ( .A(n9685), .B(n1366), .Z(n1368) );
  XOR U1499 ( .A(b[9]), .B(a[17]), .Z(n1443) );
  NANDN U1500 ( .A(n9758), .B(n1443), .Z(n1367) );
  NAND U1501 ( .A(n1368), .B(n1367), .Z(n1446) );
  XOR U1502 ( .A(n1447), .B(n1446), .Z(n1449) );
  XOR U1503 ( .A(n1448), .B(n1449), .Z(n1459) );
  NANDN U1504 ( .A(n1370), .B(n1369), .Z(n1374) );
  OR U1505 ( .A(n1372), .B(n1371), .Z(n1373) );
  AND U1506 ( .A(n1374), .B(n1373), .Z(n1458) );
  XNOR U1507 ( .A(n1459), .B(n1458), .Z(n1460) );
  NANDN U1508 ( .A(n1376), .B(n1375), .Z(n1380) );
  NANDN U1509 ( .A(n1378), .B(n1377), .Z(n1379) );
  NAND U1510 ( .A(n1380), .B(n1379), .Z(n1461) );
  XNOR U1511 ( .A(n1460), .B(n1461), .Z(n1406) );
  XOR U1512 ( .A(n1407), .B(n1406), .Z(n1465) );
  NANDN U1513 ( .A(n1382), .B(n1381), .Z(n1386) );
  NANDN U1514 ( .A(n1384), .B(n1383), .Z(n1385) );
  AND U1515 ( .A(n1386), .B(n1385), .Z(n1464) );
  XNOR U1516 ( .A(n1465), .B(n1464), .Z(n1466) );
  XOR U1517 ( .A(n1467), .B(n1466), .Z(n1399) );
  NANDN U1518 ( .A(n1388), .B(n1387), .Z(n1392) );
  NAND U1519 ( .A(n1390), .B(n1389), .Z(n1391) );
  AND U1520 ( .A(n1392), .B(n1391), .Z(n1398) );
  XNOR U1521 ( .A(n1399), .B(n1398), .Z(n1400) );
  XNOR U1522 ( .A(n1401), .B(n1400), .Z(n1470) );
  XNOR U1523 ( .A(sreg[137]), .B(n1470), .Z(n1472) );
  NANDN U1524 ( .A(sreg[136]), .B(n1393), .Z(n1397) );
  NAND U1525 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U1526 ( .A(n1397), .B(n1396), .Z(n1471) );
  XNOR U1527 ( .A(n1472), .B(n1471), .Z(c[137]) );
  NANDN U1528 ( .A(n1399), .B(n1398), .Z(n1403) );
  NANDN U1529 ( .A(n1401), .B(n1400), .Z(n1402) );
  AND U1530 ( .A(n1403), .B(n1402), .Z(n1478) );
  NANDN U1531 ( .A(n1405), .B(n1404), .Z(n1409) );
  NAND U1532 ( .A(n1407), .B(n1406), .Z(n1408) );
  AND U1533 ( .A(n1409), .B(n1408), .Z(n1544) );
  NANDN U1534 ( .A(n1411), .B(n1410), .Z(n1415) );
  NANDN U1535 ( .A(n1413), .B(n1412), .Z(n1414) );
  AND U1536 ( .A(n1415), .B(n1414), .Z(n1510) );
  NANDN U1537 ( .A(n9891), .B(n1416), .Z(n1418) );
  XOR U1538 ( .A(b[13]), .B(a[14]), .Z(n1496) );
  NANDN U1539 ( .A(n9935), .B(n1496), .Z(n1417) );
  AND U1540 ( .A(n1418), .B(n1417), .Z(n1488) );
  AND U1541 ( .A(b[15]), .B(a[10]), .Z(n1487) );
  XNOR U1542 ( .A(n1488), .B(n1487), .Z(n1489) );
  NAND U1543 ( .A(b[0]), .B(a[26]), .Z(n1419) );
  XNOR U1544 ( .A(b[1]), .B(n1419), .Z(n1421) );
  NANDN U1545 ( .A(b[0]), .B(a[25]), .Z(n1420) );
  NAND U1546 ( .A(n1421), .B(n1420), .Z(n1490) );
  XNOR U1547 ( .A(n1489), .B(n1490), .Z(n1508) );
  NANDN U1548 ( .A(n9437), .B(n1422), .Z(n1424) );
  XOR U1549 ( .A(b[5]), .B(a[22]), .Z(n1499) );
  NANDN U1550 ( .A(n9503), .B(n1499), .Z(n1423) );
  AND U1551 ( .A(n1424), .B(n1423), .Z(n1532) );
  NANDN U1552 ( .A(n9588), .B(n1425), .Z(n1427) );
  XOR U1553 ( .A(b[7]), .B(a[20]), .Z(n1502) );
  NANDN U1554 ( .A(n9639), .B(n1502), .Z(n1426) );
  AND U1555 ( .A(n1427), .B(n1426), .Z(n1530) );
  NANDN U1556 ( .A(n9374), .B(n1428), .Z(n1430) );
  XOR U1557 ( .A(b[3]), .B(a[24]), .Z(n1505) );
  NANDN U1558 ( .A(n9375), .B(n1505), .Z(n1429) );
  NAND U1559 ( .A(n1430), .B(n1429), .Z(n1529) );
  XNOR U1560 ( .A(n1530), .B(n1529), .Z(n1531) );
  XOR U1561 ( .A(n1532), .B(n1531), .Z(n1509) );
  XOR U1562 ( .A(n1508), .B(n1509), .Z(n1511) );
  XOR U1563 ( .A(n1510), .B(n1511), .Z(n1482) );
  NANDN U1564 ( .A(n1432), .B(n1431), .Z(n1436) );
  OR U1565 ( .A(n1434), .B(n1433), .Z(n1435) );
  AND U1566 ( .A(n1436), .B(n1435), .Z(n1481) );
  XNOR U1567 ( .A(n1482), .B(n1481), .Z(n1484) );
  NAND U1568 ( .A(n1437), .B(n9883), .Z(n1439) );
  XOR U1569 ( .A(b[11]), .B(a[16]), .Z(n1514) );
  NANDN U1570 ( .A(n9856), .B(n1514), .Z(n1438) );
  AND U1571 ( .A(n1439), .B(n1438), .Z(n1525) );
  NANDN U1572 ( .A(n10005), .B(n1440), .Z(n1442) );
  XOR U1573 ( .A(b[15]), .B(a[12]), .Z(n1517) );
  NANDN U1574 ( .A(n10006), .B(n1517), .Z(n1441) );
  AND U1575 ( .A(n1442), .B(n1441), .Z(n1524) );
  NANDN U1576 ( .A(n9685), .B(n1443), .Z(n1445) );
  XOR U1577 ( .A(b[9]), .B(a[18]), .Z(n1520) );
  NANDN U1578 ( .A(n9758), .B(n1520), .Z(n1444) );
  NAND U1579 ( .A(n1445), .B(n1444), .Z(n1523) );
  XOR U1580 ( .A(n1524), .B(n1523), .Z(n1526) );
  XOR U1581 ( .A(n1525), .B(n1526), .Z(n1536) );
  NANDN U1582 ( .A(n1447), .B(n1446), .Z(n1451) );
  OR U1583 ( .A(n1449), .B(n1448), .Z(n1450) );
  AND U1584 ( .A(n1451), .B(n1450), .Z(n1535) );
  XNOR U1585 ( .A(n1536), .B(n1535), .Z(n1537) );
  NANDN U1586 ( .A(n1453), .B(n1452), .Z(n1457) );
  NANDN U1587 ( .A(n1455), .B(n1454), .Z(n1456) );
  NAND U1588 ( .A(n1457), .B(n1456), .Z(n1538) );
  XNOR U1589 ( .A(n1537), .B(n1538), .Z(n1483) );
  XOR U1590 ( .A(n1484), .B(n1483), .Z(n1542) );
  NANDN U1591 ( .A(n1459), .B(n1458), .Z(n1463) );
  NANDN U1592 ( .A(n1461), .B(n1460), .Z(n1462) );
  AND U1593 ( .A(n1463), .B(n1462), .Z(n1541) );
  XNOR U1594 ( .A(n1542), .B(n1541), .Z(n1543) );
  XOR U1595 ( .A(n1544), .B(n1543), .Z(n1476) );
  NANDN U1596 ( .A(n1465), .B(n1464), .Z(n1469) );
  NAND U1597 ( .A(n1467), .B(n1466), .Z(n1468) );
  AND U1598 ( .A(n1469), .B(n1468), .Z(n1475) );
  XNOR U1599 ( .A(n1476), .B(n1475), .Z(n1477) );
  XNOR U1600 ( .A(n1478), .B(n1477), .Z(n1547) );
  XNOR U1601 ( .A(sreg[138]), .B(n1547), .Z(n1549) );
  NANDN U1602 ( .A(sreg[137]), .B(n1470), .Z(n1474) );
  NAND U1603 ( .A(n1472), .B(n1471), .Z(n1473) );
  NAND U1604 ( .A(n1474), .B(n1473), .Z(n1548) );
  XNOR U1605 ( .A(n1549), .B(n1548), .Z(c[138]) );
  NANDN U1606 ( .A(n1476), .B(n1475), .Z(n1480) );
  NANDN U1607 ( .A(n1478), .B(n1477), .Z(n1479) );
  AND U1608 ( .A(n1480), .B(n1479), .Z(n1555) );
  NANDN U1609 ( .A(n1482), .B(n1481), .Z(n1486) );
  NAND U1610 ( .A(n1484), .B(n1483), .Z(n1485) );
  AND U1611 ( .A(n1486), .B(n1485), .Z(n1621) );
  NANDN U1612 ( .A(n1488), .B(n1487), .Z(n1492) );
  NANDN U1613 ( .A(n1490), .B(n1489), .Z(n1491) );
  AND U1614 ( .A(n1492), .B(n1491), .Z(n1587) );
  NAND U1615 ( .A(b[0]), .B(a[27]), .Z(n1493) );
  XNOR U1616 ( .A(b[1]), .B(n1493), .Z(n1495) );
  NANDN U1617 ( .A(b[0]), .B(a[26]), .Z(n1494) );
  NAND U1618 ( .A(n1495), .B(n1494), .Z(n1567) );
  NANDN U1619 ( .A(n9891), .B(n1496), .Z(n1498) );
  XOR U1620 ( .A(b[13]), .B(a[15]), .Z(n1573) );
  NANDN U1621 ( .A(n9935), .B(n1573), .Z(n1497) );
  AND U1622 ( .A(n1498), .B(n1497), .Z(n1565) );
  AND U1623 ( .A(b[15]), .B(a[11]), .Z(n1564) );
  XNOR U1624 ( .A(n1565), .B(n1564), .Z(n1566) );
  XNOR U1625 ( .A(n1567), .B(n1566), .Z(n1585) );
  NANDN U1626 ( .A(n9437), .B(n1499), .Z(n1501) );
  XOR U1627 ( .A(b[5]), .B(a[23]), .Z(n1576) );
  NANDN U1628 ( .A(n9503), .B(n1576), .Z(n1500) );
  AND U1629 ( .A(n1501), .B(n1500), .Z(n1609) );
  NANDN U1630 ( .A(n9588), .B(n1502), .Z(n1504) );
  XOR U1631 ( .A(b[7]), .B(a[21]), .Z(n1579) );
  NANDN U1632 ( .A(n9639), .B(n1579), .Z(n1503) );
  AND U1633 ( .A(n1504), .B(n1503), .Z(n1607) );
  NANDN U1634 ( .A(n9374), .B(n1505), .Z(n1507) );
  XOR U1635 ( .A(b[3]), .B(a[25]), .Z(n1582) );
  NANDN U1636 ( .A(n9375), .B(n1582), .Z(n1506) );
  NAND U1637 ( .A(n1507), .B(n1506), .Z(n1606) );
  XNOR U1638 ( .A(n1607), .B(n1606), .Z(n1608) );
  XOR U1639 ( .A(n1609), .B(n1608), .Z(n1586) );
  XOR U1640 ( .A(n1585), .B(n1586), .Z(n1588) );
  XOR U1641 ( .A(n1587), .B(n1588), .Z(n1559) );
  NANDN U1642 ( .A(n1509), .B(n1508), .Z(n1513) );
  OR U1643 ( .A(n1511), .B(n1510), .Z(n1512) );
  AND U1644 ( .A(n1513), .B(n1512), .Z(n1558) );
  XNOR U1645 ( .A(n1559), .B(n1558), .Z(n1561) );
  NAND U1646 ( .A(n1514), .B(n9883), .Z(n1516) );
  XOR U1647 ( .A(b[11]), .B(a[17]), .Z(n1591) );
  NANDN U1648 ( .A(n9856), .B(n1591), .Z(n1515) );
  AND U1649 ( .A(n1516), .B(n1515), .Z(n1602) );
  NANDN U1650 ( .A(n10005), .B(n1517), .Z(n1519) );
  XOR U1651 ( .A(b[15]), .B(a[13]), .Z(n1594) );
  NANDN U1652 ( .A(n10006), .B(n1594), .Z(n1518) );
  AND U1653 ( .A(n1519), .B(n1518), .Z(n1601) );
  NANDN U1654 ( .A(n9685), .B(n1520), .Z(n1522) );
  XOR U1655 ( .A(b[9]), .B(a[19]), .Z(n1597) );
  NANDN U1656 ( .A(n9758), .B(n1597), .Z(n1521) );
  NAND U1657 ( .A(n1522), .B(n1521), .Z(n1600) );
  XOR U1658 ( .A(n1601), .B(n1600), .Z(n1603) );
  XOR U1659 ( .A(n1602), .B(n1603), .Z(n1613) );
  NANDN U1660 ( .A(n1524), .B(n1523), .Z(n1528) );
  OR U1661 ( .A(n1526), .B(n1525), .Z(n1527) );
  AND U1662 ( .A(n1528), .B(n1527), .Z(n1612) );
  XNOR U1663 ( .A(n1613), .B(n1612), .Z(n1614) );
  NANDN U1664 ( .A(n1530), .B(n1529), .Z(n1534) );
  NANDN U1665 ( .A(n1532), .B(n1531), .Z(n1533) );
  NAND U1666 ( .A(n1534), .B(n1533), .Z(n1615) );
  XNOR U1667 ( .A(n1614), .B(n1615), .Z(n1560) );
  XOR U1668 ( .A(n1561), .B(n1560), .Z(n1619) );
  NANDN U1669 ( .A(n1536), .B(n1535), .Z(n1540) );
  NANDN U1670 ( .A(n1538), .B(n1537), .Z(n1539) );
  AND U1671 ( .A(n1540), .B(n1539), .Z(n1618) );
  XNOR U1672 ( .A(n1619), .B(n1618), .Z(n1620) );
  XOR U1673 ( .A(n1621), .B(n1620), .Z(n1553) );
  NANDN U1674 ( .A(n1542), .B(n1541), .Z(n1546) );
  NAND U1675 ( .A(n1544), .B(n1543), .Z(n1545) );
  AND U1676 ( .A(n1546), .B(n1545), .Z(n1552) );
  XNOR U1677 ( .A(n1553), .B(n1552), .Z(n1554) );
  XNOR U1678 ( .A(n1555), .B(n1554), .Z(n1624) );
  XNOR U1679 ( .A(sreg[139]), .B(n1624), .Z(n1626) );
  NANDN U1680 ( .A(sreg[138]), .B(n1547), .Z(n1551) );
  NAND U1681 ( .A(n1549), .B(n1548), .Z(n1550) );
  NAND U1682 ( .A(n1551), .B(n1550), .Z(n1625) );
  XNOR U1683 ( .A(n1626), .B(n1625), .Z(c[139]) );
  NANDN U1684 ( .A(n1553), .B(n1552), .Z(n1557) );
  NANDN U1685 ( .A(n1555), .B(n1554), .Z(n1556) );
  AND U1686 ( .A(n1557), .B(n1556), .Z(n1632) );
  NANDN U1687 ( .A(n1559), .B(n1558), .Z(n1563) );
  NAND U1688 ( .A(n1561), .B(n1560), .Z(n1562) );
  AND U1689 ( .A(n1563), .B(n1562), .Z(n1698) );
  NANDN U1690 ( .A(n1565), .B(n1564), .Z(n1569) );
  NANDN U1691 ( .A(n1567), .B(n1566), .Z(n1568) );
  AND U1692 ( .A(n1569), .B(n1568), .Z(n1664) );
  NAND U1693 ( .A(b[0]), .B(a[28]), .Z(n1570) );
  XNOR U1694 ( .A(b[1]), .B(n1570), .Z(n1572) );
  NANDN U1695 ( .A(b[0]), .B(a[27]), .Z(n1571) );
  NAND U1696 ( .A(n1572), .B(n1571), .Z(n1644) );
  NANDN U1697 ( .A(n9891), .B(n1573), .Z(n1575) );
  XOR U1698 ( .A(b[13]), .B(a[16]), .Z(n1647) );
  NANDN U1699 ( .A(n9935), .B(n1647), .Z(n1574) );
  AND U1700 ( .A(n1575), .B(n1574), .Z(n1642) );
  AND U1701 ( .A(b[15]), .B(a[12]), .Z(n1641) );
  XNOR U1702 ( .A(n1642), .B(n1641), .Z(n1643) );
  XNOR U1703 ( .A(n1644), .B(n1643), .Z(n1662) );
  NANDN U1704 ( .A(n9437), .B(n1576), .Z(n1578) );
  XOR U1705 ( .A(b[5]), .B(a[24]), .Z(n1653) );
  NANDN U1706 ( .A(n9503), .B(n1653), .Z(n1577) );
  AND U1707 ( .A(n1578), .B(n1577), .Z(n1686) );
  NANDN U1708 ( .A(n9588), .B(n1579), .Z(n1581) );
  XOR U1709 ( .A(b[7]), .B(a[22]), .Z(n1656) );
  NANDN U1710 ( .A(n9639), .B(n1656), .Z(n1580) );
  AND U1711 ( .A(n1581), .B(n1580), .Z(n1684) );
  NANDN U1712 ( .A(n9374), .B(n1582), .Z(n1584) );
  XOR U1713 ( .A(b[3]), .B(a[26]), .Z(n1659) );
  NANDN U1714 ( .A(n9375), .B(n1659), .Z(n1583) );
  NAND U1715 ( .A(n1584), .B(n1583), .Z(n1683) );
  XNOR U1716 ( .A(n1684), .B(n1683), .Z(n1685) );
  XOR U1717 ( .A(n1686), .B(n1685), .Z(n1663) );
  XOR U1718 ( .A(n1662), .B(n1663), .Z(n1665) );
  XOR U1719 ( .A(n1664), .B(n1665), .Z(n1636) );
  NANDN U1720 ( .A(n1586), .B(n1585), .Z(n1590) );
  OR U1721 ( .A(n1588), .B(n1587), .Z(n1589) );
  AND U1722 ( .A(n1590), .B(n1589), .Z(n1635) );
  XNOR U1723 ( .A(n1636), .B(n1635), .Z(n1638) );
  NAND U1724 ( .A(n1591), .B(n9883), .Z(n1593) );
  XOR U1725 ( .A(b[11]), .B(a[18]), .Z(n1668) );
  NANDN U1726 ( .A(n9856), .B(n1668), .Z(n1592) );
  AND U1727 ( .A(n1593), .B(n1592), .Z(n1679) );
  NANDN U1728 ( .A(n10005), .B(n1594), .Z(n1596) );
  XOR U1729 ( .A(b[15]), .B(a[14]), .Z(n1671) );
  NANDN U1730 ( .A(n10006), .B(n1671), .Z(n1595) );
  AND U1731 ( .A(n1596), .B(n1595), .Z(n1678) );
  NANDN U1732 ( .A(n9685), .B(n1597), .Z(n1599) );
  XOR U1733 ( .A(b[9]), .B(a[20]), .Z(n1674) );
  NANDN U1734 ( .A(n9758), .B(n1674), .Z(n1598) );
  NAND U1735 ( .A(n1599), .B(n1598), .Z(n1677) );
  XOR U1736 ( .A(n1678), .B(n1677), .Z(n1680) );
  XOR U1737 ( .A(n1679), .B(n1680), .Z(n1690) );
  NANDN U1738 ( .A(n1601), .B(n1600), .Z(n1605) );
  OR U1739 ( .A(n1603), .B(n1602), .Z(n1604) );
  AND U1740 ( .A(n1605), .B(n1604), .Z(n1689) );
  XNOR U1741 ( .A(n1690), .B(n1689), .Z(n1691) );
  NANDN U1742 ( .A(n1607), .B(n1606), .Z(n1611) );
  NANDN U1743 ( .A(n1609), .B(n1608), .Z(n1610) );
  NAND U1744 ( .A(n1611), .B(n1610), .Z(n1692) );
  XNOR U1745 ( .A(n1691), .B(n1692), .Z(n1637) );
  XOR U1746 ( .A(n1638), .B(n1637), .Z(n1696) );
  NANDN U1747 ( .A(n1613), .B(n1612), .Z(n1617) );
  NANDN U1748 ( .A(n1615), .B(n1614), .Z(n1616) );
  AND U1749 ( .A(n1617), .B(n1616), .Z(n1695) );
  XNOR U1750 ( .A(n1696), .B(n1695), .Z(n1697) );
  XOR U1751 ( .A(n1698), .B(n1697), .Z(n1630) );
  NANDN U1752 ( .A(n1619), .B(n1618), .Z(n1623) );
  NAND U1753 ( .A(n1621), .B(n1620), .Z(n1622) );
  AND U1754 ( .A(n1623), .B(n1622), .Z(n1629) );
  XNOR U1755 ( .A(n1630), .B(n1629), .Z(n1631) );
  XNOR U1756 ( .A(n1632), .B(n1631), .Z(n1701) );
  XNOR U1757 ( .A(sreg[140]), .B(n1701), .Z(n1703) );
  NANDN U1758 ( .A(sreg[139]), .B(n1624), .Z(n1628) );
  NAND U1759 ( .A(n1626), .B(n1625), .Z(n1627) );
  NAND U1760 ( .A(n1628), .B(n1627), .Z(n1702) );
  XNOR U1761 ( .A(n1703), .B(n1702), .Z(c[140]) );
  NANDN U1762 ( .A(n1630), .B(n1629), .Z(n1634) );
  NANDN U1763 ( .A(n1632), .B(n1631), .Z(n1633) );
  AND U1764 ( .A(n1634), .B(n1633), .Z(n1709) );
  NANDN U1765 ( .A(n1636), .B(n1635), .Z(n1640) );
  NAND U1766 ( .A(n1638), .B(n1637), .Z(n1639) );
  AND U1767 ( .A(n1640), .B(n1639), .Z(n1775) );
  NANDN U1768 ( .A(n1642), .B(n1641), .Z(n1646) );
  NANDN U1769 ( .A(n1644), .B(n1643), .Z(n1645) );
  AND U1770 ( .A(n1646), .B(n1645), .Z(n1762) );
  NANDN U1771 ( .A(n9891), .B(n1647), .Z(n1649) );
  XOR U1772 ( .A(b[13]), .B(a[17]), .Z(n1748) );
  NANDN U1773 ( .A(n9935), .B(n1748), .Z(n1648) );
  AND U1774 ( .A(n1649), .B(n1648), .Z(n1740) );
  AND U1775 ( .A(b[15]), .B(a[13]), .Z(n1739) );
  XNOR U1776 ( .A(n1740), .B(n1739), .Z(n1741) );
  NAND U1777 ( .A(b[0]), .B(a[29]), .Z(n1650) );
  XNOR U1778 ( .A(b[1]), .B(n1650), .Z(n1652) );
  NANDN U1779 ( .A(b[0]), .B(a[28]), .Z(n1651) );
  NAND U1780 ( .A(n1652), .B(n1651), .Z(n1742) );
  XNOR U1781 ( .A(n1741), .B(n1742), .Z(n1760) );
  NANDN U1782 ( .A(n9437), .B(n1653), .Z(n1655) );
  XOR U1783 ( .A(b[5]), .B(a[25]), .Z(n1751) );
  NANDN U1784 ( .A(n9503), .B(n1751), .Z(n1654) );
  AND U1785 ( .A(n1655), .B(n1654), .Z(n1736) );
  NANDN U1786 ( .A(n9588), .B(n1656), .Z(n1658) );
  XOR U1787 ( .A(b[7]), .B(a[23]), .Z(n1754) );
  NANDN U1788 ( .A(n9639), .B(n1754), .Z(n1657) );
  AND U1789 ( .A(n1658), .B(n1657), .Z(n1734) );
  NANDN U1790 ( .A(n9374), .B(n1659), .Z(n1661) );
  XOR U1791 ( .A(b[3]), .B(a[27]), .Z(n1757) );
  NANDN U1792 ( .A(n9375), .B(n1757), .Z(n1660) );
  NAND U1793 ( .A(n1661), .B(n1660), .Z(n1733) );
  XNOR U1794 ( .A(n1734), .B(n1733), .Z(n1735) );
  XOR U1795 ( .A(n1736), .B(n1735), .Z(n1761) );
  XOR U1796 ( .A(n1760), .B(n1761), .Z(n1763) );
  XOR U1797 ( .A(n1762), .B(n1763), .Z(n1713) );
  NANDN U1798 ( .A(n1663), .B(n1662), .Z(n1667) );
  OR U1799 ( .A(n1665), .B(n1664), .Z(n1666) );
  AND U1800 ( .A(n1667), .B(n1666), .Z(n1712) );
  XNOR U1801 ( .A(n1713), .B(n1712), .Z(n1715) );
  NAND U1802 ( .A(n1668), .B(n9883), .Z(n1670) );
  XOR U1803 ( .A(b[11]), .B(a[19]), .Z(n1718) );
  NANDN U1804 ( .A(n9856), .B(n1718), .Z(n1669) );
  AND U1805 ( .A(n1670), .B(n1669), .Z(n1729) );
  NANDN U1806 ( .A(n10005), .B(n1671), .Z(n1673) );
  XOR U1807 ( .A(b[15]), .B(a[15]), .Z(n1721) );
  NANDN U1808 ( .A(n10006), .B(n1721), .Z(n1672) );
  AND U1809 ( .A(n1673), .B(n1672), .Z(n1728) );
  NANDN U1810 ( .A(n9685), .B(n1674), .Z(n1676) );
  XOR U1811 ( .A(b[9]), .B(a[21]), .Z(n1724) );
  NANDN U1812 ( .A(n9758), .B(n1724), .Z(n1675) );
  NAND U1813 ( .A(n1676), .B(n1675), .Z(n1727) );
  XOR U1814 ( .A(n1728), .B(n1727), .Z(n1730) );
  XOR U1815 ( .A(n1729), .B(n1730), .Z(n1767) );
  NANDN U1816 ( .A(n1678), .B(n1677), .Z(n1682) );
  OR U1817 ( .A(n1680), .B(n1679), .Z(n1681) );
  AND U1818 ( .A(n1682), .B(n1681), .Z(n1766) );
  XNOR U1819 ( .A(n1767), .B(n1766), .Z(n1768) );
  NANDN U1820 ( .A(n1684), .B(n1683), .Z(n1688) );
  NANDN U1821 ( .A(n1686), .B(n1685), .Z(n1687) );
  NAND U1822 ( .A(n1688), .B(n1687), .Z(n1769) );
  XNOR U1823 ( .A(n1768), .B(n1769), .Z(n1714) );
  XOR U1824 ( .A(n1715), .B(n1714), .Z(n1773) );
  NANDN U1825 ( .A(n1690), .B(n1689), .Z(n1694) );
  NANDN U1826 ( .A(n1692), .B(n1691), .Z(n1693) );
  AND U1827 ( .A(n1694), .B(n1693), .Z(n1772) );
  XNOR U1828 ( .A(n1773), .B(n1772), .Z(n1774) );
  XOR U1829 ( .A(n1775), .B(n1774), .Z(n1707) );
  NANDN U1830 ( .A(n1696), .B(n1695), .Z(n1700) );
  NAND U1831 ( .A(n1698), .B(n1697), .Z(n1699) );
  AND U1832 ( .A(n1700), .B(n1699), .Z(n1706) );
  XNOR U1833 ( .A(n1707), .B(n1706), .Z(n1708) );
  XNOR U1834 ( .A(n1709), .B(n1708), .Z(n1778) );
  XNOR U1835 ( .A(sreg[141]), .B(n1778), .Z(n1780) );
  NANDN U1836 ( .A(sreg[140]), .B(n1701), .Z(n1705) );
  NAND U1837 ( .A(n1703), .B(n1702), .Z(n1704) );
  NAND U1838 ( .A(n1705), .B(n1704), .Z(n1779) );
  XNOR U1839 ( .A(n1780), .B(n1779), .Z(c[141]) );
  NANDN U1840 ( .A(n1707), .B(n1706), .Z(n1711) );
  NANDN U1841 ( .A(n1709), .B(n1708), .Z(n1710) );
  AND U1842 ( .A(n1711), .B(n1710), .Z(n1786) );
  NANDN U1843 ( .A(n1713), .B(n1712), .Z(n1717) );
  NAND U1844 ( .A(n1715), .B(n1714), .Z(n1716) );
  AND U1845 ( .A(n1717), .B(n1716), .Z(n1852) );
  NAND U1846 ( .A(n1718), .B(n9883), .Z(n1720) );
  XOR U1847 ( .A(b[11]), .B(a[20]), .Z(n1822) );
  NANDN U1848 ( .A(n9856), .B(n1822), .Z(n1719) );
  AND U1849 ( .A(n1720), .B(n1719), .Z(n1833) );
  NANDN U1850 ( .A(n10005), .B(n1721), .Z(n1723) );
  XOR U1851 ( .A(b[15]), .B(a[16]), .Z(n1825) );
  NANDN U1852 ( .A(n10006), .B(n1825), .Z(n1722) );
  AND U1853 ( .A(n1723), .B(n1722), .Z(n1832) );
  NANDN U1854 ( .A(n9685), .B(n1724), .Z(n1726) );
  XOR U1855 ( .A(b[9]), .B(a[22]), .Z(n1828) );
  NANDN U1856 ( .A(n9758), .B(n1828), .Z(n1725) );
  NAND U1857 ( .A(n1726), .B(n1725), .Z(n1831) );
  XOR U1858 ( .A(n1832), .B(n1831), .Z(n1834) );
  XOR U1859 ( .A(n1833), .B(n1834), .Z(n1844) );
  NANDN U1860 ( .A(n1728), .B(n1727), .Z(n1732) );
  OR U1861 ( .A(n1730), .B(n1729), .Z(n1731) );
  AND U1862 ( .A(n1732), .B(n1731), .Z(n1843) );
  XNOR U1863 ( .A(n1844), .B(n1843), .Z(n1845) );
  NANDN U1864 ( .A(n1734), .B(n1733), .Z(n1738) );
  NANDN U1865 ( .A(n1736), .B(n1735), .Z(n1737) );
  NAND U1866 ( .A(n1738), .B(n1737), .Z(n1846) );
  XNOR U1867 ( .A(n1845), .B(n1846), .Z(n1792) );
  NANDN U1868 ( .A(n1740), .B(n1739), .Z(n1744) );
  NANDN U1869 ( .A(n1742), .B(n1741), .Z(n1743) );
  AND U1870 ( .A(n1744), .B(n1743), .Z(n1818) );
  NAND U1871 ( .A(b[0]), .B(a[30]), .Z(n1745) );
  XNOR U1872 ( .A(b[1]), .B(n1745), .Z(n1747) );
  NANDN U1873 ( .A(b[0]), .B(a[29]), .Z(n1746) );
  NAND U1874 ( .A(n1747), .B(n1746), .Z(n1798) );
  NANDN U1875 ( .A(n9891), .B(n1748), .Z(n1750) );
  XOR U1876 ( .A(b[13]), .B(a[18]), .Z(n1801) );
  NANDN U1877 ( .A(n9935), .B(n1801), .Z(n1749) );
  AND U1878 ( .A(n1750), .B(n1749), .Z(n1796) );
  AND U1879 ( .A(b[15]), .B(a[14]), .Z(n1795) );
  XNOR U1880 ( .A(n1796), .B(n1795), .Z(n1797) );
  XNOR U1881 ( .A(n1798), .B(n1797), .Z(n1816) );
  NANDN U1882 ( .A(n9437), .B(n1751), .Z(n1753) );
  XOR U1883 ( .A(b[5]), .B(a[26]), .Z(n1807) );
  NANDN U1884 ( .A(n9503), .B(n1807), .Z(n1752) );
  AND U1885 ( .A(n1753), .B(n1752), .Z(n1840) );
  NANDN U1886 ( .A(n9588), .B(n1754), .Z(n1756) );
  XOR U1887 ( .A(b[7]), .B(a[24]), .Z(n1810) );
  NANDN U1888 ( .A(n9639), .B(n1810), .Z(n1755) );
  AND U1889 ( .A(n1756), .B(n1755), .Z(n1838) );
  NANDN U1890 ( .A(n9374), .B(n1757), .Z(n1759) );
  XOR U1891 ( .A(b[3]), .B(a[28]), .Z(n1813) );
  NANDN U1892 ( .A(n9375), .B(n1813), .Z(n1758) );
  NAND U1893 ( .A(n1759), .B(n1758), .Z(n1837) );
  XNOR U1894 ( .A(n1838), .B(n1837), .Z(n1839) );
  XOR U1895 ( .A(n1840), .B(n1839), .Z(n1817) );
  XOR U1896 ( .A(n1816), .B(n1817), .Z(n1819) );
  XOR U1897 ( .A(n1818), .B(n1819), .Z(n1790) );
  NANDN U1898 ( .A(n1761), .B(n1760), .Z(n1765) );
  OR U1899 ( .A(n1763), .B(n1762), .Z(n1764) );
  AND U1900 ( .A(n1765), .B(n1764), .Z(n1789) );
  XNOR U1901 ( .A(n1790), .B(n1789), .Z(n1791) );
  XOR U1902 ( .A(n1792), .B(n1791), .Z(n1850) );
  NANDN U1903 ( .A(n1767), .B(n1766), .Z(n1771) );
  NANDN U1904 ( .A(n1769), .B(n1768), .Z(n1770) );
  AND U1905 ( .A(n1771), .B(n1770), .Z(n1849) );
  XNOR U1906 ( .A(n1850), .B(n1849), .Z(n1851) );
  XOR U1907 ( .A(n1852), .B(n1851), .Z(n1784) );
  NANDN U1908 ( .A(n1773), .B(n1772), .Z(n1777) );
  NAND U1909 ( .A(n1775), .B(n1774), .Z(n1776) );
  AND U1910 ( .A(n1777), .B(n1776), .Z(n1783) );
  XNOR U1911 ( .A(n1784), .B(n1783), .Z(n1785) );
  XNOR U1912 ( .A(n1786), .B(n1785), .Z(n1855) );
  XNOR U1913 ( .A(sreg[142]), .B(n1855), .Z(n1857) );
  NANDN U1914 ( .A(sreg[141]), .B(n1778), .Z(n1782) );
  NAND U1915 ( .A(n1780), .B(n1779), .Z(n1781) );
  NAND U1916 ( .A(n1782), .B(n1781), .Z(n1856) );
  XNOR U1917 ( .A(n1857), .B(n1856), .Z(c[142]) );
  NANDN U1918 ( .A(n1784), .B(n1783), .Z(n1788) );
  NANDN U1919 ( .A(n1786), .B(n1785), .Z(n1787) );
  AND U1920 ( .A(n1788), .B(n1787), .Z(n1863) );
  NANDN U1921 ( .A(n1790), .B(n1789), .Z(n1794) );
  NAND U1922 ( .A(n1792), .B(n1791), .Z(n1793) );
  AND U1923 ( .A(n1794), .B(n1793), .Z(n1929) );
  NANDN U1924 ( .A(n1796), .B(n1795), .Z(n1800) );
  NANDN U1925 ( .A(n1798), .B(n1797), .Z(n1799) );
  AND U1926 ( .A(n1800), .B(n1799), .Z(n1895) );
  NANDN U1927 ( .A(n9891), .B(n1801), .Z(n1803) );
  XOR U1928 ( .A(b[13]), .B(a[19]), .Z(n1881) );
  NANDN U1929 ( .A(n9935), .B(n1881), .Z(n1802) );
  AND U1930 ( .A(n1803), .B(n1802), .Z(n1873) );
  AND U1931 ( .A(b[15]), .B(a[15]), .Z(n1872) );
  XNOR U1932 ( .A(n1873), .B(n1872), .Z(n1874) );
  NAND U1933 ( .A(b[0]), .B(a[31]), .Z(n1804) );
  XNOR U1934 ( .A(b[1]), .B(n1804), .Z(n1806) );
  NANDN U1935 ( .A(b[0]), .B(a[30]), .Z(n1805) );
  NAND U1936 ( .A(n1806), .B(n1805), .Z(n1875) );
  XNOR U1937 ( .A(n1874), .B(n1875), .Z(n1893) );
  NANDN U1938 ( .A(n9437), .B(n1807), .Z(n1809) );
  XOR U1939 ( .A(b[5]), .B(a[27]), .Z(n1884) );
  NANDN U1940 ( .A(n9503), .B(n1884), .Z(n1808) );
  AND U1941 ( .A(n1809), .B(n1808), .Z(n1917) );
  NANDN U1942 ( .A(n9588), .B(n1810), .Z(n1812) );
  XOR U1943 ( .A(b[7]), .B(a[25]), .Z(n1887) );
  NANDN U1944 ( .A(n9639), .B(n1887), .Z(n1811) );
  AND U1945 ( .A(n1812), .B(n1811), .Z(n1915) );
  NANDN U1946 ( .A(n9374), .B(n1813), .Z(n1815) );
  XOR U1947 ( .A(b[3]), .B(a[29]), .Z(n1890) );
  NANDN U1948 ( .A(n9375), .B(n1890), .Z(n1814) );
  NAND U1949 ( .A(n1815), .B(n1814), .Z(n1914) );
  XNOR U1950 ( .A(n1915), .B(n1914), .Z(n1916) );
  XOR U1951 ( .A(n1917), .B(n1916), .Z(n1894) );
  XOR U1952 ( .A(n1893), .B(n1894), .Z(n1896) );
  XOR U1953 ( .A(n1895), .B(n1896), .Z(n1867) );
  NANDN U1954 ( .A(n1817), .B(n1816), .Z(n1821) );
  OR U1955 ( .A(n1819), .B(n1818), .Z(n1820) );
  AND U1956 ( .A(n1821), .B(n1820), .Z(n1866) );
  XNOR U1957 ( .A(n1867), .B(n1866), .Z(n1869) );
  NAND U1958 ( .A(n1822), .B(n9883), .Z(n1824) );
  XOR U1959 ( .A(b[11]), .B(a[21]), .Z(n1899) );
  NANDN U1960 ( .A(n9856), .B(n1899), .Z(n1823) );
  AND U1961 ( .A(n1824), .B(n1823), .Z(n1910) );
  NANDN U1962 ( .A(n10005), .B(n1825), .Z(n1827) );
  XOR U1963 ( .A(b[15]), .B(a[17]), .Z(n1902) );
  NANDN U1964 ( .A(n10006), .B(n1902), .Z(n1826) );
  AND U1965 ( .A(n1827), .B(n1826), .Z(n1909) );
  NANDN U1966 ( .A(n9685), .B(n1828), .Z(n1830) );
  XOR U1967 ( .A(b[9]), .B(a[23]), .Z(n1905) );
  NANDN U1968 ( .A(n9758), .B(n1905), .Z(n1829) );
  NAND U1969 ( .A(n1830), .B(n1829), .Z(n1908) );
  XOR U1970 ( .A(n1909), .B(n1908), .Z(n1911) );
  XOR U1971 ( .A(n1910), .B(n1911), .Z(n1921) );
  NANDN U1972 ( .A(n1832), .B(n1831), .Z(n1836) );
  OR U1973 ( .A(n1834), .B(n1833), .Z(n1835) );
  AND U1974 ( .A(n1836), .B(n1835), .Z(n1920) );
  XNOR U1975 ( .A(n1921), .B(n1920), .Z(n1922) );
  NANDN U1976 ( .A(n1838), .B(n1837), .Z(n1842) );
  NANDN U1977 ( .A(n1840), .B(n1839), .Z(n1841) );
  NAND U1978 ( .A(n1842), .B(n1841), .Z(n1923) );
  XNOR U1979 ( .A(n1922), .B(n1923), .Z(n1868) );
  XOR U1980 ( .A(n1869), .B(n1868), .Z(n1927) );
  NANDN U1981 ( .A(n1844), .B(n1843), .Z(n1848) );
  NANDN U1982 ( .A(n1846), .B(n1845), .Z(n1847) );
  AND U1983 ( .A(n1848), .B(n1847), .Z(n1926) );
  XNOR U1984 ( .A(n1927), .B(n1926), .Z(n1928) );
  XOR U1985 ( .A(n1929), .B(n1928), .Z(n1861) );
  NANDN U1986 ( .A(n1850), .B(n1849), .Z(n1854) );
  NAND U1987 ( .A(n1852), .B(n1851), .Z(n1853) );
  AND U1988 ( .A(n1854), .B(n1853), .Z(n1860) );
  XNOR U1989 ( .A(n1861), .B(n1860), .Z(n1862) );
  XNOR U1990 ( .A(n1863), .B(n1862), .Z(n1932) );
  XNOR U1991 ( .A(sreg[143]), .B(n1932), .Z(n1934) );
  NANDN U1992 ( .A(sreg[142]), .B(n1855), .Z(n1859) );
  NAND U1993 ( .A(n1857), .B(n1856), .Z(n1858) );
  NAND U1994 ( .A(n1859), .B(n1858), .Z(n1933) );
  XNOR U1995 ( .A(n1934), .B(n1933), .Z(c[143]) );
  NANDN U1996 ( .A(n1861), .B(n1860), .Z(n1865) );
  NANDN U1997 ( .A(n1863), .B(n1862), .Z(n1864) );
  AND U1998 ( .A(n1865), .B(n1864), .Z(n1940) );
  NANDN U1999 ( .A(n1867), .B(n1866), .Z(n1871) );
  NAND U2000 ( .A(n1869), .B(n1868), .Z(n1870) );
  AND U2001 ( .A(n1871), .B(n1870), .Z(n2006) );
  NANDN U2002 ( .A(n1873), .B(n1872), .Z(n1877) );
  NANDN U2003 ( .A(n1875), .B(n1874), .Z(n1876) );
  AND U2004 ( .A(n1877), .B(n1876), .Z(n1972) );
  NAND U2005 ( .A(b[0]), .B(a[32]), .Z(n1878) );
  XNOR U2006 ( .A(b[1]), .B(n1878), .Z(n1880) );
  NANDN U2007 ( .A(b[0]), .B(a[31]), .Z(n1879) );
  NAND U2008 ( .A(n1880), .B(n1879), .Z(n1952) );
  NANDN U2009 ( .A(n9891), .B(n1881), .Z(n1883) );
  XOR U2010 ( .A(b[13]), .B(a[20]), .Z(n1958) );
  NANDN U2011 ( .A(n9935), .B(n1958), .Z(n1882) );
  AND U2012 ( .A(n1883), .B(n1882), .Z(n1950) );
  AND U2013 ( .A(b[15]), .B(a[16]), .Z(n1949) );
  XNOR U2014 ( .A(n1950), .B(n1949), .Z(n1951) );
  XNOR U2015 ( .A(n1952), .B(n1951), .Z(n1970) );
  NANDN U2016 ( .A(n9437), .B(n1884), .Z(n1886) );
  XOR U2017 ( .A(b[5]), .B(a[28]), .Z(n1961) );
  NANDN U2018 ( .A(n9503), .B(n1961), .Z(n1885) );
  AND U2019 ( .A(n1886), .B(n1885), .Z(n1994) );
  NANDN U2020 ( .A(n9588), .B(n1887), .Z(n1889) );
  XOR U2021 ( .A(b[7]), .B(a[26]), .Z(n1964) );
  NANDN U2022 ( .A(n9639), .B(n1964), .Z(n1888) );
  AND U2023 ( .A(n1889), .B(n1888), .Z(n1992) );
  NANDN U2024 ( .A(n9374), .B(n1890), .Z(n1892) );
  XOR U2025 ( .A(b[3]), .B(a[30]), .Z(n1967) );
  NANDN U2026 ( .A(n9375), .B(n1967), .Z(n1891) );
  NAND U2027 ( .A(n1892), .B(n1891), .Z(n1991) );
  XNOR U2028 ( .A(n1992), .B(n1991), .Z(n1993) );
  XOR U2029 ( .A(n1994), .B(n1993), .Z(n1971) );
  XOR U2030 ( .A(n1970), .B(n1971), .Z(n1973) );
  XOR U2031 ( .A(n1972), .B(n1973), .Z(n1944) );
  NANDN U2032 ( .A(n1894), .B(n1893), .Z(n1898) );
  OR U2033 ( .A(n1896), .B(n1895), .Z(n1897) );
  AND U2034 ( .A(n1898), .B(n1897), .Z(n1943) );
  XNOR U2035 ( .A(n1944), .B(n1943), .Z(n1946) );
  NAND U2036 ( .A(n1899), .B(n9883), .Z(n1901) );
  XOR U2037 ( .A(b[11]), .B(a[22]), .Z(n1976) );
  NANDN U2038 ( .A(n9856), .B(n1976), .Z(n1900) );
  AND U2039 ( .A(n1901), .B(n1900), .Z(n1987) );
  NANDN U2040 ( .A(n10005), .B(n1902), .Z(n1904) );
  XOR U2041 ( .A(b[15]), .B(a[18]), .Z(n1979) );
  NANDN U2042 ( .A(n10006), .B(n1979), .Z(n1903) );
  AND U2043 ( .A(n1904), .B(n1903), .Z(n1986) );
  NANDN U2044 ( .A(n9685), .B(n1905), .Z(n1907) );
  XOR U2045 ( .A(b[9]), .B(a[24]), .Z(n1982) );
  NANDN U2046 ( .A(n9758), .B(n1982), .Z(n1906) );
  NAND U2047 ( .A(n1907), .B(n1906), .Z(n1985) );
  XOR U2048 ( .A(n1986), .B(n1985), .Z(n1988) );
  XOR U2049 ( .A(n1987), .B(n1988), .Z(n1998) );
  NANDN U2050 ( .A(n1909), .B(n1908), .Z(n1913) );
  OR U2051 ( .A(n1911), .B(n1910), .Z(n1912) );
  AND U2052 ( .A(n1913), .B(n1912), .Z(n1997) );
  XNOR U2053 ( .A(n1998), .B(n1997), .Z(n1999) );
  NANDN U2054 ( .A(n1915), .B(n1914), .Z(n1919) );
  NANDN U2055 ( .A(n1917), .B(n1916), .Z(n1918) );
  NAND U2056 ( .A(n1919), .B(n1918), .Z(n2000) );
  XNOR U2057 ( .A(n1999), .B(n2000), .Z(n1945) );
  XOR U2058 ( .A(n1946), .B(n1945), .Z(n2004) );
  NANDN U2059 ( .A(n1921), .B(n1920), .Z(n1925) );
  NANDN U2060 ( .A(n1923), .B(n1922), .Z(n1924) );
  AND U2061 ( .A(n1925), .B(n1924), .Z(n2003) );
  XNOR U2062 ( .A(n2004), .B(n2003), .Z(n2005) );
  XOR U2063 ( .A(n2006), .B(n2005), .Z(n1938) );
  NANDN U2064 ( .A(n1927), .B(n1926), .Z(n1931) );
  NAND U2065 ( .A(n1929), .B(n1928), .Z(n1930) );
  AND U2066 ( .A(n1931), .B(n1930), .Z(n1937) );
  XNOR U2067 ( .A(n1938), .B(n1937), .Z(n1939) );
  XNOR U2068 ( .A(n1940), .B(n1939), .Z(n2009) );
  XNOR U2069 ( .A(sreg[144]), .B(n2009), .Z(n2011) );
  NANDN U2070 ( .A(sreg[143]), .B(n1932), .Z(n1936) );
  NAND U2071 ( .A(n1934), .B(n1933), .Z(n1935) );
  NAND U2072 ( .A(n1936), .B(n1935), .Z(n2010) );
  XNOR U2073 ( .A(n2011), .B(n2010), .Z(c[144]) );
  NANDN U2074 ( .A(n1938), .B(n1937), .Z(n1942) );
  NANDN U2075 ( .A(n1940), .B(n1939), .Z(n1941) );
  AND U2076 ( .A(n1942), .B(n1941), .Z(n2017) );
  NANDN U2077 ( .A(n1944), .B(n1943), .Z(n1948) );
  NAND U2078 ( .A(n1946), .B(n1945), .Z(n1947) );
  AND U2079 ( .A(n1948), .B(n1947), .Z(n2083) );
  NANDN U2080 ( .A(n1950), .B(n1949), .Z(n1954) );
  NANDN U2081 ( .A(n1952), .B(n1951), .Z(n1953) );
  AND U2082 ( .A(n1954), .B(n1953), .Z(n2049) );
  NAND U2083 ( .A(b[0]), .B(a[33]), .Z(n1955) );
  XNOR U2084 ( .A(b[1]), .B(n1955), .Z(n1957) );
  NANDN U2085 ( .A(b[0]), .B(a[32]), .Z(n1956) );
  NAND U2086 ( .A(n1957), .B(n1956), .Z(n2029) );
  NANDN U2087 ( .A(n9891), .B(n1958), .Z(n1960) );
  XOR U2088 ( .A(b[13]), .B(a[21]), .Z(n2035) );
  NANDN U2089 ( .A(n9935), .B(n2035), .Z(n1959) );
  AND U2090 ( .A(n1960), .B(n1959), .Z(n2027) );
  AND U2091 ( .A(b[15]), .B(a[17]), .Z(n2026) );
  XNOR U2092 ( .A(n2027), .B(n2026), .Z(n2028) );
  XNOR U2093 ( .A(n2029), .B(n2028), .Z(n2047) );
  NANDN U2094 ( .A(n9437), .B(n1961), .Z(n1963) );
  XOR U2095 ( .A(b[5]), .B(a[29]), .Z(n2038) );
  NANDN U2096 ( .A(n9503), .B(n2038), .Z(n1962) );
  AND U2097 ( .A(n1963), .B(n1962), .Z(n2071) );
  NANDN U2098 ( .A(n9588), .B(n1964), .Z(n1966) );
  XOR U2099 ( .A(b[7]), .B(a[27]), .Z(n2041) );
  NANDN U2100 ( .A(n9639), .B(n2041), .Z(n1965) );
  AND U2101 ( .A(n1966), .B(n1965), .Z(n2069) );
  NANDN U2102 ( .A(n9374), .B(n1967), .Z(n1969) );
  XOR U2103 ( .A(b[3]), .B(a[31]), .Z(n2044) );
  NANDN U2104 ( .A(n9375), .B(n2044), .Z(n1968) );
  NAND U2105 ( .A(n1969), .B(n1968), .Z(n2068) );
  XNOR U2106 ( .A(n2069), .B(n2068), .Z(n2070) );
  XOR U2107 ( .A(n2071), .B(n2070), .Z(n2048) );
  XOR U2108 ( .A(n2047), .B(n2048), .Z(n2050) );
  XOR U2109 ( .A(n2049), .B(n2050), .Z(n2021) );
  NANDN U2110 ( .A(n1971), .B(n1970), .Z(n1975) );
  OR U2111 ( .A(n1973), .B(n1972), .Z(n1974) );
  AND U2112 ( .A(n1975), .B(n1974), .Z(n2020) );
  XNOR U2113 ( .A(n2021), .B(n2020), .Z(n2023) );
  NAND U2114 ( .A(n1976), .B(n9883), .Z(n1978) );
  XOR U2115 ( .A(b[11]), .B(a[23]), .Z(n2053) );
  NANDN U2116 ( .A(n9856), .B(n2053), .Z(n1977) );
  AND U2117 ( .A(n1978), .B(n1977), .Z(n2064) );
  NANDN U2118 ( .A(n10005), .B(n1979), .Z(n1981) );
  XOR U2119 ( .A(b[15]), .B(a[19]), .Z(n2056) );
  NANDN U2120 ( .A(n10006), .B(n2056), .Z(n1980) );
  AND U2121 ( .A(n1981), .B(n1980), .Z(n2063) );
  NANDN U2122 ( .A(n9685), .B(n1982), .Z(n1984) );
  XOR U2123 ( .A(b[9]), .B(a[25]), .Z(n2059) );
  NANDN U2124 ( .A(n9758), .B(n2059), .Z(n1983) );
  NAND U2125 ( .A(n1984), .B(n1983), .Z(n2062) );
  XOR U2126 ( .A(n2063), .B(n2062), .Z(n2065) );
  XOR U2127 ( .A(n2064), .B(n2065), .Z(n2075) );
  NANDN U2128 ( .A(n1986), .B(n1985), .Z(n1990) );
  OR U2129 ( .A(n1988), .B(n1987), .Z(n1989) );
  AND U2130 ( .A(n1990), .B(n1989), .Z(n2074) );
  XNOR U2131 ( .A(n2075), .B(n2074), .Z(n2076) );
  NANDN U2132 ( .A(n1992), .B(n1991), .Z(n1996) );
  NANDN U2133 ( .A(n1994), .B(n1993), .Z(n1995) );
  NAND U2134 ( .A(n1996), .B(n1995), .Z(n2077) );
  XNOR U2135 ( .A(n2076), .B(n2077), .Z(n2022) );
  XOR U2136 ( .A(n2023), .B(n2022), .Z(n2081) );
  NANDN U2137 ( .A(n1998), .B(n1997), .Z(n2002) );
  NANDN U2138 ( .A(n2000), .B(n1999), .Z(n2001) );
  AND U2139 ( .A(n2002), .B(n2001), .Z(n2080) );
  XNOR U2140 ( .A(n2081), .B(n2080), .Z(n2082) );
  XOR U2141 ( .A(n2083), .B(n2082), .Z(n2015) );
  NANDN U2142 ( .A(n2004), .B(n2003), .Z(n2008) );
  NAND U2143 ( .A(n2006), .B(n2005), .Z(n2007) );
  AND U2144 ( .A(n2008), .B(n2007), .Z(n2014) );
  XNOR U2145 ( .A(n2015), .B(n2014), .Z(n2016) );
  XNOR U2146 ( .A(n2017), .B(n2016), .Z(n2086) );
  XNOR U2147 ( .A(sreg[145]), .B(n2086), .Z(n2088) );
  NANDN U2148 ( .A(sreg[144]), .B(n2009), .Z(n2013) );
  NAND U2149 ( .A(n2011), .B(n2010), .Z(n2012) );
  NAND U2150 ( .A(n2013), .B(n2012), .Z(n2087) );
  XNOR U2151 ( .A(n2088), .B(n2087), .Z(c[145]) );
  NANDN U2152 ( .A(n2015), .B(n2014), .Z(n2019) );
  NANDN U2153 ( .A(n2017), .B(n2016), .Z(n2018) );
  AND U2154 ( .A(n2019), .B(n2018), .Z(n2094) );
  NANDN U2155 ( .A(n2021), .B(n2020), .Z(n2025) );
  NAND U2156 ( .A(n2023), .B(n2022), .Z(n2024) );
  AND U2157 ( .A(n2025), .B(n2024), .Z(n2160) );
  NANDN U2158 ( .A(n2027), .B(n2026), .Z(n2031) );
  NANDN U2159 ( .A(n2029), .B(n2028), .Z(n2030) );
  AND U2160 ( .A(n2031), .B(n2030), .Z(n2126) );
  NAND U2161 ( .A(b[0]), .B(a[34]), .Z(n2032) );
  XNOR U2162 ( .A(b[1]), .B(n2032), .Z(n2034) );
  NANDN U2163 ( .A(b[0]), .B(a[33]), .Z(n2033) );
  NAND U2164 ( .A(n2034), .B(n2033), .Z(n2106) );
  NANDN U2165 ( .A(n9891), .B(n2035), .Z(n2037) );
  XOR U2166 ( .A(b[13]), .B(a[22]), .Z(n2112) );
  NANDN U2167 ( .A(n9935), .B(n2112), .Z(n2036) );
  AND U2168 ( .A(n2037), .B(n2036), .Z(n2104) );
  AND U2169 ( .A(b[15]), .B(a[18]), .Z(n2103) );
  XNOR U2170 ( .A(n2104), .B(n2103), .Z(n2105) );
  XNOR U2171 ( .A(n2106), .B(n2105), .Z(n2124) );
  NANDN U2172 ( .A(n9437), .B(n2038), .Z(n2040) );
  XOR U2173 ( .A(b[5]), .B(a[30]), .Z(n2115) );
  NANDN U2174 ( .A(n9503), .B(n2115), .Z(n2039) );
  AND U2175 ( .A(n2040), .B(n2039), .Z(n2148) );
  NANDN U2176 ( .A(n9588), .B(n2041), .Z(n2043) );
  XOR U2177 ( .A(b[7]), .B(a[28]), .Z(n2118) );
  NANDN U2178 ( .A(n9639), .B(n2118), .Z(n2042) );
  AND U2179 ( .A(n2043), .B(n2042), .Z(n2146) );
  NANDN U2180 ( .A(n9374), .B(n2044), .Z(n2046) );
  XOR U2181 ( .A(b[3]), .B(a[32]), .Z(n2121) );
  NANDN U2182 ( .A(n9375), .B(n2121), .Z(n2045) );
  NAND U2183 ( .A(n2046), .B(n2045), .Z(n2145) );
  XNOR U2184 ( .A(n2146), .B(n2145), .Z(n2147) );
  XOR U2185 ( .A(n2148), .B(n2147), .Z(n2125) );
  XOR U2186 ( .A(n2124), .B(n2125), .Z(n2127) );
  XOR U2187 ( .A(n2126), .B(n2127), .Z(n2098) );
  NANDN U2188 ( .A(n2048), .B(n2047), .Z(n2052) );
  OR U2189 ( .A(n2050), .B(n2049), .Z(n2051) );
  AND U2190 ( .A(n2052), .B(n2051), .Z(n2097) );
  XNOR U2191 ( .A(n2098), .B(n2097), .Z(n2100) );
  NAND U2192 ( .A(n2053), .B(n9883), .Z(n2055) );
  XOR U2193 ( .A(b[11]), .B(a[24]), .Z(n2130) );
  NANDN U2194 ( .A(n9856), .B(n2130), .Z(n2054) );
  AND U2195 ( .A(n2055), .B(n2054), .Z(n2141) );
  NANDN U2196 ( .A(n10005), .B(n2056), .Z(n2058) );
  XOR U2197 ( .A(b[15]), .B(a[20]), .Z(n2133) );
  NANDN U2198 ( .A(n10006), .B(n2133), .Z(n2057) );
  AND U2199 ( .A(n2058), .B(n2057), .Z(n2140) );
  NANDN U2200 ( .A(n9685), .B(n2059), .Z(n2061) );
  XOR U2201 ( .A(b[9]), .B(a[26]), .Z(n2136) );
  NANDN U2202 ( .A(n9758), .B(n2136), .Z(n2060) );
  NAND U2203 ( .A(n2061), .B(n2060), .Z(n2139) );
  XOR U2204 ( .A(n2140), .B(n2139), .Z(n2142) );
  XOR U2205 ( .A(n2141), .B(n2142), .Z(n2152) );
  NANDN U2206 ( .A(n2063), .B(n2062), .Z(n2067) );
  OR U2207 ( .A(n2065), .B(n2064), .Z(n2066) );
  AND U2208 ( .A(n2067), .B(n2066), .Z(n2151) );
  XNOR U2209 ( .A(n2152), .B(n2151), .Z(n2153) );
  NANDN U2210 ( .A(n2069), .B(n2068), .Z(n2073) );
  NANDN U2211 ( .A(n2071), .B(n2070), .Z(n2072) );
  NAND U2212 ( .A(n2073), .B(n2072), .Z(n2154) );
  XNOR U2213 ( .A(n2153), .B(n2154), .Z(n2099) );
  XOR U2214 ( .A(n2100), .B(n2099), .Z(n2158) );
  NANDN U2215 ( .A(n2075), .B(n2074), .Z(n2079) );
  NANDN U2216 ( .A(n2077), .B(n2076), .Z(n2078) );
  AND U2217 ( .A(n2079), .B(n2078), .Z(n2157) );
  XNOR U2218 ( .A(n2158), .B(n2157), .Z(n2159) );
  XOR U2219 ( .A(n2160), .B(n2159), .Z(n2092) );
  NANDN U2220 ( .A(n2081), .B(n2080), .Z(n2085) );
  NAND U2221 ( .A(n2083), .B(n2082), .Z(n2084) );
  AND U2222 ( .A(n2085), .B(n2084), .Z(n2091) );
  XNOR U2223 ( .A(n2092), .B(n2091), .Z(n2093) );
  XNOR U2224 ( .A(n2094), .B(n2093), .Z(n2163) );
  XNOR U2225 ( .A(sreg[146]), .B(n2163), .Z(n2165) );
  NANDN U2226 ( .A(sreg[145]), .B(n2086), .Z(n2090) );
  NAND U2227 ( .A(n2088), .B(n2087), .Z(n2089) );
  NAND U2228 ( .A(n2090), .B(n2089), .Z(n2164) );
  XNOR U2229 ( .A(n2165), .B(n2164), .Z(c[146]) );
  NANDN U2230 ( .A(n2092), .B(n2091), .Z(n2096) );
  NANDN U2231 ( .A(n2094), .B(n2093), .Z(n2095) );
  AND U2232 ( .A(n2096), .B(n2095), .Z(n2171) );
  NANDN U2233 ( .A(n2098), .B(n2097), .Z(n2102) );
  NAND U2234 ( .A(n2100), .B(n2099), .Z(n2101) );
  AND U2235 ( .A(n2102), .B(n2101), .Z(n2237) );
  NANDN U2236 ( .A(n2104), .B(n2103), .Z(n2108) );
  NANDN U2237 ( .A(n2106), .B(n2105), .Z(n2107) );
  AND U2238 ( .A(n2108), .B(n2107), .Z(n2224) );
  NAND U2239 ( .A(b[0]), .B(a[35]), .Z(n2109) );
  XNOR U2240 ( .A(b[1]), .B(n2109), .Z(n2111) );
  NANDN U2241 ( .A(b[0]), .B(a[34]), .Z(n2110) );
  NAND U2242 ( .A(n2111), .B(n2110), .Z(n2204) );
  NANDN U2243 ( .A(n9891), .B(n2112), .Z(n2114) );
  XOR U2244 ( .A(b[13]), .B(a[23]), .Z(n2210) );
  NANDN U2245 ( .A(n9935), .B(n2210), .Z(n2113) );
  AND U2246 ( .A(n2114), .B(n2113), .Z(n2202) );
  AND U2247 ( .A(b[15]), .B(a[19]), .Z(n2201) );
  XNOR U2248 ( .A(n2202), .B(n2201), .Z(n2203) );
  XNOR U2249 ( .A(n2204), .B(n2203), .Z(n2222) );
  NANDN U2250 ( .A(n9437), .B(n2115), .Z(n2117) );
  XOR U2251 ( .A(b[5]), .B(a[31]), .Z(n2213) );
  NANDN U2252 ( .A(n9503), .B(n2213), .Z(n2116) );
  AND U2253 ( .A(n2117), .B(n2116), .Z(n2198) );
  NANDN U2254 ( .A(n9588), .B(n2118), .Z(n2120) );
  XOR U2255 ( .A(b[7]), .B(a[29]), .Z(n2216) );
  NANDN U2256 ( .A(n9639), .B(n2216), .Z(n2119) );
  AND U2257 ( .A(n2120), .B(n2119), .Z(n2196) );
  NANDN U2258 ( .A(n9374), .B(n2121), .Z(n2123) );
  XOR U2259 ( .A(b[3]), .B(a[33]), .Z(n2219) );
  NANDN U2260 ( .A(n9375), .B(n2219), .Z(n2122) );
  NAND U2261 ( .A(n2123), .B(n2122), .Z(n2195) );
  XNOR U2262 ( .A(n2196), .B(n2195), .Z(n2197) );
  XOR U2263 ( .A(n2198), .B(n2197), .Z(n2223) );
  XOR U2264 ( .A(n2222), .B(n2223), .Z(n2225) );
  XOR U2265 ( .A(n2224), .B(n2225), .Z(n2175) );
  NANDN U2266 ( .A(n2125), .B(n2124), .Z(n2129) );
  OR U2267 ( .A(n2127), .B(n2126), .Z(n2128) );
  AND U2268 ( .A(n2129), .B(n2128), .Z(n2174) );
  XNOR U2269 ( .A(n2175), .B(n2174), .Z(n2177) );
  NAND U2270 ( .A(n2130), .B(n9883), .Z(n2132) );
  XOR U2271 ( .A(b[11]), .B(a[25]), .Z(n2180) );
  NANDN U2272 ( .A(n9856), .B(n2180), .Z(n2131) );
  AND U2273 ( .A(n2132), .B(n2131), .Z(n2191) );
  NANDN U2274 ( .A(n10005), .B(n2133), .Z(n2135) );
  XOR U2275 ( .A(b[15]), .B(a[21]), .Z(n2183) );
  NANDN U2276 ( .A(n10006), .B(n2183), .Z(n2134) );
  AND U2277 ( .A(n2135), .B(n2134), .Z(n2190) );
  NANDN U2278 ( .A(n9685), .B(n2136), .Z(n2138) );
  XOR U2279 ( .A(b[9]), .B(a[27]), .Z(n2186) );
  NANDN U2280 ( .A(n9758), .B(n2186), .Z(n2137) );
  NAND U2281 ( .A(n2138), .B(n2137), .Z(n2189) );
  XOR U2282 ( .A(n2190), .B(n2189), .Z(n2192) );
  XOR U2283 ( .A(n2191), .B(n2192), .Z(n2229) );
  NANDN U2284 ( .A(n2140), .B(n2139), .Z(n2144) );
  OR U2285 ( .A(n2142), .B(n2141), .Z(n2143) );
  AND U2286 ( .A(n2144), .B(n2143), .Z(n2228) );
  XNOR U2287 ( .A(n2229), .B(n2228), .Z(n2230) );
  NANDN U2288 ( .A(n2146), .B(n2145), .Z(n2150) );
  NANDN U2289 ( .A(n2148), .B(n2147), .Z(n2149) );
  NAND U2290 ( .A(n2150), .B(n2149), .Z(n2231) );
  XNOR U2291 ( .A(n2230), .B(n2231), .Z(n2176) );
  XOR U2292 ( .A(n2177), .B(n2176), .Z(n2235) );
  NANDN U2293 ( .A(n2152), .B(n2151), .Z(n2156) );
  NANDN U2294 ( .A(n2154), .B(n2153), .Z(n2155) );
  AND U2295 ( .A(n2156), .B(n2155), .Z(n2234) );
  XNOR U2296 ( .A(n2235), .B(n2234), .Z(n2236) );
  XOR U2297 ( .A(n2237), .B(n2236), .Z(n2169) );
  NANDN U2298 ( .A(n2158), .B(n2157), .Z(n2162) );
  NAND U2299 ( .A(n2160), .B(n2159), .Z(n2161) );
  AND U2300 ( .A(n2162), .B(n2161), .Z(n2168) );
  XNOR U2301 ( .A(n2169), .B(n2168), .Z(n2170) );
  XNOR U2302 ( .A(n2171), .B(n2170), .Z(n2240) );
  XNOR U2303 ( .A(sreg[147]), .B(n2240), .Z(n2242) );
  NANDN U2304 ( .A(sreg[146]), .B(n2163), .Z(n2167) );
  NAND U2305 ( .A(n2165), .B(n2164), .Z(n2166) );
  NAND U2306 ( .A(n2167), .B(n2166), .Z(n2241) );
  XNOR U2307 ( .A(n2242), .B(n2241), .Z(c[147]) );
  NANDN U2308 ( .A(n2169), .B(n2168), .Z(n2173) );
  NANDN U2309 ( .A(n2171), .B(n2170), .Z(n2172) );
  AND U2310 ( .A(n2173), .B(n2172), .Z(n2248) );
  NANDN U2311 ( .A(n2175), .B(n2174), .Z(n2179) );
  NAND U2312 ( .A(n2177), .B(n2176), .Z(n2178) );
  AND U2313 ( .A(n2179), .B(n2178), .Z(n2314) );
  NAND U2314 ( .A(n2180), .B(n9883), .Z(n2182) );
  XOR U2315 ( .A(b[11]), .B(a[26]), .Z(n2284) );
  NANDN U2316 ( .A(n9856), .B(n2284), .Z(n2181) );
  AND U2317 ( .A(n2182), .B(n2181), .Z(n2295) );
  NANDN U2318 ( .A(n10005), .B(n2183), .Z(n2185) );
  XOR U2319 ( .A(b[15]), .B(a[22]), .Z(n2287) );
  NANDN U2320 ( .A(n10006), .B(n2287), .Z(n2184) );
  AND U2321 ( .A(n2185), .B(n2184), .Z(n2294) );
  NANDN U2322 ( .A(n9685), .B(n2186), .Z(n2188) );
  XOR U2323 ( .A(b[9]), .B(a[28]), .Z(n2290) );
  NANDN U2324 ( .A(n9758), .B(n2290), .Z(n2187) );
  NAND U2325 ( .A(n2188), .B(n2187), .Z(n2293) );
  XOR U2326 ( .A(n2294), .B(n2293), .Z(n2296) );
  XOR U2327 ( .A(n2295), .B(n2296), .Z(n2306) );
  NANDN U2328 ( .A(n2190), .B(n2189), .Z(n2194) );
  OR U2329 ( .A(n2192), .B(n2191), .Z(n2193) );
  AND U2330 ( .A(n2194), .B(n2193), .Z(n2305) );
  XNOR U2331 ( .A(n2306), .B(n2305), .Z(n2307) );
  NANDN U2332 ( .A(n2196), .B(n2195), .Z(n2200) );
  NANDN U2333 ( .A(n2198), .B(n2197), .Z(n2199) );
  NAND U2334 ( .A(n2200), .B(n2199), .Z(n2308) );
  XNOR U2335 ( .A(n2307), .B(n2308), .Z(n2254) );
  NANDN U2336 ( .A(n2202), .B(n2201), .Z(n2206) );
  NANDN U2337 ( .A(n2204), .B(n2203), .Z(n2205) );
  AND U2338 ( .A(n2206), .B(n2205), .Z(n2280) );
  NAND U2339 ( .A(b[0]), .B(a[36]), .Z(n2207) );
  XNOR U2340 ( .A(b[1]), .B(n2207), .Z(n2209) );
  NANDN U2341 ( .A(b[0]), .B(a[35]), .Z(n2208) );
  NAND U2342 ( .A(n2209), .B(n2208), .Z(n2260) );
  NANDN U2343 ( .A(n9891), .B(n2210), .Z(n2212) );
  XOR U2344 ( .A(b[13]), .B(a[24]), .Z(n2266) );
  NANDN U2345 ( .A(n9935), .B(n2266), .Z(n2211) );
  AND U2346 ( .A(n2212), .B(n2211), .Z(n2258) );
  AND U2347 ( .A(b[15]), .B(a[20]), .Z(n2257) );
  XNOR U2348 ( .A(n2258), .B(n2257), .Z(n2259) );
  XNOR U2349 ( .A(n2260), .B(n2259), .Z(n2278) );
  NANDN U2350 ( .A(n9437), .B(n2213), .Z(n2215) );
  XOR U2351 ( .A(b[5]), .B(a[32]), .Z(n2269) );
  NANDN U2352 ( .A(n9503), .B(n2269), .Z(n2214) );
  AND U2353 ( .A(n2215), .B(n2214), .Z(n2302) );
  NANDN U2354 ( .A(n9588), .B(n2216), .Z(n2218) );
  XOR U2355 ( .A(b[7]), .B(a[30]), .Z(n2272) );
  NANDN U2356 ( .A(n9639), .B(n2272), .Z(n2217) );
  AND U2357 ( .A(n2218), .B(n2217), .Z(n2300) );
  NANDN U2358 ( .A(n9374), .B(n2219), .Z(n2221) );
  XOR U2359 ( .A(b[3]), .B(a[34]), .Z(n2275) );
  NANDN U2360 ( .A(n9375), .B(n2275), .Z(n2220) );
  NAND U2361 ( .A(n2221), .B(n2220), .Z(n2299) );
  XNOR U2362 ( .A(n2300), .B(n2299), .Z(n2301) );
  XOR U2363 ( .A(n2302), .B(n2301), .Z(n2279) );
  XOR U2364 ( .A(n2278), .B(n2279), .Z(n2281) );
  XOR U2365 ( .A(n2280), .B(n2281), .Z(n2252) );
  NANDN U2366 ( .A(n2223), .B(n2222), .Z(n2227) );
  OR U2367 ( .A(n2225), .B(n2224), .Z(n2226) );
  AND U2368 ( .A(n2227), .B(n2226), .Z(n2251) );
  XNOR U2369 ( .A(n2252), .B(n2251), .Z(n2253) );
  XOR U2370 ( .A(n2254), .B(n2253), .Z(n2312) );
  NANDN U2371 ( .A(n2229), .B(n2228), .Z(n2233) );
  NANDN U2372 ( .A(n2231), .B(n2230), .Z(n2232) );
  AND U2373 ( .A(n2233), .B(n2232), .Z(n2311) );
  XNOR U2374 ( .A(n2312), .B(n2311), .Z(n2313) );
  XOR U2375 ( .A(n2314), .B(n2313), .Z(n2246) );
  NANDN U2376 ( .A(n2235), .B(n2234), .Z(n2239) );
  NAND U2377 ( .A(n2237), .B(n2236), .Z(n2238) );
  AND U2378 ( .A(n2239), .B(n2238), .Z(n2245) );
  XNOR U2379 ( .A(n2246), .B(n2245), .Z(n2247) );
  XNOR U2380 ( .A(n2248), .B(n2247), .Z(n2317) );
  XNOR U2381 ( .A(sreg[148]), .B(n2317), .Z(n2319) );
  NANDN U2382 ( .A(sreg[147]), .B(n2240), .Z(n2244) );
  NAND U2383 ( .A(n2242), .B(n2241), .Z(n2243) );
  NAND U2384 ( .A(n2244), .B(n2243), .Z(n2318) );
  XNOR U2385 ( .A(n2319), .B(n2318), .Z(c[148]) );
  NANDN U2386 ( .A(n2246), .B(n2245), .Z(n2250) );
  NANDN U2387 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U2388 ( .A(n2250), .B(n2249), .Z(n2325) );
  NANDN U2389 ( .A(n2252), .B(n2251), .Z(n2256) );
  NAND U2390 ( .A(n2254), .B(n2253), .Z(n2255) );
  AND U2391 ( .A(n2256), .B(n2255), .Z(n2391) );
  NANDN U2392 ( .A(n2258), .B(n2257), .Z(n2262) );
  NANDN U2393 ( .A(n2260), .B(n2259), .Z(n2261) );
  AND U2394 ( .A(n2262), .B(n2261), .Z(n2357) );
  NAND U2395 ( .A(b[0]), .B(a[37]), .Z(n2263) );
  XNOR U2396 ( .A(b[1]), .B(n2263), .Z(n2265) );
  NANDN U2397 ( .A(b[0]), .B(a[36]), .Z(n2264) );
  NAND U2398 ( .A(n2265), .B(n2264), .Z(n2337) );
  NANDN U2399 ( .A(n9891), .B(n2266), .Z(n2268) );
  XOR U2400 ( .A(b[13]), .B(a[25]), .Z(n2343) );
  NANDN U2401 ( .A(n9935), .B(n2343), .Z(n2267) );
  AND U2402 ( .A(n2268), .B(n2267), .Z(n2335) );
  AND U2403 ( .A(b[15]), .B(a[21]), .Z(n2334) );
  XNOR U2404 ( .A(n2335), .B(n2334), .Z(n2336) );
  XNOR U2405 ( .A(n2337), .B(n2336), .Z(n2355) );
  NANDN U2406 ( .A(n9437), .B(n2269), .Z(n2271) );
  XOR U2407 ( .A(b[5]), .B(a[33]), .Z(n2346) );
  NANDN U2408 ( .A(n9503), .B(n2346), .Z(n2270) );
  AND U2409 ( .A(n2271), .B(n2270), .Z(n2379) );
  NANDN U2410 ( .A(n9588), .B(n2272), .Z(n2274) );
  XOR U2411 ( .A(b[7]), .B(a[31]), .Z(n2349) );
  NANDN U2412 ( .A(n9639), .B(n2349), .Z(n2273) );
  AND U2413 ( .A(n2274), .B(n2273), .Z(n2377) );
  NANDN U2414 ( .A(n9374), .B(n2275), .Z(n2277) );
  XOR U2415 ( .A(b[3]), .B(a[35]), .Z(n2352) );
  NANDN U2416 ( .A(n9375), .B(n2352), .Z(n2276) );
  NAND U2417 ( .A(n2277), .B(n2276), .Z(n2376) );
  XNOR U2418 ( .A(n2377), .B(n2376), .Z(n2378) );
  XOR U2419 ( .A(n2379), .B(n2378), .Z(n2356) );
  XOR U2420 ( .A(n2355), .B(n2356), .Z(n2358) );
  XOR U2421 ( .A(n2357), .B(n2358), .Z(n2329) );
  NANDN U2422 ( .A(n2279), .B(n2278), .Z(n2283) );
  OR U2423 ( .A(n2281), .B(n2280), .Z(n2282) );
  AND U2424 ( .A(n2283), .B(n2282), .Z(n2328) );
  XNOR U2425 ( .A(n2329), .B(n2328), .Z(n2331) );
  NAND U2426 ( .A(n2284), .B(n9883), .Z(n2286) );
  XOR U2427 ( .A(b[11]), .B(a[27]), .Z(n2361) );
  NANDN U2428 ( .A(n9856), .B(n2361), .Z(n2285) );
  AND U2429 ( .A(n2286), .B(n2285), .Z(n2372) );
  NANDN U2430 ( .A(n10005), .B(n2287), .Z(n2289) );
  XOR U2431 ( .A(b[15]), .B(a[23]), .Z(n2364) );
  NANDN U2432 ( .A(n10006), .B(n2364), .Z(n2288) );
  AND U2433 ( .A(n2289), .B(n2288), .Z(n2371) );
  NANDN U2434 ( .A(n9685), .B(n2290), .Z(n2292) );
  XOR U2435 ( .A(b[9]), .B(a[29]), .Z(n2367) );
  NANDN U2436 ( .A(n9758), .B(n2367), .Z(n2291) );
  NAND U2437 ( .A(n2292), .B(n2291), .Z(n2370) );
  XOR U2438 ( .A(n2371), .B(n2370), .Z(n2373) );
  XOR U2439 ( .A(n2372), .B(n2373), .Z(n2383) );
  NANDN U2440 ( .A(n2294), .B(n2293), .Z(n2298) );
  OR U2441 ( .A(n2296), .B(n2295), .Z(n2297) );
  AND U2442 ( .A(n2298), .B(n2297), .Z(n2382) );
  XNOR U2443 ( .A(n2383), .B(n2382), .Z(n2384) );
  NANDN U2444 ( .A(n2300), .B(n2299), .Z(n2304) );
  NANDN U2445 ( .A(n2302), .B(n2301), .Z(n2303) );
  NAND U2446 ( .A(n2304), .B(n2303), .Z(n2385) );
  XNOR U2447 ( .A(n2384), .B(n2385), .Z(n2330) );
  XOR U2448 ( .A(n2331), .B(n2330), .Z(n2389) );
  NANDN U2449 ( .A(n2306), .B(n2305), .Z(n2310) );
  NANDN U2450 ( .A(n2308), .B(n2307), .Z(n2309) );
  AND U2451 ( .A(n2310), .B(n2309), .Z(n2388) );
  XNOR U2452 ( .A(n2389), .B(n2388), .Z(n2390) );
  XOR U2453 ( .A(n2391), .B(n2390), .Z(n2323) );
  NANDN U2454 ( .A(n2312), .B(n2311), .Z(n2316) );
  NAND U2455 ( .A(n2314), .B(n2313), .Z(n2315) );
  AND U2456 ( .A(n2316), .B(n2315), .Z(n2322) );
  XNOR U2457 ( .A(n2323), .B(n2322), .Z(n2324) );
  XNOR U2458 ( .A(n2325), .B(n2324), .Z(n2394) );
  XNOR U2459 ( .A(sreg[149]), .B(n2394), .Z(n2396) );
  NANDN U2460 ( .A(sreg[148]), .B(n2317), .Z(n2321) );
  NAND U2461 ( .A(n2319), .B(n2318), .Z(n2320) );
  NAND U2462 ( .A(n2321), .B(n2320), .Z(n2395) );
  XNOR U2463 ( .A(n2396), .B(n2395), .Z(c[149]) );
  NANDN U2464 ( .A(n2323), .B(n2322), .Z(n2327) );
  NANDN U2465 ( .A(n2325), .B(n2324), .Z(n2326) );
  AND U2466 ( .A(n2327), .B(n2326), .Z(n2402) );
  NANDN U2467 ( .A(n2329), .B(n2328), .Z(n2333) );
  NAND U2468 ( .A(n2331), .B(n2330), .Z(n2332) );
  AND U2469 ( .A(n2333), .B(n2332), .Z(n2468) );
  NANDN U2470 ( .A(n2335), .B(n2334), .Z(n2339) );
  NANDN U2471 ( .A(n2337), .B(n2336), .Z(n2338) );
  AND U2472 ( .A(n2339), .B(n2338), .Z(n2434) );
  NAND U2473 ( .A(b[0]), .B(a[38]), .Z(n2340) );
  XNOR U2474 ( .A(b[1]), .B(n2340), .Z(n2342) );
  NANDN U2475 ( .A(b[0]), .B(a[37]), .Z(n2341) );
  NAND U2476 ( .A(n2342), .B(n2341), .Z(n2414) );
  NANDN U2477 ( .A(n9891), .B(n2343), .Z(n2345) );
  XOR U2478 ( .A(b[13]), .B(a[26]), .Z(n2420) );
  NANDN U2479 ( .A(n9935), .B(n2420), .Z(n2344) );
  AND U2480 ( .A(n2345), .B(n2344), .Z(n2412) );
  AND U2481 ( .A(b[15]), .B(a[22]), .Z(n2411) );
  XNOR U2482 ( .A(n2412), .B(n2411), .Z(n2413) );
  XNOR U2483 ( .A(n2414), .B(n2413), .Z(n2432) );
  NANDN U2484 ( .A(n9437), .B(n2346), .Z(n2348) );
  XOR U2485 ( .A(b[5]), .B(a[34]), .Z(n2423) );
  NANDN U2486 ( .A(n9503), .B(n2423), .Z(n2347) );
  AND U2487 ( .A(n2348), .B(n2347), .Z(n2456) );
  NANDN U2488 ( .A(n9588), .B(n2349), .Z(n2351) );
  XOR U2489 ( .A(b[7]), .B(a[32]), .Z(n2426) );
  NANDN U2490 ( .A(n9639), .B(n2426), .Z(n2350) );
  AND U2491 ( .A(n2351), .B(n2350), .Z(n2454) );
  NANDN U2492 ( .A(n9374), .B(n2352), .Z(n2354) );
  XOR U2493 ( .A(b[3]), .B(a[36]), .Z(n2429) );
  NANDN U2494 ( .A(n9375), .B(n2429), .Z(n2353) );
  NAND U2495 ( .A(n2354), .B(n2353), .Z(n2453) );
  XNOR U2496 ( .A(n2454), .B(n2453), .Z(n2455) );
  XOR U2497 ( .A(n2456), .B(n2455), .Z(n2433) );
  XOR U2498 ( .A(n2432), .B(n2433), .Z(n2435) );
  XOR U2499 ( .A(n2434), .B(n2435), .Z(n2406) );
  NANDN U2500 ( .A(n2356), .B(n2355), .Z(n2360) );
  OR U2501 ( .A(n2358), .B(n2357), .Z(n2359) );
  AND U2502 ( .A(n2360), .B(n2359), .Z(n2405) );
  XNOR U2503 ( .A(n2406), .B(n2405), .Z(n2408) );
  NAND U2504 ( .A(n2361), .B(n9883), .Z(n2363) );
  XOR U2505 ( .A(b[11]), .B(a[28]), .Z(n2438) );
  NANDN U2506 ( .A(n9856), .B(n2438), .Z(n2362) );
  AND U2507 ( .A(n2363), .B(n2362), .Z(n2449) );
  NANDN U2508 ( .A(n10005), .B(n2364), .Z(n2366) );
  XOR U2509 ( .A(b[15]), .B(a[24]), .Z(n2441) );
  NANDN U2510 ( .A(n10006), .B(n2441), .Z(n2365) );
  AND U2511 ( .A(n2366), .B(n2365), .Z(n2448) );
  NANDN U2512 ( .A(n9685), .B(n2367), .Z(n2369) );
  XOR U2513 ( .A(b[9]), .B(a[30]), .Z(n2444) );
  NANDN U2514 ( .A(n9758), .B(n2444), .Z(n2368) );
  NAND U2515 ( .A(n2369), .B(n2368), .Z(n2447) );
  XOR U2516 ( .A(n2448), .B(n2447), .Z(n2450) );
  XOR U2517 ( .A(n2449), .B(n2450), .Z(n2460) );
  NANDN U2518 ( .A(n2371), .B(n2370), .Z(n2375) );
  OR U2519 ( .A(n2373), .B(n2372), .Z(n2374) );
  AND U2520 ( .A(n2375), .B(n2374), .Z(n2459) );
  XNOR U2521 ( .A(n2460), .B(n2459), .Z(n2461) );
  NANDN U2522 ( .A(n2377), .B(n2376), .Z(n2381) );
  NANDN U2523 ( .A(n2379), .B(n2378), .Z(n2380) );
  NAND U2524 ( .A(n2381), .B(n2380), .Z(n2462) );
  XNOR U2525 ( .A(n2461), .B(n2462), .Z(n2407) );
  XOR U2526 ( .A(n2408), .B(n2407), .Z(n2466) );
  NANDN U2527 ( .A(n2383), .B(n2382), .Z(n2387) );
  NANDN U2528 ( .A(n2385), .B(n2384), .Z(n2386) );
  AND U2529 ( .A(n2387), .B(n2386), .Z(n2465) );
  XNOR U2530 ( .A(n2466), .B(n2465), .Z(n2467) );
  XOR U2531 ( .A(n2468), .B(n2467), .Z(n2400) );
  NANDN U2532 ( .A(n2389), .B(n2388), .Z(n2393) );
  NAND U2533 ( .A(n2391), .B(n2390), .Z(n2392) );
  AND U2534 ( .A(n2393), .B(n2392), .Z(n2399) );
  XNOR U2535 ( .A(n2400), .B(n2399), .Z(n2401) );
  XNOR U2536 ( .A(n2402), .B(n2401), .Z(n2471) );
  XNOR U2537 ( .A(sreg[150]), .B(n2471), .Z(n2473) );
  NANDN U2538 ( .A(sreg[149]), .B(n2394), .Z(n2398) );
  NAND U2539 ( .A(n2396), .B(n2395), .Z(n2397) );
  NAND U2540 ( .A(n2398), .B(n2397), .Z(n2472) );
  XNOR U2541 ( .A(n2473), .B(n2472), .Z(c[150]) );
  NANDN U2542 ( .A(n2400), .B(n2399), .Z(n2404) );
  NANDN U2543 ( .A(n2402), .B(n2401), .Z(n2403) );
  AND U2544 ( .A(n2404), .B(n2403), .Z(n2479) );
  NANDN U2545 ( .A(n2406), .B(n2405), .Z(n2410) );
  NAND U2546 ( .A(n2408), .B(n2407), .Z(n2409) );
  AND U2547 ( .A(n2410), .B(n2409), .Z(n2545) );
  NANDN U2548 ( .A(n2412), .B(n2411), .Z(n2416) );
  NANDN U2549 ( .A(n2414), .B(n2413), .Z(n2415) );
  AND U2550 ( .A(n2416), .B(n2415), .Z(n2511) );
  NAND U2551 ( .A(b[0]), .B(a[39]), .Z(n2417) );
  XNOR U2552 ( .A(b[1]), .B(n2417), .Z(n2419) );
  NANDN U2553 ( .A(b[0]), .B(a[38]), .Z(n2418) );
  NAND U2554 ( .A(n2419), .B(n2418), .Z(n2491) );
  NANDN U2555 ( .A(n9891), .B(n2420), .Z(n2422) );
  XOR U2556 ( .A(b[13]), .B(a[27]), .Z(n2497) );
  NANDN U2557 ( .A(n9935), .B(n2497), .Z(n2421) );
  AND U2558 ( .A(n2422), .B(n2421), .Z(n2489) );
  AND U2559 ( .A(b[15]), .B(a[23]), .Z(n2488) );
  XNOR U2560 ( .A(n2489), .B(n2488), .Z(n2490) );
  XNOR U2561 ( .A(n2491), .B(n2490), .Z(n2509) );
  NANDN U2562 ( .A(n9437), .B(n2423), .Z(n2425) );
  XOR U2563 ( .A(b[5]), .B(a[35]), .Z(n2500) );
  NANDN U2564 ( .A(n9503), .B(n2500), .Z(n2424) );
  AND U2565 ( .A(n2425), .B(n2424), .Z(n2533) );
  NANDN U2566 ( .A(n9588), .B(n2426), .Z(n2428) );
  XOR U2567 ( .A(b[7]), .B(a[33]), .Z(n2503) );
  NANDN U2568 ( .A(n9639), .B(n2503), .Z(n2427) );
  AND U2569 ( .A(n2428), .B(n2427), .Z(n2531) );
  NANDN U2570 ( .A(n9374), .B(n2429), .Z(n2431) );
  XOR U2571 ( .A(b[3]), .B(a[37]), .Z(n2506) );
  NANDN U2572 ( .A(n9375), .B(n2506), .Z(n2430) );
  NAND U2573 ( .A(n2431), .B(n2430), .Z(n2530) );
  XNOR U2574 ( .A(n2531), .B(n2530), .Z(n2532) );
  XOR U2575 ( .A(n2533), .B(n2532), .Z(n2510) );
  XOR U2576 ( .A(n2509), .B(n2510), .Z(n2512) );
  XOR U2577 ( .A(n2511), .B(n2512), .Z(n2483) );
  NANDN U2578 ( .A(n2433), .B(n2432), .Z(n2437) );
  OR U2579 ( .A(n2435), .B(n2434), .Z(n2436) );
  AND U2580 ( .A(n2437), .B(n2436), .Z(n2482) );
  XNOR U2581 ( .A(n2483), .B(n2482), .Z(n2485) );
  NAND U2582 ( .A(n2438), .B(n9883), .Z(n2440) );
  XOR U2583 ( .A(b[11]), .B(a[29]), .Z(n2515) );
  NANDN U2584 ( .A(n9856), .B(n2515), .Z(n2439) );
  AND U2585 ( .A(n2440), .B(n2439), .Z(n2526) );
  NANDN U2586 ( .A(n10005), .B(n2441), .Z(n2443) );
  XOR U2587 ( .A(b[15]), .B(a[25]), .Z(n2518) );
  NANDN U2588 ( .A(n10006), .B(n2518), .Z(n2442) );
  AND U2589 ( .A(n2443), .B(n2442), .Z(n2525) );
  NANDN U2590 ( .A(n9685), .B(n2444), .Z(n2446) );
  XOR U2591 ( .A(b[9]), .B(a[31]), .Z(n2521) );
  NANDN U2592 ( .A(n9758), .B(n2521), .Z(n2445) );
  NAND U2593 ( .A(n2446), .B(n2445), .Z(n2524) );
  XOR U2594 ( .A(n2525), .B(n2524), .Z(n2527) );
  XOR U2595 ( .A(n2526), .B(n2527), .Z(n2537) );
  NANDN U2596 ( .A(n2448), .B(n2447), .Z(n2452) );
  OR U2597 ( .A(n2450), .B(n2449), .Z(n2451) );
  AND U2598 ( .A(n2452), .B(n2451), .Z(n2536) );
  XNOR U2599 ( .A(n2537), .B(n2536), .Z(n2538) );
  NANDN U2600 ( .A(n2454), .B(n2453), .Z(n2458) );
  NANDN U2601 ( .A(n2456), .B(n2455), .Z(n2457) );
  NAND U2602 ( .A(n2458), .B(n2457), .Z(n2539) );
  XNOR U2603 ( .A(n2538), .B(n2539), .Z(n2484) );
  XOR U2604 ( .A(n2485), .B(n2484), .Z(n2543) );
  NANDN U2605 ( .A(n2460), .B(n2459), .Z(n2464) );
  NANDN U2606 ( .A(n2462), .B(n2461), .Z(n2463) );
  AND U2607 ( .A(n2464), .B(n2463), .Z(n2542) );
  XNOR U2608 ( .A(n2543), .B(n2542), .Z(n2544) );
  XOR U2609 ( .A(n2545), .B(n2544), .Z(n2477) );
  NANDN U2610 ( .A(n2466), .B(n2465), .Z(n2470) );
  NAND U2611 ( .A(n2468), .B(n2467), .Z(n2469) );
  AND U2612 ( .A(n2470), .B(n2469), .Z(n2476) );
  XNOR U2613 ( .A(n2477), .B(n2476), .Z(n2478) );
  XNOR U2614 ( .A(n2479), .B(n2478), .Z(n2548) );
  XNOR U2615 ( .A(sreg[151]), .B(n2548), .Z(n2550) );
  NANDN U2616 ( .A(sreg[150]), .B(n2471), .Z(n2475) );
  NAND U2617 ( .A(n2473), .B(n2472), .Z(n2474) );
  NAND U2618 ( .A(n2475), .B(n2474), .Z(n2549) );
  XNOR U2619 ( .A(n2550), .B(n2549), .Z(c[151]) );
  NANDN U2620 ( .A(n2477), .B(n2476), .Z(n2481) );
  NANDN U2621 ( .A(n2479), .B(n2478), .Z(n2480) );
  AND U2622 ( .A(n2481), .B(n2480), .Z(n2556) );
  NANDN U2623 ( .A(n2483), .B(n2482), .Z(n2487) );
  NAND U2624 ( .A(n2485), .B(n2484), .Z(n2486) );
  AND U2625 ( .A(n2487), .B(n2486), .Z(n2622) );
  NANDN U2626 ( .A(n2489), .B(n2488), .Z(n2493) );
  NANDN U2627 ( .A(n2491), .B(n2490), .Z(n2492) );
  AND U2628 ( .A(n2493), .B(n2492), .Z(n2588) );
  NAND U2629 ( .A(b[0]), .B(a[40]), .Z(n2494) );
  XNOR U2630 ( .A(b[1]), .B(n2494), .Z(n2496) );
  NANDN U2631 ( .A(b[0]), .B(a[39]), .Z(n2495) );
  NAND U2632 ( .A(n2496), .B(n2495), .Z(n2568) );
  NANDN U2633 ( .A(n9891), .B(n2497), .Z(n2499) );
  XOR U2634 ( .A(b[13]), .B(a[28]), .Z(n2574) );
  NANDN U2635 ( .A(n9935), .B(n2574), .Z(n2498) );
  AND U2636 ( .A(n2499), .B(n2498), .Z(n2566) );
  AND U2637 ( .A(b[15]), .B(a[24]), .Z(n2565) );
  XNOR U2638 ( .A(n2566), .B(n2565), .Z(n2567) );
  XNOR U2639 ( .A(n2568), .B(n2567), .Z(n2586) );
  NANDN U2640 ( .A(n9437), .B(n2500), .Z(n2502) );
  XOR U2641 ( .A(b[5]), .B(a[36]), .Z(n2577) );
  NANDN U2642 ( .A(n9503), .B(n2577), .Z(n2501) );
  AND U2643 ( .A(n2502), .B(n2501), .Z(n2610) );
  NANDN U2644 ( .A(n9588), .B(n2503), .Z(n2505) );
  XOR U2645 ( .A(b[7]), .B(a[34]), .Z(n2580) );
  NANDN U2646 ( .A(n9639), .B(n2580), .Z(n2504) );
  AND U2647 ( .A(n2505), .B(n2504), .Z(n2608) );
  NANDN U2648 ( .A(n9374), .B(n2506), .Z(n2508) );
  XOR U2649 ( .A(b[3]), .B(a[38]), .Z(n2583) );
  NANDN U2650 ( .A(n9375), .B(n2583), .Z(n2507) );
  NAND U2651 ( .A(n2508), .B(n2507), .Z(n2607) );
  XNOR U2652 ( .A(n2608), .B(n2607), .Z(n2609) );
  XOR U2653 ( .A(n2610), .B(n2609), .Z(n2587) );
  XOR U2654 ( .A(n2586), .B(n2587), .Z(n2589) );
  XOR U2655 ( .A(n2588), .B(n2589), .Z(n2560) );
  NANDN U2656 ( .A(n2510), .B(n2509), .Z(n2514) );
  OR U2657 ( .A(n2512), .B(n2511), .Z(n2513) );
  AND U2658 ( .A(n2514), .B(n2513), .Z(n2559) );
  XNOR U2659 ( .A(n2560), .B(n2559), .Z(n2562) );
  NAND U2660 ( .A(n2515), .B(n9883), .Z(n2517) );
  XOR U2661 ( .A(b[11]), .B(a[30]), .Z(n2592) );
  NANDN U2662 ( .A(n9856), .B(n2592), .Z(n2516) );
  AND U2663 ( .A(n2517), .B(n2516), .Z(n2603) );
  NANDN U2664 ( .A(n10005), .B(n2518), .Z(n2520) );
  XOR U2665 ( .A(b[15]), .B(a[26]), .Z(n2595) );
  NANDN U2666 ( .A(n10006), .B(n2595), .Z(n2519) );
  AND U2667 ( .A(n2520), .B(n2519), .Z(n2602) );
  NANDN U2668 ( .A(n9685), .B(n2521), .Z(n2523) );
  XOR U2669 ( .A(b[9]), .B(a[32]), .Z(n2598) );
  NANDN U2670 ( .A(n9758), .B(n2598), .Z(n2522) );
  NAND U2671 ( .A(n2523), .B(n2522), .Z(n2601) );
  XOR U2672 ( .A(n2602), .B(n2601), .Z(n2604) );
  XOR U2673 ( .A(n2603), .B(n2604), .Z(n2614) );
  NANDN U2674 ( .A(n2525), .B(n2524), .Z(n2529) );
  OR U2675 ( .A(n2527), .B(n2526), .Z(n2528) );
  AND U2676 ( .A(n2529), .B(n2528), .Z(n2613) );
  XNOR U2677 ( .A(n2614), .B(n2613), .Z(n2615) );
  NANDN U2678 ( .A(n2531), .B(n2530), .Z(n2535) );
  NANDN U2679 ( .A(n2533), .B(n2532), .Z(n2534) );
  NAND U2680 ( .A(n2535), .B(n2534), .Z(n2616) );
  XNOR U2681 ( .A(n2615), .B(n2616), .Z(n2561) );
  XOR U2682 ( .A(n2562), .B(n2561), .Z(n2620) );
  NANDN U2683 ( .A(n2537), .B(n2536), .Z(n2541) );
  NANDN U2684 ( .A(n2539), .B(n2538), .Z(n2540) );
  AND U2685 ( .A(n2541), .B(n2540), .Z(n2619) );
  XNOR U2686 ( .A(n2620), .B(n2619), .Z(n2621) );
  XOR U2687 ( .A(n2622), .B(n2621), .Z(n2554) );
  NANDN U2688 ( .A(n2543), .B(n2542), .Z(n2547) );
  NAND U2689 ( .A(n2545), .B(n2544), .Z(n2546) );
  AND U2690 ( .A(n2547), .B(n2546), .Z(n2553) );
  XNOR U2691 ( .A(n2554), .B(n2553), .Z(n2555) );
  XNOR U2692 ( .A(n2556), .B(n2555), .Z(n2625) );
  XNOR U2693 ( .A(sreg[152]), .B(n2625), .Z(n2627) );
  NANDN U2694 ( .A(sreg[151]), .B(n2548), .Z(n2552) );
  NAND U2695 ( .A(n2550), .B(n2549), .Z(n2551) );
  NAND U2696 ( .A(n2552), .B(n2551), .Z(n2626) );
  XNOR U2697 ( .A(n2627), .B(n2626), .Z(c[152]) );
  NANDN U2698 ( .A(n2554), .B(n2553), .Z(n2558) );
  NANDN U2699 ( .A(n2556), .B(n2555), .Z(n2557) );
  AND U2700 ( .A(n2558), .B(n2557), .Z(n2633) );
  NANDN U2701 ( .A(n2560), .B(n2559), .Z(n2564) );
  NAND U2702 ( .A(n2562), .B(n2561), .Z(n2563) );
  AND U2703 ( .A(n2564), .B(n2563), .Z(n2699) );
  NANDN U2704 ( .A(n2566), .B(n2565), .Z(n2570) );
  NANDN U2705 ( .A(n2568), .B(n2567), .Z(n2569) );
  AND U2706 ( .A(n2570), .B(n2569), .Z(n2665) );
  NAND U2707 ( .A(b[0]), .B(a[41]), .Z(n2571) );
  XNOR U2708 ( .A(b[1]), .B(n2571), .Z(n2573) );
  NANDN U2709 ( .A(b[0]), .B(a[40]), .Z(n2572) );
  NAND U2710 ( .A(n2573), .B(n2572), .Z(n2645) );
  NANDN U2711 ( .A(n9891), .B(n2574), .Z(n2576) );
  XOR U2712 ( .A(b[13]), .B(a[29]), .Z(n2651) );
  NANDN U2713 ( .A(n9935), .B(n2651), .Z(n2575) );
  AND U2714 ( .A(n2576), .B(n2575), .Z(n2643) );
  AND U2715 ( .A(b[15]), .B(a[25]), .Z(n2642) );
  XNOR U2716 ( .A(n2643), .B(n2642), .Z(n2644) );
  XNOR U2717 ( .A(n2645), .B(n2644), .Z(n2663) );
  NANDN U2718 ( .A(n9437), .B(n2577), .Z(n2579) );
  XOR U2719 ( .A(b[5]), .B(a[37]), .Z(n2654) );
  NANDN U2720 ( .A(n9503), .B(n2654), .Z(n2578) );
  AND U2721 ( .A(n2579), .B(n2578), .Z(n2687) );
  NANDN U2722 ( .A(n9588), .B(n2580), .Z(n2582) );
  XOR U2723 ( .A(b[7]), .B(a[35]), .Z(n2657) );
  NANDN U2724 ( .A(n9639), .B(n2657), .Z(n2581) );
  AND U2725 ( .A(n2582), .B(n2581), .Z(n2685) );
  NANDN U2726 ( .A(n9374), .B(n2583), .Z(n2585) );
  XOR U2727 ( .A(b[3]), .B(a[39]), .Z(n2660) );
  NANDN U2728 ( .A(n9375), .B(n2660), .Z(n2584) );
  NAND U2729 ( .A(n2585), .B(n2584), .Z(n2684) );
  XNOR U2730 ( .A(n2685), .B(n2684), .Z(n2686) );
  XOR U2731 ( .A(n2687), .B(n2686), .Z(n2664) );
  XOR U2732 ( .A(n2663), .B(n2664), .Z(n2666) );
  XOR U2733 ( .A(n2665), .B(n2666), .Z(n2637) );
  NANDN U2734 ( .A(n2587), .B(n2586), .Z(n2591) );
  OR U2735 ( .A(n2589), .B(n2588), .Z(n2590) );
  AND U2736 ( .A(n2591), .B(n2590), .Z(n2636) );
  XNOR U2737 ( .A(n2637), .B(n2636), .Z(n2639) );
  NAND U2738 ( .A(n2592), .B(n9883), .Z(n2594) );
  XOR U2739 ( .A(b[11]), .B(a[31]), .Z(n2669) );
  NANDN U2740 ( .A(n9856), .B(n2669), .Z(n2593) );
  AND U2741 ( .A(n2594), .B(n2593), .Z(n2680) );
  NANDN U2742 ( .A(n10005), .B(n2595), .Z(n2597) );
  XOR U2743 ( .A(b[15]), .B(a[27]), .Z(n2672) );
  NANDN U2744 ( .A(n10006), .B(n2672), .Z(n2596) );
  AND U2745 ( .A(n2597), .B(n2596), .Z(n2679) );
  NANDN U2746 ( .A(n9685), .B(n2598), .Z(n2600) );
  XOR U2747 ( .A(b[9]), .B(a[33]), .Z(n2675) );
  NANDN U2748 ( .A(n9758), .B(n2675), .Z(n2599) );
  NAND U2749 ( .A(n2600), .B(n2599), .Z(n2678) );
  XOR U2750 ( .A(n2679), .B(n2678), .Z(n2681) );
  XOR U2751 ( .A(n2680), .B(n2681), .Z(n2691) );
  NANDN U2752 ( .A(n2602), .B(n2601), .Z(n2606) );
  OR U2753 ( .A(n2604), .B(n2603), .Z(n2605) );
  AND U2754 ( .A(n2606), .B(n2605), .Z(n2690) );
  XNOR U2755 ( .A(n2691), .B(n2690), .Z(n2692) );
  NANDN U2756 ( .A(n2608), .B(n2607), .Z(n2612) );
  NANDN U2757 ( .A(n2610), .B(n2609), .Z(n2611) );
  NAND U2758 ( .A(n2612), .B(n2611), .Z(n2693) );
  XNOR U2759 ( .A(n2692), .B(n2693), .Z(n2638) );
  XOR U2760 ( .A(n2639), .B(n2638), .Z(n2697) );
  NANDN U2761 ( .A(n2614), .B(n2613), .Z(n2618) );
  NANDN U2762 ( .A(n2616), .B(n2615), .Z(n2617) );
  AND U2763 ( .A(n2618), .B(n2617), .Z(n2696) );
  XNOR U2764 ( .A(n2697), .B(n2696), .Z(n2698) );
  XOR U2765 ( .A(n2699), .B(n2698), .Z(n2631) );
  NANDN U2766 ( .A(n2620), .B(n2619), .Z(n2624) );
  NAND U2767 ( .A(n2622), .B(n2621), .Z(n2623) );
  AND U2768 ( .A(n2624), .B(n2623), .Z(n2630) );
  XNOR U2769 ( .A(n2631), .B(n2630), .Z(n2632) );
  XNOR U2770 ( .A(n2633), .B(n2632), .Z(n2702) );
  XNOR U2771 ( .A(sreg[153]), .B(n2702), .Z(n2704) );
  NANDN U2772 ( .A(sreg[152]), .B(n2625), .Z(n2629) );
  NAND U2773 ( .A(n2627), .B(n2626), .Z(n2628) );
  NAND U2774 ( .A(n2629), .B(n2628), .Z(n2703) );
  XNOR U2775 ( .A(n2704), .B(n2703), .Z(c[153]) );
  NANDN U2776 ( .A(n2631), .B(n2630), .Z(n2635) );
  NANDN U2777 ( .A(n2633), .B(n2632), .Z(n2634) );
  AND U2778 ( .A(n2635), .B(n2634), .Z(n2710) );
  NANDN U2779 ( .A(n2637), .B(n2636), .Z(n2641) );
  NAND U2780 ( .A(n2639), .B(n2638), .Z(n2640) );
  AND U2781 ( .A(n2641), .B(n2640), .Z(n2776) );
  NANDN U2782 ( .A(n2643), .B(n2642), .Z(n2647) );
  NANDN U2783 ( .A(n2645), .B(n2644), .Z(n2646) );
  AND U2784 ( .A(n2647), .B(n2646), .Z(n2742) );
  NAND U2785 ( .A(b[0]), .B(a[42]), .Z(n2648) );
  XNOR U2786 ( .A(b[1]), .B(n2648), .Z(n2650) );
  NANDN U2787 ( .A(b[0]), .B(a[41]), .Z(n2649) );
  NAND U2788 ( .A(n2650), .B(n2649), .Z(n2722) );
  NANDN U2789 ( .A(n9891), .B(n2651), .Z(n2653) );
  XOR U2790 ( .A(b[13]), .B(a[30]), .Z(n2725) );
  NANDN U2791 ( .A(n9935), .B(n2725), .Z(n2652) );
  AND U2792 ( .A(n2653), .B(n2652), .Z(n2720) );
  AND U2793 ( .A(b[15]), .B(a[26]), .Z(n2719) );
  XNOR U2794 ( .A(n2720), .B(n2719), .Z(n2721) );
  XNOR U2795 ( .A(n2722), .B(n2721), .Z(n2740) );
  NANDN U2796 ( .A(n9437), .B(n2654), .Z(n2656) );
  XOR U2797 ( .A(b[5]), .B(a[38]), .Z(n2731) );
  NANDN U2798 ( .A(n9503), .B(n2731), .Z(n2655) );
  AND U2799 ( .A(n2656), .B(n2655), .Z(n2764) );
  NANDN U2800 ( .A(n9588), .B(n2657), .Z(n2659) );
  XOR U2801 ( .A(b[7]), .B(a[36]), .Z(n2734) );
  NANDN U2802 ( .A(n9639), .B(n2734), .Z(n2658) );
  AND U2803 ( .A(n2659), .B(n2658), .Z(n2762) );
  NANDN U2804 ( .A(n9374), .B(n2660), .Z(n2662) );
  XOR U2805 ( .A(b[3]), .B(a[40]), .Z(n2737) );
  NANDN U2806 ( .A(n9375), .B(n2737), .Z(n2661) );
  NAND U2807 ( .A(n2662), .B(n2661), .Z(n2761) );
  XNOR U2808 ( .A(n2762), .B(n2761), .Z(n2763) );
  XOR U2809 ( .A(n2764), .B(n2763), .Z(n2741) );
  XOR U2810 ( .A(n2740), .B(n2741), .Z(n2743) );
  XOR U2811 ( .A(n2742), .B(n2743), .Z(n2714) );
  NANDN U2812 ( .A(n2664), .B(n2663), .Z(n2668) );
  OR U2813 ( .A(n2666), .B(n2665), .Z(n2667) );
  AND U2814 ( .A(n2668), .B(n2667), .Z(n2713) );
  XNOR U2815 ( .A(n2714), .B(n2713), .Z(n2716) );
  NAND U2816 ( .A(n2669), .B(n9883), .Z(n2671) );
  XOR U2817 ( .A(b[11]), .B(a[32]), .Z(n2746) );
  NANDN U2818 ( .A(n9856), .B(n2746), .Z(n2670) );
  AND U2819 ( .A(n2671), .B(n2670), .Z(n2757) );
  NANDN U2820 ( .A(n10005), .B(n2672), .Z(n2674) );
  XOR U2821 ( .A(b[15]), .B(a[28]), .Z(n2749) );
  NANDN U2822 ( .A(n10006), .B(n2749), .Z(n2673) );
  AND U2823 ( .A(n2674), .B(n2673), .Z(n2756) );
  NANDN U2824 ( .A(n9685), .B(n2675), .Z(n2677) );
  XOR U2825 ( .A(b[9]), .B(a[34]), .Z(n2752) );
  NANDN U2826 ( .A(n9758), .B(n2752), .Z(n2676) );
  NAND U2827 ( .A(n2677), .B(n2676), .Z(n2755) );
  XOR U2828 ( .A(n2756), .B(n2755), .Z(n2758) );
  XOR U2829 ( .A(n2757), .B(n2758), .Z(n2768) );
  NANDN U2830 ( .A(n2679), .B(n2678), .Z(n2683) );
  OR U2831 ( .A(n2681), .B(n2680), .Z(n2682) );
  AND U2832 ( .A(n2683), .B(n2682), .Z(n2767) );
  XNOR U2833 ( .A(n2768), .B(n2767), .Z(n2769) );
  NANDN U2834 ( .A(n2685), .B(n2684), .Z(n2689) );
  NANDN U2835 ( .A(n2687), .B(n2686), .Z(n2688) );
  NAND U2836 ( .A(n2689), .B(n2688), .Z(n2770) );
  XNOR U2837 ( .A(n2769), .B(n2770), .Z(n2715) );
  XOR U2838 ( .A(n2716), .B(n2715), .Z(n2774) );
  NANDN U2839 ( .A(n2691), .B(n2690), .Z(n2695) );
  NANDN U2840 ( .A(n2693), .B(n2692), .Z(n2694) );
  AND U2841 ( .A(n2695), .B(n2694), .Z(n2773) );
  XNOR U2842 ( .A(n2774), .B(n2773), .Z(n2775) );
  XOR U2843 ( .A(n2776), .B(n2775), .Z(n2708) );
  NANDN U2844 ( .A(n2697), .B(n2696), .Z(n2701) );
  NAND U2845 ( .A(n2699), .B(n2698), .Z(n2700) );
  AND U2846 ( .A(n2701), .B(n2700), .Z(n2707) );
  XNOR U2847 ( .A(n2708), .B(n2707), .Z(n2709) );
  XNOR U2848 ( .A(n2710), .B(n2709), .Z(n2779) );
  XNOR U2849 ( .A(sreg[154]), .B(n2779), .Z(n2781) );
  NANDN U2850 ( .A(sreg[153]), .B(n2702), .Z(n2706) );
  NAND U2851 ( .A(n2704), .B(n2703), .Z(n2705) );
  NAND U2852 ( .A(n2706), .B(n2705), .Z(n2780) );
  XNOR U2853 ( .A(n2781), .B(n2780), .Z(c[154]) );
  NANDN U2854 ( .A(n2708), .B(n2707), .Z(n2712) );
  NANDN U2855 ( .A(n2710), .B(n2709), .Z(n2711) );
  AND U2856 ( .A(n2712), .B(n2711), .Z(n2787) );
  NANDN U2857 ( .A(n2714), .B(n2713), .Z(n2718) );
  NAND U2858 ( .A(n2716), .B(n2715), .Z(n2717) );
  AND U2859 ( .A(n2718), .B(n2717), .Z(n2853) );
  NANDN U2860 ( .A(n2720), .B(n2719), .Z(n2724) );
  NANDN U2861 ( .A(n2722), .B(n2721), .Z(n2723) );
  AND U2862 ( .A(n2724), .B(n2723), .Z(n2840) );
  NANDN U2863 ( .A(n9891), .B(n2725), .Z(n2727) );
  XOR U2864 ( .A(b[13]), .B(a[31]), .Z(n2826) );
  NANDN U2865 ( .A(n9935), .B(n2826), .Z(n2726) );
  AND U2866 ( .A(n2727), .B(n2726), .Z(n2818) );
  AND U2867 ( .A(b[15]), .B(a[27]), .Z(n2817) );
  XNOR U2868 ( .A(n2818), .B(n2817), .Z(n2819) );
  NAND U2869 ( .A(b[0]), .B(a[43]), .Z(n2728) );
  XNOR U2870 ( .A(b[1]), .B(n2728), .Z(n2730) );
  NANDN U2871 ( .A(b[0]), .B(a[42]), .Z(n2729) );
  NAND U2872 ( .A(n2730), .B(n2729), .Z(n2820) );
  XNOR U2873 ( .A(n2819), .B(n2820), .Z(n2838) );
  NANDN U2874 ( .A(n9437), .B(n2731), .Z(n2733) );
  XOR U2875 ( .A(b[5]), .B(a[39]), .Z(n2829) );
  NANDN U2876 ( .A(n9503), .B(n2829), .Z(n2732) );
  AND U2877 ( .A(n2733), .B(n2732), .Z(n2814) );
  NANDN U2878 ( .A(n9588), .B(n2734), .Z(n2736) );
  XOR U2879 ( .A(b[7]), .B(a[37]), .Z(n2832) );
  NANDN U2880 ( .A(n9639), .B(n2832), .Z(n2735) );
  AND U2881 ( .A(n2736), .B(n2735), .Z(n2812) );
  NANDN U2882 ( .A(n9374), .B(n2737), .Z(n2739) );
  XOR U2883 ( .A(b[3]), .B(a[41]), .Z(n2835) );
  NANDN U2884 ( .A(n9375), .B(n2835), .Z(n2738) );
  NAND U2885 ( .A(n2739), .B(n2738), .Z(n2811) );
  XNOR U2886 ( .A(n2812), .B(n2811), .Z(n2813) );
  XOR U2887 ( .A(n2814), .B(n2813), .Z(n2839) );
  XOR U2888 ( .A(n2838), .B(n2839), .Z(n2841) );
  XOR U2889 ( .A(n2840), .B(n2841), .Z(n2791) );
  NANDN U2890 ( .A(n2741), .B(n2740), .Z(n2745) );
  OR U2891 ( .A(n2743), .B(n2742), .Z(n2744) );
  AND U2892 ( .A(n2745), .B(n2744), .Z(n2790) );
  XNOR U2893 ( .A(n2791), .B(n2790), .Z(n2793) );
  NAND U2894 ( .A(n2746), .B(n9883), .Z(n2748) );
  XOR U2895 ( .A(b[11]), .B(a[33]), .Z(n2796) );
  NANDN U2896 ( .A(n9856), .B(n2796), .Z(n2747) );
  AND U2897 ( .A(n2748), .B(n2747), .Z(n2807) );
  NANDN U2898 ( .A(n10005), .B(n2749), .Z(n2751) );
  XOR U2899 ( .A(b[15]), .B(a[29]), .Z(n2799) );
  NANDN U2900 ( .A(n10006), .B(n2799), .Z(n2750) );
  AND U2901 ( .A(n2751), .B(n2750), .Z(n2806) );
  NANDN U2902 ( .A(n9685), .B(n2752), .Z(n2754) );
  XOR U2903 ( .A(b[9]), .B(a[35]), .Z(n2802) );
  NANDN U2904 ( .A(n9758), .B(n2802), .Z(n2753) );
  NAND U2905 ( .A(n2754), .B(n2753), .Z(n2805) );
  XOR U2906 ( .A(n2806), .B(n2805), .Z(n2808) );
  XOR U2907 ( .A(n2807), .B(n2808), .Z(n2845) );
  NANDN U2908 ( .A(n2756), .B(n2755), .Z(n2760) );
  OR U2909 ( .A(n2758), .B(n2757), .Z(n2759) );
  AND U2910 ( .A(n2760), .B(n2759), .Z(n2844) );
  XNOR U2911 ( .A(n2845), .B(n2844), .Z(n2846) );
  NANDN U2912 ( .A(n2762), .B(n2761), .Z(n2766) );
  NANDN U2913 ( .A(n2764), .B(n2763), .Z(n2765) );
  NAND U2914 ( .A(n2766), .B(n2765), .Z(n2847) );
  XNOR U2915 ( .A(n2846), .B(n2847), .Z(n2792) );
  XOR U2916 ( .A(n2793), .B(n2792), .Z(n2851) );
  NANDN U2917 ( .A(n2768), .B(n2767), .Z(n2772) );
  NANDN U2918 ( .A(n2770), .B(n2769), .Z(n2771) );
  AND U2919 ( .A(n2772), .B(n2771), .Z(n2850) );
  XNOR U2920 ( .A(n2851), .B(n2850), .Z(n2852) );
  XOR U2921 ( .A(n2853), .B(n2852), .Z(n2785) );
  NANDN U2922 ( .A(n2774), .B(n2773), .Z(n2778) );
  NAND U2923 ( .A(n2776), .B(n2775), .Z(n2777) );
  AND U2924 ( .A(n2778), .B(n2777), .Z(n2784) );
  XNOR U2925 ( .A(n2785), .B(n2784), .Z(n2786) );
  XNOR U2926 ( .A(n2787), .B(n2786), .Z(n2856) );
  XNOR U2927 ( .A(sreg[155]), .B(n2856), .Z(n2858) );
  NANDN U2928 ( .A(sreg[154]), .B(n2779), .Z(n2783) );
  NAND U2929 ( .A(n2781), .B(n2780), .Z(n2782) );
  NAND U2930 ( .A(n2783), .B(n2782), .Z(n2857) );
  XNOR U2931 ( .A(n2858), .B(n2857), .Z(c[155]) );
  NANDN U2932 ( .A(n2785), .B(n2784), .Z(n2789) );
  NANDN U2933 ( .A(n2787), .B(n2786), .Z(n2788) );
  AND U2934 ( .A(n2789), .B(n2788), .Z(n2864) );
  NANDN U2935 ( .A(n2791), .B(n2790), .Z(n2795) );
  NAND U2936 ( .A(n2793), .B(n2792), .Z(n2794) );
  AND U2937 ( .A(n2795), .B(n2794), .Z(n2930) );
  NAND U2938 ( .A(n2796), .B(n9883), .Z(n2798) );
  XOR U2939 ( .A(b[11]), .B(a[34]), .Z(n2900) );
  NANDN U2940 ( .A(n9856), .B(n2900), .Z(n2797) );
  AND U2941 ( .A(n2798), .B(n2797), .Z(n2911) );
  NANDN U2942 ( .A(n10005), .B(n2799), .Z(n2801) );
  XOR U2943 ( .A(b[15]), .B(a[30]), .Z(n2903) );
  NANDN U2944 ( .A(n10006), .B(n2903), .Z(n2800) );
  AND U2945 ( .A(n2801), .B(n2800), .Z(n2910) );
  NANDN U2946 ( .A(n9685), .B(n2802), .Z(n2804) );
  XOR U2947 ( .A(b[9]), .B(a[36]), .Z(n2906) );
  NANDN U2948 ( .A(n9758), .B(n2906), .Z(n2803) );
  NAND U2949 ( .A(n2804), .B(n2803), .Z(n2909) );
  XOR U2950 ( .A(n2910), .B(n2909), .Z(n2912) );
  XOR U2951 ( .A(n2911), .B(n2912), .Z(n2922) );
  NANDN U2952 ( .A(n2806), .B(n2805), .Z(n2810) );
  OR U2953 ( .A(n2808), .B(n2807), .Z(n2809) );
  AND U2954 ( .A(n2810), .B(n2809), .Z(n2921) );
  XNOR U2955 ( .A(n2922), .B(n2921), .Z(n2923) );
  NANDN U2956 ( .A(n2812), .B(n2811), .Z(n2816) );
  NANDN U2957 ( .A(n2814), .B(n2813), .Z(n2815) );
  NAND U2958 ( .A(n2816), .B(n2815), .Z(n2924) );
  XNOR U2959 ( .A(n2923), .B(n2924), .Z(n2870) );
  NANDN U2960 ( .A(n2818), .B(n2817), .Z(n2822) );
  NANDN U2961 ( .A(n2820), .B(n2819), .Z(n2821) );
  AND U2962 ( .A(n2822), .B(n2821), .Z(n2896) );
  NAND U2963 ( .A(b[0]), .B(a[44]), .Z(n2823) );
  XNOR U2964 ( .A(b[1]), .B(n2823), .Z(n2825) );
  NANDN U2965 ( .A(b[0]), .B(a[43]), .Z(n2824) );
  NAND U2966 ( .A(n2825), .B(n2824), .Z(n2876) );
  NANDN U2967 ( .A(n9891), .B(n2826), .Z(n2828) );
  XOR U2968 ( .A(b[13]), .B(a[32]), .Z(n2882) );
  NANDN U2969 ( .A(n9935), .B(n2882), .Z(n2827) );
  AND U2970 ( .A(n2828), .B(n2827), .Z(n2874) );
  AND U2971 ( .A(b[15]), .B(a[28]), .Z(n2873) );
  XNOR U2972 ( .A(n2874), .B(n2873), .Z(n2875) );
  XNOR U2973 ( .A(n2876), .B(n2875), .Z(n2894) );
  NANDN U2974 ( .A(n9437), .B(n2829), .Z(n2831) );
  XOR U2975 ( .A(b[5]), .B(a[40]), .Z(n2885) );
  NANDN U2976 ( .A(n9503), .B(n2885), .Z(n2830) );
  AND U2977 ( .A(n2831), .B(n2830), .Z(n2918) );
  NANDN U2978 ( .A(n9588), .B(n2832), .Z(n2834) );
  XOR U2979 ( .A(b[7]), .B(a[38]), .Z(n2888) );
  NANDN U2980 ( .A(n9639), .B(n2888), .Z(n2833) );
  AND U2981 ( .A(n2834), .B(n2833), .Z(n2916) );
  NANDN U2982 ( .A(n9374), .B(n2835), .Z(n2837) );
  XOR U2983 ( .A(b[3]), .B(a[42]), .Z(n2891) );
  NANDN U2984 ( .A(n9375), .B(n2891), .Z(n2836) );
  NAND U2985 ( .A(n2837), .B(n2836), .Z(n2915) );
  XNOR U2986 ( .A(n2916), .B(n2915), .Z(n2917) );
  XOR U2987 ( .A(n2918), .B(n2917), .Z(n2895) );
  XOR U2988 ( .A(n2894), .B(n2895), .Z(n2897) );
  XOR U2989 ( .A(n2896), .B(n2897), .Z(n2868) );
  NANDN U2990 ( .A(n2839), .B(n2838), .Z(n2843) );
  OR U2991 ( .A(n2841), .B(n2840), .Z(n2842) );
  AND U2992 ( .A(n2843), .B(n2842), .Z(n2867) );
  XNOR U2993 ( .A(n2868), .B(n2867), .Z(n2869) );
  XOR U2994 ( .A(n2870), .B(n2869), .Z(n2928) );
  NANDN U2995 ( .A(n2845), .B(n2844), .Z(n2849) );
  NANDN U2996 ( .A(n2847), .B(n2846), .Z(n2848) );
  AND U2997 ( .A(n2849), .B(n2848), .Z(n2927) );
  XNOR U2998 ( .A(n2928), .B(n2927), .Z(n2929) );
  XOR U2999 ( .A(n2930), .B(n2929), .Z(n2862) );
  NANDN U3000 ( .A(n2851), .B(n2850), .Z(n2855) );
  NAND U3001 ( .A(n2853), .B(n2852), .Z(n2854) );
  AND U3002 ( .A(n2855), .B(n2854), .Z(n2861) );
  XNOR U3003 ( .A(n2862), .B(n2861), .Z(n2863) );
  XNOR U3004 ( .A(n2864), .B(n2863), .Z(n2933) );
  XNOR U3005 ( .A(sreg[156]), .B(n2933), .Z(n2935) );
  NANDN U3006 ( .A(sreg[155]), .B(n2856), .Z(n2860) );
  NAND U3007 ( .A(n2858), .B(n2857), .Z(n2859) );
  NAND U3008 ( .A(n2860), .B(n2859), .Z(n2934) );
  XNOR U3009 ( .A(n2935), .B(n2934), .Z(c[156]) );
  NANDN U3010 ( .A(n2862), .B(n2861), .Z(n2866) );
  NANDN U3011 ( .A(n2864), .B(n2863), .Z(n2865) );
  AND U3012 ( .A(n2866), .B(n2865), .Z(n2941) );
  NANDN U3013 ( .A(n2868), .B(n2867), .Z(n2872) );
  NAND U3014 ( .A(n2870), .B(n2869), .Z(n2871) );
  AND U3015 ( .A(n2872), .B(n2871), .Z(n3007) );
  NANDN U3016 ( .A(n2874), .B(n2873), .Z(n2878) );
  NANDN U3017 ( .A(n2876), .B(n2875), .Z(n2877) );
  AND U3018 ( .A(n2878), .B(n2877), .Z(n2973) );
  NAND U3019 ( .A(b[0]), .B(a[45]), .Z(n2879) );
  XNOR U3020 ( .A(b[1]), .B(n2879), .Z(n2881) );
  NANDN U3021 ( .A(b[0]), .B(a[44]), .Z(n2880) );
  NAND U3022 ( .A(n2881), .B(n2880), .Z(n2953) );
  NANDN U3023 ( .A(n9891), .B(n2882), .Z(n2884) );
  XOR U3024 ( .A(b[13]), .B(a[33]), .Z(n2959) );
  NANDN U3025 ( .A(n9935), .B(n2959), .Z(n2883) );
  AND U3026 ( .A(n2884), .B(n2883), .Z(n2951) );
  AND U3027 ( .A(b[15]), .B(a[29]), .Z(n2950) );
  XNOR U3028 ( .A(n2951), .B(n2950), .Z(n2952) );
  XNOR U3029 ( .A(n2953), .B(n2952), .Z(n2971) );
  NANDN U3030 ( .A(n9437), .B(n2885), .Z(n2887) );
  XOR U3031 ( .A(b[5]), .B(a[41]), .Z(n2962) );
  NANDN U3032 ( .A(n9503), .B(n2962), .Z(n2886) );
  AND U3033 ( .A(n2887), .B(n2886), .Z(n2995) );
  NANDN U3034 ( .A(n9588), .B(n2888), .Z(n2890) );
  XOR U3035 ( .A(b[7]), .B(a[39]), .Z(n2965) );
  NANDN U3036 ( .A(n9639), .B(n2965), .Z(n2889) );
  AND U3037 ( .A(n2890), .B(n2889), .Z(n2993) );
  NANDN U3038 ( .A(n9374), .B(n2891), .Z(n2893) );
  XOR U3039 ( .A(b[3]), .B(a[43]), .Z(n2968) );
  NANDN U3040 ( .A(n9375), .B(n2968), .Z(n2892) );
  NAND U3041 ( .A(n2893), .B(n2892), .Z(n2992) );
  XNOR U3042 ( .A(n2993), .B(n2992), .Z(n2994) );
  XOR U3043 ( .A(n2995), .B(n2994), .Z(n2972) );
  XOR U3044 ( .A(n2971), .B(n2972), .Z(n2974) );
  XOR U3045 ( .A(n2973), .B(n2974), .Z(n2945) );
  NANDN U3046 ( .A(n2895), .B(n2894), .Z(n2899) );
  OR U3047 ( .A(n2897), .B(n2896), .Z(n2898) );
  AND U3048 ( .A(n2899), .B(n2898), .Z(n2944) );
  XNOR U3049 ( .A(n2945), .B(n2944), .Z(n2947) );
  NAND U3050 ( .A(n2900), .B(n9883), .Z(n2902) );
  XOR U3051 ( .A(b[11]), .B(a[35]), .Z(n2977) );
  NANDN U3052 ( .A(n9856), .B(n2977), .Z(n2901) );
  AND U3053 ( .A(n2902), .B(n2901), .Z(n2988) );
  NANDN U3054 ( .A(n10005), .B(n2903), .Z(n2905) );
  XOR U3055 ( .A(b[15]), .B(a[31]), .Z(n2980) );
  NANDN U3056 ( .A(n10006), .B(n2980), .Z(n2904) );
  AND U3057 ( .A(n2905), .B(n2904), .Z(n2987) );
  NANDN U3058 ( .A(n9685), .B(n2906), .Z(n2908) );
  XOR U3059 ( .A(b[9]), .B(a[37]), .Z(n2983) );
  NANDN U3060 ( .A(n9758), .B(n2983), .Z(n2907) );
  NAND U3061 ( .A(n2908), .B(n2907), .Z(n2986) );
  XOR U3062 ( .A(n2987), .B(n2986), .Z(n2989) );
  XOR U3063 ( .A(n2988), .B(n2989), .Z(n2999) );
  NANDN U3064 ( .A(n2910), .B(n2909), .Z(n2914) );
  OR U3065 ( .A(n2912), .B(n2911), .Z(n2913) );
  AND U3066 ( .A(n2914), .B(n2913), .Z(n2998) );
  XNOR U3067 ( .A(n2999), .B(n2998), .Z(n3000) );
  NANDN U3068 ( .A(n2916), .B(n2915), .Z(n2920) );
  NANDN U3069 ( .A(n2918), .B(n2917), .Z(n2919) );
  NAND U3070 ( .A(n2920), .B(n2919), .Z(n3001) );
  XNOR U3071 ( .A(n3000), .B(n3001), .Z(n2946) );
  XOR U3072 ( .A(n2947), .B(n2946), .Z(n3005) );
  NANDN U3073 ( .A(n2922), .B(n2921), .Z(n2926) );
  NANDN U3074 ( .A(n2924), .B(n2923), .Z(n2925) );
  AND U3075 ( .A(n2926), .B(n2925), .Z(n3004) );
  XNOR U3076 ( .A(n3005), .B(n3004), .Z(n3006) );
  XOR U3077 ( .A(n3007), .B(n3006), .Z(n2939) );
  NANDN U3078 ( .A(n2928), .B(n2927), .Z(n2932) );
  NAND U3079 ( .A(n2930), .B(n2929), .Z(n2931) );
  AND U3080 ( .A(n2932), .B(n2931), .Z(n2938) );
  XNOR U3081 ( .A(n2939), .B(n2938), .Z(n2940) );
  XNOR U3082 ( .A(n2941), .B(n2940), .Z(n3010) );
  XNOR U3083 ( .A(sreg[157]), .B(n3010), .Z(n3012) );
  NANDN U3084 ( .A(sreg[156]), .B(n2933), .Z(n2937) );
  NAND U3085 ( .A(n2935), .B(n2934), .Z(n2936) );
  NAND U3086 ( .A(n2937), .B(n2936), .Z(n3011) );
  XNOR U3087 ( .A(n3012), .B(n3011), .Z(c[157]) );
  NANDN U3088 ( .A(n2939), .B(n2938), .Z(n2943) );
  NANDN U3089 ( .A(n2941), .B(n2940), .Z(n2942) );
  AND U3090 ( .A(n2943), .B(n2942), .Z(n3018) );
  NANDN U3091 ( .A(n2945), .B(n2944), .Z(n2949) );
  NAND U3092 ( .A(n2947), .B(n2946), .Z(n2948) );
  AND U3093 ( .A(n2949), .B(n2948), .Z(n3084) );
  NANDN U3094 ( .A(n2951), .B(n2950), .Z(n2955) );
  NANDN U3095 ( .A(n2953), .B(n2952), .Z(n2954) );
  AND U3096 ( .A(n2955), .B(n2954), .Z(n3050) );
  NAND U3097 ( .A(b[0]), .B(a[46]), .Z(n2956) );
  XNOR U3098 ( .A(b[1]), .B(n2956), .Z(n2958) );
  NANDN U3099 ( .A(b[0]), .B(a[45]), .Z(n2957) );
  NAND U3100 ( .A(n2958), .B(n2957), .Z(n3030) );
  NANDN U3101 ( .A(n9891), .B(n2959), .Z(n2961) );
  XOR U3102 ( .A(b[13]), .B(a[34]), .Z(n3036) );
  NANDN U3103 ( .A(n9935), .B(n3036), .Z(n2960) );
  AND U3104 ( .A(n2961), .B(n2960), .Z(n3028) );
  AND U3105 ( .A(b[15]), .B(a[30]), .Z(n3027) );
  XNOR U3106 ( .A(n3028), .B(n3027), .Z(n3029) );
  XNOR U3107 ( .A(n3030), .B(n3029), .Z(n3048) );
  NANDN U3108 ( .A(n9437), .B(n2962), .Z(n2964) );
  XOR U3109 ( .A(b[5]), .B(a[42]), .Z(n3039) );
  NANDN U3110 ( .A(n9503), .B(n3039), .Z(n2963) );
  AND U3111 ( .A(n2964), .B(n2963), .Z(n3072) );
  NANDN U3112 ( .A(n9588), .B(n2965), .Z(n2967) );
  XOR U3113 ( .A(b[7]), .B(a[40]), .Z(n3042) );
  NANDN U3114 ( .A(n9639), .B(n3042), .Z(n2966) );
  AND U3115 ( .A(n2967), .B(n2966), .Z(n3070) );
  NANDN U3116 ( .A(n9374), .B(n2968), .Z(n2970) );
  XOR U3117 ( .A(b[3]), .B(a[44]), .Z(n3045) );
  NANDN U3118 ( .A(n9375), .B(n3045), .Z(n2969) );
  NAND U3119 ( .A(n2970), .B(n2969), .Z(n3069) );
  XNOR U3120 ( .A(n3070), .B(n3069), .Z(n3071) );
  XOR U3121 ( .A(n3072), .B(n3071), .Z(n3049) );
  XOR U3122 ( .A(n3048), .B(n3049), .Z(n3051) );
  XOR U3123 ( .A(n3050), .B(n3051), .Z(n3022) );
  NANDN U3124 ( .A(n2972), .B(n2971), .Z(n2976) );
  OR U3125 ( .A(n2974), .B(n2973), .Z(n2975) );
  AND U3126 ( .A(n2976), .B(n2975), .Z(n3021) );
  XNOR U3127 ( .A(n3022), .B(n3021), .Z(n3024) );
  NAND U3128 ( .A(n2977), .B(n9883), .Z(n2979) );
  XOR U3129 ( .A(b[11]), .B(a[36]), .Z(n3054) );
  NANDN U3130 ( .A(n9856), .B(n3054), .Z(n2978) );
  AND U3131 ( .A(n2979), .B(n2978), .Z(n3065) );
  NANDN U3132 ( .A(n10005), .B(n2980), .Z(n2982) );
  XOR U3133 ( .A(b[15]), .B(a[32]), .Z(n3057) );
  NANDN U3134 ( .A(n10006), .B(n3057), .Z(n2981) );
  AND U3135 ( .A(n2982), .B(n2981), .Z(n3064) );
  NANDN U3136 ( .A(n9685), .B(n2983), .Z(n2985) );
  XOR U3137 ( .A(b[9]), .B(a[38]), .Z(n3060) );
  NANDN U3138 ( .A(n9758), .B(n3060), .Z(n2984) );
  NAND U3139 ( .A(n2985), .B(n2984), .Z(n3063) );
  XOR U3140 ( .A(n3064), .B(n3063), .Z(n3066) );
  XOR U3141 ( .A(n3065), .B(n3066), .Z(n3076) );
  NANDN U3142 ( .A(n2987), .B(n2986), .Z(n2991) );
  OR U3143 ( .A(n2989), .B(n2988), .Z(n2990) );
  AND U3144 ( .A(n2991), .B(n2990), .Z(n3075) );
  XNOR U3145 ( .A(n3076), .B(n3075), .Z(n3077) );
  NANDN U3146 ( .A(n2993), .B(n2992), .Z(n2997) );
  NANDN U3147 ( .A(n2995), .B(n2994), .Z(n2996) );
  NAND U3148 ( .A(n2997), .B(n2996), .Z(n3078) );
  XNOR U3149 ( .A(n3077), .B(n3078), .Z(n3023) );
  XOR U3150 ( .A(n3024), .B(n3023), .Z(n3082) );
  NANDN U3151 ( .A(n2999), .B(n2998), .Z(n3003) );
  NANDN U3152 ( .A(n3001), .B(n3000), .Z(n3002) );
  AND U3153 ( .A(n3003), .B(n3002), .Z(n3081) );
  XNOR U3154 ( .A(n3082), .B(n3081), .Z(n3083) );
  XOR U3155 ( .A(n3084), .B(n3083), .Z(n3016) );
  NANDN U3156 ( .A(n3005), .B(n3004), .Z(n3009) );
  NAND U3157 ( .A(n3007), .B(n3006), .Z(n3008) );
  AND U3158 ( .A(n3009), .B(n3008), .Z(n3015) );
  XNOR U3159 ( .A(n3016), .B(n3015), .Z(n3017) );
  XNOR U3160 ( .A(n3018), .B(n3017), .Z(n3087) );
  XNOR U3161 ( .A(sreg[158]), .B(n3087), .Z(n3089) );
  NANDN U3162 ( .A(sreg[157]), .B(n3010), .Z(n3014) );
  NAND U3163 ( .A(n3012), .B(n3011), .Z(n3013) );
  NAND U3164 ( .A(n3014), .B(n3013), .Z(n3088) );
  XNOR U3165 ( .A(n3089), .B(n3088), .Z(c[158]) );
  NANDN U3166 ( .A(n3016), .B(n3015), .Z(n3020) );
  NANDN U3167 ( .A(n3018), .B(n3017), .Z(n3019) );
  AND U3168 ( .A(n3020), .B(n3019), .Z(n3095) );
  NANDN U3169 ( .A(n3022), .B(n3021), .Z(n3026) );
  NAND U3170 ( .A(n3024), .B(n3023), .Z(n3025) );
  AND U3171 ( .A(n3026), .B(n3025), .Z(n3161) );
  NANDN U3172 ( .A(n3028), .B(n3027), .Z(n3032) );
  NANDN U3173 ( .A(n3030), .B(n3029), .Z(n3031) );
  AND U3174 ( .A(n3032), .B(n3031), .Z(n3127) );
  NAND U3175 ( .A(b[0]), .B(a[47]), .Z(n3033) );
  XNOR U3176 ( .A(b[1]), .B(n3033), .Z(n3035) );
  NANDN U3177 ( .A(b[0]), .B(a[46]), .Z(n3034) );
  NAND U3178 ( .A(n3035), .B(n3034), .Z(n3107) );
  NANDN U3179 ( .A(n9891), .B(n3036), .Z(n3038) );
  XOR U3180 ( .A(b[13]), .B(a[35]), .Z(n3110) );
  NANDN U3181 ( .A(n9935), .B(n3110), .Z(n3037) );
  AND U3182 ( .A(n3038), .B(n3037), .Z(n3105) );
  AND U3183 ( .A(b[15]), .B(a[31]), .Z(n3104) );
  XNOR U3184 ( .A(n3105), .B(n3104), .Z(n3106) );
  XNOR U3185 ( .A(n3107), .B(n3106), .Z(n3125) );
  NANDN U3186 ( .A(n9437), .B(n3039), .Z(n3041) );
  XOR U3187 ( .A(b[5]), .B(a[43]), .Z(n3116) );
  NANDN U3188 ( .A(n9503), .B(n3116), .Z(n3040) );
  AND U3189 ( .A(n3041), .B(n3040), .Z(n3149) );
  NANDN U3190 ( .A(n9588), .B(n3042), .Z(n3044) );
  XOR U3191 ( .A(b[7]), .B(a[41]), .Z(n3119) );
  NANDN U3192 ( .A(n9639), .B(n3119), .Z(n3043) );
  AND U3193 ( .A(n3044), .B(n3043), .Z(n3147) );
  NANDN U3194 ( .A(n9374), .B(n3045), .Z(n3047) );
  XOR U3195 ( .A(b[3]), .B(a[45]), .Z(n3122) );
  NANDN U3196 ( .A(n9375), .B(n3122), .Z(n3046) );
  NAND U3197 ( .A(n3047), .B(n3046), .Z(n3146) );
  XNOR U3198 ( .A(n3147), .B(n3146), .Z(n3148) );
  XOR U3199 ( .A(n3149), .B(n3148), .Z(n3126) );
  XOR U3200 ( .A(n3125), .B(n3126), .Z(n3128) );
  XOR U3201 ( .A(n3127), .B(n3128), .Z(n3099) );
  NANDN U3202 ( .A(n3049), .B(n3048), .Z(n3053) );
  OR U3203 ( .A(n3051), .B(n3050), .Z(n3052) );
  AND U3204 ( .A(n3053), .B(n3052), .Z(n3098) );
  XNOR U3205 ( .A(n3099), .B(n3098), .Z(n3101) );
  NAND U3206 ( .A(n3054), .B(n9883), .Z(n3056) );
  XOR U3207 ( .A(b[11]), .B(a[37]), .Z(n3131) );
  NANDN U3208 ( .A(n9856), .B(n3131), .Z(n3055) );
  AND U3209 ( .A(n3056), .B(n3055), .Z(n3142) );
  NANDN U3210 ( .A(n10005), .B(n3057), .Z(n3059) );
  XOR U3211 ( .A(b[15]), .B(a[33]), .Z(n3134) );
  NANDN U3212 ( .A(n10006), .B(n3134), .Z(n3058) );
  AND U3213 ( .A(n3059), .B(n3058), .Z(n3141) );
  NANDN U3214 ( .A(n9685), .B(n3060), .Z(n3062) );
  XOR U3215 ( .A(b[9]), .B(a[39]), .Z(n3137) );
  NANDN U3216 ( .A(n9758), .B(n3137), .Z(n3061) );
  NAND U3217 ( .A(n3062), .B(n3061), .Z(n3140) );
  XOR U3218 ( .A(n3141), .B(n3140), .Z(n3143) );
  XOR U3219 ( .A(n3142), .B(n3143), .Z(n3153) );
  NANDN U3220 ( .A(n3064), .B(n3063), .Z(n3068) );
  OR U3221 ( .A(n3066), .B(n3065), .Z(n3067) );
  AND U3222 ( .A(n3068), .B(n3067), .Z(n3152) );
  XNOR U3223 ( .A(n3153), .B(n3152), .Z(n3154) );
  NANDN U3224 ( .A(n3070), .B(n3069), .Z(n3074) );
  NANDN U3225 ( .A(n3072), .B(n3071), .Z(n3073) );
  NAND U3226 ( .A(n3074), .B(n3073), .Z(n3155) );
  XNOR U3227 ( .A(n3154), .B(n3155), .Z(n3100) );
  XOR U3228 ( .A(n3101), .B(n3100), .Z(n3159) );
  NANDN U3229 ( .A(n3076), .B(n3075), .Z(n3080) );
  NANDN U3230 ( .A(n3078), .B(n3077), .Z(n3079) );
  AND U3231 ( .A(n3080), .B(n3079), .Z(n3158) );
  XNOR U3232 ( .A(n3159), .B(n3158), .Z(n3160) );
  XOR U3233 ( .A(n3161), .B(n3160), .Z(n3093) );
  NANDN U3234 ( .A(n3082), .B(n3081), .Z(n3086) );
  NAND U3235 ( .A(n3084), .B(n3083), .Z(n3085) );
  AND U3236 ( .A(n3086), .B(n3085), .Z(n3092) );
  XNOR U3237 ( .A(n3093), .B(n3092), .Z(n3094) );
  XNOR U3238 ( .A(n3095), .B(n3094), .Z(n3164) );
  XNOR U3239 ( .A(sreg[159]), .B(n3164), .Z(n3166) );
  NANDN U3240 ( .A(sreg[158]), .B(n3087), .Z(n3091) );
  NAND U3241 ( .A(n3089), .B(n3088), .Z(n3090) );
  NAND U3242 ( .A(n3091), .B(n3090), .Z(n3165) );
  XNOR U3243 ( .A(n3166), .B(n3165), .Z(c[159]) );
  NANDN U3244 ( .A(n3093), .B(n3092), .Z(n3097) );
  NANDN U3245 ( .A(n3095), .B(n3094), .Z(n3096) );
  AND U3246 ( .A(n3097), .B(n3096), .Z(n3172) );
  NANDN U3247 ( .A(n3099), .B(n3098), .Z(n3103) );
  NAND U3248 ( .A(n3101), .B(n3100), .Z(n3102) );
  AND U3249 ( .A(n3103), .B(n3102), .Z(n3238) );
  NANDN U3250 ( .A(n3105), .B(n3104), .Z(n3109) );
  NANDN U3251 ( .A(n3107), .B(n3106), .Z(n3108) );
  AND U3252 ( .A(n3109), .B(n3108), .Z(n3204) );
  NANDN U3253 ( .A(n9891), .B(n3110), .Z(n3112) );
  XOR U3254 ( .A(b[13]), .B(a[36]), .Z(n3190) );
  NANDN U3255 ( .A(n9935), .B(n3190), .Z(n3111) );
  AND U3256 ( .A(n3112), .B(n3111), .Z(n3182) );
  AND U3257 ( .A(b[15]), .B(a[32]), .Z(n3181) );
  XNOR U3258 ( .A(n3182), .B(n3181), .Z(n3183) );
  NAND U3259 ( .A(b[0]), .B(a[48]), .Z(n3113) );
  XNOR U3260 ( .A(b[1]), .B(n3113), .Z(n3115) );
  NANDN U3261 ( .A(b[0]), .B(a[47]), .Z(n3114) );
  NAND U3262 ( .A(n3115), .B(n3114), .Z(n3184) );
  XNOR U3263 ( .A(n3183), .B(n3184), .Z(n3202) );
  NANDN U3264 ( .A(n9437), .B(n3116), .Z(n3118) );
  XOR U3265 ( .A(b[5]), .B(a[44]), .Z(n3193) );
  NANDN U3266 ( .A(n9503), .B(n3193), .Z(n3117) );
  AND U3267 ( .A(n3118), .B(n3117), .Z(n3226) );
  NANDN U3268 ( .A(n9588), .B(n3119), .Z(n3121) );
  XOR U3269 ( .A(b[7]), .B(a[42]), .Z(n3196) );
  NANDN U3270 ( .A(n9639), .B(n3196), .Z(n3120) );
  AND U3271 ( .A(n3121), .B(n3120), .Z(n3224) );
  NANDN U3272 ( .A(n9374), .B(n3122), .Z(n3124) );
  XOR U3273 ( .A(b[3]), .B(a[46]), .Z(n3199) );
  NANDN U3274 ( .A(n9375), .B(n3199), .Z(n3123) );
  NAND U3275 ( .A(n3124), .B(n3123), .Z(n3223) );
  XNOR U3276 ( .A(n3224), .B(n3223), .Z(n3225) );
  XOR U3277 ( .A(n3226), .B(n3225), .Z(n3203) );
  XOR U3278 ( .A(n3202), .B(n3203), .Z(n3205) );
  XOR U3279 ( .A(n3204), .B(n3205), .Z(n3176) );
  NANDN U3280 ( .A(n3126), .B(n3125), .Z(n3130) );
  OR U3281 ( .A(n3128), .B(n3127), .Z(n3129) );
  AND U3282 ( .A(n3130), .B(n3129), .Z(n3175) );
  XNOR U3283 ( .A(n3176), .B(n3175), .Z(n3178) );
  NAND U3284 ( .A(n3131), .B(n9883), .Z(n3133) );
  XOR U3285 ( .A(b[11]), .B(a[38]), .Z(n3208) );
  NANDN U3286 ( .A(n9856), .B(n3208), .Z(n3132) );
  AND U3287 ( .A(n3133), .B(n3132), .Z(n3219) );
  NANDN U3288 ( .A(n10005), .B(n3134), .Z(n3136) );
  XOR U3289 ( .A(b[15]), .B(a[34]), .Z(n3211) );
  NANDN U3290 ( .A(n10006), .B(n3211), .Z(n3135) );
  AND U3291 ( .A(n3136), .B(n3135), .Z(n3218) );
  NANDN U3292 ( .A(n9685), .B(n3137), .Z(n3139) );
  XOR U3293 ( .A(b[9]), .B(a[40]), .Z(n3214) );
  NANDN U3294 ( .A(n9758), .B(n3214), .Z(n3138) );
  NAND U3295 ( .A(n3139), .B(n3138), .Z(n3217) );
  XOR U3296 ( .A(n3218), .B(n3217), .Z(n3220) );
  XOR U3297 ( .A(n3219), .B(n3220), .Z(n3230) );
  NANDN U3298 ( .A(n3141), .B(n3140), .Z(n3145) );
  OR U3299 ( .A(n3143), .B(n3142), .Z(n3144) );
  AND U3300 ( .A(n3145), .B(n3144), .Z(n3229) );
  XNOR U3301 ( .A(n3230), .B(n3229), .Z(n3231) );
  NANDN U3302 ( .A(n3147), .B(n3146), .Z(n3151) );
  NANDN U3303 ( .A(n3149), .B(n3148), .Z(n3150) );
  NAND U3304 ( .A(n3151), .B(n3150), .Z(n3232) );
  XNOR U3305 ( .A(n3231), .B(n3232), .Z(n3177) );
  XOR U3306 ( .A(n3178), .B(n3177), .Z(n3236) );
  NANDN U3307 ( .A(n3153), .B(n3152), .Z(n3157) );
  NANDN U3308 ( .A(n3155), .B(n3154), .Z(n3156) );
  AND U3309 ( .A(n3157), .B(n3156), .Z(n3235) );
  XNOR U3310 ( .A(n3236), .B(n3235), .Z(n3237) );
  XOR U3311 ( .A(n3238), .B(n3237), .Z(n3170) );
  NANDN U3312 ( .A(n3159), .B(n3158), .Z(n3163) );
  NAND U3313 ( .A(n3161), .B(n3160), .Z(n3162) );
  AND U3314 ( .A(n3163), .B(n3162), .Z(n3169) );
  XNOR U3315 ( .A(n3170), .B(n3169), .Z(n3171) );
  XNOR U3316 ( .A(n3172), .B(n3171), .Z(n3241) );
  XNOR U3317 ( .A(sreg[160]), .B(n3241), .Z(n3243) );
  NANDN U3318 ( .A(sreg[159]), .B(n3164), .Z(n3168) );
  NAND U3319 ( .A(n3166), .B(n3165), .Z(n3167) );
  NAND U3320 ( .A(n3168), .B(n3167), .Z(n3242) );
  XNOR U3321 ( .A(n3243), .B(n3242), .Z(c[160]) );
  NANDN U3322 ( .A(n3170), .B(n3169), .Z(n3174) );
  NANDN U3323 ( .A(n3172), .B(n3171), .Z(n3173) );
  AND U3324 ( .A(n3174), .B(n3173), .Z(n3249) );
  NANDN U3325 ( .A(n3176), .B(n3175), .Z(n3180) );
  NAND U3326 ( .A(n3178), .B(n3177), .Z(n3179) );
  AND U3327 ( .A(n3180), .B(n3179), .Z(n3315) );
  NANDN U3328 ( .A(n3182), .B(n3181), .Z(n3186) );
  NANDN U3329 ( .A(n3184), .B(n3183), .Z(n3185) );
  AND U3330 ( .A(n3186), .B(n3185), .Z(n3281) );
  NAND U3331 ( .A(b[0]), .B(a[49]), .Z(n3187) );
  XNOR U3332 ( .A(b[1]), .B(n3187), .Z(n3189) );
  NANDN U3333 ( .A(b[0]), .B(a[48]), .Z(n3188) );
  NAND U3334 ( .A(n3189), .B(n3188), .Z(n3261) );
  NANDN U3335 ( .A(n9891), .B(n3190), .Z(n3192) );
  XOR U3336 ( .A(b[13]), .B(a[37]), .Z(n3267) );
  NANDN U3337 ( .A(n9935), .B(n3267), .Z(n3191) );
  AND U3338 ( .A(n3192), .B(n3191), .Z(n3259) );
  AND U3339 ( .A(b[15]), .B(a[33]), .Z(n3258) );
  XNOR U3340 ( .A(n3259), .B(n3258), .Z(n3260) );
  XNOR U3341 ( .A(n3261), .B(n3260), .Z(n3279) );
  NANDN U3342 ( .A(n9437), .B(n3193), .Z(n3195) );
  XOR U3343 ( .A(b[5]), .B(a[45]), .Z(n3270) );
  NANDN U3344 ( .A(n9503), .B(n3270), .Z(n3194) );
  AND U3345 ( .A(n3195), .B(n3194), .Z(n3303) );
  NANDN U3346 ( .A(n9588), .B(n3196), .Z(n3198) );
  XOR U3347 ( .A(b[7]), .B(a[43]), .Z(n3273) );
  NANDN U3348 ( .A(n9639), .B(n3273), .Z(n3197) );
  AND U3349 ( .A(n3198), .B(n3197), .Z(n3301) );
  NANDN U3350 ( .A(n9374), .B(n3199), .Z(n3201) );
  XOR U3351 ( .A(b[3]), .B(a[47]), .Z(n3276) );
  NANDN U3352 ( .A(n9375), .B(n3276), .Z(n3200) );
  NAND U3353 ( .A(n3201), .B(n3200), .Z(n3300) );
  XNOR U3354 ( .A(n3301), .B(n3300), .Z(n3302) );
  XOR U3355 ( .A(n3303), .B(n3302), .Z(n3280) );
  XOR U3356 ( .A(n3279), .B(n3280), .Z(n3282) );
  XOR U3357 ( .A(n3281), .B(n3282), .Z(n3253) );
  NANDN U3358 ( .A(n3203), .B(n3202), .Z(n3207) );
  OR U3359 ( .A(n3205), .B(n3204), .Z(n3206) );
  AND U3360 ( .A(n3207), .B(n3206), .Z(n3252) );
  XNOR U3361 ( .A(n3253), .B(n3252), .Z(n3255) );
  NAND U3362 ( .A(n3208), .B(n9883), .Z(n3210) );
  XOR U3363 ( .A(b[11]), .B(a[39]), .Z(n3285) );
  NANDN U3364 ( .A(n9856), .B(n3285), .Z(n3209) );
  AND U3365 ( .A(n3210), .B(n3209), .Z(n3296) );
  NANDN U3366 ( .A(n10005), .B(n3211), .Z(n3213) );
  XOR U3367 ( .A(b[15]), .B(a[35]), .Z(n3288) );
  NANDN U3368 ( .A(n10006), .B(n3288), .Z(n3212) );
  AND U3369 ( .A(n3213), .B(n3212), .Z(n3295) );
  NANDN U3370 ( .A(n9685), .B(n3214), .Z(n3216) );
  XOR U3371 ( .A(b[9]), .B(a[41]), .Z(n3291) );
  NANDN U3372 ( .A(n9758), .B(n3291), .Z(n3215) );
  NAND U3373 ( .A(n3216), .B(n3215), .Z(n3294) );
  XOR U3374 ( .A(n3295), .B(n3294), .Z(n3297) );
  XOR U3375 ( .A(n3296), .B(n3297), .Z(n3307) );
  NANDN U3376 ( .A(n3218), .B(n3217), .Z(n3222) );
  OR U3377 ( .A(n3220), .B(n3219), .Z(n3221) );
  AND U3378 ( .A(n3222), .B(n3221), .Z(n3306) );
  XNOR U3379 ( .A(n3307), .B(n3306), .Z(n3308) );
  NANDN U3380 ( .A(n3224), .B(n3223), .Z(n3228) );
  NANDN U3381 ( .A(n3226), .B(n3225), .Z(n3227) );
  NAND U3382 ( .A(n3228), .B(n3227), .Z(n3309) );
  XNOR U3383 ( .A(n3308), .B(n3309), .Z(n3254) );
  XOR U3384 ( .A(n3255), .B(n3254), .Z(n3313) );
  NANDN U3385 ( .A(n3230), .B(n3229), .Z(n3234) );
  NANDN U3386 ( .A(n3232), .B(n3231), .Z(n3233) );
  AND U3387 ( .A(n3234), .B(n3233), .Z(n3312) );
  XNOR U3388 ( .A(n3313), .B(n3312), .Z(n3314) );
  XOR U3389 ( .A(n3315), .B(n3314), .Z(n3247) );
  NANDN U3390 ( .A(n3236), .B(n3235), .Z(n3240) );
  NAND U3391 ( .A(n3238), .B(n3237), .Z(n3239) );
  AND U3392 ( .A(n3240), .B(n3239), .Z(n3246) );
  XNOR U3393 ( .A(n3247), .B(n3246), .Z(n3248) );
  XNOR U3394 ( .A(n3249), .B(n3248), .Z(n3318) );
  XNOR U3395 ( .A(sreg[161]), .B(n3318), .Z(n3320) );
  NANDN U3396 ( .A(sreg[160]), .B(n3241), .Z(n3245) );
  NAND U3397 ( .A(n3243), .B(n3242), .Z(n3244) );
  NAND U3398 ( .A(n3245), .B(n3244), .Z(n3319) );
  XNOR U3399 ( .A(n3320), .B(n3319), .Z(c[161]) );
  NANDN U3400 ( .A(n3247), .B(n3246), .Z(n3251) );
  NANDN U3401 ( .A(n3249), .B(n3248), .Z(n3250) );
  AND U3402 ( .A(n3251), .B(n3250), .Z(n3326) );
  NANDN U3403 ( .A(n3253), .B(n3252), .Z(n3257) );
  NAND U3404 ( .A(n3255), .B(n3254), .Z(n3256) );
  AND U3405 ( .A(n3257), .B(n3256), .Z(n3392) );
  NANDN U3406 ( .A(n3259), .B(n3258), .Z(n3263) );
  NANDN U3407 ( .A(n3261), .B(n3260), .Z(n3262) );
  AND U3408 ( .A(n3263), .B(n3262), .Z(n3358) );
  NAND U3409 ( .A(b[0]), .B(a[50]), .Z(n3264) );
  XNOR U3410 ( .A(b[1]), .B(n3264), .Z(n3266) );
  NANDN U3411 ( .A(b[0]), .B(a[49]), .Z(n3265) );
  NAND U3412 ( .A(n3266), .B(n3265), .Z(n3338) );
  NANDN U3413 ( .A(n9891), .B(n3267), .Z(n3269) );
  XOR U3414 ( .A(b[13]), .B(a[38]), .Z(n3344) );
  NANDN U3415 ( .A(n9935), .B(n3344), .Z(n3268) );
  AND U3416 ( .A(n3269), .B(n3268), .Z(n3336) );
  AND U3417 ( .A(b[15]), .B(a[34]), .Z(n3335) );
  XNOR U3418 ( .A(n3336), .B(n3335), .Z(n3337) );
  XNOR U3419 ( .A(n3338), .B(n3337), .Z(n3356) );
  NANDN U3420 ( .A(n9437), .B(n3270), .Z(n3272) );
  XOR U3421 ( .A(b[5]), .B(a[46]), .Z(n3347) );
  NANDN U3422 ( .A(n9503), .B(n3347), .Z(n3271) );
  AND U3423 ( .A(n3272), .B(n3271), .Z(n3380) );
  NANDN U3424 ( .A(n9588), .B(n3273), .Z(n3275) );
  XOR U3425 ( .A(b[7]), .B(a[44]), .Z(n3350) );
  NANDN U3426 ( .A(n9639), .B(n3350), .Z(n3274) );
  AND U3427 ( .A(n3275), .B(n3274), .Z(n3378) );
  NANDN U3428 ( .A(n9374), .B(n3276), .Z(n3278) );
  XOR U3429 ( .A(b[3]), .B(a[48]), .Z(n3353) );
  NANDN U3430 ( .A(n9375), .B(n3353), .Z(n3277) );
  NAND U3431 ( .A(n3278), .B(n3277), .Z(n3377) );
  XNOR U3432 ( .A(n3378), .B(n3377), .Z(n3379) );
  XOR U3433 ( .A(n3380), .B(n3379), .Z(n3357) );
  XOR U3434 ( .A(n3356), .B(n3357), .Z(n3359) );
  XOR U3435 ( .A(n3358), .B(n3359), .Z(n3330) );
  NANDN U3436 ( .A(n3280), .B(n3279), .Z(n3284) );
  OR U3437 ( .A(n3282), .B(n3281), .Z(n3283) );
  AND U3438 ( .A(n3284), .B(n3283), .Z(n3329) );
  XNOR U3439 ( .A(n3330), .B(n3329), .Z(n3332) );
  NAND U3440 ( .A(n3285), .B(n9883), .Z(n3287) );
  XOR U3441 ( .A(b[11]), .B(a[40]), .Z(n3362) );
  NANDN U3442 ( .A(n9856), .B(n3362), .Z(n3286) );
  AND U3443 ( .A(n3287), .B(n3286), .Z(n3373) );
  NANDN U3444 ( .A(n10005), .B(n3288), .Z(n3290) );
  XOR U3445 ( .A(b[15]), .B(a[36]), .Z(n3365) );
  NANDN U3446 ( .A(n10006), .B(n3365), .Z(n3289) );
  AND U3447 ( .A(n3290), .B(n3289), .Z(n3372) );
  NANDN U3448 ( .A(n9685), .B(n3291), .Z(n3293) );
  XOR U3449 ( .A(b[9]), .B(a[42]), .Z(n3368) );
  NANDN U3450 ( .A(n9758), .B(n3368), .Z(n3292) );
  NAND U3451 ( .A(n3293), .B(n3292), .Z(n3371) );
  XOR U3452 ( .A(n3372), .B(n3371), .Z(n3374) );
  XOR U3453 ( .A(n3373), .B(n3374), .Z(n3384) );
  NANDN U3454 ( .A(n3295), .B(n3294), .Z(n3299) );
  OR U3455 ( .A(n3297), .B(n3296), .Z(n3298) );
  AND U3456 ( .A(n3299), .B(n3298), .Z(n3383) );
  XNOR U3457 ( .A(n3384), .B(n3383), .Z(n3385) );
  NANDN U3458 ( .A(n3301), .B(n3300), .Z(n3305) );
  NANDN U3459 ( .A(n3303), .B(n3302), .Z(n3304) );
  NAND U3460 ( .A(n3305), .B(n3304), .Z(n3386) );
  XNOR U3461 ( .A(n3385), .B(n3386), .Z(n3331) );
  XOR U3462 ( .A(n3332), .B(n3331), .Z(n3390) );
  NANDN U3463 ( .A(n3307), .B(n3306), .Z(n3311) );
  NANDN U3464 ( .A(n3309), .B(n3308), .Z(n3310) );
  AND U3465 ( .A(n3311), .B(n3310), .Z(n3389) );
  XNOR U3466 ( .A(n3390), .B(n3389), .Z(n3391) );
  XOR U3467 ( .A(n3392), .B(n3391), .Z(n3324) );
  NANDN U3468 ( .A(n3313), .B(n3312), .Z(n3317) );
  NAND U3469 ( .A(n3315), .B(n3314), .Z(n3316) );
  AND U3470 ( .A(n3317), .B(n3316), .Z(n3323) );
  XNOR U3471 ( .A(n3324), .B(n3323), .Z(n3325) );
  XNOR U3472 ( .A(n3326), .B(n3325), .Z(n3395) );
  XNOR U3473 ( .A(sreg[162]), .B(n3395), .Z(n3397) );
  NANDN U3474 ( .A(sreg[161]), .B(n3318), .Z(n3322) );
  NAND U3475 ( .A(n3320), .B(n3319), .Z(n3321) );
  NAND U3476 ( .A(n3322), .B(n3321), .Z(n3396) );
  XNOR U3477 ( .A(n3397), .B(n3396), .Z(c[162]) );
  NANDN U3478 ( .A(n3324), .B(n3323), .Z(n3328) );
  NANDN U3479 ( .A(n3326), .B(n3325), .Z(n3327) );
  AND U3480 ( .A(n3328), .B(n3327), .Z(n3403) );
  NANDN U3481 ( .A(n3330), .B(n3329), .Z(n3334) );
  NAND U3482 ( .A(n3332), .B(n3331), .Z(n3333) );
  AND U3483 ( .A(n3334), .B(n3333), .Z(n3469) );
  NANDN U3484 ( .A(n3336), .B(n3335), .Z(n3340) );
  NANDN U3485 ( .A(n3338), .B(n3337), .Z(n3339) );
  AND U3486 ( .A(n3340), .B(n3339), .Z(n3435) );
  NAND U3487 ( .A(b[0]), .B(a[51]), .Z(n3341) );
  XNOR U3488 ( .A(b[1]), .B(n3341), .Z(n3343) );
  NANDN U3489 ( .A(b[0]), .B(a[50]), .Z(n3342) );
  NAND U3490 ( .A(n3343), .B(n3342), .Z(n3415) );
  NANDN U3491 ( .A(n9891), .B(n3344), .Z(n3346) );
  XOR U3492 ( .A(b[13]), .B(a[39]), .Z(n3418) );
  NANDN U3493 ( .A(n9935), .B(n3418), .Z(n3345) );
  AND U3494 ( .A(n3346), .B(n3345), .Z(n3413) );
  AND U3495 ( .A(b[15]), .B(a[35]), .Z(n3412) );
  XNOR U3496 ( .A(n3413), .B(n3412), .Z(n3414) );
  XNOR U3497 ( .A(n3415), .B(n3414), .Z(n3433) );
  NANDN U3498 ( .A(n9437), .B(n3347), .Z(n3349) );
  XOR U3499 ( .A(b[5]), .B(a[47]), .Z(n3424) );
  NANDN U3500 ( .A(n9503), .B(n3424), .Z(n3348) );
  AND U3501 ( .A(n3349), .B(n3348), .Z(n3457) );
  NANDN U3502 ( .A(n9588), .B(n3350), .Z(n3352) );
  XOR U3503 ( .A(b[7]), .B(a[45]), .Z(n3427) );
  NANDN U3504 ( .A(n9639), .B(n3427), .Z(n3351) );
  AND U3505 ( .A(n3352), .B(n3351), .Z(n3455) );
  NANDN U3506 ( .A(n9374), .B(n3353), .Z(n3355) );
  XOR U3507 ( .A(b[3]), .B(a[49]), .Z(n3430) );
  NANDN U3508 ( .A(n9375), .B(n3430), .Z(n3354) );
  NAND U3509 ( .A(n3355), .B(n3354), .Z(n3454) );
  XNOR U3510 ( .A(n3455), .B(n3454), .Z(n3456) );
  XOR U3511 ( .A(n3457), .B(n3456), .Z(n3434) );
  XOR U3512 ( .A(n3433), .B(n3434), .Z(n3436) );
  XOR U3513 ( .A(n3435), .B(n3436), .Z(n3407) );
  NANDN U3514 ( .A(n3357), .B(n3356), .Z(n3361) );
  OR U3515 ( .A(n3359), .B(n3358), .Z(n3360) );
  AND U3516 ( .A(n3361), .B(n3360), .Z(n3406) );
  XNOR U3517 ( .A(n3407), .B(n3406), .Z(n3409) );
  NAND U3518 ( .A(n3362), .B(n9883), .Z(n3364) );
  XOR U3519 ( .A(b[11]), .B(a[41]), .Z(n3439) );
  NANDN U3520 ( .A(n9856), .B(n3439), .Z(n3363) );
  AND U3521 ( .A(n3364), .B(n3363), .Z(n3450) );
  NANDN U3522 ( .A(n10005), .B(n3365), .Z(n3367) );
  XOR U3523 ( .A(b[15]), .B(a[37]), .Z(n3442) );
  NANDN U3524 ( .A(n10006), .B(n3442), .Z(n3366) );
  AND U3525 ( .A(n3367), .B(n3366), .Z(n3449) );
  NANDN U3526 ( .A(n9685), .B(n3368), .Z(n3370) );
  XOR U3527 ( .A(b[9]), .B(a[43]), .Z(n3445) );
  NANDN U3528 ( .A(n9758), .B(n3445), .Z(n3369) );
  NAND U3529 ( .A(n3370), .B(n3369), .Z(n3448) );
  XOR U3530 ( .A(n3449), .B(n3448), .Z(n3451) );
  XOR U3531 ( .A(n3450), .B(n3451), .Z(n3461) );
  NANDN U3532 ( .A(n3372), .B(n3371), .Z(n3376) );
  OR U3533 ( .A(n3374), .B(n3373), .Z(n3375) );
  AND U3534 ( .A(n3376), .B(n3375), .Z(n3460) );
  XNOR U3535 ( .A(n3461), .B(n3460), .Z(n3462) );
  NANDN U3536 ( .A(n3378), .B(n3377), .Z(n3382) );
  NANDN U3537 ( .A(n3380), .B(n3379), .Z(n3381) );
  NAND U3538 ( .A(n3382), .B(n3381), .Z(n3463) );
  XNOR U3539 ( .A(n3462), .B(n3463), .Z(n3408) );
  XOR U3540 ( .A(n3409), .B(n3408), .Z(n3467) );
  NANDN U3541 ( .A(n3384), .B(n3383), .Z(n3388) );
  NANDN U3542 ( .A(n3386), .B(n3385), .Z(n3387) );
  AND U3543 ( .A(n3388), .B(n3387), .Z(n3466) );
  XNOR U3544 ( .A(n3467), .B(n3466), .Z(n3468) );
  XOR U3545 ( .A(n3469), .B(n3468), .Z(n3401) );
  NANDN U3546 ( .A(n3390), .B(n3389), .Z(n3394) );
  NAND U3547 ( .A(n3392), .B(n3391), .Z(n3393) );
  AND U3548 ( .A(n3394), .B(n3393), .Z(n3400) );
  XNOR U3549 ( .A(n3401), .B(n3400), .Z(n3402) );
  XNOR U3550 ( .A(n3403), .B(n3402), .Z(n3472) );
  XNOR U3551 ( .A(sreg[163]), .B(n3472), .Z(n3474) );
  NANDN U3552 ( .A(sreg[162]), .B(n3395), .Z(n3399) );
  NAND U3553 ( .A(n3397), .B(n3396), .Z(n3398) );
  NAND U3554 ( .A(n3399), .B(n3398), .Z(n3473) );
  XNOR U3555 ( .A(n3474), .B(n3473), .Z(c[163]) );
  NANDN U3556 ( .A(n3401), .B(n3400), .Z(n3405) );
  NANDN U3557 ( .A(n3403), .B(n3402), .Z(n3404) );
  AND U3558 ( .A(n3405), .B(n3404), .Z(n3480) );
  NANDN U3559 ( .A(n3407), .B(n3406), .Z(n3411) );
  NAND U3560 ( .A(n3409), .B(n3408), .Z(n3410) );
  AND U3561 ( .A(n3411), .B(n3410), .Z(n3546) );
  NANDN U3562 ( .A(n3413), .B(n3412), .Z(n3417) );
  NANDN U3563 ( .A(n3415), .B(n3414), .Z(n3416) );
  AND U3564 ( .A(n3417), .B(n3416), .Z(n3512) );
  NANDN U3565 ( .A(n9891), .B(n3418), .Z(n3420) );
  XOR U3566 ( .A(b[13]), .B(a[40]), .Z(n3498) );
  NANDN U3567 ( .A(n9935), .B(n3498), .Z(n3419) );
  AND U3568 ( .A(n3420), .B(n3419), .Z(n3490) );
  AND U3569 ( .A(b[15]), .B(a[36]), .Z(n3489) );
  XNOR U3570 ( .A(n3490), .B(n3489), .Z(n3491) );
  NAND U3571 ( .A(b[0]), .B(a[52]), .Z(n3421) );
  XNOR U3572 ( .A(b[1]), .B(n3421), .Z(n3423) );
  NANDN U3573 ( .A(b[0]), .B(a[51]), .Z(n3422) );
  NAND U3574 ( .A(n3423), .B(n3422), .Z(n3492) );
  XNOR U3575 ( .A(n3491), .B(n3492), .Z(n3510) );
  NANDN U3576 ( .A(n9437), .B(n3424), .Z(n3426) );
  XOR U3577 ( .A(b[5]), .B(a[48]), .Z(n3501) );
  NANDN U3578 ( .A(n9503), .B(n3501), .Z(n3425) );
  AND U3579 ( .A(n3426), .B(n3425), .Z(n3534) );
  NANDN U3580 ( .A(n9588), .B(n3427), .Z(n3429) );
  XOR U3581 ( .A(b[7]), .B(a[46]), .Z(n3504) );
  NANDN U3582 ( .A(n9639), .B(n3504), .Z(n3428) );
  AND U3583 ( .A(n3429), .B(n3428), .Z(n3532) );
  NANDN U3584 ( .A(n9374), .B(n3430), .Z(n3432) );
  XOR U3585 ( .A(b[3]), .B(a[50]), .Z(n3507) );
  NANDN U3586 ( .A(n9375), .B(n3507), .Z(n3431) );
  NAND U3587 ( .A(n3432), .B(n3431), .Z(n3531) );
  XNOR U3588 ( .A(n3532), .B(n3531), .Z(n3533) );
  XOR U3589 ( .A(n3534), .B(n3533), .Z(n3511) );
  XOR U3590 ( .A(n3510), .B(n3511), .Z(n3513) );
  XOR U3591 ( .A(n3512), .B(n3513), .Z(n3484) );
  NANDN U3592 ( .A(n3434), .B(n3433), .Z(n3438) );
  OR U3593 ( .A(n3436), .B(n3435), .Z(n3437) );
  AND U3594 ( .A(n3438), .B(n3437), .Z(n3483) );
  XNOR U3595 ( .A(n3484), .B(n3483), .Z(n3486) );
  NAND U3596 ( .A(n3439), .B(n9883), .Z(n3441) );
  XOR U3597 ( .A(b[11]), .B(a[42]), .Z(n3516) );
  NANDN U3598 ( .A(n9856), .B(n3516), .Z(n3440) );
  AND U3599 ( .A(n3441), .B(n3440), .Z(n3527) );
  NANDN U3600 ( .A(n10005), .B(n3442), .Z(n3444) );
  XOR U3601 ( .A(b[15]), .B(a[38]), .Z(n3519) );
  NANDN U3602 ( .A(n10006), .B(n3519), .Z(n3443) );
  AND U3603 ( .A(n3444), .B(n3443), .Z(n3526) );
  NANDN U3604 ( .A(n9685), .B(n3445), .Z(n3447) );
  XOR U3605 ( .A(b[9]), .B(a[44]), .Z(n3522) );
  NANDN U3606 ( .A(n9758), .B(n3522), .Z(n3446) );
  NAND U3607 ( .A(n3447), .B(n3446), .Z(n3525) );
  XOR U3608 ( .A(n3526), .B(n3525), .Z(n3528) );
  XOR U3609 ( .A(n3527), .B(n3528), .Z(n3538) );
  NANDN U3610 ( .A(n3449), .B(n3448), .Z(n3453) );
  OR U3611 ( .A(n3451), .B(n3450), .Z(n3452) );
  AND U3612 ( .A(n3453), .B(n3452), .Z(n3537) );
  XNOR U3613 ( .A(n3538), .B(n3537), .Z(n3539) );
  NANDN U3614 ( .A(n3455), .B(n3454), .Z(n3459) );
  NANDN U3615 ( .A(n3457), .B(n3456), .Z(n3458) );
  NAND U3616 ( .A(n3459), .B(n3458), .Z(n3540) );
  XNOR U3617 ( .A(n3539), .B(n3540), .Z(n3485) );
  XOR U3618 ( .A(n3486), .B(n3485), .Z(n3544) );
  NANDN U3619 ( .A(n3461), .B(n3460), .Z(n3465) );
  NANDN U3620 ( .A(n3463), .B(n3462), .Z(n3464) );
  AND U3621 ( .A(n3465), .B(n3464), .Z(n3543) );
  XNOR U3622 ( .A(n3544), .B(n3543), .Z(n3545) );
  XOR U3623 ( .A(n3546), .B(n3545), .Z(n3478) );
  NANDN U3624 ( .A(n3467), .B(n3466), .Z(n3471) );
  NAND U3625 ( .A(n3469), .B(n3468), .Z(n3470) );
  AND U3626 ( .A(n3471), .B(n3470), .Z(n3477) );
  XNOR U3627 ( .A(n3478), .B(n3477), .Z(n3479) );
  XNOR U3628 ( .A(n3480), .B(n3479), .Z(n3549) );
  XNOR U3629 ( .A(sreg[164]), .B(n3549), .Z(n3551) );
  NANDN U3630 ( .A(sreg[163]), .B(n3472), .Z(n3476) );
  NAND U3631 ( .A(n3474), .B(n3473), .Z(n3475) );
  NAND U3632 ( .A(n3476), .B(n3475), .Z(n3550) );
  XNOR U3633 ( .A(n3551), .B(n3550), .Z(c[164]) );
  NANDN U3634 ( .A(n3478), .B(n3477), .Z(n3482) );
  NANDN U3635 ( .A(n3480), .B(n3479), .Z(n3481) );
  AND U3636 ( .A(n3482), .B(n3481), .Z(n3557) );
  NANDN U3637 ( .A(n3484), .B(n3483), .Z(n3488) );
  NAND U3638 ( .A(n3486), .B(n3485), .Z(n3487) );
  AND U3639 ( .A(n3488), .B(n3487), .Z(n3623) );
  NANDN U3640 ( .A(n3490), .B(n3489), .Z(n3494) );
  NANDN U3641 ( .A(n3492), .B(n3491), .Z(n3493) );
  AND U3642 ( .A(n3494), .B(n3493), .Z(n3589) );
  NAND U3643 ( .A(b[0]), .B(a[53]), .Z(n3495) );
  XNOR U3644 ( .A(b[1]), .B(n3495), .Z(n3497) );
  NANDN U3645 ( .A(b[0]), .B(a[52]), .Z(n3496) );
  NAND U3646 ( .A(n3497), .B(n3496), .Z(n3569) );
  NANDN U3647 ( .A(n9891), .B(n3498), .Z(n3500) );
  XOR U3648 ( .A(b[13]), .B(a[41]), .Z(n3572) );
  NANDN U3649 ( .A(n9935), .B(n3572), .Z(n3499) );
  AND U3650 ( .A(n3500), .B(n3499), .Z(n3567) );
  AND U3651 ( .A(b[15]), .B(a[37]), .Z(n3566) );
  XNOR U3652 ( .A(n3567), .B(n3566), .Z(n3568) );
  XNOR U3653 ( .A(n3569), .B(n3568), .Z(n3587) );
  NANDN U3654 ( .A(n9437), .B(n3501), .Z(n3503) );
  XOR U3655 ( .A(b[5]), .B(a[49]), .Z(n3578) );
  NANDN U3656 ( .A(n9503), .B(n3578), .Z(n3502) );
  AND U3657 ( .A(n3503), .B(n3502), .Z(n3611) );
  NANDN U3658 ( .A(n9588), .B(n3504), .Z(n3506) );
  XOR U3659 ( .A(b[7]), .B(a[47]), .Z(n3581) );
  NANDN U3660 ( .A(n9639), .B(n3581), .Z(n3505) );
  AND U3661 ( .A(n3506), .B(n3505), .Z(n3609) );
  NANDN U3662 ( .A(n9374), .B(n3507), .Z(n3509) );
  XOR U3663 ( .A(b[3]), .B(a[51]), .Z(n3584) );
  NANDN U3664 ( .A(n9375), .B(n3584), .Z(n3508) );
  NAND U3665 ( .A(n3509), .B(n3508), .Z(n3608) );
  XNOR U3666 ( .A(n3609), .B(n3608), .Z(n3610) );
  XOR U3667 ( .A(n3611), .B(n3610), .Z(n3588) );
  XOR U3668 ( .A(n3587), .B(n3588), .Z(n3590) );
  XOR U3669 ( .A(n3589), .B(n3590), .Z(n3561) );
  NANDN U3670 ( .A(n3511), .B(n3510), .Z(n3515) );
  OR U3671 ( .A(n3513), .B(n3512), .Z(n3514) );
  AND U3672 ( .A(n3515), .B(n3514), .Z(n3560) );
  XNOR U3673 ( .A(n3561), .B(n3560), .Z(n3563) );
  NAND U3674 ( .A(n3516), .B(n9883), .Z(n3518) );
  XOR U3675 ( .A(b[11]), .B(a[43]), .Z(n3593) );
  NANDN U3676 ( .A(n9856), .B(n3593), .Z(n3517) );
  AND U3677 ( .A(n3518), .B(n3517), .Z(n3604) );
  NANDN U3678 ( .A(n10005), .B(n3519), .Z(n3521) );
  XOR U3679 ( .A(b[15]), .B(a[39]), .Z(n3596) );
  NANDN U3680 ( .A(n10006), .B(n3596), .Z(n3520) );
  AND U3681 ( .A(n3521), .B(n3520), .Z(n3603) );
  NANDN U3682 ( .A(n9685), .B(n3522), .Z(n3524) );
  XOR U3683 ( .A(b[9]), .B(a[45]), .Z(n3599) );
  NANDN U3684 ( .A(n9758), .B(n3599), .Z(n3523) );
  NAND U3685 ( .A(n3524), .B(n3523), .Z(n3602) );
  XOR U3686 ( .A(n3603), .B(n3602), .Z(n3605) );
  XOR U3687 ( .A(n3604), .B(n3605), .Z(n3615) );
  NANDN U3688 ( .A(n3526), .B(n3525), .Z(n3530) );
  OR U3689 ( .A(n3528), .B(n3527), .Z(n3529) );
  AND U3690 ( .A(n3530), .B(n3529), .Z(n3614) );
  XNOR U3691 ( .A(n3615), .B(n3614), .Z(n3616) );
  NANDN U3692 ( .A(n3532), .B(n3531), .Z(n3536) );
  NANDN U3693 ( .A(n3534), .B(n3533), .Z(n3535) );
  NAND U3694 ( .A(n3536), .B(n3535), .Z(n3617) );
  XNOR U3695 ( .A(n3616), .B(n3617), .Z(n3562) );
  XOR U3696 ( .A(n3563), .B(n3562), .Z(n3621) );
  NANDN U3697 ( .A(n3538), .B(n3537), .Z(n3542) );
  NANDN U3698 ( .A(n3540), .B(n3539), .Z(n3541) );
  AND U3699 ( .A(n3542), .B(n3541), .Z(n3620) );
  XNOR U3700 ( .A(n3621), .B(n3620), .Z(n3622) );
  XOR U3701 ( .A(n3623), .B(n3622), .Z(n3555) );
  NANDN U3702 ( .A(n3544), .B(n3543), .Z(n3548) );
  NAND U3703 ( .A(n3546), .B(n3545), .Z(n3547) );
  AND U3704 ( .A(n3548), .B(n3547), .Z(n3554) );
  XNOR U3705 ( .A(n3555), .B(n3554), .Z(n3556) );
  XNOR U3706 ( .A(n3557), .B(n3556), .Z(n3626) );
  XNOR U3707 ( .A(sreg[165]), .B(n3626), .Z(n3628) );
  NANDN U3708 ( .A(sreg[164]), .B(n3549), .Z(n3553) );
  NAND U3709 ( .A(n3551), .B(n3550), .Z(n3552) );
  NAND U3710 ( .A(n3553), .B(n3552), .Z(n3627) );
  XNOR U3711 ( .A(n3628), .B(n3627), .Z(c[165]) );
  NANDN U3712 ( .A(n3555), .B(n3554), .Z(n3559) );
  NANDN U3713 ( .A(n3557), .B(n3556), .Z(n3558) );
  AND U3714 ( .A(n3559), .B(n3558), .Z(n3634) );
  NANDN U3715 ( .A(n3561), .B(n3560), .Z(n3565) );
  NAND U3716 ( .A(n3563), .B(n3562), .Z(n3564) );
  AND U3717 ( .A(n3565), .B(n3564), .Z(n3700) );
  NANDN U3718 ( .A(n3567), .B(n3566), .Z(n3571) );
  NANDN U3719 ( .A(n3569), .B(n3568), .Z(n3570) );
  AND U3720 ( .A(n3571), .B(n3570), .Z(n3666) );
  NANDN U3721 ( .A(n9891), .B(n3572), .Z(n3574) );
  XOR U3722 ( .A(b[13]), .B(a[42]), .Z(n3652) );
  NANDN U3723 ( .A(n9935), .B(n3652), .Z(n3573) );
  AND U3724 ( .A(n3574), .B(n3573), .Z(n3644) );
  AND U3725 ( .A(b[15]), .B(a[38]), .Z(n3643) );
  XNOR U3726 ( .A(n3644), .B(n3643), .Z(n3645) );
  NAND U3727 ( .A(b[0]), .B(a[54]), .Z(n3575) );
  XNOR U3728 ( .A(b[1]), .B(n3575), .Z(n3577) );
  NANDN U3729 ( .A(b[0]), .B(a[53]), .Z(n3576) );
  NAND U3730 ( .A(n3577), .B(n3576), .Z(n3646) );
  XNOR U3731 ( .A(n3645), .B(n3646), .Z(n3664) );
  NANDN U3732 ( .A(n9437), .B(n3578), .Z(n3580) );
  XOR U3733 ( .A(b[5]), .B(a[50]), .Z(n3655) );
  NANDN U3734 ( .A(n9503), .B(n3655), .Z(n3579) );
  AND U3735 ( .A(n3580), .B(n3579), .Z(n3688) );
  NANDN U3736 ( .A(n9588), .B(n3581), .Z(n3583) );
  XOR U3737 ( .A(b[7]), .B(a[48]), .Z(n3658) );
  NANDN U3738 ( .A(n9639), .B(n3658), .Z(n3582) );
  AND U3739 ( .A(n3583), .B(n3582), .Z(n3686) );
  NANDN U3740 ( .A(n9374), .B(n3584), .Z(n3586) );
  XOR U3741 ( .A(b[3]), .B(a[52]), .Z(n3661) );
  NANDN U3742 ( .A(n9375), .B(n3661), .Z(n3585) );
  NAND U3743 ( .A(n3586), .B(n3585), .Z(n3685) );
  XNOR U3744 ( .A(n3686), .B(n3685), .Z(n3687) );
  XOR U3745 ( .A(n3688), .B(n3687), .Z(n3665) );
  XOR U3746 ( .A(n3664), .B(n3665), .Z(n3667) );
  XOR U3747 ( .A(n3666), .B(n3667), .Z(n3638) );
  NANDN U3748 ( .A(n3588), .B(n3587), .Z(n3592) );
  OR U3749 ( .A(n3590), .B(n3589), .Z(n3591) );
  AND U3750 ( .A(n3592), .B(n3591), .Z(n3637) );
  XNOR U3751 ( .A(n3638), .B(n3637), .Z(n3640) );
  NAND U3752 ( .A(n3593), .B(n9883), .Z(n3595) );
  XOR U3753 ( .A(b[11]), .B(a[44]), .Z(n3670) );
  NANDN U3754 ( .A(n9856), .B(n3670), .Z(n3594) );
  AND U3755 ( .A(n3595), .B(n3594), .Z(n3681) );
  NANDN U3756 ( .A(n10005), .B(n3596), .Z(n3598) );
  XOR U3757 ( .A(b[15]), .B(a[40]), .Z(n3673) );
  NANDN U3758 ( .A(n10006), .B(n3673), .Z(n3597) );
  AND U3759 ( .A(n3598), .B(n3597), .Z(n3680) );
  NANDN U3760 ( .A(n9685), .B(n3599), .Z(n3601) );
  XOR U3761 ( .A(b[9]), .B(a[46]), .Z(n3676) );
  NANDN U3762 ( .A(n9758), .B(n3676), .Z(n3600) );
  NAND U3763 ( .A(n3601), .B(n3600), .Z(n3679) );
  XOR U3764 ( .A(n3680), .B(n3679), .Z(n3682) );
  XOR U3765 ( .A(n3681), .B(n3682), .Z(n3692) );
  NANDN U3766 ( .A(n3603), .B(n3602), .Z(n3607) );
  OR U3767 ( .A(n3605), .B(n3604), .Z(n3606) );
  AND U3768 ( .A(n3607), .B(n3606), .Z(n3691) );
  XNOR U3769 ( .A(n3692), .B(n3691), .Z(n3693) );
  NANDN U3770 ( .A(n3609), .B(n3608), .Z(n3613) );
  NANDN U3771 ( .A(n3611), .B(n3610), .Z(n3612) );
  NAND U3772 ( .A(n3613), .B(n3612), .Z(n3694) );
  XNOR U3773 ( .A(n3693), .B(n3694), .Z(n3639) );
  XOR U3774 ( .A(n3640), .B(n3639), .Z(n3698) );
  NANDN U3775 ( .A(n3615), .B(n3614), .Z(n3619) );
  NANDN U3776 ( .A(n3617), .B(n3616), .Z(n3618) );
  AND U3777 ( .A(n3619), .B(n3618), .Z(n3697) );
  XNOR U3778 ( .A(n3698), .B(n3697), .Z(n3699) );
  XOR U3779 ( .A(n3700), .B(n3699), .Z(n3632) );
  NANDN U3780 ( .A(n3621), .B(n3620), .Z(n3625) );
  NAND U3781 ( .A(n3623), .B(n3622), .Z(n3624) );
  AND U3782 ( .A(n3625), .B(n3624), .Z(n3631) );
  XNOR U3783 ( .A(n3632), .B(n3631), .Z(n3633) );
  XNOR U3784 ( .A(n3634), .B(n3633), .Z(n3703) );
  XNOR U3785 ( .A(sreg[166]), .B(n3703), .Z(n3705) );
  NANDN U3786 ( .A(sreg[165]), .B(n3626), .Z(n3630) );
  NAND U3787 ( .A(n3628), .B(n3627), .Z(n3629) );
  NAND U3788 ( .A(n3630), .B(n3629), .Z(n3704) );
  XNOR U3789 ( .A(n3705), .B(n3704), .Z(c[166]) );
  NANDN U3790 ( .A(n3632), .B(n3631), .Z(n3636) );
  NANDN U3791 ( .A(n3634), .B(n3633), .Z(n3635) );
  AND U3792 ( .A(n3636), .B(n3635), .Z(n3711) );
  NANDN U3793 ( .A(n3638), .B(n3637), .Z(n3642) );
  NAND U3794 ( .A(n3640), .B(n3639), .Z(n3641) );
  AND U3795 ( .A(n3642), .B(n3641), .Z(n3777) );
  NANDN U3796 ( .A(n3644), .B(n3643), .Z(n3648) );
  NANDN U3797 ( .A(n3646), .B(n3645), .Z(n3647) );
  AND U3798 ( .A(n3648), .B(n3647), .Z(n3743) );
  NAND U3799 ( .A(b[0]), .B(a[55]), .Z(n3649) );
  XNOR U3800 ( .A(b[1]), .B(n3649), .Z(n3651) );
  NANDN U3801 ( .A(b[0]), .B(a[54]), .Z(n3650) );
  NAND U3802 ( .A(n3651), .B(n3650), .Z(n3723) );
  NANDN U3803 ( .A(n9891), .B(n3652), .Z(n3654) );
  XOR U3804 ( .A(b[13]), .B(a[43]), .Z(n3729) );
  NANDN U3805 ( .A(n9935), .B(n3729), .Z(n3653) );
  AND U3806 ( .A(n3654), .B(n3653), .Z(n3721) );
  AND U3807 ( .A(b[15]), .B(a[39]), .Z(n3720) );
  XNOR U3808 ( .A(n3721), .B(n3720), .Z(n3722) );
  XNOR U3809 ( .A(n3723), .B(n3722), .Z(n3741) );
  NANDN U3810 ( .A(n9437), .B(n3655), .Z(n3657) );
  XOR U3811 ( .A(b[5]), .B(a[51]), .Z(n3732) );
  NANDN U3812 ( .A(n9503), .B(n3732), .Z(n3656) );
  AND U3813 ( .A(n3657), .B(n3656), .Z(n3765) );
  NANDN U3814 ( .A(n9588), .B(n3658), .Z(n3660) );
  XOR U3815 ( .A(b[7]), .B(a[49]), .Z(n3735) );
  NANDN U3816 ( .A(n9639), .B(n3735), .Z(n3659) );
  AND U3817 ( .A(n3660), .B(n3659), .Z(n3763) );
  NANDN U3818 ( .A(n9374), .B(n3661), .Z(n3663) );
  XOR U3819 ( .A(b[3]), .B(a[53]), .Z(n3738) );
  NANDN U3820 ( .A(n9375), .B(n3738), .Z(n3662) );
  NAND U3821 ( .A(n3663), .B(n3662), .Z(n3762) );
  XNOR U3822 ( .A(n3763), .B(n3762), .Z(n3764) );
  XOR U3823 ( .A(n3765), .B(n3764), .Z(n3742) );
  XOR U3824 ( .A(n3741), .B(n3742), .Z(n3744) );
  XOR U3825 ( .A(n3743), .B(n3744), .Z(n3715) );
  NANDN U3826 ( .A(n3665), .B(n3664), .Z(n3669) );
  OR U3827 ( .A(n3667), .B(n3666), .Z(n3668) );
  AND U3828 ( .A(n3669), .B(n3668), .Z(n3714) );
  XNOR U3829 ( .A(n3715), .B(n3714), .Z(n3717) );
  NAND U3830 ( .A(n3670), .B(n9883), .Z(n3672) );
  XOR U3831 ( .A(b[11]), .B(a[45]), .Z(n3747) );
  NANDN U3832 ( .A(n9856), .B(n3747), .Z(n3671) );
  AND U3833 ( .A(n3672), .B(n3671), .Z(n3758) );
  NANDN U3834 ( .A(n10005), .B(n3673), .Z(n3675) );
  XOR U3835 ( .A(b[15]), .B(a[41]), .Z(n3750) );
  NANDN U3836 ( .A(n10006), .B(n3750), .Z(n3674) );
  AND U3837 ( .A(n3675), .B(n3674), .Z(n3757) );
  NANDN U3838 ( .A(n9685), .B(n3676), .Z(n3678) );
  XOR U3839 ( .A(b[9]), .B(a[47]), .Z(n3753) );
  NANDN U3840 ( .A(n9758), .B(n3753), .Z(n3677) );
  NAND U3841 ( .A(n3678), .B(n3677), .Z(n3756) );
  XOR U3842 ( .A(n3757), .B(n3756), .Z(n3759) );
  XOR U3843 ( .A(n3758), .B(n3759), .Z(n3769) );
  NANDN U3844 ( .A(n3680), .B(n3679), .Z(n3684) );
  OR U3845 ( .A(n3682), .B(n3681), .Z(n3683) );
  AND U3846 ( .A(n3684), .B(n3683), .Z(n3768) );
  XNOR U3847 ( .A(n3769), .B(n3768), .Z(n3770) );
  NANDN U3848 ( .A(n3686), .B(n3685), .Z(n3690) );
  NANDN U3849 ( .A(n3688), .B(n3687), .Z(n3689) );
  NAND U3850 ( .A(n3690), .B(n3689), .Z(n3771) );
  XNOR U3851 ( .A(n3770), .B(n3771), .Z(n3716) );
  XOR U3852 ( .A(n3717), .B(n3716), .Z(n3775) );
  NANDN U3853 ( .A(n3692), .B(n3691), .Z(n3696) );
  NANDN U3854 ( .A(n3694), .B(n3693), .Z(n3695) );
  AND U3855 ( .A(n3696), .B(n3695), .Z(n3774) );
  XNOR U3856 ( .A(n3775), .B(n3774), .Z(n3776) );
  XOR U3857 ( .A(n3777), .B(n3776), .Z(n3709) );
  NANDN U3858 ( .A(n3698), .B(n3697), .Z(n3702) );
  NAND U3859 ( .A(n3700), .B(n3699), .Z(n3701) );
  AND U3860 ( .A(n3702), .B(n3701), .Z(n3708) );
  XNOR U3861 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U3862 ( .A(n3711), .B(n3710), .Z(n3780) );
  XNOR U3863 ( .A(sreg[167]), .B(n3780), .Z(n3782) );
  NANDN U3864 ( .A(sreg[166]), .B(n3703), .Z(n3707) );
  NAND U3865 ( .A(n3705), .B(n3704), .Z(n3706) );
  NAND U3866 ( .A(n3707), .B(n3706), .Z(n3781) );
  XNOR U3867 ( .A(n3782), .B(n3781), .Z(c[167]) );
  NANDN U3868 ( .A(n3709), .B(n3708), .Z(n3713) );
  NANDN U3869 ( .A(n3711), .B(n3710), .Z(n3712) );
  AND U3870 ( .A(n3713), .B(n3712), .Z(n3788) );
  NANDN U3871 ( .A(n3715), .B(n3714), .Z(n3719) );
  NAND U3872 ( .A(n3717), .B(n3716), .Z(n3718) );
  AND U3873 ( .A(n3719), .B(n3718), .Z(n3854) );
  NANDN U3874 ( .A(n3721), .B(n3720), .Z(n3725) );
  NANDN U3875 ( .A(n3723), .B(n3722), .Z(n3724) );
  AND U3876 ( .A(n3725), .B(n3724), .Z(n3820) );
  NAND U3877 ( .A(b[0]), .B(a[56]), .Z(n3726) );
  XNOR U3878 ( .A(b[1]), .B(n3726), .Z(n3728) );
  NANDN U3879 ( .A(b[0]), .B(a[55]), .Z(n3727) );
  NAND U3880 ( .A(n3728), .B(n3727), .Z(n3800) );
  NANDN U3881 ( .A(n9891), .B(n3729), .Z(n3731) );
  XOR U3882 ( .A(b[13]), .B(a[44]), .Z(n3806) );
  NANDN U3883 ( .A(n9935), .B(n3806), .Z(n3730) );
  AND U3884 ( .A(n3731), .B(n3730), .Z(n3798) );
  AND U3885 ( .A(b[15]), .B(a[40]), .Z(n3797) );
  XNOR U3886 ( .A(n3798), .B(n3797), .Z(n3799) );
  XNOR U3887 ( .A(n3800), .B(n3799), .Z(n3818) );
  NANDN U3888 ( .A(n9437), .B(n3732), .Z(n3734) );
  XOR U3889 ( .A(b[5]), .B(a[52]), .Z(n3809) );
  NANDN U3890 ( .A(n9503), .B(n3809), .Z(n3733) );
  AND U3891 ( .A(n3734), .B(n3733), .Z(n3842) );
  NANDN U3892 ( .A(n9588), .B(n3735), .Z(n3737) );
  XOR U3893 ( .A(b[7]), .B(a[50]), .Z(n3812) );
  NANDN U3894 ( .A(n9639), .B(n3812), .Z(n3736) );
  AND U3895 ( .A(n3737), .B(n3736), .Z(n3840) );
  NANDN U3896 ( .A(n9374), .B(n3738), .Z(n3740) );
  XOR U3897 ( .A(b[3]), .B(a[54]), .Z(n3815) );
  NANDN U3898 ( .A(n9375), .B(n3815), .Z(n3739) );
  NAND U3899 ( .A(n3740), .B(n3739), .Z(n3839) );
  XNOR U3900 ( .A(n3840), .B(n3839), .Z(n3841) );
  XOR U3901 ( .A(n3842), .B(n3841), .Z(n3819) );
  XOR U3902 ( .A(n3818), .B(n3819), .Z(n3821) );
  XOR U3903 ( .A(n3820), .B(n3821), .Z(n3792) );
  NANDN U3904 ( .A(n3742), .B(n3741), .Z(n3746) );
  OR U3905 ( .A(n3744), .B(n3743), .Z(n3745) );
  AND U3906 ( .A(n3746), .B(n3745), .Z(n3791) );
  XNOR U3907 ( .A(n3792), .B(n3791), .Z(n3794) );
  NAND U3908 ( .A(n3747), .B(n9883), .Z(n3749) );
  XOR U3909 ( .A(b[11]), .B(a[46]), .Z(n3824) );
  NANDN U3910 ( .A(n9856), .B(n3824), .Z(n3748) );
  AND U3911 ( .A(n3749), .B(n3748), .Z(n3835) );
  NANDN U3912 ( .A(n10005), .B(n3750), .Z(n3752) );
  XOR U3913 ( .A(b[15]), .B(a[42]), .Z(n3827) );
  NANDN U3914 ( .A(n10006), .B(n3827), .Z(n3751) );
  AND U3915 ( .A(n3752), .B(n3751), .Z(n3834) );
  NANDN U3916 ( .A(n9685), .B(n3753), .Z(n3755) );
  XOR U3917 ( .A(b[9]), .B(a[48]), .Z(n3830) );
  NANDN U3918 ( .A(n9758), .B(n3830), .Z(n3754) );
  NAND U3919 ( .A(n3755), .B(n3754), .Z(n3833) );
  XOR U3920 ( .A(n3834), .B(n3833), .Z(n3836) );
  XOR U3921 ( .A(n3835), .B(n3836), .Z(n3846) );
  NANDN U3922 ( .A(n3757), .B(n3756), .Z(n3761) );
  OR U3923 ( .A(n3759), .B(n3758), .Z(n3760) );
  AND U3924 ( .A(n3761), .B(n3760), .Z(n3845) );
  XNOR U3925 ( .A(n3846), .B(n3845), .Z(n3847) );
  NANDN U3926 ( .A(n3763), .B(n3762), .Z(n3767) );
  NANDN U3927 ( .A(n3765), .B(n3764), .Z(n3766) );
  NAND U3928 ( .A(n3767), .B(n3766), .Z(n3848) );
  XNOR U3929 ( .A(n3847), .B(n3848), .Z(n3793) );
  XOR U3930 ( .A(n3794), .B(n3793), .Z(n3852) );
  NANDN U3931 ( .A(n3769), .B(n3768), .Z(n3773) );
  NANDN U3932 ( .A(n3771), .B(n3770), .Z(n3772) );
  AND U3933 ( .A(n3773), .B(n3772), .Z(n3851) );
  XNOR U3934 ( .A(n3852), .B(n3851), .Z(n3853) );
  XOR U3935 ( .A(n3854), .B(n3853), .Z(n3786) );
  NANDN U3936 ( .A(n3775), .B(n3774), .Z(n3779) );
  NAND U3937 ( .A(n3777), .B(n3776), .Z(n3778) );
  AND U3938 ( .A(n3779), .B(n3778), .Z(n3785) );
  XNOR U3939 ( .A(n3786), .B(n3785), .Z(n3787) );
  XNOR U3940 ( .A(n3788), .B(n3787), .Z(n3857) );
  XNOR U3941 ( .A(sreg[168]), .B(n3857), .Z(n3859) );
  NANDN U3942 ( .A(sreg[167]), .B(n3780), .Z(n3784) );
  NAND U3943 ( .A(n3782), .B(n3781), .Z(n3783) );
  NAND U3944 ( .A(n3784), .B(n3783), .Z(n3858) );
  XNOR U3945 ( .A(n3859), .B(n3858), .Z(c[168]) );
  NANDN U3946 ( .A(n3786), .B(n3785), .Z(n3790) );
  NANDN U3947 ( .A(n3788), .B(n3787), .Z(n3789) );
  AND U3948 ( .A(n3790), .B(n3789), .Z(n3865) );
  NANDN U3949 ( .A(n3792), .B(n3791), .Z(n3796) );
  NAND U3950 ( .A(n3794), .B(n3793), .Z(n3795) );
  AND U3951 ( .A(n3796), .B(n3795), .Z(n3931) );
  NANDN U3952 ( .A(n3798), .B(n3797), .Z(n3802) );
  NANDN U3953 ( .A(n3800), .B(n3799), .Z(n3801) );
  AND U3954 ( .A(n3802), .B(n3801), .Z(n3897) );
  NAND U3955 ( .A(b[0]), .B(a[57]), .Z(n3803) );
  XNOR U3956 ( .A(b[1]), .B(n3803), .Z(n3805) );
  NANDN U3957 ( .A(b[0]), .B(a[56]), .Z(n3804) );
  NAND U3958 ( .A(n3805), .B(n3804), .Z(n3877) );
  NANDN U3959 ( .A(n9891), .B(n3806), .Z(n3808) );
  XOR U3960 ( .A(b[13]), .B(a[45]), .Z(n3883) );
  NANDN U3961 ( .A(n9935), .B(n3883), .Z(n3807) );
  AND U3962 ( .A(n3808), .B(n3807), .Z(n3875) );
  AND U3963 ( .A(b[15]), .B(a[41]), .Z(n3874) );
  XNOR U3964 ( .A(n3875), .B(n3874), .Z(n3876) );
  XNOR U3965 ( .A(n3877), .B(n3876), .Z(n3895) );
  NANDN U3966 ( .A(n9437), .B(n3809), .Z(n3811) );
  XOR U3967 ( .A(b[5]), .B(a[53]), .Z(n3886) );
  NANDN U3968 ( .A(n9503), .B(n3886), .Z(n3810) );
  AND U3969 ( .A(n3811), .B(n3810), .Z(n3919) );
  NANDN U3970 ( .A(n9588), .B(n3812), .Z(n3814) );
  XOR U3971 ( .A(b[7]), .B(a[51]), .Z(n3889) );
  NANDN U3972 ( .A(n9639), .B(n3889), .Z(n3813) );
  AND U3973 ( .A(n3814), .B(n3813), .Z(n3917) );
  NANDN U3974 ( .A(n9374), .B(n3815), .Z(n3817) );
  XOR U3975 ( .A(b[3]), .B(a[55]), .Z(n3892) );
  NANDN U3976 ( .A(n9375), .B(n3892), .Z(n3816) );
  NAND U3977 ( .A(n3817), .B(n3816), .Z(n3916) );
  XNOR U3978 ( .A(n3917), .B(n3916), .Z(n3918) );
  XOR U3979 ( .A(n3919), .B(n3918), .Z(n3896) );
  XOR U3980 ( .A(n3895), .B(n3896), .Z(n3898) );
  XOR U3981 ( .A(n3897), .B(n3898), .Z(n3869) );
  NANDN U3982 ( .A(n3819), .B(n3818), .Z(n3823) );
  OR U3983 ( .A(n3821), .B(n3820), .Z(n3822) );
  AND U3984 ( .A(n3823), .B(n3822), .Z(n3868) );
  XNOR U3985 ( .A(n3869), .B(n3868), .Z(n3871) );
  NAND U3986 ( .A(n3824), .B(n9883), .Z(n3826) );
  XOR U3987 ( .A(b[11]), .B(a[47]), .Z(n3901) );
  NANDN U3988 ( .A(n9856), .B(n3901), .Z(n3825) );
  AND U3989 ( .A(n3826), .B(n3825), .Z(n3912) );
  NANDN U3990 ( .A(n10005), .B(n3827), .Z(n3829) );
  XOR U3991 ( .A(b[15]), .B(a[43]), .Z(n3904) );
  NANDN U3992 ( .A(n10006), .B(n3904), .Z(n3828) );
  AND U3993 ( .A(n3829), .B(n3828), .Z(n3911) );
  NANDN U3994 ( .A(n9685), .B(n3830), .Z(n3832) );
  XOR U3995 ( .A(b[9]), .B(a[49]), .Z(n3907) );
  NANDN U3996 ( .A(n9758), .B(n3907), .Z(n3831) );
  NAND U3997 ( .A(n3832), .B(n3831), .Z(n3910) );
  XOR U3998 ( .A(n3911), .B(n3910), .Z(n3913) );
  XOR U3999 ( .A(n3912), .B(n3913), .Z(n3923) );
  NANDN U4000 ( .A(n3834), .B(n3833), .Z(n3838) );
  OR U4001 ( .A(n3836), .B(n3835), .Z(n3837) );
  AND U4002 ( .A(n3838), .B(n3837), .Z(n3922) );
  XNOR U4003 ( .A(n3923), .B(n3922), .Z(n3924) );
  NANDN U4004 ( .A(n3840), .B(n3839), .Z(n3844) );
  NANDN U4005 ( .A(n3842), .B(n3841), .Z(n3843) );
  NAND U4006 ( .A(n3844), .B(n3843), .Z(n3925) );
  XNOR U4007 ( .A(n3924), .B(n3925), .Z(n3870) );
  XOR U4008 ( .A(n3871), .B(n3870), .Z(n3929) );
  NANDN U4009 ( .A(n3846), .B(n3845), .Z(n3850) );
  NANDN U4010 ( .A(n3848), .B(n3847), .Z(n3849) );
  AND U4011 ( .A(n3850), .B(n3849), .Z(n3928) );
  XNOR U4012 ( .A(n3929), .B(n3928), .Z(n3930) );
  XOR U4013 ( .A(n3931), .B(n3930), .Z(n3863) );
  NANDN U4014 ( .A(n3852), .B(n3851), .Z(n3856) );
  NAND U4015 ( .A(n3854), .B(n3853), .Z(n3855) );
  AND U4016 ( .A(n3856), .B(n3855), .Z(n3862) );
  XNOR U4017 ( .A(n3863), .B(n3862), .Z(n3864) );
  XNOR U4018 ( .A(n3865), .B(n3864), .Z(n3934) );
  XNOR U4019 ( .A(sreg[169]), .B(n3934), .Z(n3936) );
  NANDN U4020 ( .A(sreg[168]), .B(n3857), .Z(n3861) );
  NAND U4021 ( .A(n3859), .B(n3858), .Z(n3860) );
  NAND U4022 ( .A(n3861), .B(n3860), .Z(n3935) );
  XNOR U4023 ( .A(n3936), .B(n3935), .Z(c[169]) );
  NANDN U4024 ( .A(n3863), .B(n3862), .Z(n3867) );
  NANDN U4025 ( .A(n3865), .B(n3864), .Z(n3866) );
  AND U4026 ( .A(n3867), .B(n3866), .Z(n3942) );
  NANDN U4027 ( .A(n3869), .B(n3868), .Z(n3873) );
  NAND U4028 ( .A(n3871), .B(n3870), .Z(n3872) );
  AND U4029 ( .A(n3873), .B(n3872), .Z(n4008) );
  NANDN U4030 ( .A(n3875), .B(n3874), .Z(n3879) );
  NANDN U4031 ( .A(n3877), .B(n3876), .Z(n3878) );
  AND U4032 ( .A(n3879), .B(n3878), .Z(n3995) );
  NAND U4033 ( .A(b[0]), .B(a[58]), .Z(n3880) );
  XNOR U4034 ( .A(b[1]), .B(n3880), .Z(n3882) );
  NANDN U4035 ( .A(b[0]), .B(a[57]), .Z(n3881) );
  NAND U4036 ( .A(n3882), .B(n3881), .Z(n3975) );
  NANDN U4037 ( .A(n9891), .B(n3883), .Z(n3885) );
  XOR U4038 ( .A(b[13]), .B(a[46]), .Z(n3978) );
  NANDN U4039 ( .A(n9935), .B(n3978), .Z(n3884) );
  AND U4040 ( .A(n3885), .B(n3884), .Z(n3973) );
  AND U4041 ( .A(b[15]), .B(a[42]), .Z(n3972) );
  XNOR U4042 ( .A(n3973), .B(n3972), .Z(n3974) );
  XNOR U4043 ( .A(n3975), .B(n3974), .Z(n3993) );
  NANDN U4044 ( .A(n9437), .B(n3886), .Z(n3888) );
  XOR U4045 ( .A(b[5]), .B(a[54]), .Z(n3984) );
  NANDN U4046 ( .A(n9503), .B(n3984), .Z(n3887) );
  AND U4047 ( .A(n3888), .B(n3887), .Z(n3969) );
  NANDN U4048 ( .A(n9588), .B(n3889), .Z(n3891) );
  XOR U4049 ( .A(b[7]), .B(a[52]), .Z(n3987) );
  NANDN U4050 ( .A(n9639), .B(n3987), .Z(n3890) );
  AND U4051 ( .A(n3891), .B(n3890), .Z(n3967) );
  NANDN U4052 ( .A(n9374), .B(n3892), .Z(n3894) );
  XOR U4053 ( .A(b[3]), .B(a[56]), .Z(n3990) );
  NANDN U4054 ( .A(n9375), .B(n3990), .Z(n3893) );
  NAND U4055 ( .A(n3894), .B(n3893), .Z(n3966) );
  XNOR U4056 ( .A(n3967), .B(n3966), .Z(n3968) );
  XOR U4057 ( .A(n3969), .B(n3968), .Z(n3994) );
  XOR U4058 ( .A(n3993), .B(n3994), .Z(n3996) );
  XOR U4059 ( .A(n3995), .B(n3996), .Z(n3946) );
  NANDN U4060 ( .A(n3896), .B(n3895), .Z(n3900) );
  OR U4061 ( .A(n3898), .B(n3897), .Z(n3899) );
  AND U4062 ( .A(n3900), .B(n3899), .Z(n3945) );
  XNOR U4063 ( .A(n3946), .B(n3945), .Z(n3948) );
  NAND U4064 ( .A(n3901), .B(n9883), .Z(n3903) );
  XOR U4065 ( .A(b[11]), .B(a[48]), .Z(n3951) );
  NANDN U4066 ( .A(n9856), .B(n3951), .Z(n3902) );
  AND U4067 ( .A(n3903), .B(n3902), .Z(n3962) );
  NANDN U4068 ( .A(n10005), .B(n3904), .Z(n3906) );
  XOR U4069 ( .A(b[15]), .B(a[44]), .Z(n3954) );
  NANDN U4070 ( .A(n10006), .B(n3954), .Z(n3905) );
  AND U4071 ( .A(n3906), .B(n3905), .Z(n3961) );
  NANDN U4072 ( .A(n9685), .B(n3907), .Z(n3909) );
  XOR U4073 ( .A(b[9]), .B(a[50]), .Z(n3957) );
  NANDN U4074 ( .A(n9758), .B(n3957), .Z(n3908) );
  NAND U4075 ( .A(n3909), .B(n3908), .Z(n3960) );
  XOR U4076 ( .A(n3961), .B(n3960), .Z(n3963) );
  XOR U4077 ( .A(n3962), .B(n3963), .Z(n4000) );
  NANDN U4078 ( .A(n3911), .B(n3910), .Z(n3915) );
  OR U4079 ( .A(n3913), .B(n3912), .Z(n3914) );
  AND U4080 ( .A(n3915), .B(n3914), .Z(n3999) );
  XNOR U4081 ( .A(n4000), .B(n3999), .Z(n4001) );
  NANDN U4082 ( .A(n3917), .B(n3916), .Z(n3921) );
  NANDN U4083 ( .A(n3919), .B(n3918), .Z(n3920) );
  NAND U4084 ( .A(n3921), .B(n3920), .Z(n4002) );
  XNOR U4085 ( .A(n4001), .B(n4002), .Z(n3947) );
  XOR U4086 ( .A(n3948), .B(n3947), .Z(n4006) );
  NANDN U4087 ( .A(n3923), .B(n3922), .Z(n3927) );
  NANDN U4088 ( .A(n3925), .B(n3924), .Z(n3926) );
  AND U4089 ( .A(n3927), .B(n3926), .Z(n4005) );
  XNOR U4090 ( .A(n4006), .B(n4005), .Z(n4007) );
  XOR U4091 ( .A(n4008), .B(n4007), .Z(n3940) );
  NANDN U4092 ( .A(n3929), .B(n3928), .Z(n3933) );
  NAND U4093 ( .A(n3931), .B(n3930), .Z(n3932) );
  AND U4094 ( .A(n3933), .B(n3932), .Z(n3939) );
  XNOR U4095 ( .A(n3940), .B(n3939), .Z(n3941) );
  XNOR U4096 ( .A(n3942), .B(n3941), .Z(n4011) );
  XNOR U4097 ( .A(sreg[170]), .B(n4011), .Z(n4013) );
  NANDN U4098 ( .A(sreg[169]), .B(n3934), .Z(n3938) );
  NAND U4099 ( .A(n3936), .B(n3935), .Z(n3937) );
  NAND U4100 ( .A(n3938), .B(n3937), .Z(n4012) );
  XNOR U4101 ( .A(n4013), .B(n4012), .Z(c[170]) );
  NANDN U4102 ( .A(n3940), .B(n3939), .Z(n3944) );
  NANDN U4103 ( .A(n3942), .B(n3941), .Z(n3943) );
  AND U4104 ( .A(n3944), .B(n3943), .Z(n4019) );
  NANDN U4105 ( .A(n3946), .B(n3945), .Z(n3950) );
  NAND U4106 ( .A(n3948), .B(n3947), .Z(n3949) );
  AND U4107 ( .A(n3950), .B(n3949), .Z(n4085) );
  NAND U4108 ( .A(n3951), .B(n9883), .Z(n3953) );
  XOR U4109 ( .A(b[11]), .B(a[49]), .Z(n4028) );
  NANDN U4110 ( .A(n9856), .B(n4028), .Z(n3952) );
  AND U4111 ( .A(n3953), .B(n3952), .Z(n4039) );
  NANDN U4112 ( .A(n10005), .B(n3954), .Z(n3956) );
  XOR U4113 ( .A(b[15]), .B(a[45]), .Z(n4031) );
  NANDN U4114 ( .A(n10006), .B(n4031), .Z(n3955) );
  AND U4115 ( .A(n3956), .B(n3955), .Z(n4038) );
  NANDN U4116 ( .A(n9685), .B(n3957), .Z(n3959) );
  XOR U4117 ( .A(b[9]), .B(a[51]), .Z(n4034) );
  NANDN U4118 ( .A(n9758), .B(n4034), .Z(n3958) );
  NAND U4119 ( .A(n3959), .B(n3958), .Z(n4037) );
  XOR U4120 ( .A(n4038), .B(n4037), .Z(n4040) );
  XOR U4121 ( .A(n4039), .B(n4040), .Z(n4077) );
  NANDN U4122 ( .A(n3961), .B(n3960), .Z(n3965) );
  OR U4123 ( .A(n3963), .B(n3962), .Z(n3964) );
  AND U4124 ( .A(n3965), .B(n3964), .Z(n4076) );
  XNOR U4125 ( .A(n4077), .B(n4076), .Z(n4078) );
  NANDN U4126 ( .A(n3967), .B(n3966), .Z(n3971) );
  NANDN U4127 ( .A(n3969), .B(n3968), .Z(n3970) );
  NAND U4128 ( .A(n3971), .B(n3970), .Z(n4079) );
  XNOR U4129 ( .A(n4078), .B(n4079), .Z(n4025) );
  NANDN U4130 ( .A(n3973), .B(n3972), .Z(n3977) );
  NANDN U4131 ( .A(n3975), .B(n3974), .Z(n3976) );
  AND U4132 ( .A(n3977), .B(n3976), .Z(n4072) );
  NANDN U4133 ( .A(n9891), .B(n3978), .Z(n3980) );
  XOR U4134 ( .A(b[13]), .B(a[47]), .Z(n4058) );
  NANDN U4135 ( .A(n9935), .B(n4058), .Z(n3979) );
  AND U4136 ( .A(n3980), .B(n3979), .Z(n4050) );
  AND U4137 ( .A(b[15]), .B(a[43]), .Z(n4049) );
  XNOR U4138 ( .A(n4050), .B(n4049), .Z(n4051) );
  NAND U4139 ( .A(b[0]), .B(a[59]), .Z(n3981) );
  XNOR U4140 ( .A(b[1]), .B(n3981), .Z(n3983) );
  NANDN U4141 ( .A(b[0]), .B(a[58]), .Z(n3982) );
  NAND U4142 ( .A(n3983), .B(n3982), .Z(n4052) );
  XNOR U4143 ( .A(n4051), .B(n4052), .Z(n4070) );
  NANDN U4144 ( .A(n9437), .B(n3984), .Z(n3986) );
  XOR U4145 ( .A(b[5]), .B(a[55]), .Z(n4061) );
  NANDN U4146 ( .A(n9503), .B(n4061), .Z(n3985) );
  AND U4147 ( .A(n3986), .B(n3985), .Z(n4046) );
  NANDN U4148 ( .A(n9588), .B(n3987), .Z(n3989) );
  XOR U4149 ( .A(b[7]), .B(a[53]), .Z(n4064) );
  NANDN U4150 ( .A(n9639), .B(n4064), .Z(n3988) );
  AND U4151 ( .A(n3989), .B(n3988), .Z(n4044) );
  NANDN U4152 ( .A(n9374), .B(n3990), .Z(n3992) );
  XOR U4153 ( .A(b[3]), .B(a[57]), .Z(n4067) );
  NANDN U4154 ( .A(n9375), .B(n4067), .Z(n3991) );
  NAND U4155 ( .A(n3992), .B(n3991), .Z(n4043) );
  XNOR U4156 ( .A(n4044), .B(n4043), .Z(n4045) );
  XOR U4157 ( .A(n4046), .B(n4045), .Z(n4071) );
  XOR U4158 ( .A(n4070), .B(n4071), .Z(n4073) );
  XOR U4159 ( .A(n4072), .B(n4073), .Z(n4023) );
  NANDN U4160 ( .A(n3994), .B(n3993), .Z(n3998) );
  OR U4161 ( .A(n3996), .B(n3995), .Z(n3997) );
  AND U4162 ( .A(n3998), .B(n3997), .Z(n4022) );
  XNOR U4163 ( .A(n4023), .B(n4022), .Z(n4024) );
  XOR U4164 ( .A(n4025), .B(n4024), .Z(n4083) );
  NANDN U4165 ( .A(n4000), .B(n3999), .Z(n4004) );
  NANDN U4166 ( .A(n4002), .B(n4001), .Z(n4003) );
  AND U4167 ( .A(n4004), .B(n4003), .Z(n4082) );
  XNOR U4168 ( .A(n4083), .B(n4082), .Z(n4084) );
  XOR U4169 ( .A(n4085), .B(n4084), .Z(n4017) );
  NANDN U4170 ( .A(n4006), .B(n4005), .Z(n4010) );
  NAND U4171 ( .A(n4008), .B(n4007), .Z(n4009) );
  AND U4172 ( .A(n4010), .B(n4009), .Z(n4016) );
  XNOR U4173 ( .A(n4017), .B(n4016), .Z(n4018) );
  XNOR U4174 ( .A(n4019), .B(n4018), .Z(n4088) );
  XNOR U4175 ( .A(sreg[171]), .B(n4088), .Z(n4090) );
  NANDN U4176 ( .A(sreg[170]), .B(n4011), .Z(n4015) );
  NAND U4177 ( .A(n4013), .B(n4012), .Z(n4014) );
  NAND U4178 ( .A(n4015), .B(n4014), .Z(n4089) );
  XNOR U4179 ( .A(n4090), .B(n4089), .Z(c[171]) );
  NANDN U4180 ( .A(n4017), .B(n4016), .Z(n4021) );
  NANDN U4181 ( .A(n4019), .B(n4018), .Z(n4020) );
  AND U4182 ( .A(n4021), .B(n4020), .Z(n4096) );
  NANDN U4183 ( .A(n4023), .B(n4022), .Z(n4027) );
  NAND U4184 ( .A(n4025), .B(n4024), .Z(n4026) );
  AND U4185 ( .A(n4027), .B(n4026), .Z(n4162) );
  NAND U4186 ( .A(n4028), .B(n9883), .Z(n4030) );
  XOR U4187 ( .A(b[11]), .B(a[50]), .Z(n4132) );
  NANDN U4188 ( .A(n9856), .B(n4132), .Z(n4029) );
  AND U4189 ( .A(n4030), .B(n4029), .Z(n4143) );
  NANDN U4190 ( .A(n10005), .B(n4031), .Z(n4033) );
  XOR U4191 ( .A(b[15]), .B(a[46]), .Z(n4135) );
  NANDN U4192 ( .A(n10006), .B(n4135), .Z(n4032) );
  AND U4193 ( .A(n4033), .B(n4032), .Z(n4142) );
  NANDN U4194 ( .A(n9685), .B(n4034), .Z(n4036) );
  XOR U4195 ( .A(b[9]), .B(a[52]), .Z(n4138) );
  NANDN U4196 ( .A(n9758), .B(n4138), .Z(n4035) );
  NAND U4197 ( .A(n4036), .B(n4035), .Z(n4141) );
  XOR U4198 ( .A(n4142), .B(n4141), .Z(n4144) );
  XOR U4199 ( .A(n4143), .B(n4144), .Z(n4154) );
  NANDN U4200 ( .A(n4038), .B(n4037), .Z(n4042) );
  OR U4201 ( .A(n4040), .B(n4039), .Z(n4041) );
  AND U4202 ( .A(n4042), .B(n4041), .Z(n4153) );
  XNOR U4203 ( .A(n4154), .B(n4153), .Z(n4155) );
  NANDN U4204 ( .A(n4044), .B(n4043), .Z(n4048) );
  NANDN U4205 ( .A(n4046), .B(n4045), .Z(n4047) );
  NAND U4206 ( .A(n4048), .B(n4047), .Z(n4156) );
  XNOR U4207 ( .A(n4155), .B(n4156), .Z(n4102) );
  NANDN U4208 ( .A(n4050), .B(n4049), .Z(n4054) );
  NANDN U4209 ( .A(n4052), .B(n4051), .Z(n4053) );
  AND U4210 ( .A(n4054), .B(n4053), .Z(n4128) );
  NAND U4211 ( .A(b[0]), .B(a[60]), .Z(n4055) );
  XNOR U4212 ( .A(b[1]), .B(n4055), .Z(n4057) );
  NANDN U4213 ( .A(b[0]), .B(a[59]), .Z(n4056) );
  NAND U4214 ( .A(n4057), .B(n4056), .Z(n4108) );
  NANDN U4215 ( .A(n9891), .B(n4058), .Z(n4060) );
  XOR U4216 ( .A(b[13]), .B(a[48]), .Z(n4111) );
  NANDN U4217 ( .A(n9935), .B(n4111), .Z(n4059) );
  AND U4218 ( .A(n4060), .B(n4059), .Z(n4106) );
  AND U4219 ( .A(b[15]), .B(a[44]), .Z(n4105) );
  XNOR U4220 ( .A(n4106), .B(n4105), .Z(n4107) );
  XNOR U4221 ( .A(n4108), .B(n4107), .Z(n4126) );
  NANDN U4222 ( .A(n9437), .B(n4061), .Z(n4063) );
  XOR U4223 ( .A(b[5]), .B(a[56]), .Z(n4117) );
  NANDN U4224 ( .A(n9503), .B(n4117), .Z(n4062) );
  AND U4225 ( .A(n4063), .B(n4062), .Z(n4150) );
  NANDN U4226 ( .A(n9588), .B(n4064), .Z(n4066) );
  XOR U4227 ( .A(b[7]), .B(a[54]), .Z(n4120) );
  NANDN U4228 ( .A(n9639), .B(n4120), .Z(n4065) );
  AND U4229 ( .A(n4066), .B(n4065), .Z(n4148) );
  NANDN U4230 ( .A(n9374), .B(n4067), .Z(n4069) );
  XOR U4231 ( .A(b[3]), .B(a[58]), .Z(n4123) );
  NANDN U4232 ( .A(n9375), .B(n4123), .Z(n4068) );
  NAND U4233 ( .A(n4069), .B(n4068), .Z(n4147) );
  XNOR U4234 ( .A(n4148), .B(n4147), .Z(n4149) );
  XOR U4235 ( .A(n4150), .B(n4149), .Z(n4127) );
  XOR U4236 ( .A(n4126), .B(n4127), .Z(n4129) );
  XOR U4237 ( .A(n4128), .B(n4129), .Z(n4100) );
  NANDN U4238 ( .A(n4071), .B(n4070), .Z(n4075) );
  OR U4239 ( .A(n4073), .B(n4072), .Z(n4074) );
  AND U4240 ( .A(n4075), .B(n4074), .Z(n4099) );
  XNOR U4241 ( .A(n4100), .B(n4099), .Z(n4101) );
  XOR U4242 ( .A(n4102), .B(n4101), .Z(n4160) );
  NANDN U4243 ( .A(n4077), .B(n4076), .Z(n4081) );
  NANDN U4244 ( .A(n4079), .B(n4078), .Z(n4080) );
  AND U4245 ( .A(n4081), .B(n4080), .Z(n4159) );
  XNOR U4246 ( .A(n4160), .B(n4159), .Z(n4161) );
  XOR U4247 ( .A(n4162), .B(n4161), .Z(n4094) );
  NANDN U4248 ( .A(n4083), .B(n4082), .Z(n4087) );
  NAND U4249 ( .A(n4085), .B(n4084), .Z(n4086) );
  AND U4250 ( .A(n4087), .B(n4086), .Z(n4093) );
  XNOR U4251 ( .A(n4094), .B(n4093), .Z(n4095) );
  XNOR U4252 ( .A(n4096), .B(n4095), .Z(n4165) );
  XNOR U4253 ( .A(sreg[172]), .B(n4165), .Z(n4167) );
  NANDN U4254 ( .A(sreg[171]), .B(n4088), .Z(n4092) );
  NAND U4255 ( .A(n4090), .B(n4089), .Z(n4091) );
  NAND U4256 ( .A(n4092), .B(n4091), .Z(n4166) );
  XNOR U4257 ( .A(n4167), .B(n4166), .Z(c[172]) );
  NANDN U4258 ( .A(n4094), .B(n4093), .Z(n4098) );
  NANDN U4259 ( .A(n4096), .B(n4095), .Z(n4097) );
  AND U4260 ( .A(n4098), .B(n4097), .Z(n4173) );
  NANDN U4261 ( .A(n4100), .B(n4099), .Z(n4104) );
  NAND U4262 ( .A(n4102), .B(n4101), .Z(n4103) );
  AND U4263 ( .A(n4104), .B(n4103), .Z(n4239) );
  NANDN U4264 ( .A(n4106), .B(n4105), .Z(n4110) );
  NANDN U4265 ( .A(n4108), .B(n4107), .Z(n4109) );
  AND U4266 ( .A(n4110), .B(n4109), .Z(n4205) );
  NANDN U4267 ( .A(n9891), .B(n4111), .Z(n4113) );
  XOR U4268 ( .A(b[13]), .B(a[49]), .Z(n4191) );
  NANDN U4269 ( .A(n9935), .B(n4191), .Z(n4112) );
  AND U4270 ( .A(n4113), .B(n4112), .Z(n4183) );
  AND U4271 ( .A(b[15]), .B(a[45]), .Z(n4182) );
  XNOR U4272 ( .A(n4183), .B(n4182), .Z(n4184) );
  NAND U4273 ( .A(b[0]), .B(a[61]), .Z(n4114) );
  XNOR U4274 ( .A(b[1]), .B(n4114), .Z(n4116) );
  NANDN U4275 ( .A(b[0]), .B(a[60]), .Z(n4115) );
  NAND U4276 ( .A(n4116), .B(n4115), .Z(n4185) );
  XNOR U4277 ( .A(n4184), .B(n4185), .Z(n4203) );
  NANDN U4278 ( .A(n9437), .B(n4117), .Z(n4119) );
  XOR U4279 ( .A(b[5]), .B(a[57]), .Z(n4194) );
  NANDN U4280 ( .A(n9503), .B(n4194), .Z(n4118) );
  AND U4281 ( .A(n4119), .B(n4118), .Z(n4227) );
  NANDN U4282 ( .A(n9588), .B(n4120), .Z(n4122) );
  XOR U4283 ( .A(b[7]), .B(a[55]), .Z(n4197) );
  NANDN U4284 ( .A(n9639), .B(n4197), .Z(n4121) );
  AND U4285 ( .A(n4122), .B(n4121), .Z(n4225) );
  NANDN U4286 ( .A(n9374), .B(n4123), .Z(n4125) );
  XOR U4287 ( .A(b[3]), .B(a[59]), .Z(n4200) );
  NANDN U4288 ( .A(n9375), .B(n4200), .Z(n4124) );
  NAND U4289 ( .A(n4125), .B(n4124), .Z(n4224) );
  XNOR U4290 ( .A(n4225), .B(n4224), .Z(n4226) );
  XOR U4291 ( .A(n4227), .B(n4226), .Z(n4204) );
  XOR U4292 ( .A(n4203), .B(n4204), .Z(n4206) );
  XOR U4293 ( .A(n4205), .B(n4206), .Z(n4177) );
  NANDN U4294 ( .A(n4127), .B(n4126), .Z(n4131) );
  OR U4295 ( .A(n4129), .B(n4128), .Z(n4130) );
  AND U4296 ( .A(n4131), .B(n4130), .Z(n4176) );
  XNOR U4297 ( .A(n4177), .B(n4176), .Z(n4179) );
  NAND U4298 ( .A(n4132), .B(n9883), .Z(n4134) );
  XOR U4299 ( .A(b[11]), .B(a[51]), .Z(n4209) );
  NANDN U4300 ( .A(n9856), .B(n4209), .Z(n4133) );
  AND U4301 ( .A(n4134), .B(n4133), .Z(n4220) );
  NANDN U4302 ( .A(n10005), .B(n4135), .Z(n4137) );
  XOR U4303 ( .A(b[15]), .B(a[47]), .Z(n4212) );
  NANDN U4304 ( .A(n10006), .B(n4212), .Z(n4136) );
  AND U4305 ( .A(n4137), .B(n4136), .Z(n4219) );
  NANDN U4306 ( .A(n9685), .B(n4138), .Z(n4140) );
  XOR U4307 ( .A(b[9]), .B(a[53]), .Z(n4215) );
  NANDN U4308 ( .A(n9758), .B(n4215), .Z(n4139) );
  NAND U4309 ( .A(n4140), .B(n4139), .Z(n4218) );
  XOR U4310 ( .A(n4219), .B(n4218), .Z(n4221) );
  XOR U4311 ( .A(n4220), .B(n4221), .Z(n4231) );
  NANDN U4312 ( .A(n4142), .B(n4141), .Z(n4146) );
  OR U4313 ( .A(n4144), .B(n4143), .Z(n4145) );
  AND U4314 ( .A(n4146), .B(n4145), .Z(n4230) );
  XNOR U4315 ( .A(n4231), .B(n4230), .Z(n4232) );
  NANDN U4316 ( .A(n4148), .B(n4147), .Z(n4152) );
  NANDN U4317 ( .A(n4150), .B(n4149), .Z(n4151) );
  NAND U4318 ( .A(n4152), .B(n4151), .Z(n4233) );
  XNOR U4319 ( .A(n4232), .B(n4233), .Z(n4178) );
  XOR U4320 ( .A(n4179), .B(n4178), .Z(n4237) );
  NANDN U4321 ( .A(n4154), .B(n4153), .Z(n4158) );
  NANDN U4322 ( .A(n4156), .B(n4155), .Z(n4157) );
  AND U4323 ( .A(n4158), .B(n4157), .Z(n4236) );
  XNOR U4324 ( .A(n4237), .B(n4236), .Z(n4238) );
  XOR U4325 ( .A(n4239), .B(n4238), .Z(n4171) );
  NANDN U4326 ( .A(n4160), .B(n4159), .Z(n4164) );
  NAND U4327 ( .A(n4162), .B(n4161), .Z(n4163) );
  AND U4328 ( .A(n4164), .B(n4163), .Z(n4170) );
  XNOR U4329 ( .A(n4171), .B(n4170), .Z(n4172) );
  XNOR U4330 ( .A(n4173), .B(n4172), .Z(n4242) );
  XNOR U4331 ( .A(sreg[173]), .B(n4242), .Z(n4244) );
  NANDN U4332 ( .A(sreg[172]), .B(n4165), .Z(n4169) );
  NAND U4333 ( .A(n4167), .B(n4166), .Z(n4168) );
  NAND U4334 ( .A(n4169), .B(n4168), .Z(n4243) );
  XNOR U4335 ( .A(n4244), .B(n4243), .Z(c[173]) );
  NANDN U4336 ( .A(n4171), .B(n4170), .Z(n4175) );
  NANDN U4337 ( .A(n4173), .B(n4172), .Z(n4174) );
  AND U4338 ( .A(n4175), .B(n4174), .Z(n4250) );
  NANDN U4339 ( .A(n4177), .B(n4176), .Z(n4181) );
  NAND U4340 ( .A(n4179), .B(n4178), .Z(n4180) );
  AND U4341 ( .A(n4181), .B(n4180), .Z(n4316) );
  NANDN U4342 ( .A(n4183), .B(n4182), .Z(n4187) );
  NANDN U4343 ( .A(n4185), .B(n4184), .Z(n4186) );
  AND U4344 ( .A(n4187), .B(n4186), .Z(n4282) );
  NAND U4345 ( .A(b[0]), .B(a[62]), .Z(n4188) );
  XNOR U4346 ( .A(b[1]), .B(n4188), .Z(n4190) );
  NANDN U4347 ( .A(b[0]), .B(a[61]), .Z(n4189) );
  NAND U4348 ( .A(n4190), .B(n4189), .Z(n4262) );
  NANDN U4349 ( .A(n9891), .B(n4191), .Z(n4193) );
  XOR U4350 ( .A(b[13]), .B(a[50]), .Z(n4265) );
  NANDN U4351 ( .A(n9935), .B(n4265), .Z(n4192) );
  AND U4352 ( .A(n4193), .B(n4192), .Z(n4260) );
  AND U4353 ( .A(b[15]), .B(a[46]), .Z(n4259) );
  XNOR U4354 ( .A(n4260), .B(n4259), .Z(n4261) );
  XNOR U4355 ( .A(n4262), .B(n4261), .Z(n4280) );
  NANDN U4356 ( .A(n9437), .B(n4194), .Z(n4196) );
  XOR U4357 ( .A(b[5]), .B(a[58]), .Z(n4271) );
  NANDN U4358 ( .A(n9503), .B(n4271), .Z(n4195) );
  AND U4359 ( .A(n4196), .B(n4195), .Z(n4304) );
  NANDN U4360 ( .A(n9588), .B(n4197), .Z(n4199) );
  XOR U4361 ( .A(b[7]), .B(a[56]), .Z(n4274) );
  NANDN U4362 ( .A(n9639), .B(n4274), .Z(n4198) );
  AND U4363 ( .A(n4199), .B(n4198), .Z(n4302) );
  NANDN U4364 ( .A(n9374), .B(n4200), .Z(n4202) );
  XOR U4365 ( .A(b[3]), .B(a[60]), .Z(n4277) );
  NANDN U4366 ( .A(n9375), .B(n4277), .Z(n4201) );
  NAND U4367 ( .A(n4202), .B(n4201), .Z(n4301) );
  XNOR U4368 ( .A(n4302), .B(n4301), .Z(n4303) );
  XOR U4369 ( .A(n4304), .B(n4303), .Z(n4281) );
  XOR U4370 ( .A(n4280), .B(n4281), .Z(n4283) );
  XOR U4371 ( .A(n4282), .B(n4283), .Z(n4254) );
  NANDN U4372 ( .A(n4204), .B(n4203), .Z(n4208) );
  OR U4373 ( .A(n4206), .B(n4205), .Z(n4207) );
  AND U4374 ( .A(n4208), .B(n4207), .Z(n4253) );
  XNOR U4375 ( .A(n4254), .B(n4253), .Z(n4256) );
  NAND U4376 ( .A(n4209), .B(n9883), .Z(n4211) );
  XOR U4377 ( .A(b[11]), .B(a[52]), .Z(n4286) );
  NANDN U4378 ( .A(n9856), .B(n4286), .Z(n4210) );
  AND U4379 ( .A(n4211), .B(n4210), .Z(n4297) );
  NANDN U4380 ( .A(n10005), .B(n4212), .Z(n4214) );
  XOR U4381 ( .A(b[15]), .B(a[48]), .Z(n4289) );
  NANDN U4382 ( .A(n10006), .B(n4289), .Z(n4213) );
  AND U4383 ( .A(n4214), .B(n4213), .Z(n4296) );
  NANDN U4384 ( .A(n9685), .B(n4215), .Z(n4217) );
  XOR U4385 ( .A(b[9]), .B(a[54]), .Z(n4292) );
  NANDN U4386 ( .A(n9758), .B(n4292), .Z(n4216) );
  NAND U4387 ( .A(n4217), .B(n4216), .Z(n4295) );
  XOR U4388 ( .A(n4296), .B(n4295), .Z(n4298) );
  XOR U4389 ( .A(n4297), .B(n4298), .Z(n4308) );
  NANDN U4390 ( .A(n4219), .B(n4218), .Z(n4223) );
  OR U4391 ( .A(n4221), .B(n4220), .Z(n4222) );
  AND U4392 ( .A(n4223), .B(n4222), .Z(n4307) );
  XNOR U4393 ( .A(n4308), .B(n4307), .Z(n4309) );
  NANDN U4394 ( .A(n4225), .B(n4224), .Z(n4229) );
  NANDN U4395 ( .A(n4227), .B(n4226), .Z(n4228) );
  NAND U4396 ( .A(n4229), .B(n4228), .Z(n4310) );
  XNOR U4397 ( .A(n4309), .B(n4310), .Z(n4255) );
  XOR U4398 ( .A(n4256), .B(n4255), .Z(n4314) );
  NANDN U4399 ( .A(n4231), .B(n4230), .Z(n4235) );
  NANDN U4400 ( .A(n4233), .B(n4232), .Z(n4234) );
  AND U4401 ( .A(n4235), .B(n4234), .Z(n4313) );
  XNOR U4402 ( .A(n4314), .B(n4313), .Z(n4315) );
  XOR U4403 ( .A(n4316), .B(n4315), .Z(n4248) );
  NANDN U4404 ( .A(n4237), .B(n4236), .Z(n4241) );
  NAND U4405 ( .A(n4239), .B(n4238), .Z(n4240) );
  AND U4406 ( .A(n4241), .B(n4240), .Z(n4247) );
  XNOR U4407 ( .A(n4248), .B(n4247), .Z(n4249) );
  XNOR U4408 ( .A(n4250), .B(n4249), .Z(n4319) );
  XNOR U4409 ( .A(sreg[174]), .B(n4319), .Z(n4321) );
  NANDN U4410 ( .A(sreg[173]), .B(n4242), .Z(n4246) );
  NAND U4411 ( .A(n4244), .B(n4243), .Z(n4245) );
  NAND U4412 ( .A(n4246), .B(n4245), .Z(n4320) );
  XNOR U4413 ( .A(n4321), .B(n4320), .Z(c[174]) );
  NANDN U4414 ( .A(n4248), .B(n4247), .Z(n4252) );
  NANDN U4415 ( .A(n4250), .B(n4249), .Z(n4251) );
  AND U4416 ( .A(n4252), .B(n4251), .Z(n4327) );
  NANDN U4417 ( .A(n4254), .B(n4253), .Z(n4258) );
  NAND U4418 ( .A(n4256), .B(n4255), .Z(n4257) );
  AND U4419 ( .A(n4258), .B(n4257), .Z(n4393) );
  NANDN U4420 ( .A(n4260), .B(n4259), .Z(n4264) );
  NANDN U4421 ( .A(n4262), .B(n4261), .Z(n4263) );
  AND U4422 ( .A(n4264), .B(n4263), .Z(n4380) );
  NANDN U4423 ( .A(n9891), .B(n4265), .Z(n4267) );
  XOR U4424 ( .A(b[13]), .B(a[51]), .Z(n4366) );
  NANDN U4425 ( .A(n9935), .B(n4366), .Z(n4266) );
  AND U4426 ( .A(n4267), .B(n4266), .Z(n4358) );
  AND U4427 ( .A(b[15]), .B(a[47]), .Z(n4357) );
  XNOR U4428 ( .A(n4358), .B(n4357), .Z(n4359) );
  NAND U4429 ( .A(b[0]), .B(a[63]), .Z(n4268) );
  XNOR U4430 ( .A(b[1]), .B(n4268), .Z(n4270) );
  NANDN U4431 ( .A(b[0]), .B(a[62]), .Z(n4269) );
  NAND U4432 ( .A(n4270), .B(n4269), .Z(n4360) );
  XNOR U4433 ( .A(n4359), .B(n4360), .Z(n4378) );
  NANDN U4434 ( .A(n9437), .B(n4271), .Z(n4273) );
  XOR U4435 ( .A(b[5]), .B(a[59]), .Z(n4369) );
  NANDN U4436 ( .A(n9503), .B(n4369), .Z(n4272) );
  AND U4437 ( .A(n4273), .B(n4272), .Z(n4354) );
  NANDN U4438 ( .A(n9588), .B(n4274), .Z(n4276) );
  XOR U4439 ( .A(b[7]), .B(a[57]), .Z(n4372) );
  NANDN U4440 ( .A(n9639), .B(n4372), .Z(n4275) );
  AND U4441 ( .A(n4276), .B(n4275), .Z(n4352) );
  NANDN U4442 ( .A(n9374), .B(n4277), .Z(n4279) );
  XOR U4443 ( .A(b[3]), .B(a[61]), .Z(n4375) );
  NANDN U4444 ( .A(n9375), .B(n4375), .Z(n4278) );
  NAND U4445 ( .A(n4279), .B(n4278), .Z(n4351) );
  XNOR U4446 ( .A(n4352), .B(n4351), .Z(n4353) );
  XOR U4447 ( .A(n4354), .B(n4353), .Z(n4379) );
  XOR U4448 ( .A(n4378), .B(n4379), .Z(n4381) );
  XOR U4449 ( .A(n4380), .B(n4381), .Z(n4331) );
  NANDN U4450 ( .A(n4281), .B(n4280), .Z(n4285) );
  OR U4451 ( .A(n4283), .B(n4282), .Z(n4284) );
  AND U4452 ( .A(n4285), .B(n4284), .Z(n4330) );
  XNOR U4453 ( .A(n4331), .B(n4330), .Z(n4333) );
  NAND U4454 ( .A(n4286), .B(n9883), .Z(n4288) );
  XOR U4455 ( .A(b[11]), .B(a[53]), .Z(n4336) );
  NANDN U4456 ( .A(n9856), .B(n4336), .Z(n4287) );
  AND U4457 ( .A(n4288), .B(n4287), .Z(n4347) );
  NANDN U4458 ( .A(n10005), .B(n4289), .Z(n4291) );
  XOR U4459 ( .A(b[15]), .B(a[49]), .Z(n4339) );
  NANDN U4460 ( .A(n10006), .B(n4339), .Z(n4290) );
  AND U4461 ( .A(n4291), .B(n4290), .Z(n4346) );
  NANDN U4462 ( .A(n9685), .B(n4292), .Z(n4294) );
  XOR U4463 ( .A(b[9]), .B(a[55]), .Z(n4342) );
  NANDN U4464 ( .A(n9758), .B(n4342), .Z(n4293) );
  NAND U4465 ( .A(n4294), .B(n4293), .Z(n4345) );
  XOR U4466 ( .A(n4346), .B(n4345), .Z(n4348) );
  XOR U4467 ( .A(n4347), .B(n4348), .Z(n4385) );
  NANDN U4468 ( .A(n4296), .B(n4295), .Z(n4300) );
  OR U4469 ( .A(n4298), .B(n4297), .Z(n4299) );
  AND U4470 ( .A(n4300), .B(n4299), .Z(n4384) );
  XNOR U4471 ( .A(n4385), .B(n4384), .Z(n4386) );
  NANDN U4472 ( .A(n4302), .B(n4301), .Z(n4306) );
  NANDN U4473 ( .A(n4304), .B(n4303), .Z(n4305) );
  NAND U4474 ( .A(n4306), .B(n4305), .Z(n4387) );
  XNOR U4475 ( .A(n4386), .B(n4387), .Z(n4332) );
  XOR U4476 ( .A(n4333), .B(n4332), .Z(n4391) );
  NANDN U4477 ( .A(n4308), .B(n4307), .Z(n4312) );
  NANDN U4478 ( .A(n4310), .B(n4309), .Z(n4311) );
  AND U4479 ( .A(n4312), .B(n4311), .Z(n4390) );
  XNOR U4480 ( .A(n4391), .B(n4390), .Z(n4392) );
  XOR U4481 ( .A(n4393), .B(n4392), .Z(n4325) );
  NANDN U4482 ( .A(n4314), .B(n4313), .Z(n4318) );
  NAND U4483 ( .A(n4316), .B(n4315), .Z(n4317) );
  AND U4484 ( .A(n4318), .B(n4317), .Z(n4324) );
  XNOR U4485 ( .A(n4325), .B(n4324), .Z(n4326) );
  XNOR U4486 ( .A(n4327), .B(n4326), .Z(n4396) );
  XNOR U4487 ( .A(sreg[175]), .B(n4396), .Z(n4398) );
  NANDN U4488 ( .A(sreg[174]), .B(n4319), .Z(n4323) );
  NAND U4489 ( .A(n4321), .B(n4320), .Z(n4322) );
  NAND U4490 ( .A(n4323), .B(n4322), .Z(n4397) );
  XNOR U4491 ( .A(n4398), .B(n4397), .Z(c[175]) );
  NANDN U4492 ( .A(n4325), .B(n4324), .Z(n4329) );
  NANDN U4493 ( .A(n4327), .B(n4326), .Z(n4328) );
  AND U4494 ( .A(n4329), .B(n4328), .Z(n4404) );
  NANDN U4495 ( .A(n4331), .B(n4330), .Z(n4335) );
  NAND U4496 ( .A(n4333), .B(n4332), .Z(n4334) );
  AND U4497 ( .A(n4335), .B(n4334), .Z(n4470) );
  NAND U4498 ( .A(n4336), .B(n9883), .Z(n4338) );
  XOR U4499 ( .A(b[11]), .B(a[54]), .Z(n4440) );
  NANDN U4500 ( .A(n9856), .B(n4440), .Z(n4337) );
  AND U4501 ( .A(n4338), .B(n4337), .Z(n4451) );
  NANDN U4502 ( .A(n10005), .B(n4339), .Z(n4341) );
  XOR U4503 ( .A(b[15]), .B(a[50]), .Z(n4443) );
  NANDN U4504 ( .A(n10006), .B(n4443), .Z(n4340) );
  AND U4505 ( .A(n4341), .B(n4340), .Z(n4450) );
  NANDN U4506 ( .A(n9685), .B(n4342), .Z(n4344) );
  XOR U4507 ( .A(b[9]), .B(a[56]), .Z(n4446) );
  NANDN U4508 ( .A(n9758), .B(n4446), .Z(n4343) );
  NAND U4509 ( .A(n4344), .B(n4343), .Z(n4449) );
  XOR U4510 ( .A(n4450), .B(n4449), .Z(n4452) );
  XOR U4511 ( .A(n4451), .B(n4452), .Z(n4462) );
  NANDN U4512 ( .A(n4346), .B(n4345), .Z(n4350) );
  OR U4513 ( .A(n4348), .B(n4347), .Z(n4349) );
  AND U4514 ( .A(n4350), .B(n4349), .Z(n4461) );
  XNOR U4515 ( .A(n4462), .B(n4461), .Z(n4463) );
  NANDN U4516 ( .A(n4352), .B(n4351), .Z(n4356) );
  NANDN U4517 ( .A(n4354), .B(n4353), .Z(n4355) );
  NAND U4518 ( .A(n4356), .B(n4355), .Z(n4464) );
  XNOR U4519 ( .A(n4463), .B(n4464), .Z(n4410) );
  NANDN U4520 ( .A(n4358), .B(n4357), .Z(n4362) );
  NANDN U4521 ( .A(n4360), .B(n4359), .Z(n4361) );
  AND U4522 ( .A(n4362), .B(n4361), .Z(n4436) );
  NAND U4523 ( .A(b[0]), .B(a[64]), .Z(n4363) );
  XNOR U4524 ( .A(b[1]), .B(n4363), .Z(n4365) );
  NANDN U4525 ( .A(b[0]), .B(a[63]), .Z(n4364) );
  NAND U4526 ( .A(n4365), .B(n4364), .Z(n4416) );
  NANDN U4527 ( .A(n9891), .B(n4366), .Z(n4368) );
  XOR U4528 ( .A(b[13]), .B(a[52]), .Z(n4422) );
  NANDN U4529 ( .A(n9935), .B(n4422), .Z(n4367) );
  AND U4530 ( .A(n4368), .B(n4367), .Z(n4414) );
  AND U4531 ( .A(b[15]), .B(a[48]), .Z(n4413) );
  XNOR U4532 ( .A(n4414), .B(n4413), .Z(n4415) );
  XNOR U4533 ( .A(n4416), .B(n4415), .Z(n4434) );
  NANDN U4534 ( .A(n9437), .B(n4369), .Z(n4371) );
  XOR U4535 ( .A(b[5]), .B(a[60]), .Z(n4425) );
  NANDN U4536 ( .A(n9503), .B(n4425), .Z(n4370) );
  AND U4537 ( .A(n4371), .B(n4370), .Z(n4458) );
  NANDN U4538 ( .A(n9588), .B(n4372), .Z(n4374) );
  XOR U4539 ( .A(b[7]), .B(a[58]), .Z(n4428) );
  NANDN U4540 ( .A(n9639), .B(n4428), .Z(n4373) );
  AND U4541 ( .A(n4374), .B(n4373), .Z(n4456) );
  NANDN U4542 ( .A(n9374), .B(n4375), .Z(n4377) );
  XOR U4543 ( .A(b[3]), .B(a[62]), .Z(n4431) );
  NANDN U4544 ( .A(n9375), .B(n4431), .Z(n4376) );
  NAND U4545 ( .A(n4377), .B(n4376), .Z(n4455) );
  XNOR U4546 ( .A(n4456), .B(n4455), .Z(n4457) );
  XOR U4547 ( .A(n4458), .B(n4457), .Z(n4435) );
  XOR U4548 ( .A(n4434), .B(n4435), .Z(n4437) );
  XOR U4549 ( .A(n4436), .B(n4437), .Z(n4408) );
  NANDN U4550 ( .A(n4379), .B(n4378), .Z(n4383) );
  OR U4551 ( .A(n4381), .B(n4380), .Z(n4382) );
  AND U4552 ( .A(n4383), .B(n4382), .Z(n4407) );
  XNOR U4553 ( .A(n4408), .B(n4407), .Z(n4409) );
  XOR U4554 ( .A(n4410), .B(n4409), .Z(n4468) );
  NANDN U4555 ( .A(n4385), .B(n4384), .Z(n4389) );
  NANDN U4556 ( .A(n4387), .B(n4386), .Z(n4388) );
  AND U4557 ( .A(n4389), .B(n4388), .Z(n4467) );
  XNOR U4558 ( .A(n4468), .B(n4467), .Z(n4469) );
  XOR U4559 ( .A(n4470), .B(n4469), .Z(n4402) );
  NANDN U4560 ( .A(n4391), .B(n4390), .Z(n4395) );
  NAND U4561 ( .A(n4393), .B(n4392), .Z(n4394) );
  AND U4562 ( .A(n4395), .B(n4394), .Z(n4401) );
  XNOR U4563 ( .A(n4402), .B(n4401), .Z(n4403) );
  XNOR U4564 ( .A(n4404), .B(n4403), .Z(n4473) );
  XNOR U4565 ( .A(sreg[176]), .B(n4473), .Z(n4475) );
  NANDN U4566 ( .A(sreg[175]), .B(n4396), .Z(n4400) );
  NAND U4567 ( .A(n4398), .B(n4397), .Z(n4399) );
  NAND U4568 ( .A(n4400), .B(n4399), .Z(n4474) );
  XNOR U4569 ( .A(n4475), .B(n4474), .Z(c[176]) );
  NANDN U4570 ( .A(n4402), .B(n4401), .Z(n4406) );
  NANDN U4571 ( .A(n4404), .B(n4403), .Z(n4405) );
  AND U4572 ( .A(n4406), .B(n4405), .Z(n4481) );
  NANDN U4573 ( .A(n4408), .B(n4407), .Z(n4412) );
  NAND U4574 ( .A(n4410), .B(n4409), .Z(n4411) );
  AND U4575 ( .A(n4412), .B(n4411), .Z(n4547) );
  NANDN U4576 ( .A(n4414), .B(n4413), .Z(n4418) );
  NANDN U4577 ( .A(n4416), .B(n4415), .Z(n4417) );
  AND U4578 ( .A(n4418), .B(n4417), .Z(n4513) );
  AND U4579 ( .A(b[0]), .B(a[65]), .Z(n4419) );
  XOR U4580 ( .A(b[1]), .B(n4419), .Z(n4421) );
  NANDN U4581 ( .A(b[0]), .B(a[64]), .Z(n4420) );
  AND U4582 ( .A(n4421), .B(n4420), .Z(n4492) );
  NANDN U4583 ( .A(n9891), .B(n4422), .Z(n4424) );
  XOR U4584 ( .A(b[13]), .B(a[53]), .Z(n4499) );
  NANDN U4585 ( .A(n9935), .B(n4499), .Z(n4423) );
  AND U4586 ( .A(n4424), .B(n4423), .Z(n4491) );
  AND U4587 ( .A(b[15]), .B(a[49]), .Z(n4490) );
  XOR U4588 ( .A(n4491), .B(n4490), .Z(n4493) );
  XNOR U4589 ( .A(n4492), .B(n4493), .Z(n4511) );
  NANDN U4590 ( .A(n9437), .B(n4425), .Z(n4427) );
  XOR U4591 ( .A(b[5]), .B(a[61]), .Z(n4502) );
  NANDN U4592 ( .A(n9503), .B(n4502), .Z(n4426) );
  AND U4593 ( .A(n4427), .B(n4426), .Z(n4535) );
  NANDN U4594 ( .A(n9588), .B(n4428), .Z(n4430) );
  XOR U4595 ( .A(b[7]), .B(a[59]), .Z(n4505) );
  NANDN U4596 ( .A(n9639), .B(n4505), .Z(n4429) );
  AND U4597 ( .A(n4430), .B(n4429), .Z(n4533) );
  NANDN U4598 ( .A(n9374), .B(n4431), .Z(n4433) );
  XOR U4599 ( .A(b[3]), .B(a[63]), .Z(n4508) );
  NANDN U4600 ( .A(n9375), .B(n4508), .Z(n4432) );
  NAND U4601 ( .A(n4433), .B(n4432), .Z(n4532) );
  XNOR U4602 ( .A(n4533), .B(n4532), .Z(n4534) );
  XOR U4603 ( .A(n4535), .B(n4534), .Z(n4512) );
  XOR U4604 ( .A(n4511), .B(n4512), .Z(n4514) );
  XOR U4605 ( .A(n4513), .B(n4514), .Z(n4485) );
  NANDN U4606 ( .A(n4435), .B(n4434), .Z(n4439) );
  OR U4607 ( .A(n4437), .B(n4436), .Z(n4438) );
  AND U4608 ( .A(n4439), .B(n4438), .Z(n4484) );
  XNOR U4609 ( .A(n4485), .B(n4484), .Z(n4487) );
  NAND U4610 ( .A(n4440), .B(n9883), .Z(n4442) );
  XOR U4611 ( .A(b[11]), .B(a[55]), .Z(n4517) );
  NANDN U4612 ( .A(n9856), .B(n4517), .Z(n4441) );
  AND U4613 ( .A(n4442), .B(n4441), .Z(n4528) );
  NANDN U4614 ( .A(n10005), .B(n4443), .Z(n4445) );
  XOR U4615 ( .A(b[15]), .B(a[51]), .Z(n4520) );
  NANDN U4616 ( .A(n10006), .B(n4520), .Z(n4444) );
  AND U4617 ( .A(n4445), .B(n4444), .Z(n4527) );
  NANDN U4618 ( .A(n9685), .B(n4446), .Z(n4448) );
  XOR U4619 ( .A(b[9]), .B(a[57]), .Z(n4523) );
  NANDN U4620 ( .A(n9758), .B(n4523), .Z(n4447) );
  NAND U4621 ( .A(n4448), .B(n4447), .Z(n4526) );
  XOR U4622 ( .A(n4527), .B(n4526), .Z(n4529) );
  XOR U4623 ( .A(n4528), .B(n4529), .Z(n4539) );
  NANDN U4624 ( .A(n4450), .B(n4449), .Z(n4454) );
  OR U4625 ( .A(n4452), .B(n4451), .Z(n4453) );
  AND U4626 ( .A(n4454), .B(n4453), .Z(n4538) );
  XNOR U4627 ( .A(n4539), .B(n4538), .Z(n4540) );
  NANDN U4628 ( .A(n4456), .B(n4455), .Z(n4460) );
  NANDN U4629 ( .A(n4458), .B(n4457), .Z(n4459) );
  NAND U4630 ( .A(n4460), .B(n4459), .Z(n4541) );
  XNOR U4631 ( .A(n4540), .B(n4541), .Z(n4486) );
  XOR U4632 ( .A(n4487), .B(n4486), .Z(n4545) );
  NANDN U4633 ( .A(n4462), .B(n4461), .Z(n4466) );
  NANDN U4634 ( .A(n4464), .B(n4463), .Z(n4465) );
  AND U4635 ( .A(n4466), .B(n4465), .Z(n4544) );
  XNOR U4636 ( .A(n4545), .B(n4544), .Z(n4546) );
  XOR U4637 ( .A(n4547), .B(n4546), .Z(n4479) );
  NANDN U4638 ( .A(n4468), .B(n4467), .Z(n4472) );
  NAND U4639 ( .A(n4470), .B(n4469), .Z(n4471) );
  AND U4640 ( .A(n4472), .B(n4471), .Z(n4478) );
  XNOR U4641 ( .A(n4479), .B(n4478), .Z(n4480) );
  XNOR U4642 ( .A(n4481), .B(n4480), .Z(n4550) );
  XNOR U4643 ( .A(sreg[177]), .B(n4550), .Z(n4552) );
  NANDN U4644 ( .A(sreg[176]), .B(n4473), .Z(n4477) );
  NAND U4645 ( .A(n4475), .B(n4474), .Z(n4476) );
  NAND U4646 ( .A(n4477), .B(n4476), .Z(n4551) );
  XNOR U4647 ( .A(n4552), .B(n4551), .Z(c[177]) );
  NANDN U4648 ( .A(n4479), .B(n4478), .Z(n4483) );
  NANDN U4649 ( .A(n4481), .B(n4480), .Z(n4482) );
  AND U4650 ( .A(n4483), .B(n4482), .Z(n4558) );
  NANDN U4651 ( .A(n4485), .B(n4484), .Z(n4489) );
  NAND U4652 ( .A(n4487), .B(n4486), .Z(n4488) );
  AND U4653 ( .A(n4489), .B(n4488), .Z(n4624) );
  NANDN U4654 ( .A(n4491), .B(n4490), .Z(n4495) );
  NANDN U4655 ( .A(n4493), .B(n4492), .Z(n4494) );
  AND U4656 ( .A(n4495), .B(n4494), .Z(n4590) );
  NAND U4657 ( .A(b[0]), .B(a[66]), .Z(n4496) );
  XNOR U4658 ( .A(b[1]), .B(n4496), .Z(n4498) );
  NANDN U4659 ( .A(b[0]), .B(a[65]), .Z(n4497) );
  NAND U4660 ( .A(n4498), .B(n4497), .Z(n4570) );
  NANDN U4661 ( .A(n9891), .B(n4499), .Z(n4501) );
  XOR U4662 ( .A(b[13]), .B(a[54]), .Z(n4573) );
  NANDN U4663 ( .A(n9935), .B(n4573), .Z(n4500) );
  AND U4664 ( .A(n4501), .B(n4500), .Z(n4568) );
  AND U4665 ( .A(b[15]), .B(a[50]), .Z(n4567) );
  XNOR U4666 ( .A(n4568), .B(n4567), .Z(n4569) );
  XNOR U4667 ( .A(n4570), .B(n4569), .Z(n4588) );
  NANDN U4668 ( .A(n9437), .B(n4502), .Z(n4504) );
  XOR U4669 ( .A(b[5]), .B(a[62]), .Z(n4579) );
  NANDN U4670 ( .A(n9503), .B(n4579), .Z(n4503) );
  AND U4671 ( .A(n4504), .B(n4503), .Z(n4612) );
  NANDN U4672 ( .A(n9588), .B(n4505), .Z(n4507) );
  XOR U4673 ( .A(b[7]), .B(a[60]), .Z(n4582) );
  NANDN U4674 ( .A(n9639), .B(n4582), .Z(n4506) );
  AND U4675 ( .A(n4507), .B(n4506), .Z(n4610) );
  NANDN U4676 ( .A(n9374), .B(n4508), .Z(n4510) );
  XOR U4677 ( .A(b[3]), .B(a[64]), .Z(n4585) );
  NANDN U4678 ( .A(n9375), .B(n4585), .Z(n4509) );
  NAND U4679 ( .A(n4510), .B(n4509), .Z(n4609) );
  XNOR U4680 ( .A(n4610), .B(n4609), .Z(n4611) );
  XOR U4681 ( .A(n4612), .B(n4611), .Z(n4589) );
  XOR U4682 ( .A(n4588), .B(n4589), .Z(n4591) );
  XOR U4683 ( .A(n4590), .B(n4591), .Z(n4562) );
  NANDN U4684 ( .A(n4512), .B(n4511), .Z(n4516) );
  OR U4685 ( .A(n4514), .B(n4513), .Z(n4515) );
  AND U4686 ( .A(n4516), .B(n4515), .Z(n4561) );
  XNOR U4687 ( .A(n4562), .B(n4561), .Z(n4564) );
  NAND U4688 ( .A(n4517), .B(n9883), .Z(n4519) );
  XOR U4689 ( .A(b[11]), .B(a[56]), .Z(n4594) );
  NANDN U4690 ( .A(n9856), .B(n4594), .Z(n4518) );
  AND U4691 ( .A(n4519), .B(n4518), .Z(n4605) );
  NANDN U4692 ( .A(n10005), .B(n4520), .Z(n4522) );
  XOR U4693 ( .A(b[15]), .B(a[52]), .Z(n4597) );
  NANDN U4694 ( .A(n10006), .B(n4597), .Z(n4521) );
  AND U4695 ( .A(n4522), .B(n4521), .Z(n4604) );
  NANDN U4696 ( .A(n9685), .B(n4523), .Z(n4525) );
  XOR U4697 ( .A(b[9]), .B(a[58]), .Z(n4600) );
  NANDN U4698 ( .A(n9758), .B(n4600), .Z(n4524) );
  NAND U4699 ( .A(n4525), .B(n4524), .Z(n4603) );
  XOR U4700 ( .A(n4604), .B(n4603), .Z(n4606) );
  XOR U4701 ( .A(n4605), .B(n4606), .Z(n4616) );
  NANDN U4702 ( .A(n4527), .B(n4526), .Z(n4531) );
  OR U4703 ( .A(n4529), .B(n4528), .Z(n4530) );
  AND U4704 ( .A(n4531), .B(n4530), .Z(n4615) );
  XNOR U4705 ( .A(n4616), .B(n4615), .Z(n4617) );
  NANDN U4706 ( .A(n4533), .B(n4532), .Z(n4537) );
  NANDN U4707 ( .A(n4535), .B(n4534), .Z(n4536) );
  NAND U4708 ( .A(n4537), .B(n4536), .Z(n4618) );
  XNOR U4709 ( .A(n4617), .B(n4618), .Z(n4563) );
  XOR U4710 ( .A(n4564), .B(n4563), .Z(n4622) );
  NANDN U4711 ( .A(n4539), .B(n4538), .Z(n4543) );
  NANDN U4712 ( .A(n4541), .B(n4540), .Z(n4542) );
  AND U4713 ( .A(n4543), .B(n4542), .Z(n4621) );
  XNOR U4714 ( .A(n4622), .B(n4621), .Z(n4623) );
  XOR U4715 ( .A(n4624), .B(n4623), .Z(n4556) );
  NANDN U4716 ( .A(n4545), .B(n4544), .Z(n4549) );
  NAND U4717 ( .A(n4547), .B(n4546), .Z(n4548) );
  AND U4718 ( .A(n4549), .B(n4548), .Z(n4555) );
  XNOR U4719 ( .A(n4556), .B(n4555), .Z(n4557) );
  XNOR U4720 ( .A(n4558), .B(n4557), .Z(n4627) );
  XNOR U4721 ( .A(sreg[178]), .B(n4627), .Z(n4629) );
  NANDN U4722 ( .A(sreg[177]), .B(n4550), .Z(n4554) );
  NAND U4723 ( .A(n4552), .B(n4551), .Z(n4553) );
  NAND U4724 ( .A(n4554), .B(n4553), .Z(n4628) );
  XNOR U4725 ( .A(n4629), .B(n4628), .Z(c[178]) );
  NANDN U4726 ( .A(n4556), .B(n4555), .Z(n4560) );
  NANDN U4727 ( .A(n4558), .B(n4557), .Z(n4559) );
  AND U4728 ( .A(n4560), .B(n4559), .Z(n4635) );
  NANDN U4729 ( .A(n4562), .B(n4561), .Z(n4566) );
  NAND U4730 ( .A(n4564), .B(n4563), .Z(n4565) );
  AND U4731 ( .A(n4566), .B(n4565), .Z(n4701) );
  NANDN U4732 ( .A(n4568), .B(n4567), .Z(n4572) );
  NANDN U4733 ( .A(n4570), .B(n4569), .Z(n4571) );
  AND U4734 ( .A(n4572), .B(n4571), .Z(n4667) );
  NANDN U4735 ( .A(n9891), .B(n4573), .Z(n4575) );
  XOR U4736 ( .A(b[13]), .B(a[55]), .Z(n4653) );
  NANDN U4737 ( .A(n9935), .B(n4653), .Z(n4574) );
  AND U4738 ( .A(n4575), .B(n4574), .Z(n4645) );
  AND U4739 ( .A(b[15]), .B(a[51]), .Z(n4644) );
  XNOR U4740 ( .A(n4645), .B(n4644), .Z(n4646) );
  NAND U4741 ( .A(b[0]), .B(a[67]), .Z(n4576) );
  XNOR U4742 ( .A(b[1]), .B(n4576), .Z(n4578) );
  NANDN U4743 ( .A(b[0]), .B(a[66]), .Z(n4577) );
  NAND U4744 ( .A(n4578), .B(n4577), .Z(n4647) );
  XNOR U4745 ( .A(n4646), .B(n4647), .Z(n4665) );
  NANDN U4746 ( .A(n9437), .B(n4579), .Z(n4581) );
  XOR U4747 ( .A(b[5]), .B(a[63]), .Z(n4656) );
  NANDN U4748 ( .A(n9503), .B(n4656), .Z(n4580) );
  AND U4749 ( .A(n4581), .B(n4580), .Z(n4689) );
  NANDN U4750 ( .A(n9588), .B(n4582), .Z(n4584) );
  XOR U4751 ( .A(b[7]), .B(a[61]), .Z(n4659) );
  NANDN U4752 ( .A(n9639), .B(n4659), .Z(n4583) );
  AND U4753 ( .A(n4584), .B(n4583), .Z(n4687) );
  NANDN U4754 ( .A(n9374), .B(n4585), .Z(n4587) );
  XOR U4755 ( .A(b[3]), .B(a[65]), .Z(n4662) );
  NANDN U4756 ( .A(n9375), .B(n4662), .Z(n4586) );
  NAND U4757 ( .A(n4587), .B(n4586), .Z(n4686) );
  XNOR U4758 ( .A(n4687), .B(n4686), .Z(n4688) );
  XOR U4759 ( .A(n4689), .B(n4688), .Z(n4666) );
  XOR U4760 ( .A(n4665), .B(n4666), .Z(n4668) );
  XOR U4761 ( .A(n4667), .B(n4668), .Z(n4639) );
  NANDN U4762 ( .A(n4589), .B(n4588), .Z(n4593) );
  OR U4763 ( .A(n4591), .B(n4590), .Z(n4592) );
  AND U4764 ( .A(n4593), .B(n4592), .Z(n4638) );
  XNOR U4765 ( .A(n4639), .B(n4638), .Z(n4641) );
  NAND U4766 ( .A(n4594), .B(n9883), .Z(n4596) );
  XOR U4767 ( .A(b[11]), .B(a[57]), .Z(n4671) );
  NANDN U4768 ( .A(n9856), .B(n4671), .Z(n4595) );
  AND U4769 ( .A(n4596), .B(n4595), .Z(n4682) );
  NANDN U4770 ( .A(n10005), .B(n4597), .Z(n4599) );
  XOR U4771 ( .A(b[15]), .B(a[53]), .Z(n4674) );
  NANDN U4772 ( .A(n10006), .B(n4674), .Z(n4598) );
  AND U4773 ( .A(n4599), .B(n4598), .Z(n4681) );
  NANDN U4774 ( .A(n9685), .B(n4600), .Z(n4602) );
  XOR U4775 ( .A(b[9]), .B(a[59]), .Z(n4677) );
  NANDN U4776 ( .A(n9758), .B(n4677), .Z(n4601) );
  NAND U4777 ( .A(n4602), .B(n4601), .Z(n4680) );
  XOR U4778 ( .A(n4681), .B(n4680), .Z(n4683) );
  XOR U4779 ( .A(n4682), .B(n4683), .Z(n4693) );
  NANDN U4780 ( .A(n4604), .B(n4603), .Z(n4608) );
  OR U4781 ( .A(n4606), .B(n4605), .Z(n4607) );
  AND U4782 ( .A(n4608), .B(n4607), .Z(n4692) );
  XNOR U4783 ( .A(n4693), .B(n4692), .Z(n4694) );
  NANDN U4784 ( .A(n4610), .B(n4609), .Z(n4614) );
  NANDN U4785 ( .A(n4612), .B(n4611), .Z(n4613) );
  NAND U4786 ( .A(n4614), .B(n4613), .Z(n4695) );
  XNOR U4787 ( .A(n4694), .B(n4695), .Z(n4640) );
  XOR U4788 ( .A(n4641), .B(n4640), .Z(n4699) );
  NANDN U4789 ( .A(n4616), .B(n4615), .Z(n4620) );
  NANDN U4790 ( .A(n4618), .B(n4617), .Z(n4619) );
  AND U4791 ( .A(n4620), .B(n4619), .Z(n4698) );
  XNOR U4792 ( .A(n4699), .B(n4698), .Z(n4700) );
  XOR U4793 ( .A(n4701), .B(n4700), .Z(n4633) );
  NANDN U4794 ( .A(n4622), .B(n4621), .Z(n4626) );
  NAND U4795 ( .A(n4624), .B(n4623), .Z(n4625) );
  AND U4796 ( .A(n4626), .B(n4625), .Z(n4632) );
  XNOR U4797 ( .A(n4633), .B(n4632), .Z(n4634) );
  XNOR U4798 ( .A(n4635), .B(n4634), .Z(n4704) );
  XNOR U4799 ( .A(sreg[179]), .B(n4704), .Z(n4706) );
  NANDN U4800 ( .A(sreg[178]), .B(n4627), .Z(n4631) );
  NAND U4801 ( .A(n4629), .B(n4628), .Z(n4630) );
  NAND U4802 ( .A(n4631), .B(n4630), .Z(n4705) );
  XNOR U4803 ( .A(n4706), .B(n4705), .Z(c[179]) );
  NANDN U4804 ( .A(n4633), .B(n4632), .Z(n4637) );
  NANDN U4805 ( .A(n4635), .B(n4634), .Z(n4636) );
  AND U4806 ( .A(n4637), .B(n4636), .Z(n4712) );
  NANDN U4807 ( .A(n4639), .B(n4638), .Z(n4643) );
  NAND U4808 ( .A(n4641), .B(n4640), .Z(n4642) );
  AND U4809 ( .A(n4643), .B(n4642), .Z(n4778) );
  NANDN U4810 ( .A(n4645), .B(n4644), .Z(n4649) );
  NANDN U4811 ( .A(n4647), .B(n4646), .Z(n4648) );
  AND U4812 ( .A(n4649), .B(n4648), .Z(n4744) );
  NAND U4813 ( .A(b[0]), .B(a[68]), .Z(n4650) );
  XNOR U4814 ( .A(b[1]), .B(n4650), .Z(n4652) );
  NANDN U4815 ( .A(b[0]), .B(a[67]), .Z(n4651) );
  NAND U4816 ( .A(n4652), .B(n4651), .Z(n4724) );
  NANDN U4817 ( .A(n9891), .B(n4653), .Z(n4655) );
  XOR U4818 ( .A(b[13]), .B(a[56]), .Z(n4730) );
  NANDN U4819 ( .A(n9935), .B(n4730), .Z(n4654) );
  AND U4820 ( .A(n4655), .B(n4654), .Z(n4722) );
  AND U4821 ( .A(b[15]), .B(a[52]), .Z(n4721) );
  XNOR U4822 ( .A(n4722), .B(n4721), .Z(n4723) );
  XNOR U4823 ( .A(n4724), .B(n4723), .Z(n4742) );
  NANDN U4824 ( .A(n9437), .B(n4656), .Z(n4658) );
  XOR U4825 ( .A(b[5]), .B(a[64]), .Z(n4733) );
  NANDN U4826 ( .A(n9503), .B(n4733), .Z(n4657) );
  AND U4827 ( .A(n4658), .B(n4657), .Z(n4766) );
  NANDN U4828 ( .A(n9588), .B(n4659), .Z(n4661) );
  XOR U4829 ( .A(b[7]), .B(a[62]), .Z(n4736) );
  NANDN U4830 ( .A(n9639), .B(n4736), .Z(n4660) );
  AND U4831 ( .A(n4661), .B(n4660), .Z(n4764) );
  NANDN U4832 ( .A(n9374), .B(n4662), .Z(n4664) );
  XOR U4833 ( .A(b[3]), .B(a[66]), .Z(n4739) );
  NANDN U4834 ( .A(n9375), .B(n4739), .Z(n4663) );
  NAND U4835 ( .A(n4664), .B(n4663), .Z(n4763) );
  XNOR U4836 ( .A(n4764), .B(n4763), .Z(n4765) );
  XOR U4837 ( .A(n4766), .B(n4765), .Z(n4743) );
  XOR U4838 ( .A(n4742), .B(n4743), .Z(n4745) );
  XOR U4839 ( .A(n4744), .B(n4745), .Z(n4716) );
  NANDN U4840 ( .A(n4666), .B(n4665), .Z(n4670) );
  OR U4841 ( .A(n4668), .B(n4667), .Z(n4669) );
  AND U4842 ( .A(n4670), .B(n4669), .Z(n4715) );
  XNOR U4843 ( .A(n4716), .B(n4715), .Z(n4718) );
  NAND U4844 ( .A(n4671), .B(n9883), .Z(n4673) );
  XOR U4845 ( .A(b[11]), .B(a[58]), .Z(n4748) );
  NANDN U4846 ( .A(n9856), .B(n4748), .Z(n4672) );
  AND U4847 ( .A(n4673), .B(n4672), .Z(n4759) );
  NANDN U4848 ( .A(n10005), .B(n4674), .Z(n4676) );
  XOR U4849 ( .A(b[15]), .B(a[54]), .Z(n4751) );
  NANDN U4850 ( .A(n10006), .B(n4751), .Z(n4675) );
  AND U4851 ( .A(n4676), .B(n4675), .Z(n4758) );
  NANDN U4852 ( .A(n9685), .B(n4677), .Z(n4679) );
  XOR U4853 ( .A(b[9]), .B(a[60]), .Z(n4754) );
  NANDN U4854 ( .A(n9758), .B(n4754), .Z(n4678) );
  NAND U4855 ( .A(n4679), .B(n4678), .Z(n4757) );
  XOR U4856 ( .A(n4758), .B(n4757), .Z(n4760) );
  XOR U4857 ( .A(n4759), .B(n4760), .Z(n4770) );
  NANDN U4858 ( .A(n4681), .B(n4680), .Z(n4685) );
  OR U4859 ( .A(n4683), .B(n4682), .Z(n4684) );
  AND U4860 ( .A(n4685), .B(n4684), .Z(n4769) );
  XNOR U4861 ( .A(n4770), .B(n4769), .Z(n4771) );
  NANDN U4862 ( .A(n4687), .B(n4686), .Z(n4691) );
  NANDN U4863 ( .A(n4689), .B(n4688), .Z(n4690) );
  NAND U4864 ( .A(n4691), .B(n4690), .Z(n4772) );
  XNOR U4865 ( .A(n4771), .B(n4772), .Z(n4717) );
  XOR U4866 ( .A(n4718), .B(n4717), .Z(n4776) );
  NANDN U4867 ( .A(n4693), .B(n4692), .Z(n4697) );
  NANDN U4868 ( .A(n4695), .B(n4694), .Z(n4696) );
  AND U4869 ( .A(n4697), .B(n4696), .Z(n4775) );
  XNOR U4870 ( .A(n4776), .B(n4775), .Z(n4777) );
  XOR U4871 ( .A(n4778), .B(n4777), .Z(n4710) );
  NANDN U4872 ( .A(n4699), .B(n4698), .Z(n4703) );
  NAND U4873 ( .A(n4701), .B(n4700), .Z(n4702) );
  AND U4874 ( .A(n4703), .B(n4702), .Z(n4709) );
  XNOR U4875 ( .A(n4710), .B(n4709), .Z(n4711) );
  XNOR U4876 ( .A(n4712), .B(n4711), .Z(n4781) );
  XNOR U4877 ( .A(sreg[180]), .B(n4781), .Z(n4783) );
  NANDN U4878 ( .A(sreg[179]), .B(n4704), .Z(n4708) );
  NAND U4879 ( .A(n4706), .B(n4705), .Z(n4707) );
  NAND U4880 ( .A(n4708), .B(n4707), .Z(n4782) );
  XNOR U4881 ( .A(n4783), .B(n4782), .Z(c[180]) );
  NANDN U4882 ( .A(n4710), .B(n4709), .Z(n4714) );
  NANDN U4883 ( .A(n4712), .B(n4711), .Z(n4713) );
  AND U4884 ( .A(n4714), .B(n4713), .Z(n4789) );
  NANDN U4885 ( .A(n4716), .B(n4715), .Z(n4720) );
  NAND U4886 ( .A(n4718), .B(n4717), .Z(n4719) );
  AND U4887 ( .A(n4720), .B(n4719), .Z(n4855) );
  NANDN U4888 ( .A(n4722), .B(n4721), .Z(n4726) );
  NANDN U4889 ( .A(n4724), .B(n4723), .Z(n4725) );
  AND U4890 ( .A(n4726), .B(n4725), .Z(n4821) );
  NAND U4891 ( .A(b[0]), .B(a[69]), .Z(n4727) );
  XNOR U4892 ( .A(b[1]), .B(n4727), .Z(n4729) );
  NANDN U4893 ( .A(b[0]), .B(a[68]), .Z(n4728) );
  NAND U4894 ( .A(n4729), .B(n4728), .Z(n4801) );
  NANDN U4895 ( .A(n9891), .B(n4730), .Z(n4732) );
  XOR U4896 ( .A(b[13]), .B(a[57]), .Z(n4807) );
  NANDN U4897 ( .A(n9935), .B(n4807), .Z(n4731) );
  AND U4898 ( .A(n4732), .B(n4731), .Z(n4799) );
  AND U4899 ( .A(b[15]), .B(a[53]), .Z(n4798) );
  XNOR U4900 ( .A(n4799), .B(n4798), .Z(n4800) );
  XNOR U4901 ( .A(n4801), .B(n4800), .Z(n4819) );
  NANDN U4902 ( .A(n9437), .B(n4733), .Z(n4735) );
  XOR U4903 ( .A(b[5]), .B(a[65]), .Z(n4810) );
  NANDN U4904 ( .A(n9503), .B(n4810), .Z(n4734) );
  AND U4905 ( .A(n4735), .B(n4734), .Z(n4843) );
  NANDN U4906 ( .A(n9588), .B(n4736), .Z(n4738) );
  XOR U4907 ( .A(b[7]), .B(a[63]), .Z(n4813) );
  NANDN U4908 ( .A(n9639), .B(n4813), .Z(n4737) );
  AND U4909 ( .A(n4738), .B(n4737), .Z(n4841) );
  NANDN U4910 ( .A(n9374), .B(n4739), .Z(n4741) );
  XOR U4911 ( .A(b[3]), .B(a[67]), .Z(n4816) );
  NANDN U4912 ( .A(n9375), .B(n4816), .Z(n4740) );
  NAND U4913 ( .A(n4741), .B(n4740), .Z(n4840) );
  XNOR U4914 ( .A(n4841), .B(n4840), .Z(n4842) );
  XOR U4915 ( .A(n4843), .B(n4842), .Z(n4820) );
  XOR U4916 ( .A(n4819), .B(n4820), .Z(n4822) );
  XOR U4917 ( .A(n4821), .B(n4822), .Z(n4793) );
  NANDN U4918 ( .A(n4743), .B(n4742), .Z(n4747) );
  OR U4919 ( .A(n4745), .B(n4744), .Z(n4746) );
  AND U4920 ( .A(n4747), .B(n4746), .Z(n4792) );
  XNOR U4921 ( .A(n4793), .B(n4792), .Z(n4795) );
  NAND U4922 ( .A(n4748), .B(n9883), .Z(n4750) );
  XOR U4923 ( .A(b[11]), .B(a[59]), .Z(n4825) );
  NANDN U4924 ( .A(n9856), .B(n4825), .Z(n4749) );
  AND U4925 ( .A(n4750), .B(n4749), .Z(n4836) );
  NANDN U4926 ( .A(n10005), .B(n4751), .Z(n4753) );
  XOR U4927 ( .A(b[15]), .B(a[55]), .Z(n4828) );
  NANDN U4928 ( .A(n10006), .B(n4828), .Z(n4752) );
  AND U4929 ( .A(n4753), .B(n4752), .Z(n4835) );
  NANDN U4930 ( .A(n9685), .B(n4754), .Z(n4756) );
  XOR U4931 ( .A(b[9]), .B(a[61]), .Z(n4831) );
  NANDN U4932 ( .A(n9758), .B(n4831), .Z(n4755) );
  NAND U4933 ( .A(n4756), .B(n4755), .Z(n4834) );
  XOR U4934 ( .A(n4835), .B(n4834), .Z(n4837) );
  XOR U4935 ( .A(n4836), .B(n4837), .Z(n4847) );
  NANDN U4936 ( .A(n4758), .B(n4757), .Z(n4762) );
  OR U4937 ( .A(n4760), .B(n4759), .Z(n4761) );
  AND U4938 ( .A(n4762), .B(n4761), .Z(n4846) );
  XNOR U4939 ( .A(n4847), .B(n4846), .Z(n4848) );
  NANDN U4940 ( .A(n4764), .B(n4763), .Z(n4768) );
  NANDN U4941 ( .A(n4766), .B(n4765), .Z(n4767) );
  NAND U4942 ( .A(n4768), .B(n4767), .Z(n4849) );
  XNOR U4943 ( .A(n4848), .B(n4849), .Z(n4794) );
  XOR U4944 ( .A(n4795), .B(n4794), .Z(n4853) );
  NANDN U4945 ( .A(n4770), .B(n4769), .Z(n4774) );
  NANDN U4946 ( .A(n4772), .B(n4771), .Z(n4773) );
  AND U4947 ( .A(n4774), .B(n4773), .Z(n4852) );
  XNOR U4948 ( .A(n4853), .B(n4852), .Z(n4854) );
  XOR U4949 ( .A(n4855), .B(n4854), .Z(n4787) );
  NANDN U4950 ( .A(n4776), .B(n4775), .Z(n4780) );
  NAND U4951 ( .A(n4778), .B(n4777), .Z(n4779) );
  AND U4952 ( .A(n4780), .B(n4779), .Z(n4786) );
  XNOR U4953 ( .A(n4787), .B(n4786), .Z(n4788) );
  XNOR U4954 ( .A(n4789), .B(n4788), .Z(n4858) );
  XNOR U4955 ( .A(sreg[181]), .B(n4858), .Z(n4860) );
  NANDN U4956 ( .A(sreg[180]), .B(n4781), .Z(n4785) );
  NAND U4957 ( .A(n4783), .B(n4782), .Z(n4784) );
  NAND U4958 ( .A(n4785), .B(n4784), .Z(n4859) );
  XNOR U4959 ( .A(n4860), .B(n4859), .Z(c[181]) );
  NANDN U4960 ( .A(n4787), .B(n4786), .Z(n4791) );
  NANDN U4961 ( .A(n4789), .B(n4788), .Z(n4790) );
  AND U4962 ( .A(n4791), .B(n4790), .Z(n4866) );
  NANDN U4963 ( .A(n4793), .B(n4792), .Z(n4797) );
  NAND U4964 ( .A(n4795), .B(n4794), .Z(n4796) );
  AND U4965 ( .A(n4797), .B(n4796), .Z(n4932) );
  NANDN U4966 ( .A(n4799), .B(n4798), .Z(n4803) );
  NANDN U4967 ( .A(n4801), .B(n4800), .Z(n4802) );
  AND U4968 ( .A(n4803), .B(n4802), .Z(n4898) );
  NAND U4969 ( .A(b[0]), .B(a[70]), .Z(n4804) );
  XNOR U4970 ( .A(b[1]), .B(n4804), .Z(n4806) );
  NANDN U4971 ( .A(b[0]), .B(a[69]), .Z(n4805) );
  NAND U4972 ( .A(n4806), .B(n4805), .Z(n4878) );
  NANDN U4973 ( .A(n9891), .B(n4807), .Z(n4809) );
  XOR U4974 ( .A(b[13]), .B(a[58]), .Z(n4881) );
  NANDN U4975 ( .A(n9935), .B(n4881), .Z(n4808) );
  AND U4976 ( .A(n4809), .B(n4808), .Z(n4876) );
  AND U4977 ( .A(b[15]), .B(a[54]), .Z(n4875) );
  XNOR U4978 ( .A(n4876), .B(n4875), .Z(n4877) );
  XNOR U4979 ( .A(n4878), .B(n4877), .Z(n4896) );
  NANDN U4980 ( .A(n9437), .B(n4810), .Z(n4812) );
  XOR U4981 ( .A(b[5]), .B(a[66]), .Z(n4887) );
  NANDN U4982 ( .A(n9503), .B(n4887), .Z(n4811) );
  AND U4983 ( .A(n4812), .B(n4811), .Z(n4920) );
  NANDN U4984 ( .A(n9588), .B(n4813), .Z(n4815) );
  XOR U4985 ( .A(b[7]), .B(a[64]), .Z(n4890) );
  NANDN U4986 ( .A(n9639), .B(n4890), .Z(n4814) );
  AND U4987 ( .A(n4815), .B(n4814), .Z(n4918) );
  NANDN U4988 ( .A(n9374), .B(n4816), .Z(n4818) );
  XOR U4989 ( .A(b[3]), .B(a[68]), .Z(n4893) );
  NANDN U4990 ( .A(n9375), .B(n4893), .Z(n4817) );
  NAND U4991 ( .A(n4818), .B(n4817), .Z(n4917) );
  XNOR U4992 ( .A(n4918), .B(n4917), .Z(n4919) );
  XOR U4993 ( .A(n4920), .B(n4919), .Z(n4897) );
  XOR U4994 ( .A(n4896), .B(n4897), .Z(n4899) );
  XOR U4995 ( .A(n4898), .B(n4899), .Z(n4870) );
  NANDN U4996 ( .A(n4820), .B(n4819), .Z(n4824) );
  OR U4997 ( .A(n4822), .B(n4821), .Z(n4823) );
  AND U4998 ( .A(n4824), .B(n4823), .Z(n4869) );
  XNOR U4999 ( .A(n4870), .B(n4869), .Z(n4872) );
  NAND U5000 ( .A(n4825), .B(n9883), .Z(n4827) );
  XOR U5001 ( .A(b[11]), .B(a[60]), .Z(n4902) );
  NANDN U5002 ( .A(n9856), .B(n4902), .Z(n4826) );
  AND U5003 ( .A(n4827), .B(n4826), .Z(n4913) );
  NANDN U5004 ( .A(n10005), .B(n4828), .Z(n4830) );
  XOR U5005 ( .A(b[15]), .B(a[56]), .Z(n4905) );
  NANDN U5006 ( .A(n10006), .B(n4905), .Z(n4829) );
  AND U5007 ( .A(n4830), .B(n4829), .Z(n4912) );
  NANDN U5008 ( .A(n9685), .B(n4831), .Z(n4833) );
  XOR U5009 ( .A(b[9]), .B(a[62]), .Z(n4908) );
  NANDN U5010 ( .A(n9758), .B(n4908), .Z(n4832) );
  NAND U5011 ( .A(n4833), .B(n4832), .Z(n4911) );
  XOR U5012 ( .A(n4912), .B(n4911), .Z(n4914) );
  XOR U5013 ( .A(n4913), .B(n4914), .Z(n4924) );
  NANDN U5014 ( .A(n4835), .B(n4834), .Z(n4839) );
  OR U5015 ( .A(n4837), .B(n4836), .Z(n4838) );
  AND U5016 ( .A(n4839), .B(n4838), .Z(n4923) );
  XNOR U5017 ( .A(n4924), .B(n4923), .Z(n4925) );
  NANDN U5018 ( .A(n4841), .B(n4840), .Z(n4845) );
  NANDN U5019 ( .A(n4843), .B(n4842), .Z(n4844) );
  NAND U5020 ( .A(n4845), .B(n4844), .Z(n4926) );
  XNOR U5021 ( .A(n4925), .B(n4926), .Z(n4871) );
  XOR U5022 ( .A(n4872), .B(n4871), .Z(n4930) );
  NANDN U5023 ( .A(n4847), .B(n4846), .Z(n4851) );
  NANDN U5024 ( .A(n4849), .B(n4848), .Z(n4850) );
  AND U5025 ( .A(n4851), .B(n4850), .Z(n4929) );
  XNOR U5026 ( .A(n4930), .B(n4929), .Z(n4931) );
  XOR U5027 ( .A(n4932), .B(n4931), .Z(n4864) );
  NANDN U5028 ( .A(n4853), .B(n4852), .Z(n4857) );
  NAND U5029 ( .A(n4855), .B(n4854), .Z(n4856) );
  AND U5030 ( .A(n4857), .B(n4856), .Z(n4863) );
  XNOR U5031 ( .A(n4864), .B(n4863), .Z(n4865) );
  XNOR U5032 ( .A(n4866), .B(n4865), .Z(n4935) );
  XNOR U5033 ( .A(sreg[182]), .B(n4935), .Z(n4937) );
  NANDN U5034 ( .A(sreg[181]), .B(n4858), .Z(n4862) );
  NAND U5035 ( .A(n4860), .B(n4859), .Z(n4861) );
  NAND U5036 ( .A(n4862), .B(n4861), .Z(n4936) );
  XNOR U5037 ( .A(n4937), .B(n4936), .Z(c[182]) );
  NANDN U5038 ( .A(n4864), .B(n4863), .Z(n4868) );
  NANDN U5039 ( .A(n4866), .B(n4865), .Z(n4867) );
  AND U5040 ( .A(n4868), .B(n4867), .Z(n4943) );
  NANDN U5041 ( .A(n4870), .B(n4869), .Z(n4874) );
  NAND U5042 ( .A(n4872), .B(n4871), .Z(n4873) );
  AND U5043 ( .A(n4874), .B(n4873), .Z(n5009) );
  NANDN U5044 ( .A(n4876), .B(n4875), .Z(n4880) );
  NANDN U5045 ( .A(n4878), .B(n4877), .Z(n4879) );
  AND U5046 ( .A(n4880), .B(n4879), .Z(n4975) );
  NANDN U5047 ( .A(n9891), .B(n4881), .Z(n4883) );
  XOR U5048 ( .A(b[13]), .B(a[59]), .Z(n4961) );
  NANDN U5049 ( .A(n9935), .B(n4961), .Z(n4882) );
  AND U5050 ( .A(n4883), .B(n4882), .Z(n4953) );
  AND U5051 ( .A(b[15]), .B(a[55]), .Z(n4952) );
  XNOR U5052 ( .A(n4953), .B(n4952), .Z(n4954) );
  NAND U5053 ( .A(b[0]), .B(a[71]), .Z(n4884) );
  XNOR U5054 ( .A(b[1]), .B(n4884), .Z(n4886) );
  NANDN U5055 ( .A(b[0]), .B(a[70]), .Z(n4885) );
  NAND U5056 ( .A(n4886), .B(n4885), .Z(n4955) );
  XNOR U5057 ( .A(n4954), .B(n4955), .Z(n4973) );
  NANDN U5058 ( .A(n9437), .B(n4887), .Z(n4889) );
  XOR U5059 ( .A(b[5]), .B(a[67]), .Z(n4964) );
  NANDN U5060 ( .A(n9503), .B(n4964), .Z(n4888) );
  AND U5061 ( .A(n4889), .B(n4888), .Z(n4997) );
  NANDN U5062 ( .A(n9588), .B(n4890), .Z(n4892) );
  XOR U5063 ( .A(b[7]), .B(a[65]), .Z(n4967) );
  NANDN U5064 ( .A(n9639), .B(n4967), .Z(n4891) );
  AND U5065 ( .A(n4892), .B(n4891), .Z(n4995) );
  NANDN U5066 ( .A(n9374), .B(n4893), .Z(n4895) );
  XOR U5067 ( .A(b[3]), .B(a[69]), .Z(n4970) );
  NANDN U5068 ( .A(n9375), .B(n4970), .Z(n4894) );
  NAND U5069 ( .A(n4895), .B(n4894), .Z(n4994) );
  XNOR U5070 ( .A(n4995), .B(n4994), .Z(n4996) );
  XOR U5071 ( .A(n4997), .B(n4996), .Z(n4974) );
  XOR U5072 ( .A(n4973), .B(n4974), .Z(n4976) );
  XOR U5073 ( .A(n4975), .B(n4976), .Z(n4947) );
  NANDN U5074 ( .A(n4897), .B(n4896), .Z(n4901) );
  OR U5075 ( .A(n4899), .B(n4898), .Z(n4900) );
  AND U5076 ( .A(n4901), .B(n4900), .Z(n4946) );
  XNOR U5077 ( .A(n4947), .B(n4946), .Z(n4949) );
  NAND U5078 ( .A(n4902), .B(n9883), .Z(n4904) );
  XOR U5079 ( .A(b[11]), .B(a[61]), .Z(n4979) );
  NANDN U5080 ( .A(n9856), .B(n4979), .Z(n4903) );
  AND U5081 ( .A(n4904), .B(n4903), .Z(n4990) );
  NANDN U5082 ( .A(n10005), .B(n4905), .Z(n4907) );
  XOR U5083 ( .A(b[15]), .B(a[57]), .Z(n4982) );
  NANDN U5084 ( .A(n10006), .B(n4982), .Z(n4906) );
  AND U5085 ( .A(n4907), .B(n4906), .Z(n4989) );
  NANDN U5086 ( .A(n9685), .B(n4908), .Z(n4910) );
  XOR U5087 ( .A(b[9]), .B(a[63]), .Z(n4985) );
  NANDN U5088 ( .A(n9758), .B(n4985), .Z(n4909) );
  NAND U5089 ( .A(n4910), .B(n4909), .Z(n4988) );
  XOR U5090 ( .A(n4989), .B(n4988), .Z(n4991) );
  XOR U5091 ( .A(n4990), .B(n4991), .Z(n5001) );
  NANDN U5092 ( .A(n4912), .B(n4911), .Z(n4916) );
  OR U5093 ( .A(n4914), .B(n4913), .Z(n4915) );
  AND U5094 ( .A(n4916), .B(n4915), .Z(n5000) );
  XNOR U5095 ( .A(n5001), .B(n5000), .Z(n5002) );
  NANDN U5096 ( .A(n4918), .B(n4917), .Z(n4922) );
  NANDN U5097 ( .A(n4920), .B(n4919), .Z(n4921) );
  NAND U5098 ( .A(n4922), .B(n4921), .Z(n5003) );
  XNOR U5099 ( .A(n5002), .B(n5003), .Z(n4948) );
  XOR U5100 ( .A(n4949), .B(n4948), .Z(n5007) );
  NANDN U5101 ( .A(n4924), .B(n4923), .Z(n4928) );
  NANDN U5102 ( .A(n4926), .B(n4925), .Z(n4927) );
  AND U5103 ( .A(n4928), .B(n4927), .Z(n5006) );
  XNOR U5104 ( .A(n5007), .B(n5006), .Z(n5008) );
  XOR U5105 ( .A(n5009), .B(n5008), .Z(n4941) );
  NANDN U5106 ( .A(n4930), .B(n4929), .Z(n4934) );
  NAND U5107 ( .A(n4932), .B(n4931), .Z(n4933) );
  AND U5108 ( .A(n4934), .B(n4933), .Z(n4940) );
  XNOR U5109 ( .A(n4941), .B(n4940), .Z(n4942) );
  XNOR U5110 ( .A(n4943), .B(n4942), .Z(n5012) );
  XNOR U5111 ( .A(sreg[183]), .B(n5012), .Z(n5014) );
  NANDN U5112 ( .A(sreg[182]), .B(n4935), .Z(n4939) );
  NAND U5113 ( .A(n4937), .B(n4936), .Z(n4938) );
  NAND U5114 ( .A(n4939), .B(n4938), .Z(n5013) );
  XNOR U5115 ( .A(n5014), .B(n5013), .Z(c[183]) );
  NANDN U5116 ( .A(n4941), .B(n4940), .Z(n4945) );
  NANDN U5117 ( .A(n4943), .B(n4942), .Z(n4944) );
  AND U5118 ( .A(n4945), .B(n4944), .Z(n5020) );
  NANDN U5119 ( .A(n4947), .B(n4946), .Z(n4951) );
  NAND U5120 ( .A(n4949), .B(n4948), .Z(n4950) );
  AND U5121 ( .A(n4951), .B(n4950), .Z(n5086) );
  NANDN U5122 ( .A(n4953), .B(n4952), .Z(n4957) );
  NANDN U5123 ( .A(n4955), .B(n4954), .Z(n4956) );
  AND U5124 ( .A(n4957), .B(n4956), .Z(n5052) );
  NAND U5125 ( .A(b[0]), .B(a[72]), .Z(n4958) );
  XNOR U5126 ( .A(b[1]), .B(n4958), .Z(n4960) );
  NANDN U5127 ( .A(b[0]), .B(a[71]), .Z(n4959) );
  NAND U5128 ( .A(n4960), .B(n4959), .Z(n5032) );
  NANDN U5129 ( .A(n9891), .B(n4961), .Z(n4963) );
  XOR U5130 ( .A(b[13]), .B(a[60]), .Z(n5038) );
  NANDN U5131 ( .A(n9935), .B(n5038), .Z(n4962) );
  AND U5132 ( .A(n4963), .B(n4962), .Z(n5030) );
  AND U5133 ( .A(b[15]), .B(a[56]), .Z(n5029) );
  XNOR U5134 ( .A(n5030), .B(n5029), .Z(n5031) );
  XNOR U5135 ( .A(n5032), .B(n5031), .Z(n5050) );
  NANDN U5136 ( .A(n9437), .B(n4964), .Z(n4966) );
  XOR U5137 ( .A(b[5]), .B(a[68]), .Z(n5041) );
  NANDN U5138 ( .A(n9503), .B(n5041), .Z(n4965) );
  AND U5139 ( .A(n4966), .B(n4965), .Z(n5074) );
  NANDN U5140 ( .A(n9588), .B(n4967), .Z(n4969) );
  XOR U5141 ( .A(b[7]), .B(a[66]), .Z(n5044) );
  NANDN U5142 ( .A(n9639), .B(n5044), .Z(n4968) );
  AND U5143 ( .A(n4969), .B(n4968), .Z(n5072) );
  NANDN U5144 ( .A(n9374), .B(n4970), .Z(n4972) );
  XOR U5145 ( .A(b[3]), .B(a[70]), .Z(n5047) );
  NANDN U5146 ( .A(n9375), .B(n5047), .Z(n4971) );
  NAND U5147 ( .A(n4972), .B(n4971), .Z(n5071) );
  XNOR U5148 ( .A(n5072), .B(n5071), .Z(n5073) );
  XOR U5149 ( .A(n5074), .B(n5073), .Z(n5051) );
  XOR U5150 ( .A(n5050), .B(n5051), .Z(n5053) );
  XOR U5151 ( .A(n5052), .B(n5053), .Z(n5024) );
  NANDN U5152 ( .A(n4974), .B(n4973), .Z(n4978) );
  OR U5153 ( .A(n4976), .B(n4975), .Z(n4977) );
  AND U5154 ( .A(n4978), .B(n4977), .Z(n5023) );
  XNOR U5155 ( .A(n5024), .B(n5023), .Z(n5026) );
  NAND U5156 ( .A(n4979), .B(n9883), .Z(n4981) );
  XOR U5157 ( .A(b[11]), .B(a[62]), .Z(n5056) );
  NANDN U5158 ( .A(n9856), .B(n5056), .Z(n4980) );
  AND U5159 ( .A(n4981), .B(n4980), .Z(n5067) );
  NANDN U5160 ( .A(n10005), .B(n4982), .Z(n4984) );
  XOR U5161 ( .A(b[15]), .B(a[58]), .Z(n5059) );
  NANDN U5162 ( .A(n10006), .B(n5059), .Z(n4983) );
  AND U5163 ( .A(n4984), .B(n4983), .Z(n5066) );
  NANDN U5164 ( .A(n9685), .B(n4985), .Z(n4987) );
  XOR U5165 ( .A(b[9]), .B(a[64]), .Z(n5062) );
  NANDN U5166 ( .A(n9758), .B(n5062), .Z(n4986) );
  NAND U5167 ( .A(n4987), .B(n4986), .Z(n5065) );
  XOR U5168 ( .A(n5066), .B(n5065), .Z(n5068) );
  XOR U5169 ( .A(n5067), .B(n5068), .Z(n5078) );
  NANDN U5170 ( .A(n4989), .B(n4988), .Z(n4993) );
  OR U5171 ( .A(n4991), .B(n4990), .Z(n4992) );
  AND U5172 ( .A(n4993), .B(n4992), .Z(n5077) );
  XNOR U5173 ( .A(n5078), .B(n5077), .Z(n5079) );
  NANDN U5174 ( .A(n4995), .B(n4994), .Z(n4999) );
  NANDN U5175 ( .A(n4997), .B(n4996), .Z(n4998) );
  NAND U5176 ( .A(n4999), .B(n4998), .Z(n5080) );
  XNOR U5177 ( .A(n5079), .B(n5080), .Z(n5025) );
  XOR U5178 ( .A(n5026), .B(n5025), .Z(n5084) );
  NANDN U5179 ( .A(n5001), .B(n5000), .Z(n5005) );
  NANDN U5180 ( .A(n5003), .B(n5002), .Z(n5004) );
  AND U5181 ( .A(n5005), .B(n5004), .Z(n5083) );
  XNOR U5182 ( .A(n5084), .B(n5083), .Z(n5085) );
  XOR U5183 ( .A(n5086), .B(n5085), .Z(n5018) );
  NANDN U5184 ( .A(n5007), .B(n5006), .Z(n5011) );
  NAND U5185 ( .A(n5009), .B(n5008), .Z(n5010) );
  AND U5186 ( .A(n5011), .B(n5010), .Z(n5017) );
  XNOR U5187 ( .A(n5018), .B(n5017), .Z(n5019) );
  XNOR U5188 ( .A(n5020), .B(n5019), .Z(n5089) );
  XNOR U5189 ( .A(sreg[184]), .B(n5089), .Z(n5091) );
  NANDN U5190 ( .A(sreg[183]), .B(n5012), .Z(n5016) );
  NAND U5191 ( .A(n5014), .B(n5013), .Z(n5015) );
  NAND U5192 ( .A(n5016), .B(n5015), .Z(n5090) );
  XNOR U5193 ( .A(n5091), .B(n5090), .Z(c[184]) );
  NANDN U5194 ( .A(n5018), .B(n5017), .Z(n5022) );
  NANDN U5195 ( .A(n5020), .B(n5019), .Z(n5021) );
  AND U5196 ( .A(n5022), .B(n5021), .Z(n5097) );
  NANDN U5197 ( .A(n5024), .B(n5023), .Z(n5028) );
  NAND U5198 ( .A(n5026), .B(n5025), .Z(n5027) );
  AND U5199 ( .A(n5028), .B(n5027), .Z(n5163) );
  NANDN U5200 ( .A(n5030), .B(n5029), .Z(n5034) );
  NANDN U5201 ( .A(n5032), .B(n5031), .Z(n5033) );
  AND U5202 ( .A(n5034), .B(n5033), .Z(n5129) );
  NAND U5203 ( .A(b[0]), .B(a[73]), .Z(n5035) );
  XNOR U5204 ( .A(b[1]), .B(n5035), .Z(n5037) );
  NANDN U5205 ( .A(b[0]), .B(a[72]), .Z(n5036) );
  NAND U5206 ( .A(n5037), .B(n5036), .Z(n5109) );
  NANDN U5207 ( .A(n9891), .B(n5038), .Z(n5040) );
  XOR U5208 ( .A(b[13]), .B(a[61]), .Z(n5115) );
  NANDN U5209 ( .A(n9935), .B(n5115), .Z(n5039) );
  AND U5210 ( .A(n5040), .B(n5039), .Z(n5107) );
  AND U5211 ( .A(b[15]), .B(a[57]), .Z(n5106) );
  XNOR U5212 ( .A(n5107), .B(n5106), .Z(n5108) );
  XNOR U5213 ( .A(n5109), .B(n5108), .Z(n5127) );
  NANDN U5214 ( .A(n9437), .B(n5041), .Z(n5043) );
  XOR U5215 ( .A(b[5]), .B(a[69]), .Z(n5118) );
  NANDN U5216 ( .A(n9503), .B(n5118), .Z(n5042) );
  AND U5217 ( .A(n5043), .B(n5042), .Z(n5151) );
  NANDN U5218 ( .A(n9588), .B(n5044), .Z(n5046) );
  XOR U5219 ( .A(b[7]), .B(a[67]), .Z(n5121) );
  NANDN U5220 ( .A(n9639), .B(n5121), .Z(n5045) );
  AND U5221 ( .A(n5046), .B(n5045), .Z(n5149) );
  NANDN U5222 ( .A(n9374), .B(n5047), .Z(n5049) );
  XOR U5223 ( .A(b[3]), .B(a[71]), .Z(n5124) );
  NANDN U5224 ( .A(n9375), .B(n5124), .Z(n5048) );
  NAND U5225 ( .A(n5049), .B(n5048), .Z(n5148) );
  XNOR U5226 ( .A(n5149), .B(n5148), .Z(n5150) );
  XOR U5227 ( .A(n5151), .B(n5150), .Z(n5128) );
  XOR U5228 ( .A(n5127), .B(n5128), .Z(n5130) );
  XOR U5229 ( .A(n5129), .B(n5130), .Z(n5101) );
  NANDN U5230 ( .A(n5051), .B(n5050), .Z(n5055) );
  OR U5231 ( .A(n5053), .B(n5052), .Z(n5054) );
  AND U5232 ( .A(n5055), .B(n5054), .Z(n5100) );
  XNOR U5233 ( .A(n5101), .B(n5100), .Z(n5103) );
  NAND U5234 ( .A(n5056), .B(n9883), .Z(n5058) );
  XOR U5235 ( .A(b[11]), .B(a[63]), .Z(n5133) );
  NANDN U5236 ( .A(n9856), .B(n5133), .Z(n5057) );
  AND U5237 ( .A(n5058), .B(n5057), .Z(n5144) );
  NANDN U5238 ( .A(n10005), .B(n5059), .Z(n5061) );
  XOR U5239 ( .A(b[15]), .B(a[59]), .Z(n5136) );
  NANDN U5240 ( .A(n10006), .B(n5136), .Z(n5060) );
  AND U5241 ( .A(n5061), .B(n5060), .Z(n5143) );
  NANDN U5242 ( .A(n9685), .B(n5062), .Z(n5064) );
  XOR U5243 ( .A(b[9]), .B(a[65]), .Z(n5139) );
  NANDN U5244 ( .A(n9758), .B(n5139), .Z(n5063) );
  NAND U5245 ( .A(n5064), .B(n5063), .Z(n5142) );
  XOR U5246 ( .A(n5143), .B(n5142), .Z(n5145) );
  XOR U5247 ( .A(n5144), .B(n5145), .Z(n5155) );
  NANDN U5248 ( .A(n5066), .B(n5065), .Z(n5070) );
  OR U5249 ( .A(n5068), .B(n5067), .Z(n5069) );
  AND U5250 ( .A(n5070), .B(n5069), .Z(n5154) );
  XNOR U5251 ( .A(n5155), .B(n5154), .Z(n5156) );
  NANDN U5252 ( .A(n5072), .B(n5071), .Z(n5076) );
  NANDN U5253 ( .A(n5074), .B(n5073), .Z(n5075) );
  NAND U5254 ( .A(n5076), .B(n5075), .Z(n5157) );
  XNOR U5255 ( .A(n5156), .B(n5157), .Z(n5102) );
  XOR U5256 ( .A(n5103), .B(n5102), .Z(n5161) );
  NANDN U5257 ( .A(n5078), .B(n5077), .Z(n5082) );
  NANDN U5258 ( .A(n5080), .B(n5079), .Z(n5081) );
  AND U5259 ( .A(n5082), .B(n5081), .Z(n5160) );
  XNOR U5260 ( .A(n5161), .B(n5160), .Z(n5162) );
  XOR U5261 ( .A(n5163), .B(n5162), .Z(n5095) );
  NANDN U5262 ( .A(n5084), .B(n5083), .Z(n5088) );
  NAND U5263 ( .A(n5086), .B(n5085), .Z(n5087) );
  AND U5264 ( .A(n5088), .B(n5087), .Z(n5094) );
  XNOR U5265 ( .A(n5095), .B(n5094), .Z(n5096) );
  XNOR U5266 ( .A(n5097), .B(n5096), .Z(n5166) );
  XNOR U5267 ( .A(sreg[185]), .B(n5166), .Z(n5168) );
  NANDN U5268 ( .A(sreg[184]), .B(n5089), .Z(n5093) );
  NAND U5269 ( .A(n5091), .B(n5090), .Z(n5092) );
  NAND U5270 ( .A(n5093), .B(n5092), .Z(n5167) );
  XNOR U5271 ( .A(n5168), .B(n5167), .Z(c[185]) );
  NANDN U5272 ( .A(n5095), .B(n5094), .Z(n5099) );
  NANDN U5273 ( .A(n5097), .B(n5096), .Z(n5098) );
  AND U5274 ( .A(n5099), .B(n5098), .Z(n5174) );
  NANDN U5275 ( .A(n5101), .B(n5100), .Z(n5105) );
  NAND U5276 ( .A(n5103), .B(n5102), .Z(n5104) );
  AND U5277 ( .A(n5105), .B(n5104), .Z(n5240) );
  NANDN U5278 ( .A(n5107), .B(n5106), .Z(n5111) );
  NANDN U5279 ( .A(n5109), .B(n5108), .Z(n5110) );
  AND U5280 ( .A(n5111), .B(n5110), .Z(n5206) );
  NAND U5281 ( .A(b[0]), .B(a[74]), .Z(n5112) );
  XNOR U5282 ( .A(b[1]), .B(n5112), .Z(n5114) );
  NANDN U5283 ( .A(b[0]), .B(a[73]), .Z(n5113) );
  NAND U5284 ( .A(n5114), .B(n5113), .Z(n5186) );
  NANDN U5285 ( .A(n9891), .B(n5115), .Z(n5117) );
  XOR U5286 ( .A(b[13]), .B(a[62]), .Z(n5192) );
  NANDN U5287 ( .A(n9935), .B(n5192), .Z(n5116) );
  AND U5288 ( .A(n5117), .B(n5116), .Z(n5184) );
  AND U5289 ( .A(b[15]), .B(a[58]), .Z(n5183) );
  XNOR U5290 ( .A(n5184), .B(n5183), .Z(n5185) );
  XNOR U5291 ( .A(n5186), .B(n5185), .Z(n5204) );
  NANDN U5292 ( .A(n9437), .B(n5118), .Z(n5120) );
  XOR U5293 ( .A(b[5]), .B(a[70]), .Z(n5195) );
  NANDN U5294 ( .A(n9503), .B(n5195), .Z(n5119) );
  AND U5295 ( .A(n5120), .B(n5119), .Z(n5228) );
  NANDN U5296 ( .A(n9588), .B(n5121), .Z(n5123) );
  XOR U5297 ( .A(b[7]), .B(a[68]), .Z(n5198) );
  NANDN U5298 ( .A(n9639), .B(n5198), .Z(n5122) );
  AND U5299 ( .A(n5123), .B(n5122), .Z(n5226) );
  NANDN U5300 ( .A(n9374), .B(n5124), .Z(n5126) );
  XOR U5301 ( .A(b[3]), .B(a[72]), .Z(n5201) );
  NANDN U5302 ( .A(n9375), .B(n5201), .Z(n5125) );
  NAND U5303 ( .A(n5126), .B(n5125), .Z(n5225) );
  XNOR U5304 ( .A(n5226), .B(n5225), .Z(n5227) );
  XOR U5305 ( .A(n5228), .B(n5227), .Z(n5205) );
  XOR U5306 ( .A(n5204), .B(n5205), .Z(n5207) );
  XOR U5307 ( .A(n5206), .B(n5207), .Z(n5178) );
  NANDN U5308 ( .A(n5128), .B(n5127), .Z(n5132) );
  OR U5309 ( .A(n5130), .B(n5129), .Z(n5131) );
  AND U5310 ( .A(n5132), .B(n5131), .Z(n5177) );
  XNOR U5311 ( .A(n5178), .B(n5177), .Z(n5180) );
  NAND U5312 ( .A(n5133), .B(n9883), .Z(n5135) );
  XOR U5313 ( .A(b[11]), .B(a[64]), .Z(n5210) );
  NANDN U5314 ( .A(n9856), .B(n5210), .Z(n5134) );
  AND U5315 ( .A(n5135), .B(n5134), .Z(n5221) );
  NANDN U5316 ( .A(n10005), .B(n5136), .Z(n5138) );
  XOR U5317 ( .A(b[15]), .B(a[60]), .Z(n5213) );
  NANDN U5318 ( .A(n10006), .B(n5213), .Z(n5137) );
  AND U5319 ( .A(n5138), .B(n5137), .Z(n5220) );
  NANDN U5320 ( .A(n9685), .B(n5139), .Z(n5141) );
  XOR U5321 ( .A(b[9]), .B(a[66]), .Z(n5216) );
  NANDN U5322 ( .A(n9758), .B(n5216), .Z(n5140) );
  NAND U5323 ( .A(n5141), .B(n5140), .Z(n5219) );
  XOR U5324 ( .A(n5220), .B(n5219), .Z(n5222) );
  XOR U5325 ( .A(n5221), .B(n5222), .Z(n5232) );
  NANDN U5326 ( .A(n5143), .B(n5142), .Z(n5147) );
  OR U5327 ( .A(n5145), .B(n5144), .Z(n5146) );
  AND U5328 ( .A(n5147), .B(n5146), .Z(n5231) );
  XNOR U5329 ( .A(n5232), .B(n5231), .Z(n5233) );
  NANDN U5330 ( .A(n5149), .B(n5148), .Z(n5153) );
  NANDN U5331 ( .A(n5151), .B(n5150), .Z(n5152) );
  NAND U5332 ( .A(n5153), .B(n5152), .Z(n5234) );
  XNOR U5333 ( .A(n5233), .B(n5234), .Z(n5179) );
  XOR U5334 ( .A(n5180), .B(n5179), .Z(n5238) );
  NANDN U5335 ( .A(n5155), .B(n5154), .Z(n5159) );
  NANDN U5336 ( .A(n5157), .B(n5156), .Z(n5158) );
  AND U5337 ( .A(n5159), .B(n5158), .Z(n5237) );
  XNOR U5338 ( .A(n5238), .B(n5237), .Z(n5239) );
  XOR U5339 ( .A(n5240), .B(n5239), .Z(n5172) );
  NANDN U5340 ( .A(n5161), .B(n5160), .Z(n5165) );
  NAND U5341 ( .A(n5163), .B(n5162), .Z(n5164) );
  AND U5342 ( .A(n5165), .B(n5164), .Z(n5171) );
  XNOR U5343 ( .A(n5172), .B(n5171), .Z(n5173) );
  XNOR U5344 ( .A(n5174), .B(n5173), .Z(n5243) );
  XNOR U5345 ( .A(sreg[186]), .B(n5243), .Z(n5245) );
  NANDN U5346 ( .A(sreg[185]), .B(n5166), .Z(n5170) );
  NAND U5347 ( .A(n5168), .B(n5167), .Z(n5169) );
  NAND U5348 ( .A(n5170), .B(n5169), .Z(n5244) );
  XNOR U5349 ( .A(n5245), .B(n5244), .Z(c[186]) );
  NANDN U5350 ( .A(n5172), .B(n5171), .Z(n5176) );
  NANDN U5351 ( .A(n5174), .B(n5173), .Z(n5175) );
  AND U5352 ( .A(n5176), .B(n5175), .Z(n5251) );
  NANDN U5353 ( .A(n5178), .B(n5177), .Z(n5182) );
  NAND U5354 ( .A(n5180), .B(n5179), .Z(n5181) );
  AND U5355 ( .A(n5182), .B(n5181), .Z(n5317) );
  NANDN U5356 ( .A(n5184), .B(n5183), .Z(n5188) );
  NANDN U5357 ( .A(n5186), .B(n5185), .Z(n5187) );
  AND U5358 ( .A(n5188), .B(n5187), .Z(n5283) );
  NAND U5359 ( .A(b[0]), .B(a[75]), .Z(n5189) );
  XNOR U5360 ( .A(b[1]), .B(n5189), .Z(n5191) );
  NANDN U5361 ( .A(b[0]), .B(a[74]), .Z(n5190) );
  NAND U5362 ( .A(n5191), .B(n5190), .Z(n5263) );
  NANDN U5363 ( .A(n9891), .B(n5192), .Z(n5194) );
  XOR U5364 ( .A(b[13]), .B(a[63]), .Z(n5269) );
  NANDN U5365 ( .A(n9935), .B(n5269), .Z(n5193) );
  AND U5366 ( .A(n5194), .B(n5193), .Z(n5261) );
  AND U5367 ( .A(b[15]), .B(a[59]), .Z(n5260) );
  XNOR U5368 ( .A(n5261), .B(n5260), .Z(n5262) );
  XNOR U5369 ( .A(n5263), .B(n5262), .Z(n5281) );
  NANDN U5370 ( .A(n9437), .B(n5195), .Z(n5197) );
  XOR U5371 ( .A(b[5]), .B(a[71]), .Z(n5272) );
  NANDN U5372 ( .A(n9503), .B(n5272), .Z(n5196) );
  AND U5373 ( .A(n5197), .B(n5196), .Z(n5305) );
  NANDN U5374 ( .A(n9588), .B(n5198), .Z(n5200) );
  XOR U5375 ( .A(b[7]), .B(a[69]), .Z(n5275) );
  NANDN U5376 ( .A(n9639), .B(n5275), .Z(n5199) );
  AND U5377 ( .A(n5200), .B(n5199), .Z(n5303) );
  NANDN U5378 ( .A(n9374), .B(n5201), .Z(n5203) );
  XOR U5379 ( .A(b[3]), .B(a[73]), .Z(n5278) );
  NANDN U5380 ( .A(n9375), .B(n5278), .Z(n5202) );
  NAND U5381 ( .A(n5203), .B(n5202), .Z(n5302) );
  XNOR U5382 ( .A(n5303), .B(n5302), .Z(n5304) );
  XOR U5383 ( .A(n5305), .B(n5304), .Z(n5282) );
  XOR U5384 ( .A(n5281), .B(n5282), .Z(n5284) );
  XOR U5385 ( .A(n5283), .B(n5284), .Z(n5255) );
  NANDN U5386 ( .A(n5205), .B(n5204), .Z(n5209) );
  OR U5387 ( .A(n5207), .B(n5206), .Z(n5208) );
  AND U5388 ( .A(n5209), .B(n5208), .Z(n5254) );
  XNOR U5389 ( .A(n5255), .B(n5254), .Z(n5257) );
  NAND U5390 ( .A(n5210), .B(n9883), .Z(n5212) );
  XOR U5391 ( .A(b[11]), .B(a[65]), .Z(n5287) );
  NANDN U5392 ( .A(n9856), .B(n5287), .Z(n5211) );
  AND U5393 ( .A(n5212), .B(n5211), .Z(n5298) );
  NANDN U5394 ( .A(n10005), .B(n5213), .Z(n5215) );
  XOR U5395 ( .A(b[15]), .B(a[61]), .Z(n5290) );
  NANDN U5396 ( .A(n10006), .B(n5290), .Z(n5214) );
  AND U5397 ( .A(n5215), .B(n5214), .Z(n5297) );
  NANDN U5398 ( .A(n9685), .B(n5216), .Z(n5218) );
  XOR U5399 ( .A(b[9]), .B(a[67]), .Z(n5293) );
  NANDN U5400 ( .A(n9758), .B(n5293), .Z(n5217) );
  NAND U5401 ( .A(n5218), .B(n5217), .Z(n5296) );
  XOR U5402 ( .A(n5297), .B(n5296), .Z(n5299) );
  XOR U5403 ( .A(n5298), .B(n5299), .Z(n5309) );
  NANDN U5404 ( .A(n5220), .B(n5219), .Z(n5224) );
  OR U5405 ( .A(n5222), .B(n5221), .Z(n5223) );
  AND U5406 ( .A(n5224), .B(n5223), .Z(n5308) );
  XNOR U5407 ( .A(n5309), .B(n5308), .Z(n5310) );
  NANDN U5408 ( .A(n5226), .B(n5225), .Z(n5230) );
  NANDN U5409 ( .A(n5228), .B(n5227), .Z(n5229) );
  NAND U5410 ( .A(n5230), .B(n5229), .Z(n5311) );
  XNOR U5411 ( .A(n5310), .B(n5311), .Z(n5256) );
  XOR U5412 ( .A(n5257), .B(n5256), .Z(n5315) );
  NANDN U5413 ( .A(n5232), .B(n5231), .Z(n5236) );
  NANDN U5414 ( .A(n5234), .B(n5233), .Z(n5235) );
  AND U5415 ( .A(n5236), .B(n5235), .Z(n5314) );
  XNOR U5416 ( .A(n5315), .B(n5314), .Z(n5316) );
  XOR U5417 ( .A(n5317), .B(n5316), .Z(n5249) );
  NANDN U5418 ( .A(n5238), .B(n5237), .Z(n5242) );
  NAND U5419 ( .A(n5240), .B(n5239), .Z(n5241) );
  AND U5420 ( .A(n5242), .B(n5241), .Z(n5248) );
  XNOR U5421 ( .A(n5249), .B(n5248), .Z(n5250) );
  XNOR U5422 ( .A(n5251), .B(n5250), .Z(n5320) );
  XNOR U5423 ( .A(sreg[187]), .B(n5320), .Z(n5322) );
  NANDN U5424 ( .A(sreg[186]), .B(n5243), .Z(n5247) );
  NAND U5425 ( .A(n5245), .B(n5244), .Z(n5246) );
  NAND U5426 ( .A(n5247), .B(n5246), .Z(n5321) );
  XNOR U5427 ( .A(n5322), .B(n5321), .Z(c[187]) );
  NANDN U5428 ( .A(n5249), .B(n5248), .Z(n5253) );
  NANDN U5429 ( .A(n5251), .B(n5250), .Z(n5252) );
  AND U5430 ( .A(n5253), .B(n5252), .Z(n5328) );
  NANDN U5431 ( .A(n5255), .B(n5254), .Z(n5259) );
  NAND U5432 ( .A(n5257), .B(n5256), .Z(n5258) );
  AND U5433 ( .A(n5259), .B(n5258), .Z(n5394) );
  NANDN U5434 ( .A(n5261), .B(n5260), .Z(n5265) );
  NANDN U5435 ( .A(n5263), .B(n5262), .Z(n5264) );
  AND U5436 ( .A(n5265), .B(n5264), .Z(n5381) );
  NAND U5437 ( .A(b[0]), .B(a[76]), .Z(n5266) );
  XNOR U5438 ( .A(b[1]), .B(n5266), .Z(n5268) );
  NANDN U5439 ( .A(b[0]), .B(a[75]), .Z(n5267) );
  NAND U5440 ( .A(n5268), .B(n5267), .Z(n5361) );
  NANDN U5441 ( .A(n9891), .B(n5269), .Z(n5271) );
  XOR U5442 ( .A(b[13]), .B(a[64]), .Z(n5367) );
  NANDN U5443 ( .A(n9935), .B(n5367), .Z(n5270) );
  AND U5444 ( .A(n5271), .B(n5270), .Z(n5359) );
  AND U5445 ( .A(b[15]), .B(a[60]), .Z(n5358) );
  XNOR U5446 ( .A(n5359), .B(n5358), .Z(n5360) );
  XNOR U5447 ( .A(n5361), .B(n5360), .Z(n5379) );
  NANDN U5448 ( .A(n9437), .B(n5272), .Z(n5274) );
  XOR U5449 ( .A(b[5]), .B(a[72]), .Z(n5370) );
  NANDN U5450 ( .A(n9503), .B(n5370), .Z(n5273) );
  AND U5451 ( .A(n5274), .B(n5273), .Z(n5355) );
  NANDN U5452 ( .A(n9588), .B(n5275), .Z(n5277) );
  XOR U5453 ( .A(b[7]), .B(a[70]), .Z(n5373) );
  NANDN U5454 ( .A(n9639), .B(n5373), .Z(n5276) );
  AND U5455 ( .A(n5277), .B(n5276), .Z(n5353) );
  NANDN U5456 ( .A(n9374), .B(n5278), .Z(n5280) );
  XOR U5457 ( .A(b[3]), .B(a[74]), .Z(n5376) );
  NANDN U5458 ( .A(n9375), .B(n5376), .Z(n5279) );
  NAND U5459 ( .A(n5280), .B(n5279), .Z(n5352) );
  XNOR U5460 ( .A(n5353), .B(n5352), .Z(n5354) );
  XOR U5461 ( .A(n5355), .B(n5354), .Z(n5380) );
  XOR U5462 ( .A(n5379), .B(n5380), .Z(n5382) );
  XOR U5463 ( .A(n5381), .B(n5382), .Z(n5332) );
  NANDN U5464 ( .A(n5282), .B(n5281), .Z(n5286) );
  OR U5465 ( .A(n5284), .B(n5283), .Z(n5285) );
  AND U5466 ( .A(n5286), .B(n5285), .Z(n5331) );
  XNOR U5467 ( .A(n5332), .B(n5331), .Z(n5334) );
  NAND U5468 ( .A(n5287), .B(n9883), .Z(n5289) );
  XOR U5469 ( .A(b[11]), .B(a[66]), .Z(n5337) );
  NANDN U5470 ( .A(n9856), .B(n5337), .Z(n5288) );
  AND U5471 ( .A(n5289), .B(n5288), .Z(n5348) );
  NANDN U5472 ( .A(n10005), .B(n5290), .Z(n5292) );
  XOR U5473 ( .A(b[15]), .B(a[62]), .Z(n5340) );
  NANDN U5474 ( .A(n10006), .B(n5340), .Z(n5291) );
  AND U5475 ( .A(n5292), .B(n5291), .Z(n5347) );
  NANDN U5476 ( .A(n9685), .B(n5293), .Z(n5295) );
  XOR U5477 ( .A(b[9]), .B(a[68]), .Z(n5343) );
  NANDN U5478 ( .A(n9758), .B(n5343), .Z(n5294) );
  NAND U5479 ( .A(n5295), .B(n5294), .Z(n5346) );
  XOR U5480 ( .A(n5347), .B(n5346), .Z(n5349) );
  XOR U5481 ( .A(n5348), .B(n5349), .Z(n5386) );
  NANDN U5482 ( .A(n5297), .B(n5296), .Z(n5301) );
  OR U5483 ( .A(n5299), .B(n5298), .Z(n5300) );
  AND U5484 ( .A(n5301), .B(n5300), .Z(n5385) );
  XNOR U5485 ( .A(n5386), .B(n5385), .Z(n5387) );
  NANDN U5486 ( .A(n5303), .B(n5302), .Z(n5307) );
  NANDN U5487 ( .A(n5305), .B(n5304), .Z(n5306) );
  NAND U5488 ( .A(n5307), .B(n5306), .Z(n5388) );
  XNOR U5489 ( .A(n5387), .B(n5388), .Z(n5333) );
  XOR U5490 ( .A(n5334), .B(n5333), .Z(n5392) );
  NANDN U5491 ( .A(n5309), .B(n5308), .Z(n5313) );
  NANDN U5492 ( .A(n5311), .B(n5310), .Z(n5312) );
  AND U5493 ( .A(n5313), .B(n5312), .Z(n5391) );
  XNOR U5494 ( .A(n5392), .B(n5391), .Z(n5393) );
  XOR U5495 ( .A(n5394), .B(n5393), .Z(n5326) );
  NANDN U5496 ( .A(n5315), .B(n5314), .Z(n5319) );
  NAND U5497 ( .A(n5317), .B(n5316), .Z(n5318) );
  AND U5498 ( .A(n5319), .B(n5318), .Z(n5325) );
  XNOR U5499 ( .A(n5326), .B(n5325), .Z(n5327) );
  XNOR U5500 ( .A(n5328), .B(n5327), .Z(n5397) );
  XNOR U5501 ( .A(sreg[188]), .B(n5397), .Z(n5399) );
  NANDN U5502 ( .A(sreg[187]), .B(n5320), .Z(n5324) );
  NAND U5503 ( .A(n5322), .B(n5321), .Z(n5323) );
  NAND U5504 ( .A(n5324), .B(n5323), .Z(n5398) );
  XNOR U5505 ( .A(n5399), .B(n5398), .Z(c[188]) );
  NANDN U5506 ( .A(n5326), .B(n5325), .Z(n5330) );
  NANDN U5507 ( .A(n5328), .B(n5327), .Z(n5329) );
  AND U5508 ( .A(n5330), .B(n5329), .Z(n5405) );
  NANDN U5509 ( .A(n5332), .B(n5331), .Z(n5336) );
  NAND U5510 ( .A(n5334), .B(n5333), .Z(n5335) );
  AND U5511 ( .A(n5336), .B(n5335), .Z(n5471) );
  NAND U5512 ( .A(n5337), .B(n9883), .Z(n5339) );
  XOR U5513 ( .A(b[11]), .B(a[67]), .Z(n5441) );
  NANDN U5514 ( .A(n9856), .B(n5441), .Z(n5338) );
  AND U5515 ( .A(n5339), .B(n5338), .Z(n5452) );
  NANDN U5516 ( .A(n10005), .B(n5340), .Z(n5342) );
  XOR U5517 ( .A(b[15]), .B(a[63]), .Z(n5444) );
  NANDN U5518 ( .A(n10006), .B(n5444), .Z(n5341) );
  AND U5519 ( .A(n5342), .B(n5341), .Z(n5451) );
  NANDN U5520 ( .A(n9685), .B(n5343), .Z(n5345) );
  XOR U5521 ( .A(b[9]), .B(a[69]), .Z(n5447) );
  NANDN U5522 ( .A(n9758), .B(n5447), .Z(n5344) );
  NAND U5523 ( .A(n5345), .B(n5344), .Z(n5450) );
  XOR U5524 ( .A(n5451), .B(n5450), .Z(n5453) );
  XOR U5525 ( .A(n5452), .B(n5453), .Z(n5463) );
  NANDN U5526 ( .A(n5347), .B(n5346), .Z(n5351) );
  OR U5527 ( .A(n5349), .B(n5348), .Z(n5350) );
  AND U5528 ( .A(n5351), .B(n5350), .Z(n5462) );
  XNOR U5529 ( .A(n5463), .B(n5462), .Z(n5464) );
  NANDN U5530 ( .A(n5353), .B(n5352), .Z(n5357) );
  NANDN U5531 ( .A(n5355), .B(n5354), .Z(n5356) );
  NAND U5532 ( .A(n5357), .B(n5356), .Z(n5465) );
  XNOR U5533 ( .A(n5464), .B(n5465), .Z(n5411) );
  NANDN U5534 ( .A(n5359), .B(n5358), .Z(n5363) );
  NANDN U5535 ( .A(n5361), .B(n5360), .Z(n5362) );
  AND U5536 ( .A(n5363), .B(n5362), .Z(n5437) );
  NAND U5537 ( .A(b[0]), .B(a[77]), .Z(n5364) );
  XNOR U5538 ( .A(b[1]), .B(n5364), .Z(n5366) );
  NANDN U5539 ( .A(b[0]), .B(a[76]), .Z(n5365) );
  NAND U5540 ( .A(n5366), .B(n5365), .Z(n5417) );
  NANDN U5541 ( .A(n9891), .B(n5367), .Z(n5369) );
  XOR U5542 ( .A(b[13]), .B(a[65]), .Z(n5423) );
  NANDN U5543 ( .A(n9935), .B(n5423), .Z(n5368) );
  AND U5544 ( .A(n5369), .B(n5368), .Z(n5415) );
  AND U5545 ( .A(b[15]), .B(a[61]), .Z(n5414) );
  XNOR U5546 ( .A(n5415), .B(n5414), .Z(n5416) );
  XNOR U5547 ( .A(n5417), .B(n5416), .Z(n5435) );
  NANDN U5548 ( .A(n9437), .B(n5370), .Z(n5372) );
  XOR U5549 ( .A(b[5]), .B(a[73]), .Z(n5426) );
  NANDN U5550 ( .A(n9503), .B(n5426), .Z(n5371) );
  AND U5551 ( .A(n5372), .B(n5371), .Z(n5459) );
  NANDN U5552 ( .A(n9588), .B(n5373), .Z(n5375) );
  XOR U5553 ( .A(b[7]), .B(a[71]), .Z(n5429) );
  NANDN U5554 ( .A(n9639), .B(n5429), .Z(n5374) );
  AND U5555 ( .A(n5375), .B(n5374), .Z(n5457) );
  NANDN U5556 ( .A(n9374), .B(n5376), .Z(n5378) );
  XOR U5557 ( .A(b[3]), .B(a[75]), .Z(n5432) );
  NANDN U5558 ( .A(n9375), .B(n5432), .Z(n5377) );
  NAND U5559 ( .A(n5378), .B(n5377), .Z(n5456) );
  XNOR U5560 ( .A(n5457), .B(n5456), .Z(n5458) );
  XOR U5561 ( .A(n5459), .B(n5458), .Z(n5436) );
  XOR U5562 ( .A(n5435), .B(n5436), .Z(n5438) );
  XOR U5563 ( .A(n5437), .B(n5438), .Z(n5409) );
  NANDN U5564 ( .A(n5380), .B(n5379), .Z(n5384) );
  OR U5565 ( .A(n5382), .B(n5381), .Z(n5383) );
  AND U5566 ( .A(n5384), .B(n5383), .Z(n5408) );
  XNOR U5567 ( .A(n5409), .B(n5408), .Z(n5410) );
  XOR U5568 ( .A(n5411), .B(n5410), .Z(n5469) );
  NANDN U5569 ( .A(n5386), .B(n5385), .Z(n5390) );
  NANDN U5570 ( .A(n5388), .B(n5387), .Z(n5389) );
  AND U5571 ( .A(n5390), .B(n5389), .Z(n5468) );
  XNOR U5572 ( .A(n5469), .B(n5468), .Z(n5470) );
  XOR U5573 ( .A(n5471), .B(n5470), .Z(n5403) );
  NANDN U5574 ( .A(n5392), .B(n5391), .Z(n5396) );
  NAND U5575 ( .A(n5394), .B(n5393), .Z(n5395) );
  AND U5576 ( .A(n5396), .B(n5395), .Z(n5402) );
  XNOR U5577 ( .A(n5403), .B(n5402), .Z(n5404) );
  XNOR U5578 ( .A(n5405), .B(n5404), .Z(n5474) );
  XNOR U5579 ( .A(sreg[189]), .B(n5474), .Z(n5476) );
  NANDN U5580 ( .A(sreg[188]), .B(n5397), .Z(n5401) );
  NAND U5581 ( .A(n5399), .B(n5398), .Z(n5400) );
  NAND U5582 ( .A(n5401), .B(n5400), .Z(n5475) );
  XNOR U5583 ( .A(n5476), .B(n5475), .Z(c[189]) );
  NANDN U5584 ( .A(n5403), .B(n5402), .Z(n5407) );
  NANDN U5585 ( .A(n5405), .B(n5404), .Z(n5406) );
  AND U5586 ( .A(n5407), .B(n5406), .Z(n5482) );
  NANDN U5587 ( .A(n5409), .B(n5408), .Z(n5413) );
  NAND U5588 ( .A(n5411), .B(n5410), .Z(n5412) );
  AND U5589 ( .A(n5413), .B(n5412), .Z(n5548) );
  NANDN U5590 ( .A(n5415), .B(n5414), .Z(n5419) );
  NANDN U5591 ( .A(n5417), .B(n5416), .Z(n5418) );
  AND U5592 ( .A(n5419), .B(n5418), .Z(n5514) );
  NAND U5593 ( .A(b[0]), .B(a[78]), .Z(n5420) );
  XNOR U5594 ( .A(b[1]), .B(n5420), .Z(n5422) );
  NANDN U5595 ( .A(b[0]), .B(a[77]), .Z(n5421) );
  NAND U5596 ( .A(n5422), .B(n5421), .Z(n5494) );
  NANDN U5597 ( .A(n9891), .B(n5423), .Z(n5425) );
  XOR U5598 ( .A(b[13]), .B(a[66]), .Z(n5500) );
  NANDN U5599 ( .A(n9935), .B(n5500), .Z(n5424) );
  AND U5600 ( .A(n5425), .B(n5424), .Z(n5492) );
  AND U5601 ( .A(b[15]), .B(a[62]), .Z(n5491) );
  XNOR U5602 ( .A(n5492), .B(n5491), .Z(n5493) );
  XNOR U5603 ( .A(n5494), .B(n5493), .Z(n5512) );
  NANDN U5604 ( .A(n9437), .B(n5426), .Z(n5428) );
  XOR U5605 ( .A(b[5]), .B(a[74]), .Z(n5503) );
  NANDN U5606 ( .A(n9503), .B(n5503), .Z(n5427) );
  AND U5607 ( .A(n5428), .B(n5427), .Z(n5536) );
  NANDN U5608 ( .A(n9588), .B(n5429), .Z(n5431) );
  XOR U5609 ( .A(b[7]), .B(a[72]), .Z(n5506) );
  NANDN U5610 ( .A(n9639), .B(n5506), .Z(n5430) );
  AND U5611 ( .A(n5431), .B(n5430), .Z(n5534) );
  NANDN U5612 ( .A(n9374), .B(n5432), .Z(n5434) );
  XOR U5613 ( .A(b[3]), .B(a[76]), .Z(n5509) );
  NANDN U5614 ( .A(n9375), .B(n5509), .Z(n5433) );
  NAND U5615 ( .A(n5434), .B(n5433), .Z(n5533) );
  XNOR U5616 ( .A(n5534), .B(n5533), .Z(n5535) );
  XOR U5617 ( .A(n5536), .B(n5535), .Z(n5513) );
  XOR U5618 ( .A(n5512), .B(n5513), .Z(n5515) );
  XOR U5619 ( .A(n5514), .B(n5515), .Z(n5486) );
  NANDN U5620 ( .A(n5436), .B(n5435), .Z(n5440) );
  OR U5621 ( .A(n5438), .B(n5437), .Z(n5439) );
  AND U5622 ( .A(n5440), .B(n5439), .Z(n5485) );
  XNOR U5623 ( .A(n5486), .B(n5485), .Z(n5488) );
  NAND U5624 ( .A(n5441), .B(n9883), .Z(n5443) );
  XOR U5625 ( .A(b[11]), .B(a[68]), .Z(n5518) );
  NANDN U5626 ( .A(n9856), .B(n5518), .Z(n5442) );
  AND U5627 ( .A(n5443), .B(n5442), .Z(n5529) );
  NANDN U5628 ( .A(n10005), .B(n5444), .Z(n5446) );
  XOR U5629 ( .A(b[15]), .B(a[64]), .Z(n5521) );
  NANDN U5630 ( .A(n10006), .B(n5521), .Z(n5445) );
  AND U5631 ( .A(n5446), .B(n5445), .Z(n5528) );
  NANDN U5632 ( .A(n9685), .B(n5447), .Z(n5449) );
  XOR U5633 ( .A(b[9]), .B(a[70]), .Z(n5524) );
  NANDN U5634 ( .A(n9758), .B(n5524), .Z(n5448) );
  NAND U5635 ( .A(n5449), .B(n5448), .Z(n5527) );
  XOR U5636 ( .A(n5528), .B(n5527), .Z(n5530) );
  XOR U5637 ( .A(n5529), .B(n5530), .Z(n5540) );
  NANDN U5638 ( .A(n5451), .B(n5450), .Z(n5455) );
  OR U5639 ( .A(n5453), .B(n5452), .Z(n5454) );
  AND U5640 ( .A(n5455), .B(n5454), .Z(n5539) );
  XNOR U5641 ( .A(n5540), .B(n5539), .Z(n5541) );
  NANDN U5642 ( .A(n5457), .B(n5456), .Z(n5461) );
  NANDN U5643 ( .A(n5459), .B(n5458), .Z(n5460) );
  NAND U5644 ( .A(n5461), .B(n5460), .Z(n5542) );
  XNOR U5645 ( .A(n5541), .B(n5542), .Z(n5487) );
  XOR U5646 ( .A(n5488), .B(n5487), .Z(n5546) );
  NANDN U5647 ( .A(n5463), .B(n5462), .Z(n5467) );
  NANDN U5648 ( .A(n5465), .B(n5464), .Z(n5466) );
  AND U5649 ( .A(n5467), .B(n5466), .Z(n5545) );
  XNOR U5650 ( .A(n5546), .B(n5545), .Z(n5547) );
  XOR U5651 ( .A(n5548), .B(n5547), .Z(n5480) );
  NANDN U5652 ( .A(n5469), .B(n5468), .Z(n5473) );
  NAND U5653 ( .A(n5471), .B(n5470), .Z(n5472) );
  AND U5654 ( .A(n5473), .B(n5472), .Z(n5479) );
  XNOR U5655 ( .A(n5480), .B(n5479), .Z(n5481) );
  XNOR U5656 ( .A(n5482), .B(n5481), .Z(n5551) );
  XNOR U5657 ( .A(sreg[190]), .B(n5551), .Z(n5553) );
  NANDN U5658 ( .A(sreg[189]), .B(n5474), .Z(n5478) );
  NAND U5659 ( .A(n5476), .B(n5475), .Z(n5477) );
  NAND U5660 ( .A(n5478), .B(n5477), .Z(n5552) );
  XNOR U5661 ( .A(n5553), .B(n5552), .Z(c[190]) );
  NANDN U5662 ( .A(n5480), .B(n5479), .Z(n5484) );
  NANDN U5663 ( .A(n5482), .B(n5481), .Z(n5483) );
  AND U5664 ( .A(n5484), .B(n5483), .Z(n5559) );
  NANDN U5665 ( .A(n5486), .B(n5485), .Z(n5490) );
  NAND U5666 ( .A(n5488), .B(n5487), .Z(n5489) );
  AND U5667 ( .A(n5490), .B(n5489), .Z(n5625) );
  NANDN U5668 ( .A(n5492), .B(n5491), .Z(n5496) );
  NANDN U5669 ( .A(n5494), .B(n5493), .Z(n5495) );
  AND U5670 ( .A(n5496), .B(n5495), .Z(n5591) );
  NAND U5671 ( .A(b[0]), .B(a[79]), .Z(n5497) );
  XNOR U5672 ( .A(b[1]), .B(n5497), .Z(n5499) );
  NANDN U5673 ( .A(b[0]), .B(a[78]), .Z(n5498) );
  NAND U5674 ( .A(n5499), .B(n5498), .Z(n5571) );
  NANDN U5675 ( .A(n9891), .B(n5500), .Z(n5502) );
  XOR U5676 ( .A(b[13]), .B(a[67]), .Z(n5574) );
  NANDN U5677 ( .A(n9935), .B(n5574), .Z(n5501) );
  AND U5678 ( .A(n5502), .B(n5501), .Z(n5569) );
  AND U5679 ( .A(b[15]), .B(a[63]), .Z(n5568) );
  XNOR U5680 ( .A(n5569), .B(n5568), .Z(n5570) );
  XNOR U5681 ( .A(n5571), .B(n5570), .Z(n5589) );
  NANDN U5682 ( .A(n9437), .B(n5503), .Z(n5505) );
  XOR U5683 ( .A(b[5]), .B(a[75]), .Z(n5580) );
  NANDN U5684 ( .A(n9503), .B(n5580), .Z(n5504) );
  AND U5685 ( .A(n5505), .B(n5504), .Z(n5613) );
  NANDN U5686 ( .A(n9588), .B(n5506), .Z(n5508) );
  XOR U5687 ( .A(b[7]), .B(a[73]), .Z(n5583) );
  NANDN U5688 ( .A(n9639), .B(n5583), .Z(n5507) );
  AND U5689 ( .A(n5508), .B(n5507), .Z(n5611) );
  NANDN U5690 ( .A(n9374), .B(n5509), .Z(n5511) );
  XOR U5691 ( .A(b[3]), .B(a[77]), .Z(n5586) );
  NANDN U5692 ( .A(n9375), .B(n5586), .Z(n5510) );
  NAND U5693 ( .A(n5511), .B(n5510), .Z(n5610) );
  XNOR U5694 ( .A(n5611), .B(n5610), .Z(n5612) );
  XOR U5695 ( .A(n5613), .B(n5612), .Z(n5590) );
  XOR U5696 ( .A(n5589), .B(n5590), .Z(n5592) );
  XOR U5697 ( .A(n5591), .B(n5592), .Z(n5563) );
  NANDN U5698 ( .A(n5513), .B(n5512), .Z(n5517) );
  OR U5699 ( .A(n5515), .B(n5514), .Z(n5516) );
  AND U5700 ( .A(n5517), .B(n5516), .Z(n5562) );
  XNOR U5701 ( .A(n5563), .B(n5562), .Z(n5565) );
  NAND U5702 ( .A(n5518), .B(n9883), .Z(n5520) );
  XOR U5703 ( .A(b[11]), .B(a[69]), .Z(n5595) );
  NANDN U5704 ( .A(n9856), .B(n5595), .Z(n5519) );
  AND U5705 ( .A(n5520), .B(n5519), .Z(n5606) );
  NANDN U5706 ( .A(n10005), .B(n5521), .Z(n5523) );
  XOR U5707 ( .A(b[15]), .B(a[65]), .Z(n5598) );
  NANDN U5708 ( .A(n10006), .B(n5598), .Z(n5522) );
  AND U5709 ( .A(n5523), .B(n5522), .Z(n5605) );
  NANDN U5710 ( .A(n9685), .B(n5524), .Z(n5526) );
  XOR U5711 ( .A(b[9]), .B(a[71]), .Z(n5601) );
  NANDN U5712 ( .A(n9758), .B(n5601), .Z(n5525) );
  NAND U5713 ( .A(n5526), .B(n5525), .Z(n5604) );
  XOR U5714 ( .A(n5605), .B(n5604), .Z(n5607) );
  XOR U5715 ( .A(n5606), .B(n5607), .Z(n5617) );
  NANDN U5716 ( .A(n5528), .B(n5527), .Z(n5532) );
  OR U5717 ( .A(n5530), .B(n5529), .Z(n5531) );
  AND U5718 ( .A(n5532), .B(n5531), .Z(n5616) );
  XNOR U5719 ( .A(n5617), .B(n5616), .Z(n5618) );
  NANDN U5720 ( .A(n5534), .B(n5533), .Z(n5538) );
  NANDN U5721 ( .A(n5536), .B(n5535), .Z(n5537) );
  NAND U5722 ( .A(n5538), .B(n5537), .Z(n5619) );
  XNOR U5723 ( .A(n5618), .B(n5619), .Z(n5564) );
  XOR U5724 ( .A(n5565), .B(n5564), .Z(n5623) );
  NANDN U5725 ( .A(n5540), .B(n5539), .Z(n5544) );
  NANDN U5726 ( .A(n5542), .B(n5541), .Z(n5543) );
  AND U5727 ( .A(n5544), .B(n5543), .Z(n5622) );
  XNOR U5728 ( .A(n5623), .B(n5622), .Z(n5624) );
  XOR U5729 ( .A(n5625), .B(n5624), .Z(n5557) );
  NANDN U5730 ( .A(n5546), .B(n5545), .Z(n5550) );
  NAND U5731 ( .A(n5548), .B(n5547), .Z(n5549) );
  AND U5732 ( .A(n5550), .B(n5549), .Z(n5556) );
  XNOR U5733 ( .A(n5557), .B(n5556), .Z(n5558) );
  XNOR U5734 ( .A(n5559), .B(n5558), .Z(n5628) );
  XNOR U5735 ( .A(sreg[191]), .B(n5628), .Z(n5630) );
  NANDN U5736 ( .A(sreg[190]), .B(n5551), .Z(n5555) );
  NAND U5737 ( .A(n5553), .B(n5552), .Z(n5554) );
  NAND U5738 ( .A(n5555), .B(n5554), .Z(n5629) );
  XNOR U5739 ( .A(n5630), .B(n5629), .Z(c[191]) );
  NANDN U5740 ( .A(n5557), .B(n5556), .Z(n5561) );
  NANDN U5741 ( .A(n5559), .B(n5558), .Z(n5560) );
  AND U5742 ( .A(n5561), .B(n5560), .Z(n5636) );
  NANDN U5743 ( .A(n5563), .B(n5562), .Z(n5567) );
  NAND U5744 ( .A(n5565), .B(n5564), .Z(n5566) );
  AND U5745 ( .A(n5567), .B(n5566), .Z(n5702) );
  NANDN U5746 ( .A(n5569), .B(n5568), .Z(n5573) );
  NANDN U5747 ( .A(n5571), .B(n5570), .Z(n5572) );
  AND U5748 ( .A(n5573), .B(n5572), .Z(n5668) );
  NANDN U5749 ( .A(n9891), .B(n5574), .Z(n5576) );
  XOR U5750 ( .A(b[13]), .B(a[68]), .Z(n5654) );
  NANDN U5751 ( .A(n9935), .B(n5654), .Z(n5575) );
  AND U5752 ( .A(n5576), .B(n5575), .Z(n5646) );
  AND U5753 ( .A(b[15]), .B(a[64]), .Z(n5645) );
  XNOR U5754 ( .A(n5646), .B(n5645), .Z(n5647) );
  NAND U5755 ( .A(b[0]), .B(a[80]), .Z(n5577) );
  XNOR U5756 ( .A(b[1]), .B(n5577), .Z(n5579) );
  NANDN U5757 ( .A(b[0]), .B(a[79]), .Z(n5578) );
  NAND U5758 ( .A(n5579), .B(n5578), .Z(n5648) );
  XNOR U5759 ( .A(n5647), .B(n5648), .Z(n5666) );
  NANDN U5760 ( .A(n9437), .B(n5580), .Z(n5582) );
  XOR U5761 ( .A(b[5]), .B(a[76]), .Z(n5657) );
  NANDN U5762 ( .A(n9503), .B(n5657), .Z(n5581) );
  AND U5763 ( .A(n5582), .B(n5581), .Z(n5690) );
  NANDN U5764 ( .A(n9588), .B(n5583), .Z(n5585) );
  XOR U5765 ( .A(b[7]), .B(a[74]), .Z(n5660) );
  NANDN U5766 ( .A(n9639), .B(n5660), .Z(n5584) );
  AND U5767 ( .A(n5585), .B(n5584), .Z(n5688) );
  NANDN U5768 ( .A(n9374), .B(n5586), .Z(n5588) );
  XOR U5769 ( .A(b[3]), .B(a[78]), .Z(n5663) );
  NANDN U5770 ( .A(n9375), .B(n5663), .Z(n5587) );
  NAND U5771 ( .A(n5588), .B(n5587), .Z(n5687) );
  XNOR U5772 ( .A(n5688), .B(n5687), .Z(n5689) );
  XOR U5773 ( .A(n5690), .B(n5689), .Z(n5667) );
  XOR U5774 ( .A(n5666), .B(n5667), .Z(n5669) );
  XOR U5775 ( .A(n5668), .B(n5669), .Z(n5640) );
  NANDN U5776 ( .A(n5590), .B(n5589), .Z(n5594) );
  OR U5777 ( .A(n5592), .B(n5591), .Z(n5593) );
  AND U5778 ( .A(n5594), .B(n5593), .Z(n5639) );
  XNOR U5779 ( .A(n5640), .B(n5639), .Z(n5642) );
  NAND U5780 ( .A(n5595), .B(n9883), .Z(n5597) );
  XOR U5781 ( .A(b[11]), .B(a[70]), .Z(n5672) );
  NANDN U5782 ( .A(n9856), .B(n5672), .Z(n5596) );
  AND U5783 ( .A(n5597), .B(n5596), .Z(n5683) );
  NANDN U5784 ( .A(n10005), .B(n5598), .Z(n5600) );
  XOR U5785 ( .A(b[15]), .B(a[66]), .Z(n5675) );
  NANDN U5786 ( .A(n10006), .B(n5675), .Z(n5599) );
  AND U5787 ( .A(n5600), .B(n5599), .Z(n5682) );
  NANDN U5788 ( .A(n9685), .B(n5601), .Z(n5603) );
  XOR U5789 ( .A(b[9]), .B(a[72]), .Z(n5678) );
  NANDN U5790 ( .A(n9758), .B(n5678), .Z(n5602) );
  NAND U5791 ( .A(n5603), .B(n5602), .Z(n5681) );
  XOR U5792 ( .A(n5682), .B(n5681), .Z(n5684) );
  XOR U5793 ( .A(n5683), .B(n5684), .Z(n5694) );
  NANDN U5794 ( .A(n5605), .B(n5604), .Z(n5609) );
  OR U5795 ( .A(n5607), .B(n5606), .Z(n5608) );
  AND U5796 ( .A(n5609), .B(n5608), .Z(n5693) );
  XNOR U5797 ( .A(n5694), .B(n5693), .Z(n5695) );
  NANDN U5798 ( .A(n5611), .B(n5610), .Z(n5615) );
  NANDN U5799 ( .A(n5613), .B(n5612), .Z(n5614) );
  NAND U5800 ( .A(n5615), .B(n5614), .Z(n5696) );
  XNOR U5801 ( .A(n5695), .B(n5696), .Z(n5641) );
  XOR U5802 ( .A(n5642), .B(n5641), .Z(n5700) );
  NANDN U5803 ( .A(n5617), .B(n5616), .Z(n5621) );
  NANDN U5804 ( .A(n5619), .B(n5618), .Z(n5620) );
  AND U5805 ( .A(n5621), .B(n5620), .Z(n5699) );
  XNOR U5806 ( .A(n5700), .B(n5699), .Z(n5701) );
  XOR U5807 ( .A(n5702), .B(n5701), .Z(n5634) );
  NANDN U5808 ( .A(n5623), .B(n5622), .Z(n5627) );
  NAND U5809 ( .A(n5625), .B(n5624), .Z(n5626) );
  AND U5810 ( .A(n5627), .B(n5626), .Z(n5633) );
  XNOR U5811 ( .A(n5634), .B(n5633), .Z(n5635) );
  XNOR U5812 ( .A(n5636), .B(n5635), .Z(n5705) );
  XNOR U5813 ( .A(sreg[192]), .B(n5705), .Z(n5707) );
  NANDN U5814 ( .A(sreg[191]), .B(n5628), .Z(n5632) );
  NAND U5815 ( .A(n5630), .B(n5629), .Z(n5631) );
  NAND U5816 ( .A(n5632), .B(n5631), .Z(n5706) );
  XNOR U5817 ( .A(n5707), .B(n5706), .Z(c[192]) );
  NANDN U5818 ( .A(n5634), .B(n5633), .Z(n5638) );
  NANDN U5819 ( .A(n5636), .B(n5635), .Z(n5637) );
  AND U5820 ( .A(n5638), .B(n5637), .Z(n5713) );
  NANDN U5821 ( .A(n5640), .B(n5639), .Z(n5644) );
  NAND U5822 ( .A(n5642), .B(n5641), .Z(n5643) );
  AND U5823 ( .A(n5644), .B(n5643), .Z(n5779) );
  NANDN U5824 ( .A(n5646), .B(n5645), .Z(n5650) );
  NANDN U5825 ( .A(n5648), .B(n5647), .Z(n5649) );
  AND U5826 ( .A(n5650), .B(n5649), .Z(n5745) );
  NAND U5827 ( .A(b[0]), .B(a[81]), .Z(n5651) );
  XNOR U5828 ( .A(b[1]), .B(n5651), .Z(n5653) );
  NANDN U5829 ( .A(b[0]), .B(a[80]), .Z(n5652) );
  NAND U5830 ( .A(n5653), .B(n5652), .Z(n5725) );
  NANDN U5831 ( .A(n9891), .B(n5654), .Z(n5656) );
  XOR U5832 ( .A(b[13]), .B(a[69]), .Z(n5731) );
  NANDN U5833 ( .A(n9935), .B(n5731), .Z(n5655) );
  AND U5834 ( .A(n5656), .B(n5655), .Z(n5723) );
  AND U5835 ( .A(b[15]), .B(a[65]), .Z(n5722) );
  XNOR U5836 ( .A(n5723), .B(n5722), .Z(n5724) );
  XNOR U5837 ( .A(n5725), .B(n5724), .Z(n5743) );
  NANDN U5838 ( .A(n9437), .B(n5657), .Z(n5659) );
  XOR U5839 ( .A(b[5]), .B(a[77]), .Z(n5734) );
  NANDN U5840 ( .A(n9503), .B(n5734), .Z(n5658) );
  AND U5841 ( .A(n5659), .B(n5658), .Z(n5767) );
  NANDN U5842 ( .A(n9588), .B(n5660), .Z(n5662) );
  XOR U5843 ( .A(b[7]), .B(a[75]), .Z(n5737) );
  NANDN U5844 ( .A(n9639), .B(n5737), .Z(n5661) );
  AND U5845 ( .A(n5662), .B(n5661), .Z(n5765) );
  NANDN U5846 ( .A(n9374), .B(n5663), .Z(n5665) );
  XOR U5847 ( .A(b[3]), .B(a[79]), .Z(n5740) );
  NANDN U5848 ( .A(n9375), .B(n5740), .Z(n5664) );
  NAND U5849 ( .A(n5665), .B(n5664), .Z(n5764) );
  XNOR U5850 ( .A(n5765), .B(n5764), .Z(n5766) );
  XOR U5851 ( .A(n5767), .B(n5766), .Z(n5744) );
  XOR U5852 ( .A(n5743), .B(n5744), .Z(n5746) );
  XOR U5853 ( .A(n5745), .B(n5746), .Z(n5717) );
  NANDN U5854 ( .A(n5667), .B(n5666), .Z(n5671) );
  OR U5855 ( .A(n5669), .B(n5668), .Z(n5670) );
  AND U5856 ( .A(n5671), .B(n5670), .Z(n5716) );
  XNOR U5857 ( .A(n5717), .B(n5716), .Z(n5719) );
  NAND U5858 ( .A(n5672), .B(n9883), .Z(n5674) );
  XOR U5859 ( .A(b[11]), .B(a[71]), .Z(n5749) );
  NANDN U5860 ( .A(n9856), .B(n5749), .Z(n5673) );
  AND U5861 ( .A(n5674), .B(n5673), .Z(n5760) );
  NANDN U5862 ( .A(n10005), .B(n5675), .Z(n5677) );
  XOR U5863 ( .A(b[15]), .B(a[67]), .Z(n5752) );
  NANDN U5864 ( .A(n10006), .B(n5752), .Z(n5676) );
  AND U5865 ( .A(n5677), .B(n5676), .Z(n5759) );
  NANDN U5866 ( .A(n9685), .B(n5678), .Z(n5680) );
  XOR U5867 ( .A(b[9]), .B(a[73]), .Z(n5755) );
  NANDN U5868 ( .A(n9758), .B(n5755), .Z(n5679) );
  NAND U5869 ( .A(n5680), .B(n5679), .Z(n5758) );
  XOR U5870 ( .A(n5759), .B(n5758), .Z(n5761) );
  XOR U5871 ( .A(n5760), .B(n5761), .Z(n5771) );
  NANDN U5872 ( .A(n5682), .B(n5681), .Z(n5686) );
  OR U5873 ( .A(n5684), .B(n5683), .Z(n5685) );
  AND U5874 ( .A(n5686), .B(n5685), .Z(n5770) );
  XNOR U5875 ( .A(n5771), .B(n5770), .Z(n5772) );
  NANDN U5876 ( .A(n5688), .B(n5687), .Z(n5692) );
  NANDN U5877 ( .A(n5690), .B(n5689), .Z(n5691) );
  NAND U5878 ( .A(n5692), .B(n5691), .Z(n5773) );
  XNOR U5879 ( .A(n5772), .B(n5773), .Z(n5718) );
  XOR U5880 ( .A(n5719), .B(n5718), .Z(n5777) );
  NANDN U5881 ( .A(n5694), .B(n5693), .Z(n5698) );
  NANDN U5882 ( .A(n5696), .B(n5695), .Z(n5697) );
  AND U5883 ( .A(n5698), .B(n5697), .Z(n5776) );
  XNOR U5884 ( .A(n5777), .B(n5776), .Z(n5778) );
  XOR U5885 ( .A(n5779), .B(n5778), .Z(n5711) );
  NANDN U5886 ( .A(n5700), .B(n5699), .Z(n5704) );
  NAND U5887 ( .A(n5702), .B(n5701), .Z(n5703) );
  AND U5888 ( .A(n5704), .B(n5703), .Z(n5710) );
  XNOR U5889 ( .A(n5711), .B(n5710), .Z(n5712) );
  XNOR U5890 ( .A(n5713), .B(n5712), .Z(n5782) );
  XNOR U5891 ( .A(sreg[193]), .B(n5782), .Z(n5784) );
  NANDN U5892 ( .A(sreg[192]), .B(n5705), .Z(n5709) );
  NAND U5893 ( .A(n5707), .B(n5706), .Z(n5708) );
  NAND U5894 ( .A(n5709), .B(n5708), .Z(n5783) );
  XNOR U5895 ( .A(n5784), .B(n5783), .Z(c[193]) );
  NANDN U5896 ( .A(n5711), .B(n5710), .Z(n5715) );
  NANDN U5897 ( .A(n5713), .B(n5712), .Z(n5714) );
  AND U5898 ( .A(n5715), .B(n5714), .Z(n5790) );
  NANDN U5899 ( .A(n5717), .B(n5716), .Z(n5721) );
  NAND U5900 ( .A(n5719), .B(n5718), .Z(n5720) );
  AND U5901 ( .A(n5721), .B(n5720), .Z(n5856) );
  NANDN U5902 ( .A(n5723), .B(n5722), .Z(n5727) );
  NANDN U5903 ( .A(n5725), .B(n5724), .Z(n5726) );
  AND U5904 ( .A(n5727), .B(n5726), .Z(n5822) );
  NAND U5905 ( .A(b[0]), .B(a[82]), .Z(n5728) );
  XNOR U5906 ( .A(b[1]), .B(n5728), .Z(n5730) );
  NANDN U5907 ( .A(b[0]), .B(a[81]), .Z(n5729) );
  NAND U5908 ( .A(n5730), .B(n5729), .Z(n5802) );
  NANDN U5909 ( .A(n9891), .B(n5731), .Z(n5733) );
  XOR U5910 ( .A(b[13]), .B(a[70]), .Z(n5808) );
  NANDN U5911 ( .A(n9935), .B(n5808), .Z(n5732) );
  AND U5912 ( .A(n5733), .B(n5732), .Z(n5800) );
  AND U5913 ( .A(b[15]), .B(a[66]), .Z(n5799) );
  XNOR U5914 ( .A(n5800), .B(n5799), .Z(n5801) );
  XNOR U5915 ( .A(n5802), .B(n5801), .Z(n5820) );
  NANDN U5916 ( .A(n9437), .B(n5734), .Z(n5736) );
  XOR U5917 ( .A(b[5]), .B(a[78]), .Z(n5811) );
  NANDN U5918 ( .A(n9503), .B(n5811), .Z(n5735) );
  AND U5919 ( .A(n5736), .B(n5735), .Z(n5844) );
  NANDN U5920 ( .A(n9588), .B(n5737), .Z(n5739) );
  XOR U5921 ( .A(b[7]), .B(a[76]), .Z(n5814) );
  NANDN U5922 ( .A(n9639), .B(n5814), .Z(n5738) );
  AND U5923 ( .A(n5739), .B(n5738), .Z(n5842) );
  NANDN U5924 ( .A(n9374), .B(n5740), .Z(n5742) );
  XOR U5925 ( .A(b[3]), .B(a[80]), .Z(n5817) );
  NANDN U5926 ( .A(n9375), .B(n5817), .Z(n5741) );
  NAND U5927 ( .A(n5742), .B(n5741), .Z(n5841) );
  XNOR U5928 ( .A(n5842), .B(n5841), .Z(n5843) );
  XOR U5929 ( .A(n5844), .B(n5843), .Z(n5821) );
  XOR U5930 ( .A(n5820), .B(n5821), .Z(n5823) );
  XOR U5931 ( .A(n5822), .B(n5823), .Z(n5794) );
  NANDN U5932 ( .A(n5744), .B(n5743), .Z(n5748) );
  OR U5933 ( .A(n5746), .B(n5745), .Z(n5747) );
  AND U5934 ( .A(n5748), .B(n5747), .Z(n5793) );
  XNOR U5935 ( .A(n5794), .B(n5793), .Z(n5796) );
  NAND U5936 ( .A(n5749), .B(n9883), .Z(n5751) );
  XOR U5937 ( .A(b[11]), .B(a[72]), .Z(n5826) );
  NANDN U5938 ( .A(n9856), .B(n5826), .Z(n5750) );
  AND U5939 ( .A(n5751), .B(n5750), .Z(n5837) );
  NANDN U5940 ( .A(n10005), .B(n5752), .Z(n5754) );
  XOR U5941 ( .A(b[15]), .B(a[68]), .Z(n5829) );
  NANDN U5942 ( .A(n10006), .B(n5829), .Z(n5753) );
  AND U5943 ( .A(n5754), .B(n5753), .Z(n5836) );
  NANDN U5944 ( .A(n9685), .B(n5755), .Z(n5757) );
  XOR U5945 ( .A(b[9]), .B(a[74]), .Z(n5832) );
  NANDN U5946 ( .A(n9758), .B(n5832), .Z(n5756) );
  NAND U5947 ( .A(n5757), .B(n5756), .Z(n5835) );
  XOR U5948 ( .A(n5836), .B(n5835), .Z(n5838) );
  XOR U5949 ( .A(n5837), .B(n5838), .Z(n5848) );
  NANDN U5950 ( .A(n5759), .B(n5758), .Z(n5763) );
  OR U5951 ( .A(n5761), .B(n5760), .Z(n5762) );
  AND U5952 ( .A(n5763), .B(n5762), .Z(n5847) );
  XNOR U5953 ( .A(n5848), .B(n5847), .Z(n5849) );
  NANDN U5954 ( .A(n5765), .B(n5764), .Z(n5769) );
  NANDN U5955 ( .A(n5767), .B(n5766), .Z(n5768) );
  NAND U5956 ( .A(n5769), .B(n5768), .Z(n5850) );
  XNOR U5957 ( .A(n5849), .B(n5850), .Z(n5795) );
  XOR U5958 ( .A(n5796), .B(n5795), .Z(n5854) );
  NANDN U5959 ( .A(n5771), .B(n5770), .Z(n5775) );
  NANDN U5960 ( .A(n5773), .B(n5772), .Z(n5774) );
  AND U5961 ( .A(n5775), .B(n5774), .Z(n5853) );
  XNOR U5962 ( .A(n5854), .B(n5853), .Z(n5855) );
  XOR U5963 ( .A(n5856), .B(n5855), .Z(n5788) );
  NANDN U5964 ( .A(n5777), .B(n5776), .Z(n5781) );
  NAND U5965 ( .A(n5779), .B(n5778), .Z(n5780) );
  AND U5966 ( .A(n5781), .B(n5780), .Z(n5787) );
  XNOR U5967 ( .A(n5788), .B(n5787), .Z(n5789) );
  XNOR U5968 ( .A(n5790), .B(n5789), .Z(n5859) );
  XNOR U5969 ( .A(sreg[194]), .B(n5859), .Z(n5861) );
  NANDN U5970 ( .A(sreg[193]), .B(n5782), .Z(n5786) );
  NAND U5971 ( .A(n5784), .B(n5783), .Z(n5785) );
  NAND U5972 ( .A(n5786), .B(n5785), .Z(n5860) );
  XNOR U5973 ( .A(n5861), .B(n5860), .Z(c[194]) );
  NANDN U5974 ( .A(n5788), .B(n5787), .Z(n5792) );
  NANDN U5975 ( .A(n5790), .B(n5789), .Z(n5791) );
  AND U5976 ( .A(n5792), .B(n5791), .Z(n5867) );
  NANDN U5977 ( .A(n5794), .B(n5793), .Z(n5798) );
  NAND U5978 ( .A(n5796), .B(n5795), .Z(n5797) );
  AND U5979 ( .A(n5798), .B(n5797), .Z(n5933) );
  NANDN U5980 ( .A(n5800), .B(n5799), .Z(n5804) );
  NANDN U5981 ( .A(n5802), .B(n5801), .Z(n5803) );
  AND U5982 ( .A(n5804), .B(n5803), .Z(n5899) );
  NAND U5983 ( .A(b[0]), .B(a[83]), .Z(n5805) );
  XNOR U5984 ( .A(b[1]), .B(n5805), .Z(n5807) );
  NANDN U5985 ( .A(b[0]), .B(a[82]), .Z(n5806) );
  NAND U5986 ( .A(n5807), .B(n5806), .Z(n5879) );
  NANDN U5987 ( .A(n9891), .B(n5808), .Z(n5810) );
  XOR U5988 ( .A(b[13]), .B(a[71]), .Z(n5882) );
  NANDN U5989 ( .A(n9935), .B(n5882), .Z(n5809) );
  AND U5990 ( .A(n5810), .B(n5809), .Z(n5877) );
  AND U5991 ( .A(b[15]), .B(a[67]), .Z(n5876) );
  XNOR U5992 ( .A(n5877), .B(n5876), .Z(n5878) );
  XNOR U5993 ( .A(n5879), .B(n5878), .Z(n5897) );
  NANDN U5994 ( .A(n9437), .B(n5811), .Z(n5813) );
  XOR U5995 ( .A(b[5]), .B(a[79]), .Z(n5888) );
  NANDN U5996 ( .A(n9503), .B(n5888), .Z(n5812) );
  AND U5997 ( .A(n5813), .B(n5812), .Z(n5921) );
  NANDN U5998 ( .A(n9588), .B(n5814), .Z(n5816) );
  XOR U5999 ( .A(b[7]), .B(a[77]), .Z(n5891) );
  NANDN U6000 ( .A(n9639), .B(n5891), .Z(n5815) );
  AND U6001 ( .A(n5816), .B(n5815), .Z(n5919) );
  NANDN U6002 ( .A(n9374), .B(n5817), .Z(n5819) );
  XOR U6003 ( .A(b[3]), .B(a[81]), .Z(n5894) );
  NANDN U6004 ( .A(n9375), .B(n5894), .Z(n5818) );
  NAND U6005 ( .A(n5819), .B(n5818), .Z(n5918) );
  XNOR U6006 ( .A(n5919), .B(n5918), .Z(n5920) );
  XOR U6007 ( .A(n5921), .B(n5920), .Z(n5898) );
  XOR U6008 ( .A(n5897), .B(n5898), .Z(n5900) );
  XOR U6009 ( .A(n5899), .B(n5900), .Z(n5871) );
  NANDN U6010 ( .A(n5821), .B(n5820), .Z(n5825) );
  OR U6011 ( .A(n5823), .B(n5822), .Z(n5824) );
  AND U6012 ( .A(n5825), .B(n5824), .Z(n5870) );
  XNOR U6013 ( .A(n5871), .B(n5870), .Z(n5873) );
  NAND U6014 ( .A(n5826), .B(n9883), .Z(n5828) );
  XOR U6015 ( .A(b[11]), .B(a[73]), .Z(n5903) );
  NANDN U6016 ( .A(n9856), .B(n5903), .Z(n5827) );
  AND U6017 ( .A(n5828), .B(n5827), .Z(n5914) );
  NANDN U6018 ( .A(n10005), .B(n5829), .Z(n5831) );
  XOR U6019 ( .A(b[15]), .B(a[69]), .Z(n5906) );
  NANDN U6020 ( .A(n10006), .B(n5906), .Z(n5830) );
  AND U6021 ( .A(n5831), .B(n5830), .Z(n5913) );
  NANDN U6022 ( .A(n9685), .B(n5832), .Z(n5834) );
  XOR U6023 ( .A(b[9]), .B(a[75]), .Z(n5909) );
  NANDN U6024 ( .A(n9758), .B(n5909), .Z(n5833) );
  NAND U6025 ( .A(n5834), .B(n5833), .Z(n5912) );
  XOR U6026 ( .A(n5913), .B(n5912), .Z(n5915) );
  XOR U6027 ( .A(n5914), .B(n5915), .Z(n5925) );
  NANDN U6028 ( .A(n5836), .B(n5835), .Z(n5840) );
  OR U6029 ( .A(n5838), .B(n5837), .Z(n5839) );
  AND U6030 ( .A(n5840), .B(n5839), .Z(n5924) );
  XNOR U6031 ( .A(n5925), .B(n5924), .Z(n5926) );
  NANDN U6032 ( .A(n5842), .B(n5841), .Z(n5846) );
  NANDN U6033 ( .A(n5844), .B(n5843), .Z(n5845) );
  NAND U6034 ( .A(n5846), .B(n5845), .Z(n5927) );
  XNOR U6035 ( .A(n5926), .B(n5927), .Z(n5872) );
  XOR U6036 ( .A(n5873), .B(n5872), .Z(n5931) );
  NANDN U6037 ( .A(n5848), .B(n5847), .Z(n5852) );
  NANDN U6038 ( .A(n5850), .B(n5849), .Z(n5851) );
  AND U6039 ( .A(n5852), .B(n5851), .Z(n5930) );
  XNOR U6040 ( .A(n5931), .B(n5930), .Z(n5932) );
  XOR U6041 ( .A(n5933), .B(n5932), .Z(n5865) );
  NANDN U6042 ( .A(n5854), .B(n5853), .Z(n5858) );
  NAND U6043 ( .A(n5856), .B(n5855), .Z(n5857) );
  AND U6044 ( .A(n5858), .B(n5857), .Z(n5864) );
  XNOR U6045 ( .A(n5865), .B(n5864), .Z(n5866) );
  XNOR U6046 ( .A(n5867), .B(n5866), .Z(n5936) );
  XNOR U6047 ( .A(sreg[195]), .B(n5936), .Z(n5938) );
  NANDN U6048 ( .A(sreg[194]), .B(n5859), .Z(n5863) );
  NAND U6049 ( .A(n5861), .B(n5860), .Z(n5862) );
  NAND U6050 ( .A(n5863), .B(n5862), .Z(n5937) );
  XNOR U6051 ( .A(n5938), .B(n5937), .Z(c[195]) );
  NANDN U6052 ( .A(n5865), .B(n5864), .Z(n5869) );
  NANDN U6053 ( .A(n5867), .B(n5866), .Z(n5868) );
  AND U6054 ( .A(n5869), .B(n5868), .Z(n5944) );
  NANDN U6055 ( .A(n5871), .B(n5870), .Z(n5875) );
  NAND U6056 ( .A(n5873), .B(n5872), .Z(n5874) );
  AND U6057 ( .A(n5875), .B(n5874), .Z(n6010) );
  NANDN U6058 ( .A(n5877), .B(n5876), .Z(n5881) );
  NANDN U6059 ( .A(n5879), .B(n5878), .Z(n5880) );
  AND U6060 ( .A(n5881), .B(n5880), .Z(n5997) );
  NANDN U6061 ( .A(n9891), .B(n5882), .Z(n5884) );
  XOR U6062 ( .A(b[13]), .B(a[72]), .Z(n5983) );
  NANDN U6063 ( .A(n9935), .B(n5983), .Z(n5883) );
  AND U6064 ( .A(n5884), .B(n5883), .Z(n5975) );
  AND U6065 ( .A(b[15]), .B(a[68]), .Z(n5974) );
  XNOR U6066 ( .A(n5975), .B(n5974), .Z(n5976) );
  NAND U6067 ( .A(b[0]), .B(a[84]), .Z(n5885) );
  XNOR U6068 ( .A(b[1]), .B(n5885), .Z(n5887) );
  NANDN U6069 ( .A(b[0]), .B(a[83]), .Z(n5886) );
  NAND U6070 ( .A(n5887), .B(n5886), .Z(n5977) );
  XNOR U6071 ( .A(n5976), .B(n5977), .Z(n5995) );
  NANDN U6072 ( .A(n9437), .B(n5888), .Z(n5890) );
  XOR U6073 ( .A(b[5]), .B(a[80]), .Z(n5986) );
  NANDN U6074 ( .A(n9503), .B(n5986), .Z(n5889) );
  AND U6075 ( .A(n5890), .B(n5889), .Z(n5971) );
  NANDN U6076 ( .A(n9588), .B(n5891), .Z(n5893) );
  XOR U6077 ( .A(b[7]), .B(a[78]), .Z(n5989) );
  NANDN U6078 ( .A(n9639), .B(n5989), .Z(n5892) );
  AND U6079 ( .A(n5893), .B(n5892), .Z(n5969) );
  NANDN U6080 ( .A(n9374), .B(n5894), .Z(n5896) );
  XOR U6081 ( .A(b[3]), .B(a[82]), .Z(n5992) );
  NANDN U6082 ( .A(n9375), .B(n5992), .Z(n5895) );
  NAND U6083 ( .A(n5896), .B(n5895), .Z(n5968) );
  XNOR U6084 ( .A(n5969), .B(n5968), .Z(n5970) );
  XOR U6085 ( .A(n5971), .B(n5970), .Z(n5996) );
  XOR U6086 ( .A(n5995), .B(n5996), .Z(n5998) );
  XOR U6087 ( .A(n5997), .B(n5998), .Z(n5948) );
  NANDN U6088 ( .A(n5898), .B(n5897), .Z(n5902) );
  OR U6089 ( .A(n5900), .B(n5899), .Z(n5901) );
  AND U6090 ( .A(n5902), .B(n5901), .Z(n5947) );
  XNOR U6091 ( .A(n5948), .B(n5947), .Z(n5950) );
  NAND U6092 ( .A(n5903), .B(n9883), .Z(n5905) );
  XOR U6093 ( .A(b[11]), .B(a[74]), .Z(n5953) );
  NANDN U6094 ( .A(n9856), .B(n5953), .Z(n5904) );
  AND U6095 ( .A(n5905), .B(n5904), .Z(n5964) );
  NANDN U6096 ( .A(n10005), .B(n5906), .Z(n5908) );
  XOR U6097 ( .A(b[15]), .B(a[70]), .Z(n5956) );
  NANDN U6098 ( .A(n10006), .B(n5956), .Z(n5907) );
  AND U6099 ( .A(n5908), .B(n5907), .Z(n5963) );
  NANDN U6100 ( .A(n9685), .B(n5909), .Z(n5911) );
  XOR U6101 ( .A(b[9]), .B(a[76]), .Z(n5959) );
  NANDN U6102 ( .A(n9758), .B(n5959), .Z(n5910) );
  NAND U6103 ( .A(n5911), .B(n5910), .Z(n5962) );
  XOR U6104 ( .A(n5963), .B(n5962), .Z(n5965) );
  XOR U6105 ( .A(n5964), .B(n5965), .Z(n6002) );
  NANDN U6106 ( .A(n5913), .B(n5912), .Z(n5917) );
  OR U6107 ( .A(n5915), .B(n5914), .Z(n5916) );
  AND U6108 ( .A(n5917), .B(n5916), .Z(n6001) );
  XNOR U6109 ( .A(n6002), .B(n6001), .Z(n6003) );
  NANDN U6110 ( .A(n5919), .B(n5918), .Z(n5923) );
  NANDN U6111 ( .A(n5921), .B(n5920), .Z(n5922) );
  NAND U6112 ( .A(n5923), .B(n5922), .Z(n6004) );
  XNOR U6113 ( .A(n6003), .B(n6004), .Z(n5949) );
  XOR U6114 ( .A(n5950), .B(n5949), .Z(n6008) );
  NANDN U6115 ( .A(n5925), .B(n5924), .Z(n5929) );
  NANDN U6116 ( .A(n5927), .B(n5926), .Z(n5928) );
  AND U6117 ( .A(n5929), .B(n5928), .Z(n6007) );
  XNOR U6118 ( .A(n6008), .B(n6007), .Z(n6009) );
  XOR U6119 ( .A(n6010), .B(n6009), .Z(n5942) );
  NANDN U6120 ( .A(n5931), .B(n5930), .Z(n5935) );
  NAND U6121 ( .A(n5933), .B(n5932), .Z(n5934) );
  AND U6122 ( .A(n5935), .B(n5934), .Z(n5941) );
  XNOR U6123 ( .A(n5942), .B(n5941), .Z(n5943) );
  XNOR U6124 ( .A(n5944), .B(n5943), .Z(n6013) );
  XNOR U6125 ( .A(sreg[196]), .B(n6013), .Z(n6015) );
  NANDN U6126 ( .A(sreg[195]), .B(n5936), .Z(n5940) );
  NAND U6127 ( .A(n5938), .B(n5937), .Z(n5939) );
  NAND U6128 ( .A(n5940), .B(n5939), .Z(n6014) );
  XNOR U6129 ( .A(n6015), .B(n6014), .Z(c[196]) );
  NANDN U6130 ( .A(n5942), .B(n5941), .Z(n5946) );
  NANDN U6131 ( .A(n5944), .B(n5943), .Z(n5945) );
  AND U6132 ( .A(n5946), .B(n5945), .Z(n6021) );
  NANDN U6133 ( .A(n5948), .B(n5947), .Z(n5952) );
  NAND U6134 ( .A(n5950), .B(n5949), .Z(n5951) );
  AND U6135 ( .A(n5952), .B(n5951), .Z(n6087) );
  NAND U6136 ( .A(n5953), .B(n9883), .Z(n5955) );
  XOR U6137 ( .A(b[11]), .B(a[75]), .Z(n6057) );
  NANDN U6138 ( .A(n9856), .B(n6057), .Z(n5954) );
  AND U6139 ( .A(n5955), .B(n5954), .Z(n6068) );
  NANDN U6140 ( .A(n10005), .B(n5956), .Z(n5958) );
  XOR U6141 ( .A(b[15]), .B(a[71]), .Z(n6060) );
  NANDN U6142 ( .A(n10006), .B(n6060), .Z(n5957) );
  AND U6143 ( .A(n5958), .B(n5957), .Z(n6067) );
  NANDN U6144 ( .A(n9685), .B(n5959), .Z(n5961) );
  XOR U6145 ( .A(b[9]), .B(a[77]), .Z(n6063) );
  NANDN U6146 ( .A(n9758), .B(n6063), .Z(n5960) );
  NAND U6147 ( .A(n5961), .B(n5960), .Z(n6066) );
  XOR U6148 ( .A(n6067), .B(n6066), .Z(n6069) );
  XOR U6149 ( .A(n6068), .B(n6069), .Z(n6079) );
  NANDN U6150 ( .A(n5963), .B(n5962), .Z(n5967) );
  OR U6151 ( .A(n5965), .B(n5964), .Z(n5966) );
  AND U6152 ( .A(n5967), .B(n5966), .Z(n6078) );
  XNOR U6153 ( .A(n6079), .B(n6078), .Z(n6080) );
  NANDN U6154 ( .A(n5969), .B(n5968), .Z(n5973) );
  NANDN U6155 ( .A(n5971), .B(n5970), .Z(n5972) );
  NAND U6156 ( .A(n5973), .B(n5972), .Z(n6081) );
  XNOR U6157 ( .A(n6080), .B(n6081), .Z(n6027) );
  NANDN U6158 ( .A(n5975), .B(n5974), .Z(n5979) );
  NANDN U6159 ( .A(n5977), .B(n5976), .Z(n5978) );
  AND U6160 ( .A(n5979), .B(n5978), .Z(n6053) );
  NAND U6161 ( .A(b[0]), .B(a[85]), .Z(n5980) );
  XNOR U6162 ( .A(b[1]), .B(n5980), .Z(n5982) );
  NANDN U6163 ( .A(b[0]), .B(a[84]), .Z(n5981) );
  NAND U6164 ( .A(n5982), .B(n5981), .Z(n6033) );
  NANDN U6165 ( .A(n9891), .B(n5983), .Z(n5985) );
  XOR U6166 ( .A(b[13]), .B(a[73]), .Z(n6039) );
  NANDN U6167 ( .A(n9935), .B(n6039), .Z(n5984) );
  AND U6168 ( .A(n5985), .B(n5984), .Z(n6031) );
  AND U6169 ( .A(b[15]), .B(a[69]), .Z(n6030) );
  XNOR U6170 ( .A(n6031), .B(n6030), .Z(n6032) );
  XNOR U6171 ( .A(n6033), .B(n6032), .Z(n6051) );
  NANDN U6172 ( .A(n9437), .B(n5986), .Z(n5988) );
  XOR U6173 ( .A(b[5]), .B(a[81]), .Z(n6042) );
  NANDN U6174 ( .A(n9503), .B(n6042), .Z(n5987) );
  AND U6175 ( .A(n5988), .B(n5987), .Z(n6075) );
  NANDN U6176 ( .A(n9588), .B(n5989), .Z(n5991) );
  XOR U6177 ( .A(b[7]), .B(a[79]), .Z(n6045) );
  NANDN U6178 ( .A(n9639), .B(n6045), .Z(n5990) );
  AND U6179 ( .A(n5991), .B(n5990), .Z(n6073) );
  NANDN U6180 ( .A(n9374), .B(n5992), .Z(n5994) );
  XOR U6181 ( .A(b[3]), .B(a[83]), .Z(n6048) );
  NANDN U6182 ( .A(n9375), .B(n6048), .Z(n5993) );
  NAND U6183 ( .A(n5994), .B(n5993), .Z(n6072) );
  XNOR U6184 ( .A(n6073), .B(n6072), .Z(n6074) );
  XOR U6185 ( .A(n6075), .B(n6074), .Z(n6052) );
  XOR U6186 ( .A(n6051), .B(n6052), .Z(n6054) );
  XOR U6187 ( .A(n6053), .B(n6054), .Z(n6025) );
  NANDN U6188 ( .A(n5996), .B(n5995), .Z(n6000) );
  OR U6189 ( .A(n5998), .B(n5997), .Z(n5999) );
  AND U6190 ( .A(n6000), .B(n5999), .Z(n6024) );
  XNOR U6191 ( .A(n6025), .B(n6024), .Z(n6026) );
  XOR U6192 ( .A(n6027), .B(n6026), .Z(n6085) );
  NANDN U6193 ( .A(n6002), .B(n6001), .Z(n6006) );
  NANDN U6194 ( .A(n6004), .B(n6003), .Z(n6005) );
  AND U6195 ( .A(n6006), .B(n6005), .Z(n6084) );
  XNOR U6196 ( .A(n6085), .B(n6084), .Z(n6086) );
  XOR U6197 ( .A(n6087), .B(n6086), .Z(n6019) );
  NANDN U6198 ( .A(n6008), .B(n6007), .Z(n6012) );
  NAND U6199 ( .A(n6010), .B(n6009), .Z(n6011) );
  AND U6200 ( .A(n6012), .B(n6011), .Z(n6018) );
  XNOR U6201 ( .A(n6019), .B(n6018), .Z(n6020) );
  XNOR U6202 ( .A(n6021), .B(n6020), .Z(n6090) );
  XNOR U6203 ( .A(sreg[197]), .B(n6090), .Z(n6092) );
  NANDN U6204 ( .A(sreg[196]), .B(n6013), .Z(n6017) );
  NAND U6205 ( .A(n6015), .B(n6014), .Z(n6016) );
  NAND U6206 ( .A(n6017), .B(n6016), .Z(n6091) );
  XNOR U6207 ( .A(n6092), .B(n6091), .Z(c[197]) );
  NANDN U6208 ( .A(n6019), .B(n6018), .Z(n6023) );
  NANDN U6209 ( .A(n6021), .B(n6020), .Z(n6022) );
  AND U6210 ( .A(n6023), .B(n6022), .Z(n6098) );
  NANDN U6211 ( .A(n6025), .B(n6024), .Z(n6029) );
  NAND U6212 ( .A(n6027), .B(n6026), .Z(n6028) );
  AND U6213 ( .A(n6029), .B(n6028), .Z(n6164) );
  NANDN U6214 ( .A(n6031), .B(n6030), .Z(n6035) );
  NANDN U6215 ( .A(n6033), .B(n6032), .Z(n6034) );
  AND U6216 ( .A(n6035), .B(n6034), .Z(n6130) );
  NAND U6217 ( .A(b[0]), .B(a[86]), .Z(n6036) );
  XNOR U6218 ( .A(b[1]), .B(n6036), .Z(n6038) );
  NANDN U6219 ( .A(b[0]), .B(a[85]), .Z(n6037) );
  NAND U6220 ( .A(n6038), .B(n6037), .Z(n6110) );
  NANDN U6221 ( .A(n9891), .B(n6039), .Z(n6041) );
  XOR U6222 ( .A(b[13]), .B(a[74]), .Z(n6113) );
  NANDN U6223 ( .A(n9935), .B(n6113), .Z(n6040) );
  AND U6224 ( .A(n6041), .B(n6040), .Z(n6108) );
  AND U6225 ( .A(b[15]), .B(a[70]), .Z(n6107) );
  XNOR U6226 ( .A(n6108), .B(n6107), .Z(n6109) );
  XNOR U6227 ( .A(n6110), .B(n6109), .Z(n6128) );
  NANDN U6228 ( .A(n9437), .B(n6042), .Z(n6044) );
  XOR U6229 ( .A(b[5]), .B(a[82]), .Z(n6119) );
  NANDN U6230 ( .A(n9503), .B(n6119), .Z(n6043) );
  AND U6231 ( .A(n6044), .B(n6043), .Z(n6152) );
  NANDN U6232 ( .A(n9588), .B(n6045), .Z(n6047) );
  XOR U6233 ( .A(b[7]), .B(a[80]), .Z(n6122) );
  NANDN U6234 ( .A(n9639), .B(n6122), .Z(n6046) );
  AND U6235 ( .A(n6047), .B(n6046), .Z(n6150) );
  NANDN U6236 ( .A(n9374), .B(n6048), .Z(n6050) );
  XOR U6237 ( .A(b[3]), .B(a[84]), .Z(n6125) );
  NANDN U6238 ( .A(n9375), .B(n6125), .Z(n6049) );
  NAND U6239 ( .A(n6050), .B(n6049), .Z(n6149) );
  XNOR U6240 ( .A(n6150), .B(n6149), .Z(n6151) );
  XOR U6241 ( .A(n6152), .B(n6151), .Z(n6129) );
  XOR U6242 ( .A(n6128), .B(n6129), .Z(n6131) );
  XOR U6243 ( .A(n6130), .B(n6131), .Z(n6102) );
  NANDN U6244 ( .A(n6052), .B(n6051), .Z(n6056) );
  OR U6245 ( .A(n6054), .B(n6053), .Z(n6055) );
  AND U6246 ( .A(n6056), .B(n6055), .Z(n6101) );
  XNOR U6247 ( .A(n6102), .B(n6101), .Z(n6104) );
  NAND U6248 ( .A(n6057), .B(n9883), .Z(n6059) );
  XOR U6249 ( .A(b[11]), .B(a[76]), .Z(n6134) );
  NANDN U6250 ( .A(n9856), .B(n6134), .Z(n6058) );
  AND U6251 ( .A(n6059), .B(n6058), .Z(n6145) );
  NANDN U6252 ( .A(n10005), .B(n6060), .Z(n6062) );
  XOR U6253 ( .A(b[15]), .B(a[72]), .Z(n6137) );
  NANDN U6254 ( .A(n10006), .B(n6137), .Z(n6061) );
  AND U6255 ( .A(n6062), .B(n6061), .Z(n6144) );
  NANDN U6256 ( .A(n9685), .B(n6063), .Z(n6065) );
  XOR U6257 ( .A(b[9]), .B(a[78]), .Z(n6140) );
  NANDN U6258 ( .A(n9758), .B(n6140), .Z(n6064) );
  NAND U6259 ( .A(n6065), .B(n6064), .Z(n6143) );
  XOR U6260 ( .A(n6144), .B(n6143), .Z(n6146) );
  XOR U6261 ( .A(n6145), .B(n6146), .Z(n6156) );
  NANDN U6262 ( .A(n6067), .B(n6066), .Z(n6071) );
  OR U6263 ( .A(n6069), .B(n6068), .Z(n6070) );
  AND U6264 ( .A(n6071), .B(n6070), .Z(n6155) );
  XNOR U6265 ( .A(n6156), .B(n6155), .Z(n6157) );
  NANDN U6266 ( .A(n6073), .B(n6072), .Z(n6077) );
  NANDN U6267 ( .A(n6075), .B(n6074), .Z(n6076) );
  NAND U6268 ( .A(n6077), .B(n6076), .Z(n6158) );
  XNOR U6269 ( .A(n6157), .B(n6158), .Z(n6103) );
  XOR U6270 ( .A(n6104), .B(n6103), .Z(n6162) );
  NANDN U6271 ( .A(n6079), .B(n6078), .Z(n6083) );
  NANDN U6272 ( .A(n6081), .B(n6080), .Z(n6082) );
  AND U6273 ( .A(n6083), .B(n6082), .Z(n6161) );
  XNOR U6274 ( .A(n6162), .B(n6161), .Z(n6163) );
  XOR U6275 ( .A(n6164), .B(n6163), .Z(n6096) );
  NANDN U6276 ( .A(n6085), .B(n6084), .Z(n6089) );
  NAND U6277 ( .A(n6087), .B(n6086), .Z(n6088) );
  AND U6278 ( .A(n6089), .B(n6088), .Z(n6095) );
  XNOR U6279 ( .A(n6096), .B(n6095), .Z(n6097) );
  XNOR U6280 ( .A(n6098), .B(n6097), .Z(n6167) );
  XNOR U6281 ( .A(sreg[198]), .B(n6167), .Z(n6169) );
  NANDN U6282 ( .A(sreg[197]), .B(n6090), .Z(n6094) );
  NAND U6283 ( .A(n6092), .B(n6091), .Z(n6093) );
  NAND U6284 ( .A(n6094), .B(n6093), .Z(n6168) );
  XNOR U6285 ( .A(n6169), .B(n6168), .Z(c[198]) );
  NANDN U6286 ( .A(n6096), .B(n6095), .Z(n6100) );
  NANDN U6287 ( .A(n6098), .B(n6097), .Z(n6099) );
  AND U6288 ( .A(n6100), .B(n6099), .Z(n6175) );
  NANDN U6289 ( .A(n6102), .B(n6101), .Z(n6106) );
  NAND U6290 ( .A(n6104), .B(n6103), .Z(n6105) );
  AND U6291 ( .A(n6106), .B(n6105), .Z(n6241) );
  NANDN U6292 ( .A(n6108), .B(n6107), .Z(n6112) );
  NANDN U6293 ( .A(n6110), .B(n6109), .Z(n6111) );
  AND U6294 ( .A(n6112), .B(n6111), .Z(n6207) );
  NANDN U6295 ( .A(n9891), .B(n6113), .Z(n6115) );
  XOR U6296 ( .A(b[13]), .B(a[75]), .Z(n6190) );
  NANDN U6297 ( .A(n9935), .B(n6190), .Z(n6114) );
  AND U6298 ( .A(n6115), .B(n6114), .Z(n6185) );
  AND U6299 ( .A(b[15]), .B(a[71]), .Z(n6184) );
  XNOR U6300 ( .A(n6185), .B(n6184), .Z(n6186) );
  NAND U6301 ( .A(b[0]), .B(a[87]), .Z(n6116) );
  XNOR U6302 ( .A(b[1]), .B(n6116), .Z(n6118) );
  NANDN U6303 ( .A(b[0]), .B(a[86]), .Z(n6117) );
  NAND U6304 ( .A(n6118), .B(n6117), .Z(n6187) );
  XNOR U6305 ( .A(n6186), .B(n6187), .Z(n6205) );
  NANDN U6306 ( .A(n9437), .B(n6119), .Z(n6121) );
  XOR U6307 ( .A(b[5]), .B(a[83]), .Z(n6196) );
  NANDN U6308 ( .A(n9503), .B(n6196), .Z(n6120) );
  AND U6309 ( .A(n6121), .B(n6120), .Z(n6229) );
  NANDN U6310 ( .A(n9588), .B(n6122), .Z(n6124) );
  XOR U6311 ( .A(b[7]), .B(a[81]), .Z(n6199) );
  NANDN U6312 ( .A(n9639), .B(n6199), .Z(n6123) );
  AND U6313 ( .A(n6124), .B(n6123), .Z(n6227) );
  NANDN U6314 ( .A(n9374), .B(n6125), .Z(n6127) );
  XOR U6315 ( .A(b[3]), .B(a[85]), .Z(n6202) );
  NANDN U6316 ( .A(n9375), .B(n6202), .Z(n6126) );
  NAND U6317 ( .A(n6127), .B(n6126), .Z(n6226) );
  XNOR U6318 ( .A(n6227), .B(n6226), .Z(n6228) );
  XOR U6319 ( .A(n6229), .B(n6228), .Z(n6206) );
  XOR U6320 ( .A(n6205), .B(n6206), .Z(n6208) );
  XOR U6321 ( .A(n6207), .B(n6208), .Z(n6179) );
  NANDN U6322 ( .A(n6129), .B(n6128), .Z(n6133) );
  OR U6323 ( .A(n6131), .B(n6130), .Z(n6132) );
  AND U6324 ( .A(n6133), .B(n6132), .Z(n6178) );
  XNOR U6325 ( .A(n6179), .B(n6178), .Z(n6181) );
  NAND U6326 ( .A(n6134), .B(n9883), .Z(n6136) );
  XOR U6327 ( .A(b[11]), .B(a[77]), .Z(n6211) );
  NANDN U6328 ( .A(n9856), .B(n6211), .Z(n6135) );
  AND U6329 ( .A(n6136), .B(n6135), .Z(n6222) );
  NANDN U6330 ( .A(n10005), .B(n6137), .Z(n6139) );
  XOR U6331 ( .A(b[15]), .B(a[73]), .Z(n6214) );
  NANDN U6332 ( .A(n10006), .B(n6214), .Z(n6138) );
  AND U6333 ( .A(n6139), .B(n6138), .Z(n6221) );
  NANDN U6334 ( .A(n9685), .B(n6140), .Z(n6142) );
  XOR U6335 ( .A(b[9]), .B(a[79]), .Z(n6217) );
  NANDN U6336 ( .A(n9758), .B(n6217), .Z(n6141) );
  NAND U6337 ( .A(n6142), .B(n6141), .Z(n6220) );
  XOR U6338 ( .A(n6221), .B(n6220), .Z(n6223) );
  XOR U6339 ( .A(n6222), .B(n6223), .Z(n6233) );
  NANDN U6340 ( .A(n6144), .B(n6143), .Z(n6148) );
  OR U6341 ( .A(n6146), .B(n6145), .Z(n6147) );
  AND U6342 ( .A(n6148), .B(n6147), .Z(n6232) );
  XNOR U6343 ( .A(n6233), .B(n6232), .Z(n6234) );
  NANDN U6344 ( .A(n6150), .B(n6149), .Z(n6154) );
  NANDN U6345 ( .A(n6152), .B(n6151), .Z(n6153) );
  NAND U6346 ( .A(n6154), .B(n6153), .Z(n6235) );
  XNOR U6347 ( .A(n6234), .B(n6235), .Z(n6180) );
  XOR U6348 ( .A(n6181), .B(n6180), .Z(n6239) );
  NANDN U6349 ( .A(n6156), .B(n6155), .Z(n6160) );
  NANDN U6350 ( .A(n6158), .B(n6157), .Z(n6159) );
  AND U6351 ( .A(n6160), .B(n6159), .Z(n6238) );
  XNOR U6352 ( .A(n6239), .B(n6238), .Z(n6240) );
  XOR U6353 ( .A(n6241), .B(n6240), .Z(n6173) );
  NANDN U6354 ( .A(n6162), .B(n6161), .Z(n6166) );
  NAND U6355 ( .A(n6164), .B(n6163), .Z(n6165) );
  AND U6356 ( .A(n6166), .B(n6165), .Z(n6172) );
  XNOR U6357 ( .A(n6173), .B(n6172), .Z(n6174) );
  XNOR U6358 ( .A(n6175), .B(n6174), .Z(n6244) );
  XNOR U6359 ( .A(sreg[199]), .B(n6244), .Z(n6246) );
  NANDN U6360 ( .A(sreg[198]), .B(n6167), .Z(n6171) );
  NAND U6361 ( .A(n6169), .B(n6168), .Z(n6170) );
  NAND U6362 ( .A(n6171), .B(n6170), .Z(n6245) );
  XNOR U6363 ( .A(n6246), .B(n6245), .Z(c[199]) );
  NANDN U6364 ( .A(n6173), .B(n6172), .Z(n6177) );
  NANDN U6365 ( .A(n6175), .B(n6174), .Z(n6176) );
  AND U6366 ( .A(n6177), .B(n6176), .Z(n6252) );
  NANDN U6367 ( .A(n6179), .B(n6178), .Z(n6183) );
  NAND U6368 ( .A(n6181), .B(n6180), .Z(n6182) );
  AND U6369 ( .A(n6183), .B(n6182), .Z(n6318) );
  NANDN U6370 ( .A(n6185), .B(n6184), .Z(n6189) );
  NANDN U6371 ( .A(n6187), .B(n6186), .Z(n6188) );
  AND U6372 ( .A(n6189), .B(n6188), .Z(n6284) );
  NANDN U6373 ( .A(n9891), .B(n6190), .Z(n6192) );
  XOR U6374 ( .A(b[13]), .B(a[76]), .Z(n6270) );
  NANDN U6375 ( .A(n9935), .B(n6270), .Z(n6191) );
  AND U6376 ( .A(n6192), .B(n6191), .Z(n6262) );
  AND U6377 ( .A(b[15]), .B(a[72]), .Z(n6261) );
  XNOR U6378 ( .A(n6262), .B(n6261), .Z(n6263) );
  NAND U6379 ( .A(b[0]), .B(a[88]), .Z(n6193) );
  XNOR U6380 ( .A(b[1]), .B(n6193), .Z(n6195) );
  NANDN U6381 ( .A(b[0]), .B(a[87]), .Z(n6194) );
  NAND U6382 ( .A(n6195), .B(n6194), .Z(n6264) );
  XNOR U6383 ( .A(n6263), .B(n6264), .Z(n6282) );
  NANDN U6384 ( .A(n9437), .B(n6196), .Z(n6198) );
  XOR U6385 ( .A(b[5]), .B(a[84]), .Z(n6273) );
  NANDN U6386 ( .A(n9503), .B(n6273), .Z(n6197) );
  AND U6387 ( .A(n6198), .B(n6197), .Z(n6306) );
  NANDN U6388 ( .A(n9588), .B(n6199), .Z(n6201) );
  XOR U6389 ( .A(b[7]), .B(a[82]), .Z(n6276) );
  NANDN U6390 ( .A(n9639), .B(n6276), .Z(n6200) );
  AND U6391 ( .A(n6201), .B(n6200), .Z(n6304) );
  NANDN U6392 ( .A(n9374), .B(n6202), .Z(n6204) );
  XOR U6393 ( .A(b[3]), .B(a[86]), .Z(n6279) );
  NANDN U6394 ( .A(n9375), .B(n6279), .Z(n6203) );
  NAND U6395 ( .A(n6204), .B(n6203), .Z(n6303) );
  XNOR U6396 ( .A(n6304), .B(n6303), .Z(n6305) );
  XOR U6397 ( .A(n6306), .B(n6305), .Z(n6283) );
  XOR U6398 ( .A(n6282), .B(n6283), .Z(n6285) );
  XOR U6399 ( .A(n6284), .B(n6285), .Z(n6256) );
  NANDN U6400 ( .A(n6206), .B(n6205), .Z(n6210) );
  OR U6401 ( .A(n6208), .B(n6207), .Z(n6209) );
  AND U6402 ( .A(n6210), .B(n6209), .Z(n6255) );
  XNOR U6403 ( .A(n6256), .B(n6255), .Z(n6258) );
  NAND U6404 ( .A(n6211), .B(n9883), .Z(n6213) );
  XOR U6405 ( .A(b[11]), .B(a[78]), .Z(n6288) );
  NANDN U6406 ( .A(n9856), .B(n6288), .Z(n6212) );
  AND U6407 ( .A(n6213), .B(n6212), .Z(n6299) );
  NANDN U6408 ( .A(n10005), .B(n6214), .Z(n6216) );
  XOR U6409 ( .A(b[15]), .B(a[74]), .Z(n6291) );
  NANDN U6410 ( .A(n10006), .B(n6291), .Z(n6215) );
  AND U6411 ( .A(n6216), .B(n6215), .Z(n6298) );
  NANDN U6412 ( .A(n9685), .B(n6217), .Z(n6219) );
  XOR U6413 ( .A(b[9]), .B(a[80]), .Z(n6294) );
  NANDN U6414 ( .A(n9758), .B(n6294), .Z(n6218) );
  NAND U6415 ( .A(n6219), .B(n6218), .Z(n6297) );
  XOR U6416 ( .A(n6298), .B(n6297), .Z(n6300) );
  XOR U6417 ( .A(n6299), .B(n6300), .Z(n6310) );
  NANDN U6418 ( .A(n6221), .B(n6220), .Z(n6225) );
  OR U6419 ( .A(n6223), .B(n6222), .Z(n6224) );
  AND U6420 ( .A(n6225), .B(n6224), .Z(n6309) );
  XNOR U6421 ( .A(n6310), .B(n6309), .Z(n6311) );
  NANDN U6422 ( .A(n6227), .B(n6226), .Z(n6231) );
  NANDN U6423 ( .A(n6229), .B(n6228), .Z(n6230) );
  NAND U6424 ( .A(n6231), .B(n6230), .Z(n6312) );
  XNOR U6425 ( .A(n6311), .B(n6312), .Z(n6257) );
  XOR U6426 ( .A(n6258), .B(n6257), .Z(n6316) );
  NANDN U6427 ( .A(n6233), .B(n6232), .Z(n6237) );
  NANDN U6428 ( .A(n6235), .B(n6234), .Z(n6236) );
  AND U6429 ( .A(n6237), .B(n6236), .Z(n6315) );
  XNOR U6430 ( .A(n6316), .B(n6315), .Z(n6317) );
  XOR U6431 ( .A(n6318), .B(n6317), .Z(n6250) );
  NANDN U6432 ( .A(n6239), .B(n6238), .Z(n6243) );
  NAND U6433 ( .A(n6241), .B(n6240), .Z(n6242) );
  AND U6434 ( .A(n6243), .B(n6242), .Z(n6249) );
  XNOR U6435 ( .A(n6250), .B(n6249), .Z(n6251) );
  XNOR U6436 ( .A(n6252), .B(n6251), .Z(n6321) );
  XNOR U6437 ( .A(sreg[200]), .B(n6321), .Z(n6323) );
  NANDN U6438 ( .A(sreg[199]), .B(n6244), .Z(n6248) );
  NAND U6439 ( .A(n6246), .B(n6245), .Z(n6247) );
  NAND U6440 ( .A(n6248), .B(n6247), .Z(n6322) );
  XNOR U6441 ( .A(n6323), .B(n6322), .Z(c[200]) );
  NANDN U6442 ( .A(n6250), .B(n6249), .Z(n6254) );
  NANDN U6443 ( .A(n6252), .B(n6251), .Z(n6253) );
  AND U6444 ( .A(n6254), .B(n6253), .Z(n6329) );
  NANDN U6445 ( .A(n6256), .B(n6255), .Z(n6260) );
  NAND U6446 ( .A(n6258), .B(n6257), .Z(n6259) );
  AND U6447 ( .A(n6260), .B(n6259), .Z(n6395) );
  NANDN U6448 ( .A(n6262), .B(n6261), .Z(n6266) );
  NANDN U6449 ( .A(n6264), .B(n6263), .Z(n6265) );
  AND U6450 ( .A(n6266), .B(n6265), .Z(n6361) );
  NAND U6451 ( .A(b[0]), .B(a[89]), .Z(n6267) );
  XNOR U6452 ( .A(b[1]), .B(n6267), .Z(n6269) );
  NANDN U6453 ( .A(b[0]), .B(a[88]), .Z(n6268) );
  NAND U6454 ( .A(n6269), .B(n6268), .Z(n6341) );
  NANDN U6455 ( .A(n9891), .B(n6270), .Z(n6272) );
  XOR U6456 ( .A(b[13]), .B(a[77]), .Z(n6344) );
  NANDN U6457 ( .A(n9935), .B(n6344), .Z(n6271) );
  AND U6458 ( .A(n6272), .B(n6271), .Z(n6339) );
  AND U6459 ( .A(b[15]), .B(a[73]), .Z(n6338) );
  XNOR U6460 ( .A(n6339), .B(n6338), .Z(n6340) );
  XNOR U6461 ( .A(n6341), .B(n6340), .Z(n6359) );
  NANDN U6462 ( .A(n9437), .B(n6273), .Z(n6275) );
  XOR U6463 ( .A(b[5]), .B(a[85]), .Z(n6350) );
  NANDN U6464 ( .A(n9503), .B(n6350), .Z(n6274) );
  AND U6465 ( .A(n6275), .B(n6274), .Z(n6383) );
  NANDN U6466 ( .A(n9588), .B(n6276), .Z(n6278) );
  XOR U6467 ( .A(b[7]), .B(a[83]), .Z(n6353) );
  NANDN U6468 ( .A(n9639), .B(n6353), .Z(n6277) );
  AND U6469 ( .A(n6278), .B(n6277), .Z(n6381) );
  NANDN U6470 ( .A(n9374), .B(n6279), .Z(n6281) );
  XOR U6471 ( .A(b[3]), .B(a[87]), .Z(n6356) );
  NANDN U6472 ( .A(n9375), .B(n6356), .Z(n6280) );
  NAND U6473 ( .A(n6281), .B(n6280), .Z(n6380) );
  XNOR U6474 ( .A(n6381), .B(n6380), .Z(n6382) );
  XOR U6475 ( .A(n6383), .B(n6382), .Z(n6360) );
  XOR U6476 ( .A(n6359), .B(n6360), .Z(n6362) );
  XOR U6477 ( .A(n6361), .B(n6362), .Z(n6333) );
  NANDN U6478 ( .A(n6283), .B(n6282), .Z(n6287) );
  OR U6479 ( .A(n6285), .B(n6284), .Z(n6286) );
  AND U6480 ( .A(n6287), .B(n6286), .Z(n6332) );
  XNOR U6481 ( .A(n6333), .B(n6332), .Z(n6335) );
  NAND U6482 ( .A(n6288), .B(n9883), .Z(n6290) );
  XOR U6483 ( .A(b[11]), .B(a[79]), .Z(n6365) );
  NANDN U6484 ( .A(n9856), .B(n6365), .Z(n6289) );
  AND U6485 ( .A(n6290), .B(n6289), .Z(n6376) );
  NANDN U6486 ( .A(n10005), .B(n6291), .Z(n6293) );
  XOR U6487 ( .A(b[15]), .B(a[75]), .Z(n6368) );
  NANDN U6488 ( .A(n10006), .B(n6368), .Z(n6292) );
  AND U6489 ( .A(n6293), .B(n6292), .Z(n6375) );
  NANDN U6490 ( .A(n9685), .B(n6294), .Z(n6296) );
  XOR U6491 ( .A(b[9]), .B(a[81]), .Z(n6371) );
  NANDN U6492 ( .A(n9758), .B(n6371), .Z(n6295) );
  NAND U6493 ( .A(n6296), .B(n6295), .Z(n6374) );
  XOR U6494 ( .A(n6375), .B(n6374), .Z(n6377) );
  XOR U6495 ( .A(n6376), .B(n6377), .Z(n6387) );
  NANDN U6496 ( .A(n6298), .B(n6297), .Z(n6302) );
  OR U6497 ( .A(n6300), .B(n6299), .Z(n6301) );
  AND U6498 ( .A(n6302), .B(n6301), .Z(n6386) );
  XNOR U6499 ( .A(n6387), .B(n6386), .Z(n6388) );
  NANDN U6500 ( .A(n6304), .B(n6303), .Z(n6308) );
  NANDN U6501 ( .A(n6306), .B(n6305), .Z(n6307) );
  NAND U6502 ( .A(n6308), .B(n6307), .Z(n6389) );
  XNOR U6503 ( .A(n6388), .B(n6389), .Z(n6334) );
  XOR U6504 ( .A(n6335), .B(n6334), .Z(n6393) );
  NANDN U6505 ( .A(n6310), .B(n6309), .Z(n6314) );
  NANDN U6506 ( .A(n6312), .B(n6311), .Z(n6313) );
  AND U6507 ( .A(n6314), .B(n6313), .Z(n6392) );
  XNOR U6508 ( .A(n6393), .B(n6392), .Z(n6394) );
  XOR U6509 ( .A(n6395), .B(n6394), .Z(n6327) );
  NANDN U6510 ( .A(n6316), .B(n6315), .Z(n6320) );
  NAND U6511 ( .A(n6318), .B(n6317), .Z(n6319) );
  AND U6512 ( .A(n6320), .B(n6319), .Z(n6326) );
  XNOR U6513 ( .A(n6327), .B(n6326), .Z(n6328) );
  XNOR U6514 ( .A(n6329), .B(n6328), .Z(n6398) );
  XNOR U6515 ( .A(sreg[201]), .B(n6398), .Z(n6400) );
  NANDN U6516 ( .A(sreg[200]), .B(n6321), .Z(n6325) );
  NAND U6517 ( .A(n6323), .B(n6322), .Z(n6324) );
  NAND U6518 ( .A(n6325), .B(n6324), .Z(n6399) );
  XNOR U6519 ( .A(n6400), .B(n6399), .Z(c[201]) );
  NANDN U6520 ( .A(n6327), .B(n6326), .Z(n6331) );
  NANDN U6521 ( .A(n6329), .B(n6328), .Z(n6330) );
  AND U6522 ( .A(n6331), .B(n6330), .Z(n6406) );
  NANDN U6523 ( .A(n6333), .B(n6332), .Z(n6337) );
  NAND U6524 ( .A(n6335), .B(n6334), .Z(n6336) );
  AND U6525 ( .A(n6337), .B(n6336), .Z(n6472) );
  NANDN U6526 ( .A(n6339), .B(n6338), .Z(n6343) );
  NANDN U6527 ( .A(n6341), .B(n6340), .Z(n6342) );
  AND U6528 ( .A(n6343), .B(n6342), .Z(n6438) );
  NANDN U6529 ( .A(n9891), .B(n6344), .Z(n6346) );
  XOR U6530 ( .A(b[13]), .B(a[78]), .Z(n6424) );
  NANDN U6531 ( .A(n9935), .B(n6424), .Z(n6345) );
  AND U6532 ( .A(n6346), .B(n6345), .Z(n6416) );
  AND U6533 ( .A(b[15]), .B(a[74]), .Z(n6415) );
  XNOR U6534 ( .A(n6416), .B(n6415), .Z(n6417) );
  NAND U6535 ( .A(b[0]), .B(a[90]), .Z(n6347) );
  XNOR U6536 ( .A(b[1]), .B(n6347), .Z(n6349) );
  NANDN U6537 ( .A(b[0]), .B(a[89]), .Z(n6348) );
  NAND U6538 ( .A(n6349), .B(n6348), .Z(n6418) );
  XNOR U6539 ( .A(n6417), .B(n6418), .Z(n6436) );
  NANDN U6540 ( .A(n9437), .B(n6350), .Z(n6352) );
  XOR U6541 ( .A(b[5]), .B(a[86]), .Z(n6427) );
  NANDN U6542 ( .A(n9503), .B(n6427), .Z(n6351) );
  AND U6543 ( .A(n6352), .B(n6351), .Z(n6460) );
  NANDN U6544 ( .A(n9588), .B(n6353), .Z(n6355) );
  XOR U6545 ( .A(b[7]), .B(a[84]), .Z(n6430) );
  NANDN U6546 ( .A(n9639), .B(n6430), .Z(n6354) );
  AND U6547 ( .A(n6355), .B(n6354), .Z(n6458) );
  NANDN U6548 ( .A(n9374), .B(n6356), .Z(n6358) );
  XOR U6549 ( .A(b[3]), .B(a[88]), .Z(n6433) );
  NANDN U6550 ( .A(n9375), .B(n6433), .Z(n6357) );
  NAND U6551 ( .A(n6358), .B(n6357), .Z(n6457) );
  XNOR U6552 ( .A(n6458), .B(n6457), .Z(n6459) );
  XOR U6553 ( .A(n6460), .B(n6459), .Z(n6437) );
  XOR U6554 ( .A(n6436), .B(n6437), .Z(n6439) );
  XOR U6555 ( .A(n6438), .B(n6439), .Z(n6410) );
  NANDN U6556 ( .A(n6360), .B(n6359), .Z(n6364) );
  OR U6557 ( .A(n6362), .B(n6361), .Z(n6363) );
  AND U6558 ( .A(n6364), .B(n6363), .Z(n6409) );
  XNOR U6559 ( .A(n6410), .B(n6409), .Z(n6412) );
  NAND U6560 ( .A(n6365), .B(n9883), .Z(n6367) );
  XOR U6561 ( .A(b[11]), .B(a[80]), .Z(n6442) );
  NANDN U6562 ( .A(n9856), .B(n6442), .Z(n6366) );
  AND U6563 ( .A(n6367), .B(n6366), .Z(n6453) );
  NANDN U6564 ( .A(n10005), .B(n6368), .Z(n6370) );
  XOR U6565 ( .A(b[15]), .B(a[76]), .Z(n6445) );
  NANDN U6566 ( .A(n10006), .B(n6445), .Z(n6369) );
  AND U6567 ( .A(n6370), .B(n6369), .Z(n6452) );
  NANDN U6568 ( .A(n9685), .B(n6371), .Z(n6373) );
  XOR U6569 ( .A(b[9]), .B(a[82]), .Z(n6448) );
  NANDN U6570 ( .A(n9758), .B(n6448), .Z(n6372) );
  NAND U6571 ( .A(n6373), .B(n6372), .Z(n6451) );
  XOR U6572 ( .A(n6452), .B(n6451), .Z(n6454) );
  XOR U6573 ( .A(n6453), .B(n6454), .Z(n6464) );
  NANDN U6574 ( .A(n6375), .B(n6374), .Z(n6379) );
  OR U6575 ( .A(n6377), .B(n6376), .Z(n6378) );
  AND U6576 ( .A(n6379), .B(n6378), .Z(n6463) );
  XNOR U6577 ( .A(n6464), .B(n6463), .Z(n6465) );
  NANDN U6578 ( .A(n6381), .B(n6380), .Z(n6385) );
  NANDN U6579 ( .A(n6383), .B(n6382), .Z(n6384) );
  NAND U6580 ( .A(n6385), .B(n6384), .Z(n6466) );
  XNOR U6581 ( .A(n6465), .B(n6466), .Z(n6411) );
  XOR U6582 ( .A(n6412), .B(n6411), .Z(n6470) );
  NANDN U6583 ( .A(n6387), .B(n6386), .Z(n6391) );
  NANDN U6584 ( .A(n6389), .B(n6388), .Z(n6390) );
  AND U6585 ( .A(n6391), .B(n6390), .Z(n6469) );
  XNOR U6586 ( .A(n6470), .B(n6469), .Z(n6471) );
  XOR U6587 ( .A(n6472), .B(n6471), .Z(n6404) );
  NANDN U6588 ( .A(n6393), .B(n6392), .Z(n6397) );
  NAND U6589 ( .A(n6395), .B(n6394), .Z(n6396) );
  AND U6590 ( .A(n6397), .B(n6396), .Z(n6403) );
  XNOR U6591 ( .A(n6404), .B(n6403), .Z(n6405) );
  XNOR U6592 ( .A(n6406), .B(n6405), .Z(n6475) );
  XNOR U6593 ( .A(sreg[202]), .B(n6475), .Z(n6477) );
  NANDN U6594 ( .A(sreg[201]), .B(n6398), .Z(n6402) );
  NAND U6595 ( .A(n6400), .B(n6399), .Z(n6401) );
  NAND U6596 ( .A(n6402), .B(n6401), .Z(n6476) );
  XNOR U6597 ( .A(n6477), .B(n6476), .Z(c[202]) );
  NANDN U6598 ( .A(n6404), .B(n6403), .Z(n6408) );
  NANDN U6599 ( .A(n6406), .B(n6405), .Z(n6407) );
  AND U6600 ( .A(n6408), .B(n6407), .Z(n6483) );
  NANDN U6601 ( .A(n6410), .B(n6409), .Z(n6414) );
  NAND U6602 ( .A(n6412), .B(n6411), .Z(n6413) );
  AND U6603 ( .A(n6414), .B(n6413), .Z(n6549) );
  NANDN U6604 ( .A(n6416), .B(n6415), .Z(n6420) );
  NANDN U6605 ( .A(n6418), .B(n6417), .Z(n6419) );
  AND U6606 ( .A(n6420), .B(n6419), .Z(n6536) );
  NAND U6607 ( .A(b[0]), .B(a[91]), .Z(n6421) );
  XNOR U6608 ( .A(b[1]), .B(n6421), .Z(n6423) );
  NANDN U6609 ( .A(b[0]), .B(a[90]), .Z(n6422) );
  NAND U6610 ( .A(n6423), .B(n6422), .Z(n6516) );
  NANDN U6611 ( .A(n9891), .B(n6424), .Z(n6426) );
  XOR U6612 ( .A(b[13]), .B(a[79]), .Z(n6522) );
  NANDN U6613 ( .A(n9935), .B(n6522), .Z(n6425) );
  AND U6614 ( .A(n6426), .B(n6425), .Z(n6514) );
  AND U6615 ( .A(b[15]), .B(a[75]), .Z(n6513) );
  XNOR U6616 ( .A(n6514), .B(n6513), .Z(n6515) );
  XNOR U6617 ( .A(n6516), .B(n6515), .Z(n6534) );
  NANDN U6618 ( .A(n9437), .B(n6427), .Z(n6429) );
  XOR U6619 ( .A(b[5]), .B(a[87]), .Z(n6525) );
  NANDN U6620 ( .A(n9503), .B(n6525), .Z(n6428) );
  AND U6621 ( .A(n6429), .B(n6428), .Z(n6510) );
  NANDN U6622 ( .A(n9588), .B(n6430), .Z(n6432) );
  XOR U6623 ( .A(b[7]), .B(a[85]), .Z(n6528) );
  NANDN U6624 ( .A(n9639), .B(n6528), .Z(n6431) );
  AND U6625 ( .A(n6432), .B(n6431), .Z(n6508) );
  NANDN U6626 ( .A(n9374), .B(n6433), .Z(n6435) );
  XOR U6627 ( .A(b[3]), .B(a[89]), .Z(n6531) );
  NANDN U6628 ( .A(n9375), .B(n6531), .Z(n6434) );
  NAND U6629 ( .A(n6435), .B(n6434), .Z(n6507) );
  XNOR U6630 ( .A(n6508), .B(n6507), .Z(n6509) );
  XOR U6631 ( .A(n6510), .B(n6509), .Z(n6535) );
  XOR U6632 ( .A(n6534), .B(n6535), .Z(n6537) );
  XOR U6633 ( .A(n6536), .B(n6537), .Z(n6487) );
  NANDN U6634 ( .A(n6437), .B(n6436), .Z(n6441) );
  OR U6635 ( .A(n6439), .B(n6438), .Z(n6440) );
  AND U6636 ( .A(n6441), .B(n6440), .Z(n6486) );
  XNOR U6637 ( .A(n6487), .B(n6486), .Z(n6489) );
  NAND U6638 ( .A(n6442), .B(n9883), .Z(n6444) );
  XOR U6639 ( .A(b[11]), .B(a[81]), .Z(n6492) );
  NANDN U6640 ( .A(n9856), .B(n6492), .Z(n6443) );
  AND U6641 ( .A(n6444), .B(n6443), .Z(n6503) );
  NANDN U6642 ( .A(n10005), .B(n6445), .Z(n6447) );
  XOR U6643 ( .A(b[15]), .B(a[77]), .Z(n6495) );
  NANDN U6644 ( .A(n10006), .B(n6495), .Z(n6446) );
  AND U6645 ( .A(n6447), .B(n6446), .Z(n6502) );
  NANDN U6646 ( .A(n9685), .B(n6448), .Z(n6450) );
  XOR U6647 ( .A(b[9]), .B(a[83]), .Z(n6498) );
  NANDN U6648 ( .A(n9758), .B(n6498), .Z(n6449) );
  NAND U6649 ( .A(n6450), .B(n6449), .Z(n6501) );
  XOR U6650 ( .A(n6502), .B(n6501), .Z(n6504) );
  XOR U6651 ( .A(n6503), .B(n6504), .Z(n6541) );
  NANDN U6652 ( .A(n6452), .B(n6451), .Z(n6456) );
  OR U6653 ( .A(n6454), .B(n6453), .Z(n6455) );
  AND U6654 ( .A(n6456), .B(n6455), .Z(n6540) );
  XNOR U6655 ( .A(n6541), .B(n6540), .Z(n6542) );
  NANDN U6656 ( .A(n6458), .B(n6457), .Z(n6462) );
  NANDN U6657 ( .A(n6460), .B(n6459), .Z(n6461) );
  NAND U6658 ( .A(n6462), .B(n6461), .Z(n6543) );
  XNOR U6659 ( .A(n6542), .B(n6543), .Z(n6488) );
  XOR U6660 ( .A(n6489), .B(n6488), .Z(n6547) );
  NANDN U6661 ( .A(n6464), .B(n6463), .Z(n6468) );
  NANDN U6662 ( .A(n6466), .B(n6465), .Z(n6467) );
  AND U6663 ( .A(n6468), .B(n6467), .Z(n6546) );
  XNOR U6664 ( .A(n6547), .B(n6546), .Z(n6548) );
  XOR U6665 ( .A(n6549), .B(n6548), .Z(n6481) );
  NANDN U6666 ( .A(n6470), .B(n6469), .Z(n6474) );
  NAND U6667 ( .A(n6472), .B(n6471), .Z(n6473) );
  AND U6668 ( .A(n6474), .B(n6473), .Z(n6480) );
  XNOR U6669 ( .A(n6481), .B(n6480), .Z(n6482) );
  XNOR U6670 ( .A(n6483), .B(n6482), .Z(n6552) );
  XNOR U6671 ( .A(sreg[203]), .B(n6552), .Z(n6554) );
  NANDN U6672 ( .A(sreg[202]), .B(n6475), .Z(n6479) );
  NAND U6673 ( .A(n6477), .B(n6476), .Z(n6478) );
  NAND U6674 ( .A(n6479), .B(n6478), .Z(n6553) );
  XNOR U6675 ( .A(n6554), .B(n6553), .Z(c[203]) );
  NANDN U6676 ( .A(n6481), .B(n6480), .Z(n6485) );
  NANDN U6677 ( .A(n6483), .B(n6482), .Z(n6484) );
  AND U6678 ( .A(n6485), .B(n6484), .Z(n6560) );
  NANDN U6679 ( .A(n6487), .B(n6486), .Z(n6491) );
  NAND U6680 ( .A(n6489), .B(n6488), .Z(n6490) );
  AND U6681 ( .A(n6491), .B(n6490), .Z(n6626) );
  NAND U6682 ( .A(n6492), .B(n9883), .Z(n6494) );
  XOR U6683 ( .A(b[11]), .B(a[82]), .Z(n6596) );
  NANDN U6684 ( .A(n9856), .B(n6596), .Z(n6493) );
  AND U6685 ( .A(n6494), .B(n6493), .Z(n6607) );
  NANDN U6686 ( .A(n10005), .B(n6495), .Z(n6497) );
  XOR U6687 ( .A(b[15]), .B(a[78]), .Z(n6599) );
  NANDN U6688 ( .A(n10006), .B(n6599), .Z(n6496) );
  AND U6689 ( .A(n6497), .B(n6496), .Z(n6606) );
  NANDN U6690 ( .A(n9685), .B(n6498), .Z(n6500) );
  XOR U6691 ( .A(b[9]), .B(a[84]), .Z(n6602) );
  NANDN U6692 ( .A(n9758), .B(n6602), .Z(n6499) );
  NAND U6693 ( .A(n6500), .B(n6499), .Z(n6605) );
  XOR U6694 ( .A(n6606), .B(n6605), .Z(n6608) );
  XOR U6695 ( .A(n6607), .B(n6608), .Z(n6618) );
  NANDN U6696 ( .A(n6502), .B(n6501), .Z(n6506) );
  OR U6697 ( .A(n6504), .B(n6503), .Z(n6505) );
  AND U6698 ( .A(n6506), .B(n6505), .Z(n6617) );
  XNOR U6699 ( .A(n6618), .B(n6617), .Z(n6619) );
  NANDN U6700 ( .A(n6508), .B(n6507), .Z(n6512) );
  NANDN U6701 ( .A(n6510), .B(n6509), .Z(n6511) );
  NAND U6702 ( .A(n6512), .B(n6511), .Z(n6620) );
  XNOR U6703 ( .A(n6619), .B(n6620), .Z(n6566) );
  NANDN U6704 ( .A(n6514), .B(n6513), .Z(n6518) );
  NANDN U6705 ( .A(n6516), .B(n6515), .Z(n6517) );
  AND U6706 ( .A(n6518), .B(n6517), .Z(n6592) );
  NAND U6707 ( .A(b[0]), .B(a[92]), .Z(n6519) );
  XNOR U6708 ( .A(b[1]), .B(n6519), .Z(n6521) );
  NANDN U6709 ( .A(b[0]), .B(a[91]), .Z(n6520) );
  NAND U6710 ( .A(n6521), .B(n6520), .Z(n6572) );
  NANDN U6711 ( .A(n9891), .B(n6522), .Z(n6524) );
  XOR U6712 ( .A(b[13]), .B(a[80]), .Z(n6575) );
  NANDN U6713 ( .A(n9935), .B(n6575), .Z(n6523) );
  AND U6714 ( .A(n6524), .B(n6523), .Z(n6570) );
  AND U6715 ( .A(b[15]), .B(a[76]), .Z(n6569) );
  XNOR U6716 ( .A(n6570), .B(n6569), .Z(n6571) );
  XNOR U6717 ( .A(n6572), .B(n6571), .Z(n6590) );
  NANDN U6718 ( .A(n9437), .B(n6525), .Z(n6527) );
  XOR U6719 ( .A(b[5]), .B(a[88]), .Z(n6581) );
  NANDN U6720 ( .A(n9503), .B(n6581), .Z(n6526) );
  AND U6721 ( .A(n6527), .B(n6526), .Z(n6614) );
  NANDN U6722 ( .A(n9588), .B(n6528), .Z(n6530) );
  XOR U6723 ( .A(b[7]), .B(a[86]), .Z(n6584) );
  NANDN U6724 ( .A(n9639), .B(n6584), .Z(n6529) );
  AND U6725 ( .A(n6530), .B(n6529), .Z(n6612) );
  NANDN U6726 ( .A(n9374), .B(n6531), .Z(n6533) );
  XOR U6727 ( .A(b[3]), .B(a[90]), .Z(n6587) );
  NANDN U6728 ( .A(n9375), .B(n6587), .Z(n6532) );
  NAND U6729 ( .A(n6533), .B(n6532), .Z(n6611) );
  XNOR U6730 ( .A(n6612), .B(n6611), .Z(n6613) );
  XOR U6731 ( .A(n6614), .B(n6613), .Z(n6591) );
  XOR U6732 ( .A(n6590), .B(n6591), .Z(n6593) );
  XOR U6733 ( .A(n6592), .B(n6593), .Z(n6564) );
  NANDN U6734 ( .A(n6535), .B(n6534), .Z(n6539) );
  OR U6735 ( .A(n6537), .B(n6536), .Z(n6538) );
  AND U6736 ( .A(n6539), .B(n6538), .Z(n6563) );
  XNOR U6737 ( .A(n6564), .B(n6563), .Z(n6565) );
  XOR U6738 ( .A(n6566), .B(n6565), .Z(n6624) );
  NANDN U6739 ( .A(n6541), .B(n6540), .Z(n6545) );
  NANDN U6740 ( .A(n6543), .B(n6542), .Z(n6544) );
  AND U6741 ( .A(n6545), .B(n6544), .Z(n6623) );
  XNOR U6742 ( .A(n6624), .B(n6623), .Z(n6625) );
  XOR U6743 ( .A(n6626), .B(n6625), .Z(n6558) );
  NANDN U6744 ( .A(n6547), .B(n6546), .Z(n6551) );
  NAND U6745 ( .A(n6549), .B(n6548), .Z(n6550) );
  AND U6746 ( .A(n6551), .B(n6550), .Z(n6557) );
  XNOR U6747 ( .A(n6558), .B(n6557), .Z(n6559) );
  XNOR U6748 ( .A(n6560), .B(n6559), .Z(n6629) );
  XNOR U6749 ( .A(sreg[204]), .B(n6629), .Z(n6631) );
  NANDN U6750 ( .A(sreg[203]), .B(n6552), .Z(n6556) );
  NAND U6751 ( .A(n6554), .B(n6553), .Z(n6555) );
  NAND U6752 ( .A(n6556), .B(n6555), .Z(n6630) );
  XNOR U6753 ( .A(n6631), .B(n6630), .Z(c[204]) );
  NANDN U6754 ( .A(n6558), .B(n6557), .Z(n6562) );
  NANDN U6755 ( .A(n6560), .B(n6559), .Z(n6561) );
  AND U6756 ( .A(n6562), .B(n6561), .Z(n6637) );
  NANDN U6757 ( .A(n6564), .B(n6563), .Z(n6568) );
  NAND U6758 ( .A(n6566), .B(n6565), .Z(n6567) );
  AND U6759 ( .A(n6568), .B(n6567), .Z(n6703) );
  NANDN U6760 ( .A(n6570), .B(n6569), .Z(n6574) );
  NANDN U6761 ( .A(n6572), .B(n6571), .Z(n6573) );
  AND U6762 ( .A(n6574), .B(n6573), .Z(n6669) );
  NANDN U6763 ( .A(n9891), .B(n6575), .Z(n6577) );
  XOR U6764 ( .A(b[13]), .B(a[81]), .Z(n6655) );
  NANDN U6765 ( .A(n9935), .B(n6655), .Z(n6576) );
  AND U6766 ( .A(n6577), .B(n6576), .Z(n6647) );
  AND U6767 ( .A(b[15]), .B(a[77]), .Z(n6646) );
  XNOR U6768 ( .A(n6647), .B(n6646), .Z(n6648) );
  NAND U6769 ( .A(b[0]), .B(a[93]), .Z(n6578) );
  XNOR U6770 ( .A(b[1]), .B(n6578), .Z(n6580) );
  NANDN U6771 ( .A(b[0]), .B(a[92]), .Z(n6579) );
  NAND U6772 ( .A(n6580), .B(n6579), .Z(n6649) );
  XNOR U6773 ( .A(n6648), .B(n6649), .Z(n6667) );
  NANDN U6774 ( .A(n9437), .B(n6581), .Z(n6583) );
  XOR U6775 ( .A(b[5]), .B(a[89]), .Z(n6658) );
  NANDN U6776 ( .A(n9503), .B(n6658), .Z(n6582) );
  AND U6777 ( .A(n6583), .B(n6582), .Z(n6691) );
  NANDN U6778 ( .A(n9588), .B(n6584), .Z(n6586) );
  XOR U6779 ( .A(b[7]), .B(a[87]), .Z(n6661) );
  NANDN U6780 ( .A(n9639), .B(n6661), .Z(n6585) );
  AND U6781 ( .A(n6586), .B(n6585), .Z(n6689) );
  NANDN U6782 ( .A(n9374), .B(n6587), .Z(n6589) );
  XOR U6783 ( .A(b[3]), .B(a[91]), .Z(n6664) );
  NANDN U6784 ( .A(n9375), .B(n6664), .Z(n6588) );
  NAND U6785 ( .A(n6589), .B(n6588), .Z(n6688) );
  XNOR U6786 ( .A(n6689), .B(n6688), .Z(n6690) );
  XOR U6787 ( .A(n6691), .B(n6690), .Z(n6668) );
  XOR U6788 ( .A(n6667), .B(n6668), .Z(n6670) );
  XOR U6789 ( .A(n6669), .B(n6670), .Z(n6641) );
  NANDN U6790 ( .A(n6591), .B(n6590), .Z(n6595) );
  OR U6791 ( .A(n6593), .B(n6592), .Z(n6594) );
  AND U6792 ( .A(n6595), .B(n6594), .Z(n6640) );
  XNOR U6793 ( .A(n6641), .B(n6640), .Z(n6643) );
  NAND U6794 ( .A(n6596), .B(n9883), .Z(n6598) );
  XOR U6795 ( .A(b[11]), .B(a[83]), .Z(n6673) );
  NANDN U6796 ( .A(n9856), .B(n6673), .Z(n6597) );
  AND U6797 ( .A(n6598), .B(n6597), .Z(n6684) );
  NANDN U6798 ( .A(n10005), .B(n6599), .Z(n6601) );
  XOR U6799 ( .A(b[15]), .B(a[79]), .Z(n6676) );
  NANDN U6800 ( .A(n10006), .B(n6676), .Z(n6600) );
  AND U6801 ( .A(n6601), .B(n6600), .Z(n6683) );
  NANDN U6802 ( .A(n9685), .B(n6602), .Z(n6604) );
  XOR U6803 ( .A(b[9]), .B(a[85]), .Z(n6679) );
  NANDN U6804 ( .A(n9758), .B(n6679), .Z(n6603) );
  NAND U6805 ( .A(n6604), .B(n6603), .Z(n6682) );
  XOR U6806 ( .A(n6683), .B(n6682), .Z(n6685) );
  XOR U6807 ( .A(n6684), .B(n6685), .Z(n6695) );
  NANDN U6808 ( .A(n6606), .B(n6605), .Z(n6610) );
  OR U6809 ( .A(n6608), .B(n6607), .Z(n6609) );
  AND U6810 ( .A(n6610), .B(n6609), .Z(n6694) );
  XNOR U6811 ( .A(n6695), .B(n6694), .Z(n6696) );
  NANDN U6812 ( .A(n6612), .B(n6611), .Z(n6616) );
  NANDN U6813 ( .A(n6614), .B(n6613), .Z(n6615) );
  NAND U6814 ( .A(n6616), .B(n6615), .Z(n6697) );
  XNOR U6815 ( .A(n6696), .B(n6697), .Z(n6642) );
  XOR U6816 ( .A(n6643), .B(n6642), .Z(n6701) );
  NANDN U6817 ( .A(n6618), .B(n6617), .Z(n6622) );
  NANDN U6818 ( .A(n6620), .B(n6619), .Z(n6621) );
  AND U6819 ( .A(n6622), .B(n6621), .Z(n6700) );
  XNOR U6820 ( .A(n6701), .B(n6700), .Z(n6702) );
  XOR U6821 ( .A(n6703), .B(n6702), .Z(n6635) );
  NANDN U6822 ( .A(n6624), .B(n6623), .Z(n6628) );
  NAND U6823 ( .A(n6626), .B(n6625), .Z(n6627) );
  AND U6824 ( .A(n6628), .B(n6627), .Z(n6634) );
  XNOR U6825 ( .A(n6635), .B(n6634), .Z(n6636) );
  XNOR U6826 ( .A(n6637), .B(n6636), .Z(n6706) );
  XNOR U6827 ( .A(sreg[205]), .B(n6706), .Z(n6708) );
  NANDN U6828 ( .A(sreg[204]), .B(n6629), .Z(n6633) );
  NAND U6829 ( .A(n6631), .B(n6630), .Z(n6632) );
  NAND U6830 ( .A(n6633), .B(n6632), .Z(n6707) );
  XNOR U6831 ( .A(n6708), .B(n6707), .Z(c[205]) );
  NANDN U6832 ( .A(n6635), .B(n6634), .Z(n6639) );
  NANDN U6833 ( .A(n6637), .B(n6636), .Z(n6638) );
  AND U6834 ( .A(n6639), .B(n6638), .Z(n6714) );
  NANDN U6835 ( .A(n6641), .B(n6640), .Z(n6645) );
  NAND U6836 ( .A(n6643), .B(n6642), .Z(n6644) );
  AND U6837 ( .A(n6645), .B(n6644), .Z(n6780) );
  NANDN U6838 ( .A(n6647), .B(n6646), .Z(n6651) );
  NANDN U6839 ( .A(n6649), .B(n6648), .Z(n6650) );
  AND U6840 ( .A(n6651), .B(n6650), .Z(n6746) );
  NAND U6841 ( .A(b[0]), .B(a[94]), .Z(n6652) );
  XNOR U6842 ( .A(b[1]), .B(n6652), .Z(n6654) );
  NANDN U6843 ( .A(b[0]), .B(a[93]), .Z(n6653) );
  NAND U6844 ( .A(n6654), .B(n6653), .Z(n6726) );
  NANDN U6845 ( .A(n9891), .B(n6655), .Z(n6657) );
  XOR U6846 ( .A(b[13]), .B(a[82]), .Z(n6729) );
  NANDN U6847 ( .A(n9935), .B(n6729), .Z(n6656) );
  AND U6848 ( .A(n6657), .B(n6656), .Z(n6724) );
  AND U6849 ( .A(b[15]), .B(a[78]), .Z(n6723) );
  XNOR U6850 ( .A(n6724), .B(n6723), .Z(n6725) );
  XNOR U6851 ( .A(n6726), .B(n6725), .Z(n6744) );
  NANDN U6852 ( .A(n9437), .B(n6658), .Z(n6660) );
  XOR U6853 ( .A(b[5]), .B(a[90]), .Z(n6735) );
  NANDN U6854 ( .A(n9503), .B(n6735), .Z(n6659) );
  AND U6855 ( .A(n6660), .B(n6659), .Z(n6768) );
  NANDN U6856 ( .A(n9588), .B(n6661), .Z(n6663) );
  XOR U6857 ( .A(b[7]), .B(a[88]), .Z(n6738) );
  NANDN U6858 ( .A(n9639), .B(n6738), .Z(n6662) );
  AND U6859 ( .A(n6663), .B(n6662), .Z(n6766) );
  NANDN U6860 ( .A(n9374), .B(n6664), .Z(n6666) );
  XOR U6861 ( .A(b[3]), .B(a[92]), .Z(n6741) );
  NANDN U6862 ( .A(n9375), .B(n6741), .Z(n6665) );
  NAND U6863 ( .A(n6666), .B(n6665), .Z(n6765) );
  XNOR U6864 ( .A(n6766), .B(n6765), .Z(n6767) );
  XOR U6865 ( .A(n6768), .B(n6767), .Z(n6745) );
  XOR U6866 ( .A(n6744), .B(n6745), .Z(n6747) );
  XOR U6867 ( .A(n6746), .B(n6747), .Z(n6718) );
  NANDN U6868 ( .A(n6668), .B(n6667), .Z(n6672) );
  OR U6869 ( .A(n6670), .B(n6669), .Z(n6671) );
  AND U6870 ( .A(n6672), .B(n6671), .Z(n6717) );
  XNOR U6871 ( .A(n6718), .B(n6717), .Z(n6720) );
  NAND U6872 ( .A(n6673), .B(n9883), .Z(n6675) );
  XOR U6873 ( .A(b[11]), .B(a[84]), .Z(n6750) );
  NANDN U6874 ( .A(n9856), .B(n6750), .Z(n6674) );
  AND U6875 ( .A(n6675), .B(n6674), .Z(n6761) );
  NANDN U6876 ( .A(n10005), .B(n6676), .Z(n6678) );
  XOR U6877 ( .A(b[15]), .B(a[80]), .Z(n6753) );
  NANDN U6878 ( .A(n10006), .B(n6753), .Z(n6677) );
  AND U6879 ( .A(n6678), .B(n6677), .Z(n6760) );
  NANDN U6880 ( .A(n9685), .B(n6679), .Z(n6681) );
  XOR U6881 ( .A(b[9]), .B(a[86]), .Z(n6756) );
  NANDN U6882 ( .A(n9758), .B(n6756), .Z(n6680) );
  NAND U6883 ( .A(n6681), .B(n6680), .Z(n6759) );
  XOR U6884 ( .A(n6760), .B(n6759), .Z(n6762) );
  XOR U6885 ( .A(n6761), .B(n6762), .Z(n6772) );
  NANDN U6886 ( .A(n6683), .B(n6682), .Z(n6687) );
  OR U6887 ( .A(n6685), .B(n6684), .Z(n6686) );
  AND U6888 ( .A(n6687), .B(n6686), .Z(n6771) );
  XNOR U6889 ( .A(n6772), .B(n6771), .Z(n6773) );
  NANDN U6890 ( .A(n6689), .B(n6688), .Z(n6693) );
  NANDN U6891 ( .A(n6691), .B(n6690), .Z(n6692) );
  NAND U6892 ( .A(n6693), .B(n6692), .Z(n6774) );
  XNOR U6893 ( .A(n6773), .B(n6774), .Z(n6719) );
  XOR U6894 ( .A(n6720), .B(n6719), .Z(n6778) );
  NANDN U6895 ( .A(n6695), .B(n6694), .Z(n6699) );
  NANDN U6896 ( .A(n6697), .B(n6696), .Z(n6698) );
  AND U6897 ( .A(n6699), .B(n6698), .Z(n6777) );
  XNOR U6898 ( .A(n6778), .B(n6777), .Z(n6779) );
  XOR U6899 ( .A(n6780), .B(n6779), .Z(n6712) );
  NANDN U6900 ( .A(n6701), .B(n6700), .Z(n6705) );
  NAND U6901 ( .A(n6703), .B(n6702), .Z(n6704) );
  AND U6902 ( .A(n6705), .B(n6704), .Z(n6711) );
  XNOR U6903 ( .A(n6712), .B(n6711), .Z(n6713) );
  XNOR U6904 ( .A(n6714), .B(n6713), .Z(n6783) );
  XNOR U6905 ( .A(sreg[206]), .B(n6783), .Z(n6785) );
  NANDN U6906 ( .A(sreg[205]), .B(n6706), .Z(n6710) );
  NAND U6907 ( .A(n6708), .B(n6707), .Z(n6709) );
  NAND U6908 ( .A(n6710), .B(n6709), .Z(n6784) );
  XNOR U6909 ( .A(n6785), .B(n6784), .Z(c[206]) );
  NANDN U6910 ( .A(n6712), .B(n6711), .Z(n6716) );
  NANDN U6911 ( .A(n6714), .B(n6713), .Z(n6715) );
  AND U6912 ( .A(n6716), .B(n6715), .Z(n6791) );
  NANDN U6913 ( .A(n6718), .B(n6717), .Z(n6722) );
  NAND U6914 ( .A(n6720), .B(n6719), .Z(n6721) );
  AND U6915 ( .A(n6722), .B(n6721), .Z(n6857) );
  NANDN U6916 ( .A(n6724), .B(n6723), .Z(n6728) );
  NANDN U6917 ( .A(n6726), .B(n6725), .Z(n6727) );
  AND U6918 ( .A(n6728), .B(n6727), .Z(n6823) );
  NANDN U6919 ( .A(n9891), .B(n6729), .Z(n6731) );
  XOR U6920 ( .A(b[13]), .B(a[83]), .Z(n6806) );
  NANDN U6921 ( .A(n9935), .B(n6806), .Z(n6730) );
  AND U6922 ( .A(n6731), .B(n6730), .Z(n6801) );
  AND U6923 ( .A(b[15]), .B(a[79]), .Z(n6800) );
  XNOR U6924 ( .A(n6801), .B(n6800), .Z(n6802) );
  NAND U6925 ( .A(b[0]), .B(a[95]), .Z(n6732) );
  XNOR U6926 ( .A(b[1]), .B(n6732), .Z(n6734) );
  NANDN U6927 ( .A(b[0]), .B(a[94]), .Z(n6733) );
  NAND U6928 ( .A(n6734), .B(n6733), .Z(n6803) );
  XNOR U6929 ( .A(n6802), .B(n6803), .Z(n6821) );
  NANDN U6930 ( .A(n9437), .B(n6735), .Z(n6737) );
  XOR U6931 ( .A(b[5]), .B(a[91]), .Z(n6812) );
  NANDN U6932 ( .A(n9503), .B(n6812), .Z(n6736) );
  AND U6933 ( .A(n6737), .B(n6736), .Z(n6845) );
  NANDN U6934 ( .A(n9588), .B(n6738), .Z(n6740) );
  XOR U6935 ( .A(b[7]), .B(a[89]), .Z(n6815) );
  NANDN U6936 ( .A(n9639), .B(n6815), .Z(n6739) );
  AND U6937 ( .A(n6740), .B(n6739), .Z(n6843) );
  NANDN U6938 ( .A(n9374), .B(n6741), .Z(n6743) );
  XOR U6939 ( .A(b[3]), .B(a[93]), .Z(n6818) );
  NANDN U6940 ( .A(n9375), .B(n6818), .Z(n6742) );
  NAND U6941 ( .A(n6743), .B(n6742), .Z(n6842) );
  XNOR U6942 ( .A(n6843), .B(n6842), .Z(n6844) );
  XOR U6943 ( .A(n6845), .B(n6844), .Z(n6822) );
  XOR U6944 ( .A(n6821), .B(n6822), .Z(n6824) );
  XOR U6945 ( .A(n6823), .B(n6824), .Z(n6795) );
  NANDN U6946 ( .A(n6745), .B(n6744), .Z(n6749) );
  OR U6947 ( .A(n6747), .B(n6746), .Z(n6748) );
  AND U6948 ( .A(n6749), .B(n6748), .Z(n6794) );
  XNOR U6949 ( .A(n6795), .B(n6794), .Z(n6797) );
  NAND U6950 ( .A(n6750), .B(n9883), .Z(n6752) );
  XOR U6951 ( .A(b[11]), .B(a[85]), .Z(n6827) );
  NANDN U6952 ( .A(n9856), .B(n6827), .Z(n6751) );
  AND U6953 ( .A(n6752), .B(n6751), .Z(n6838) );
  NANDN U6954 ( .A(n10005), .B(n6753), .Z(n6755) );
  XOR U6955 ( .A(b[15]), .B(a[81]), .Z(n6830) );
  NANDN U6956 ( .A(n10006), .B(n6830), .Z(n6754) );
  AND U6957 ( .A(n6755), .B(n6754), .Z(n6837) );
  NANDN U6958 ( .A(n9685), .B(n6756), .Z(n6758) );
  XOR U6959 ( .A(b[9]), .B(a[87]), .Z(n6833) );
  NANDN U6960 ( .A(n9758), .B(n6833), .Z(n6757) );
  NAND U6961 ( .A(n6758), .B(n6757), .Z(n6836) );
  XOR U6962 ( .A(n6837), .B(n6836), .Z(n6839) );
  XOR U6963 ( .A(n6838), .B(n6839), .Z(n6849) );
  NANDN U6964 ( .A(n6760), .B(n6759), .Z(n6764) );
  OR U6965 ( .A(n6762), .B(n6761), .Z(n6763) );
  AND U6966 ( .A(n6764), .B(n6763), .Z(n6848) );
  XNOR U6967 ( .A(n6849), .B(n6848), .Z(n6850) );
  NANDN U6968 ( .A(n6766), .B(n6765), .Z(n6770) );
  NANDN U6969 ( .A(n6768), .B(n6767), .Z(n6769) );
  NAND U6970 ( .A(n6770), .B(n6769), .Z(n6851) );
  XNOR U6971 ( .A(n6850), .B(n6851), .Z(n6796) );
  XOR U6972 ( .A(n6797), .B(n6796), .Z(n6855) );
  NANDN U6973 ( .A(n6772), .B(n6771), .Z(n6776) );
  NANDN U6974 ( .A(n6774), .B(n6773), .Z(n6775) );
  AND U6975 ( .A(n6776), .B(n6775), .Z(n6854) );
  XNOR U6976 ( .A(n6855), .B(n6854), .Z(n6856) );
  XOR U6977 ( .A(n6857), .B(n6856), .Z(n6789) );
  NANDN U6978 ( .A(n6778), .B(n6777), .Z(n6782) );
  NAND U6979 ( .A(n6780), .B(n6779), .Z(n6781) );
  AND U6980 ( .A(n6782), .B(n6781), .Z(n6788) );
  XNOR U6981 ( .A(n6789), .B(n6788), .Z(n6790) );
  XNOR U6982 ( .A(n6791), .B(n6790), .Z(n6860) );
  XNOR U6983 ( .A(sreg[207]), .B(n6860), .Z(n6862) );
  NANDN U6984 ( .A(sreg[206]), .B(n6783), .Z(n6787) );
  NAND U6985 ( .A(n6785), .B(n6784), .Z(n6786) );
  NAND U6986 ( .A(n6787), .B(n6786), .Z(n6861) );
  XNOR U6987 ( .A(n6862), .B(n6861), .Z(c[207]) );
  NANDN U6988 ( .A(n6789), .B(n6788), .Z(n6793) );
  NANDN U6989 ( .A(n6791), .B(n6790), .Z(n6792) );
  AND U6990 ( .A(n6793), .B(n6792), .Z(n6868) );
  NANDN U6991 ( .A(n6795), .B(n6794), .Z(n6799) );
  NAND U6992 ( .A(n6797), .B(n6796), .Z(n6798) );
  AND U6993 ( .A(n6799), .B(n6798), .Z(n6934) );
  NANDN U6994 ( .A(n6801), .B(n6800), .Z(n6805) );
  NANDN U6995 ( .A(n6803), .B(n6802), .Z(n6804) );
  AND U6996 ( .A(n6805), .B(n6804), .Z(n6900) );
  NANDN U6997 ( .A(n9891), .B(n6806), .Z(n6808) );
  XOR U6998 ( .A(b[13]), .B(a[84]), .Z(n6883) );
  NANDN U6999 ( .A(n9935), .B(n6883), .Z(n6807) );
  AND U7000 ( .A(n6808), .B(n6807), .Z(n6878) );
  AND U7001 ( .A(b[15]), .B(a[80]), .Z(n6877) );
  XNOR U7002 ( .A(n6878), .B(n6877), .Z(n6879) );
  NAND U7003 ( .A(b[0]), .B(a[96]), .Z(n6809) );
  XNOR U7004 ( .A(b[1]), .B(n6809), .Z(n6811) );
  NANDN U7005 ( .A(b[0]), .B(a[95]), .Z(n6810) );
  NAND U7006 ( .A(n6811), .B(n6810), .Z(n6880) );
  XNOR U7007 ( .A(n6879), .B(n6880), .Z(n6898) );
  NANDN U7008 ( .A(n9437), .B(n6812), .Z(n6814) );
  XOR U7009 ( .A(b[5]), .B(a[92]), .Z(n6889) );
  NANDN U7010 ( .A(n9503), .B(n6889), .Z(n6813) );
  AND U7011 ( .A(n6814), .B(n6813), .Z(n6922) );
  NANDN U7012 ( .A(n9588), .B(n6815), .Z(n6817) );
  XOR U7013 ( .A(b[7]), .B(a[90]), .Z(n6892) );
  NANDN U7014 ( .A(n9639), .B(n6892), .Z(n6816) );
  AND U7015 ( .A(n6817), .B(n6816), .Z(n6920) );
  NANDN U7016 ( .A(n9374), .B(n6818), .Z(n6820) );
  XOR U7017 ( .A(b[3]), .B(a[94]), .Z(n6895) );
  NANDN U7018 ( .A(n9375), .B(n6895), .Z(n6819) );
  NAND U7019 ( .A(n6820), .B(n6819), .Z(n6919) );
  XNOR U7020 ( .A(n6920), .B(n6919), .Z(n6921) );
  XOR U7021 ( .A(n6922), .B(n6921), .Z(n6899) );
  XOR U7022 ( .A(n6898), .B(n6899), .Z(n6901) );
  XOR U7023 ( .A(n6900), .B(n6901), .Z(n6872) );
  NANDN U7024 ( .A(n6822), .B(n6821), .Z(n6826) );
  OR U7025 ( .A(n6824), .B(n6823), .Z(n6825) );
  AND U7026 ( .A(n6826), .B(n6825), .Z(n6871) );
  XNOR U7027 ( .A(n6872), .B(n6871), .Z(n6874) );
  NAND U7028 ( .A(n6827), .B(n9883), .Z(n6829) );
  XOR U7029 ( .A(b[11]), .B(a[86]), .Z(n6904) );
  NANDN U7030 ( .A(n9856), .B(n6904), .Z(n6828) );
  AND U7031 ( .A(n6829), .B(n6828), .Z(n6915) );
  NANDN U7032 ( .A(n10005), .B(n6830), .Z(n6832) );
  XOR U7033 ( .A(b[15]), .B(a[82]), .Z(n6907) );
  NANDN U7034 ( .A(n10006), .B(n6907), .Z(n6831) );
  AND U7035 ( .A(n6832), .B(n6831), .Z(n6914) );
  NANDN U7036 ( .A(n9685), .B(n6833), .Z(n6835) );
  XOR U7037 ( .A(b[9]), .B(a[88]), .Z(n6910) );
  NANDN U7038 ( .A(n9758), .B(n6910), .Z(n6834) );
  NAND U7039 ( .A(n6835), .B(n6834), .Z(n6913) );
  XOR U7040 ( .A(n6914), .B(n6913), .Z(n6916) );
  XOR U7041 ( .A(n6915), .B(n6916), .Z(n6926) );
  NANDN U7042 ( .A(n6837), .B(n6836), .Z(n6841) );
  OR U7043 ( .A(n6839), .B(n6838), .Z(n6840) );
  AND U7044 ( .A(n6841), .B(n6840), .Z(n6925) );
  XNOR U7045 ( .A(n6926), .B(n6925), .Z(n6927) );
  NANDN U7046 ( .A(n6843), .B(n6842), .Z(n6847) );
  NANDN U7047 ( .A(n6845), .B(n6844), .Z(n6846) );
  NAND U7048 ( .A(n6847), .B(n6846), .Z(n6928) );
  XNOR U7049 ( .A(n6927), .B(n6928), .Z(n6873) );
  XOR U7050 ( .A(n6874), .B(n6873), .Z(n6932) );
  NANDN U7051 ( .A(n6849), .B(n6848), .Z(n6853) );
  NANDN U7052 ( .A(n6851), .B(n6850), .Z(n6852) );
  AND U7053 ( .A(n6853), .B(n6852), .Z(n6931) );
  XNOR U7054 ( .A(n6932), .B(n6931), .Z(n6933) );
  XOR U7055 ( .A(n6934), .B(n6933), .Z(n6866) );
  NANDN U7056 ( .A(n6855), .B(n6854), .Z(n6859) );
  NAND U7057 ( .A(n6857), .B(n6856), .Z(n6858) );
  AND U7058 ( .A(n6859), .B(n6858), .Z(n6865) );
  XNOR U7059 ( .A(n6866), .B(n6865), .Z(n6867) );
  XNOR U7060 ( .A(n6868), .B(n6867), .Z(n6937) );
  XNOR U7061 ( .A(sreg[208]), .B(n6937), .Z(n6939) );
  NANDN U7062 ( .A(sreg[207]), .B(n6860), .Z(n6864) );
  NAND U7063 ( .A(n6862), .B(n6861), .Z(n6863) );
  NAND U7064 ( .A(n6864), .B(n6863), .Z(n6938) );
  XNOR U7065 ( .A(n6939), .B(n6938), .Z(c[208]) );
  NANDN U7066 ( .A(n6866), .B(n6865), .Z(n6870) );
  NANDN U7067 ( .A(n6868), .B(n6867), .Z(n6869) );
  AND U7068 ( .A(n6870), .B(n6869), .Z(n6945) );
  NANDN U7069 ( .A(n6872), .B(n6871), .Z(n6876) );
  NAND U7070 ( .A(n6874), .B(n6873), .Z(n6875) );
  AND U7071 ( .A(n6876), .B(n6875), .Z(n7011) );
  NANDN U7072 ( .A(n6878), .B(n6877), .Z(n6882) );
  NANDN U7073 ( .A(n6880), .B(n6879), .Z(n6881) );
  AND U7074 ( .A(n6882), .B(n6881), .Z(n6977) );
  NANDN U7075 ( .A(n9891), .B(n6883), .Z(n6885) );
  XOR U7076 ( .A(b[13]), .B(a[85]), .Z(n6963) );
  NANDN U7077 ( .A(n9935), .B(n6963), .Z(n6884) );
  AND U7078 ( .A(n6885), .B(n6884), .Z(n6955) );
  AND U7079 ( .A(b[15]), .B(a[81]), .Z(n6954) );
  XNOR U7080 ( .A(n6955), .B(n6954), .Z(n6956) );
  NAND U7081 ( .A(b[0]), .B(a[97]), .Z(n6886) );
  XNOR U7082 ( .A(b[1]), .B(n6886), .Z(n6888) );
  NANDN U7083 ( .A(b[0]), .B(a[96]), .Z(n6887) );
  NAND U7084 ( .A(n6888), .B(n6887), .Z(n6957) );
  XNOR U7085 ( .A(n6956), .B(n6957), .Z(n6975) );
  NANDN U7086 ( .A(n9437), .B(n6889), .Z(n6891) );
  XOR U7087 ( .A(b[5]), .B(a[93]), .Z(n6966) );
  NANDN U7088 ( .A(n9503), .B(n6966), .Z(n6890) );
  AND U7089 ( .A(n6891), .B(n6890), .Z(n6999) );
  NANDN U7090 ( .A(n9588), .B(n6892), .Z(n6894) );
  XOR U7091 ( .A(b[7]), .B(a[91]), .Z(n6969) );
  NANDN U7092 ( .A(n9639), .B(n6969), .Z(n6893) );
  AND U7093 ( .A(n6894), .B(n6893), .Z(n6997) );
  NANDN U7094 ( .A(n9374), .B(n6895), .Z(n6897) );
  XOR U7095 ( .A(b[3]), .B(a[95]), .Z(n6972) );
  NANDN U7096 ( .A(n9375), .B(n6972), .Z(n6896) );
  NAND U7097 ( .A(n6897), .B(n6896), .Z(n6996) );
  XNOR U7098 ( .A(n6997), .B(n6996), .Z(n6998) );
  XOR U7099 ( .A(n6999), .B(n6998), .Z(n6976) );
  XOR U7100 ( .A(n6975), .B(n6976), .Z(n6978) );
  XOR U7101 ( .A(n6977), .B(n6978), .Z(n6949) );
  NANDN U7102 ( .A(n6899), .B(n6898), .Z(n6903) );
  OR U7103 ( .A(n6901), .B(n6900), .Z(n6902) );
  AND U7104 ( .A(n6903), .B(n6902), .Z(n6948) );
  XNOR U7105 ( .A(n6949), .B(n6948), .Z(n6951) );
  NAND U7106 ( .A(n6904), .B(n9883), .Z(n6906) );
  XOR U7107 ( .A(b[11]), .B(a[87]), .Z(n6981) );
  NANDN U7108 ( .A(n9856), .B(n6981), .Z(n6905) );
  AND U7109 ( .A(n6906), .B(n6905), .Z(n6992) );
  NANDN U7110 ( .A(n10005), .B(n6907), .Z(n6909) );
  XOR U7111 ( .A(b[15]), .B(a[83]), .Z(n6984) );
  NANDN U7112 ( .A(n10006), .B(n6984), .Z(n6908) );
  AND U7113 ( .A(n6909), .B(n6908), .Z(n6991) );
  NANDN U7114 ( .A(n9685), .B(n6910), .Z(n6912) );
  XOR U7115 ( .A(b[9]), .B(a[89]), .Z(n6987) );
  NANDN U7116 ( .A(n9758), .B(n6987), .Z(n6911) );
  NAND U7117 ( .A(n6912), .B(n6911), .Z(n6990) );
  XOR U7118 ( .A(n6991), .B(n6990), .Z(n6993) );
  XOR U7119 ( .A(n6992), .B(n6993), .Z(n7003) );
  NANDN U7120 ( .A(n6914), .B(n6913), .Z(n6918) );
  OR U7121 ( .A(n6916), .B(n6915), .Z(n6917) );
  AND U7122 ( .A(n6918), .B(n6917), .Z(n7002) );
  XNOR U7123 ( .A(n7003), .B(n7002), .Z(n7004) );
  NANDN U7124 ( .A(n6920), .B(n6919), .Z(n6924) );
  NANDN U7125 ( .A(n6922), .B(n6921), .Z(n6923) );
  NAND U7126 ( .A(n6924), .B(n6923), .Z(n7005) );
  XNOR U7127 ( .A(n7004), .B(n7005), .Z(n6950) );
  XOR U7128 ( .A(n6951), .B(n6950), .Z(n7009) );
  NANDN U7129 ( .A(n6926), .B(n6925), .Z(n6930) );
  NANDN U7130 ( .A(n6928), .B(n6927), .Z(n6929) );
  AND U7131 ( .A(n6930), .B(n6929), .Z(n7008) );
  XNOR U7132 ( .A(n7009), .B(n7008), .Z(n7010) );
  XOR U7133 ( .A(n7011), .B(n7010), .Z(n6943) );
  NANDN U7134 ( .A(n6932), .B(n6931), .Z(n6936) );
  NAND U7135 ( .A(n6934), .B(n6933), .Z(n6935) );
  AND U7136 ( .A(n6936), .B(n6935), .Z(n6942) );
  XNOR U7137 ( .A(n6943), .B(n6942), .Z(n6944) );
  XNOR U7138 ( .A(n6945), .B(n6944), .Z(n7014) );
  XNOR U7139 ( .A(sreg[209]), .B(n7014), .Z(n7016) );
  NANDN U7140 ( .A(sreg[208]), .B(n6937), .Z(n6941) );
  NAND U7141 ( .A(n6939), .B(n6938), .Z(n6940) );
  NAND U7142 ( .A(n6941), .B(n6940), .Z(n7015) );
  XNOR U7143 ( .A(n7016), .B(n7015), .Z(c[209]) );
  NANDN U7144 ( .A(n6943), .B(n6942), .Z(n6947) );
  NANDN U7145 ( .A(n6945), .B(n6944), .Z(n6946) );
  AND U7146 ( .A(n6947), .B(n6946), .Z(n7022) );
  NANDN U7147 ( .A(n6949), .B(n6948), .Z(n6953) );
  NAND U7148 ( .A(n6951), .B(n6950), .Z(n6952) );
  AND U7149 ( .A(n6953), .B(n6952), .Z(n7088) );
  NANDN U7150 ( .A(n6955), .B(n6954), .Z(n6959) );
  NANDN U7151 ( .A(n6957), .B(n6956), .Z(n6958) );
  AND U7152 ( .A(n6959), .B(n6958), .Z(n7075) );
  NAND U7153 ( .A(b[0]), .B(a[98]), .Z(n6960) );
  XNOR U7154 ( .A(b[1]), .B(n6960), .Z(n6962) );
  NANDN U7155 ( .A(b[0]), .B(a[97]), .Z(n6961) );
  NAND U7156 ( .A(n6962), .B(n6961), .Z(n7055) );
  NANDN U7157 ( .A(n9891), .B(n6963), .Z(n6965) );
  XOR U7158 ( .A(b[13]), .B(a[86]), .Z(n7058) );
  NANDN U7159 ( .A(n9935), .B(n7058), .Z(n6964) );
  AND U7160 ( .A(n6965), .B(n6964), .Z(n7053) );
  AND U7161 ( .A(b[15]), .B(a[82]), .Z(n7052) );
  XNOR U7162 ( .A(n7053), .B(n7052), .Z(n7054) );
  XNOR U7163 ( .A(n7055), .B(n7054), .Z(n7073) );
  NANDN U7164 ( .A(n9437), .B(n6966), .Z(n6968) );
  XOR U7165 ( .A(b[5]), .B(a[94]), .Z(n7064) );
  NANDN U7166 ( .A(n9503), .B(n7064), .Z(n6967) );
  AND U7167 ( .A(n6968), .B(n6967), .Z(n7049) );
  NANDN U7168 ( .A(n9588), .B(n6969), .Z(n6971) );
  XOR U7169 ( .A(b[7]), .B(a[92]), .Z(n7067) );
  NANDN U7170 ( .A(n9639), .B(n7067), .Z(n6970) );
  AND U7171 ( .A(n6971), .B(n6970), .Z(n7047) );
  NANDN U7172 ( .A(n9374), .B(n6972), .Z(n6974) );
  XOR U7173 ( .A(b[3]), .B(a[96]), .Z(n7070) );
  NANDN U7174 ( .A(n9375), .B(n7070), .Z(n6973) );
  NAND U7175 ( .A(n6974), .B(n6973), .Z(n7046) );
  XNOR U7176 ( .A(n7047), .B(n7046), .Z(n7048) );
  XOR U7177 ( .A(n7049), .B(n7048), .Z(n7074) );
  XOR U7178 ( .A(n7073), .B(n7074), .Z(n7076) );
  XOR U7179 ( .A(n7075), .B(n7076), .Z(n7026) );
  NANDN U7180 ( .A(n6976), .B(n6975), .Z(n6980) );
  OR U7181 ( .A(n6978), .B(n6977), .Z(n6979) );
  AND U7182 ( .A(n6980), .B(n6979), .Z(n7025) );
  XNOR U7183 ( .A(n7026), .B(n7025), .Z(n7028) );
  NAND U7184 ( .A(n6981), .B(n9883), .Z(n6983) );
  XOR U7185 ( .A(b[11]), .B(a[88]), .Z(n7031) );
  NANDN U7186 ( .A(n9856), .B(n7031), .Z(n6982) );
  AND U7187 ( .A(n6983), .B(n6982), .Z(n7042) );
  NANDN U7188 ( .A(n10005), .B(n6984), .Z(n6986) );
  XOR U7189 ( .A(b[15]), .B(a[84]), .Z(n7034) );
  NANDN U7190 ( .A(n10006), .B(n7034), .Z(n6985) );
  AND U7191 ( .A(n6986), .B(n6985), .Z(n7041) );
  NANDN U7192 ( .A(n9685), .B(n6987), .Z(n6989) );
  XOR U7193 ( .A(b[9]), .B(a[90]), .Z(n7037) );
  NANDN U7194 ( .A(n9758), .B(n7037), .Z(n6988) );
  NAND U7195 ( .A(n6989), .B(n6988), .Z(n7040) );
  XOR U7196 ( .A(n7041), .B(n7040), .Z(n7043) );
  XOR U7197 ( .A(n7042), .B(n7043), .Z(n7080) );
  NANDN U7198 ( .A(n6991), .B(n6990), .Z(n6995) );
  OR U7199 ( .A(n6993), .B(n6992), .Z(n6994) );
  AND U7200 ( .A(n6995), .B(n6994), .Z(n7079) );
  XNOR U7201 ( .A(n7080), .B(n7079), .Z(n7081) );
  NANDN U7202 ( .A(n6997), .B(n6996), .Z(n7001) );
  NANDN U7203 ( .A(n6999), .B(n6998), .Z(n7000) );
  NAND U7204 ( .A(n7001), .B(n7000), .Z(n7082) );
  XNOR U7205 ( .A(n7081), .B(n7082), .Z(n7027) );
  XOR U7206 ( .A(n7028), .B(n7027), .Z(n7086) );
  NANDN U7207 ( .A(n7003), .B(n7002), .Z(n7007) );
  NANDN U7208 ( .A(n7005), .B(n7004), .Z(n7006) );
  AND U7209 ( .A(n7007), .B(n7006), .Z(n7085) );
  XNOR U7210 ( .A(n7086), .B(n7085), .Z(n7087) );
  XOR U7211 ( .A(n7088), .B(n7087), .Z(n7020) );
  NANDN U7212 ( .A(n7009), .B(n7008), .Z(n7013) );
  NAND U7213 ( .A(n7011), .B(n7010), .Z(n7012) );
  AND U7214 ( .A(n7013), .B(n7012), .Z(n7019) );
  XNOR U7215 ( .A(n7020), .B(n7019), .Z(n7021) );
  XNOR U7216 ( .A(n7022), .B(n7021), .Z(n7091) );
  XNOR U7217 ( .A(sreg[210]), .B(n7091), .Z(n7093) );
  NANDN U7218 ( .A(sreg[209]), .B(n7014), .Z(n7018) );
  NAND U7219 ( .A(n7016), .B(n7015), .Z(n7017) );
  NAND U7220 ( .A(n7018), .B(n7017), .Z(n7092) );
  XNOR U7221 ( .A(n7093), .B(n7092), .Z(c[210]) );
  NANDN U7222 ( .A(n7020), .B(n7019), .Z(n7024) );
  NANDN U7223 ( .A(n7022), .B(n7021), .Z(n7023) );
  AND U7224 ( .A(n7024), .B(n7023), .Z(n7099) );
  NANDN U7225 ( .A(n7026), .B(n7025), .Z(n7030) );
  NAND U7226 ( .A(n7028), .B(n7027), .Z(n7029) );
  AND U7227 ( .A(n7030), .B(n7029), .Z(n7165) );
  NAND U7228 ( .A(n7031), .B(n9883), .Z(n7033) );
  XOR U7229 ( .A(b[11]), .B(a[89]), .Z(n7135) );
  NANDN U7230 ( .A(n9856), .B(n7135), .Z(n7032) );
  AND U7231 ( .A(n7033), .B(n7032), .Z(n7146) );
  NANDN U7232 ( .A(n10005), .B(n7034), .Z(n7036) );
  XOR U7233 ( .A(b[15]), .B(a[85]), .Z(n7138) );
  NANDN U7234 ( .A(n10006), .B(n7138), .Z(n7035) );
  AND U7235 ( .A(n7036), .B(n7035), .Z(n7145) );
  NANDN U7236 ( .A(n9685), .B(n7037), .Z(n7039) );
  XOR U7237 ( .A(b[9]), .B(a[91]), .Z(n7141) );
  NANDN U7238 ( .A(n9758), .B(n7141), .Z(n7038) );
  NAND U7239 ( .A(n7039), .B(n7038), .Z(n7144) );
  XOR U7240 ( .A(n7145), .B(n7144), .Z(n7147) );
  XOR U7241 ( .A(n7146), .B(n7147), .Z(n7157) );
  NANDN U7242 ( .A(n7041), .B(n7040), .Z(n7045) );
  OR U7243 ( .A(n7043), .B(n7042), .Z(n7044) );
  AND U7244 ( .A(n7045), .B(n7044), .Z(n7156) );
  XNOR U7245 ( .A(n7157), .B(n7156), .Z(n7158) );
  NANDN U7246 ( .A(n7047), .B(n7046), .Z(n7051) );
  NANDN U7247 ( .A(n7049), .B(n7048), .Z(n7050) );
  NAND U7248 ( .A(n7051), .B(n7050), .Z(n7159) );
  XNOR U7249 ( .A(n7158), .B(n7159), .Z(n7105) );
  NANDN U7250 ( .A(n7053), .B(n7052), .Z(n7057) );
  NANDN U7251 ( .A(n7055), .B(n7054), .Z(n7056) );
  AND U7252 ( .A(n7057), .B(n7056), .Z(n7131) );
  NANDN U7253 ( .A(n9891), .B(n7058), .Z(n7060) );
  XOR U7254 ( .A(b[13]), .B(a[87]), .Z(n7117) );
  NANDN U7255 ( .A(n9935), .B(n7117), .Z(n7059) );
  AND U7256 ( .A(n7060), .B(n7059), .Z(n7109) );
  AND U7257 ( .A(b[15]), .B(a[83]), .Z(n7108) );
  XNOR U7258 ( .A(n7109), .B(n7108), .Z(n7110) );
  NAND U7259 ( .A(b[0]), .B(a[99]), .Z(n7061) );
  XNOR U7260 ( .A(b[1]), .B(n7061), .Z(n7063) );
  NANDN U7261 ( .A(b[0]), .B(a[98]), .Z(n7062) );
  NAND U7262 ( .A(n7063), .B(n7062), .Z(n7111) );
  XNOR U7263 ( .A(n7110), .B(n7111), .Z(n7129) );
  NANDN U7264 ( .A(n9437), .B(n7064), .Z(n7066) );
  XOR U7265 ( .A(b[5]), .B(a[95]), .Z(n7120) );
  NANDN U7266 ( .A(n9503), .B(n7120), .Z(n7065) );
  AND U7267 ( .A(n7066), .B(n7065), .Z(n7153) );
  NANDN U7268 ( .A(n9588), .B(n7067), .Z(n7069) );
  XOR U7269 ( .A(b[7]), .B(a[93]), .Z(n7123) );
  NANDN U7270 ( .A(n9639), .B(n7123), .Z(n7068) );
  AND U7271 ( .A(n7069), .B(n7068), .Z(n7151) );
  NANDN U7272 ( .A(n9374), .B(n7070), .Z(n7072) );
  XOR U7273 ( .A(b[3]), .B(a[97]), .Z(n7126) );
  NANDN U7274 ( .A(n9375), .B(n7126), .Z(n7071) );
  NAND U7275 ( .A(n7072), .B(n7071), .Z(n7150) );
  XNOR U7276 ( .A(n7151), .B(n7150), .Z(n7152) );
  XOR U7277 ( .A(n7153), .B(n7152), .Z(n7130) );
  XOR U7278 ( .A(n7129), .B(n7130), .Z(n7132) );
  XOR U7279 ( .A(n7131), .B(n7132), .Z(n7103) );
  NANDN U7280 ( .A(n7074), .B(n7073), .Z(n7078) );
  OR U7281 ( .A(n7076), .B(n7075), .Z(n7077) );
  AND U7282 ( .A(n7078), .B(n7077), .Z(n7102) );
  XNOR U7283 ( .A(n7103), .B(n7102), .Z(n7104) );
  XOR U7284 ( .A(n7105), .B(n7104), .Z(n7163) );
  NANDN U7285 ( .A(n7080), .B(n7079), .Z(n7084) );
  NANDN U7286 ( .A(n7082), .B(n7081), .Z(n7083) );
  AND U7287 ( .A(n7084), .B(n7083), .Z(n7162) );
  XNOR U7288 ( .A(n7163), .B(n7162), .Z(n7164) );
  XOR U7289 ( .A(n7165), .B(n7164), .Z(n7097) );
  NANDN U7290 ( .A(n7086), .B(n7085), .Z(n7090) );
  NAND U7291 ( .A(n7088), .B(n7087), .Z(n7089) );
  AND U7292 ( .A(n7090), .B(n7089), .Z(n7096) );
  XNOR U7293 ( .A(n7097), .B(n7096), .Z(n7098) );
  XNOR U7294 ( .A(n7099), .B(n7098), .Z(n7168) );
  XNOR U7295 ( .A(sreg[211]), .B(n7168), .Z(n7170) );
  NANDN U7296 ( .A(sreg[210]), .B(n7091), .Z(n7095) );
  NAND U7297 ( .A(n7093), .B(n7092), .Z(n7094) );
  NAND U7298 ( .A(n7095), .B(n7094), .Z(n7169) );
  XNOR U7299 ( .A(n7170), .B(n7169), .Z(c[211]) );
  NANDN U7300 ( .A(n7097), .B(n7096), .Z(n7101) );
  NANDN U7301 ( .A(n7099), .B(n7098), .Z(n7100) );
  AND U7302 ( .A(n7101), .B(n7100), .Z(n7176) );
  NANDN U7303 ( .A(n7103), .B(n7102), .Z(n7107) );
  NAND U7304 ( .A(n7105), .B(n7104), .Z(n7106) );
  AND U7305 ( .A(n7107), .B(n7106), .Z(n7242) );
  NANDN U7306 ( .A(n7109), .B(n7108), .Z(n7113) );
  NANDN U7307 ( .A(n7111), .B(n7110), .Z(n7112) );
  AND U7308 ( .A(n7113), .B(n7112), .Z(n7208) );
  NAND U7309 ( .A(b[0]), .B(a[100]), .Z(n7114) );
  XNOR U7310 ( .A(b[1]), .B(n7114), .Z(n7116) );
  NANDN U7311 ( .A(b[0]), .B(a[99]), .Z(n7115) );
  NAND U7312 ( .A(n7116), .B(n7115), .Z(n7188) );
  NANDN U7313 ( .A(n9891), .B(n7117), .Z(n7119) );
  XOR U7314 ( .A(b[13]), .B(a[88]), .Z(n7194) );
  NANDN U7315 ( .A(n9935), .B(n7194), .Z(n7118) );
  AND U7316 ( .A(n7119), .B(n7118), .Z(n7186) );
  AND U7317 ( .A(b[15]), .B(a[84]), .Z(n7185) );
  XNOR U7318 ( .A(n7186), .B(n7185), .Z(n7187) );
  XNOR U7319 ( .A(n7188), .B(n7187), .Z(n7206) );
  NANDN U7320 ( .A(n9437), .B(n7120), .Z(n7122) );
  XOR U7321 ( .A(b[5]), .B(a[96]), .Z(n7197) );
  NANDN U7322 ( .A(n9503), .B(n7197), .Z(n7121) );
  AND U7323 ( .A(n7122), .B(n7121), .Z(n7230) );
  NANDN U7324 ( .A(n9588), .B(n7123), .Z(n7125) );
  XOR U7325 ( .A(b[7]), .B(a[94]), .Z(n7200) );
  NANDN U7326 ( .A(n9639), .B(n7200), .Z(n7124) );
  AND U7327 ( .A(n7125), .B(n7124), .Z(n7228) );
  NANDN U7328 ( .A(n9374), .B(n7126), .Z(n7128) );
  XOR U7329 ( .A(b[3]), .B(a[98]), .Z(n7203) );
  NANDN U7330 ( .A(n9375), .B(n7203), .Z(n7127) );
  NAND U7331 ( .A(n7128), .B(n7127), .Z(n7227) );
  XNOR U7332 ( .A(n7228), .B(n7227), .Z(n7229) );
  XOR U7333 ( .A(n7230), .B(n7229), .Z(n7207) );
  XOR U7334 ( .A(n7206), .B(n7207), .Z(n7209) );
  XOR U7335 ( .A(n7208), .B(n7209), .Z(n7180) );
  NANDN U7336 ( .A(n7130), .B(n7129), .Z(n7134) );
  OR U7337 ( .A(n7132), .B(n7131), .Z(n7133) );
  AND U7338 ( .A(n7134), .B(n7133), .Z(n7179) );
  XNOR U7339 ( .A(n7180), .B(n7179), .Z(n7182) );
  NAND U7340 ( .A(n7135), .B(n9883), .Z(n7137) );
  XOR U7341 ( .A(b[11]), .B(a[90]), .Z(n7212) );
  NANDN U7342 ( .A(n9856), .B(n7212), .Z(n7136) );
  AND U7343 ( .A(n7137), .B(n7136), .Z(n7223) );
  NANDN U7344 ( .A(n10005), .B(n7138), .Z(n7140) );
  XOR U7345 ( .A(b[15]), .B(a[86]), .Z(n7215) );
  NANDN U7346 ( .A(n10006), .B(n7215), .Z(n7139) );
  AND U7347 ( .A(n7140), .B(n7139), .Z(n7222) );
  NANDN U7348 ( .A(n9685), .B(n7141), .Z(n7143) );
  XOR U7349 ( .A(b[9]), .B(a[92]), .Z(n7218) );
  NANDN U7350 ( .A(n9758), .B(n7218), .Z(n7142) );
  NAND U7351 ( .A(n7143), .B(n7142), .Z(n7221) );
  XOR U7352 ( .A(n7222), .B(n7221), .Z(n7224) );
  XOR U7353 ( .A(n7223), .B(n7224), .Z(n7234) );
  NANDN U7354 ( .A(n7145), .B(n7144), .Z(n7149) );
  OR U7355 ( .A(n7147), .B(n7146), .Z(n7148) );
  AND U7356 ( .A(n7149), .B(n7148), .Z(n7233) );
  XNOR U7357 ( .A(n7234), .B(n7233), .Z(n7235) );
  NANDN U7358 ( .A(n7151), .B(n7150), .Z(n7155) );
  NANDN U7359 ( .A(n7153), .B(n7152), .Z(n7154) );
  NAND U7360 ( .A(n7155), .B(n7154), .Z(n7236) );
  XNOR U7361 ( .A(n7235), .B(n7236), .Z(n7181) );
  XOR U7362 ( .A(n7182), .B(n7181), .Z(n7240) );
  NANDN U7363 ( .A(n7157), .B(n7156), .Z(n7161) );
  NANDN U7364 ( .A(n7159), .B(n7158), .Z(n7160) );
  AND U7365 ( .A(n7161), .B(n7160), .Z(n7239) );
  XNOR U7366 ( .A(n7240), .B(n7239), .Z(n7241) );
  XOR U7367 ( .A(n7242), .B(n7241), .Z(n7174) );
  NANDN U7368 ( .A(n7163), .B(n7162), .Z(n7167) );
  NAND U7369 ( .A(n7165), .B(n7164), .Z(n7166) );
  AND U7370 ( .A(n7167), .B(n7166), .Z(n7173) );
  XNOR U7371 ( .A(n7174), .B(n7173), .Z(n7175) );
  XNOR U7372 ( .A(n7176), .B(n7175), .Z(n7245) );
  XNOR U7373 ( .A(sreg[212]), .B(n7245), .Z(n7247) );
  NANDN U7374 ( .A(sreg[211]), .B(n7168), .Z(n7172) );
  NAND U7375 ( .A(n7170), .B(n7169), .Z(n7171) );
  NAND U7376 ( .A(n7172), .B(n7171), .Z(n7246) );
  XNOR U7377 ( .A(n7247), .B(n7246), .Z(c[212]) );
  NANDN U7378 ( .A(n7174), .B(n7173), .Z(n7178) );
  NANDN U7379 ( .A(n7176), .B(n7175), .Z(n7177) );
  AND U7380 ( .A(n7178), .B(n7177), .Z(n7253) );
  NANDN U7381 ( .A(n7180), .B(n7179), .Z(n7184) );
  NAND U7382 ( .A(n7182), .B(n7181), .Z(n7183) );
  AND U7383 ( .A(n7184), .B(n7183), .Z(n7319) );
  NANDN U7384 ( .A(n7186), .B(n7185), .Z(n7190) );
  NANDN U7385 ( .A(n7188), .B(n7187), .Z(n7189) );
  AND U7386 ( .A(n7190), .B(n7189), .Z(n7285) );
  NAND U7387 ( .A(b[0]), .B(a[101]), .Z(n7191) );
  XNOR U7388 ( .A(b[1]), .B(n7191), .Z(n7193) );
  NANDN U7389 ( .A(b[0]), .B(a[100]), .Z(n7192) );
  NAND U7390 ( .A(n7193), .B(n7192), .Z(n7265) );
  NANDN U7391 ( .A(n9891), .B(n7194), .Z(n7196) );
  XOR U7392 ( .A(b[13]), .B(a[89]), .Z(n7268) );
  NANDN U7393 ( .A(n9935), .B(n7268), .Z(n7195) );
  AND U7394 ( .A(n7196), .B(n7195), .Z(n7263) );
  AND U7395 ( .A(b[15]), .B(a[85]), .Z(n7262) );
  XNOR U7396 ( .A(n7263), .B(n7262), .Z(n7264) );
  XNOR U7397 ( .A(n7265), .B(n7264), .Z(n7283) );
  NANDN U7398 ( .A(n9437), .B(n7197), .Z(n7199) );
  XOR U7399 ( .A(b[5]), .B(a[97]), .Z(n7274) );
  NANDN U7400 ( .A(n9503), .B(n7274), .Z(n7198) );
  AND U7401 ( .A(n7199), .B(n7198), .Z(n7307) );
  NANDN U7402 ( .A(n9588), .B(n7200), .Z(n7202) );
  XOR U7403 ( .A(b[7]), .B(a[95]), .Z(n7277) );
  NANDN U7404 ( .A(n9639), .B(n7277), .Z(n7201) );
  AND U7405 ( .A(n7202), .B(n7201), .Z(n7305) );
  NANDN U7406 ( .A(n9374), .B(n7203), .Z(n7205) );
  XOR U7407 ( .A(b[3]), .B(a[99]), .Z(n7280) );
  NANDN U7408 ( .A(n9375), .B(n7280), .Z(n7204) );
  NAND U7409 ( .A(n7205), .B(n7204), .Z(n7304) );
  XNOR U7410 ( .A(n7305), .B(n7304), .Z(n7306) );
  XOR U7411 ( .A(n7307), .B(n7306), .Z(n7284) );
  XOR U7412 ( .A(n7283), .B(n7284), .Z(n7286) );
  XOR U7413 ( .A(n7285), .B(n7286), .Z(n7257) );
  NANDN U7414 ( .A(n7207), .B(n7206), .Z(n7211) );
  OR U7415 ( .A(n7209), .B(n7208), .Z(n7210) );
  AND U7416 ( .A(n7211), .B(n7210), .Z(n7256) );
  XNOR U7417 ( .A(n7257), .B(n7256), .Z(n7259) );
  NAND U7418 ( .A(n7212), .B(n9883), .Z(n7214) );
  XOR U7419 ( .A(b[11]), .B(a[91]), .Z(n7289) );
  NANDN U7420 ( .A(n9856), .B(n7289), .Z(n7213) );
  AND U7421 ( .A(n7214), .B(n7213), .Z(n7300) );
  NANDN U7422 ( .A(n10005), .B(n7215), .Z(n7217) );
  XOR U7423 ( .A(b[15]), .B(a[87]), .Z(n7292) );
  NANDN U7424 ( .A(n10006), .B(n7292), .Z(n7216) );
  AND U7425 ( .A(n7217), .B(n7216), .Z(n7299) );
  NANDN U7426 ( .A(n9685), .B(n7218), .Z(n7220) );
  XOR U7427 ( .A(b[9]), .B(a[93]), .Z(n7295) );
  NANDN U7428 ( .A(n9758), .B(n7295), .Z(n7219) );
  NAND U7429 ( .A(n7220), .B(n7219), .Z(n7298) );
  XOR U7430 ( .A(n7299), .B(n7298), .Z(n7301) );
  XOR U7431 ( .A(n7300), .B(n7301), .Z(n7311) );
  NANDN U7432 ( .A(n7222), .B(n7221), .Z(n7226) );
  OR U7433 ( .A(n7224), .B(n7223), .Z(n7225) );
  AND U7434 ( .A(n7226), .B(n7225), .Z(n7310) );
  XNOR U7435 ( .A(n7311), .B(n7310), .Z(n7312) );
  NANDN U7436 ( .A(n7228), .B(n7227), .Z(n7232) );
  NANDN U7437 ( .A(n7230), .B(n7229), .Z(n7231) );
  NAND U7438 ( .A(n7232), .B(n7231), .Z(n7313) );
  XNOR U7439 ( .A(n7312), .B(n7313), .Z(n7258) );
  XOR U7440 ( .A(n7259), .B(n7258), .Z(n7317) );
  NANDN U7441 ( .A(n7234), .B(n7233), .Z(n7238) );
  NANDN U7442 ( .A(n7236), .B(n7235), .Z(n7237) );
  AND U7443 ( .A(n7238), .B(n7237), .Z(n7316) );
  XNOR U7444 ( .A(n7317), .B(n7316), .Z(n7318) );
  XOR U7445 ( .A(n7319), .B(n7318), .Z(n7251) );
  NANDN U7446 ( .A(n7240), .B(n7239), .Z(n7244) );
  NAND U7447 ( .A(n7242), .B(n7241), .Z(n7243) );
  AND U7448 ( .A(n7244), .B(n7243), .Z(n7250) );
  XNOR U7449 ( .A(n7251), .B(n7250), .Z(n7252) );
  XNOR U7450 ( .A(n7253), .B(n7252), .Z(n7322) );
  XNOR U7451 ( .A(sreg[213]), .B(n7322), .Z(n7324) );
  NANDN U7452 ( .A(sreg[212]), .B(n7245), .Z(n7249) );
  NAND U7453 ( .A(n7247), .B(n7246), .Z(n7248) );
  NAND U7454 ( .A(n7249), .B(n7248), .Z(n7323) );
  XNOR U7455 ( .A(n7324), .B(n7323), .Z(c[213]) );
  NANDN U7456 ( .A(n7251), .B(n7250), .Z(n7255) );
  NANDN U7457 ( .A(n7253), .B(n7252), .Z(n7254) );
  AND U7458 ( .A(n7255), .B(n7254), .Z(n7330) );
  NANDN U7459 ( .A(n7257), .B(n7256), .Z(n7261) );
  NAND U7460 ( .A(n7259), .B(n7258), .Z(n7260) );
  AND U7461 ( .A(n7261), .B(n7260), .Z(n7396) );
  NANDN U7462 ( .A(n7263), .B(n7262), .Z(n7267) );
  NANDN U7463 ( .A(n7265), .B(n7264), .Z(n7266) );
  AND U7464 ( .A(n7267), .B(n7266), .Z(n7362) );
  NANDN U7465 ( .A(n9891), .B(n7268), .Z(n7270) );
  XOR U7466 ( .A(b[13]), .B(a[90]), .Z(n7348) );
  NANDN U7467 ( .A(n9935), .B(n7348), .Z(n7269) );
  AND U7468 ( .A(n7270), .B(n7269), .Z(n7340) );
  AND U7469 ( .A(b[15]), .B(a[86]), .Z(n7339) );
  XNOR U7470 ( .A(n7340), .B(n7339), .Z(n7341) );
  NAND U7471 ( .A(b[0]), .B(a[102]), .Z(n7271) );
  XNOR U7472 ( .A(b[1]), .B(n7271), .Z(n7273) );
  NANDN U7473 ( .A(b[0]), .B(a[101]), .Z(n7272) );
  NAND U7474 ( .A(n7273), .B(n7272), .Z(n7342) );
  XNOR U7475 ( .A(n7341), .B(n7342), .Z(n7360) );
  NANDN U7476 ( .A(n9437), .B(n7274), .Z(n7276) );
  XOR U7477 ( .A(b[5]), .B(a[98]), .Z(n7351) );
  NANDN U7478 ( .A(n9503), .B(n7351), .Z(n7275) );
  AND U7479 ( .A(n7276), .B(n7275), .Z(n7384) );
  NANDN U7480 ( .A(n9588), .B(n7277), .Z(n7279) );
  XOR U7481 ( .A(b[7]), .B(a[96]), .Z(n7354) );
  NANDN U7482 ( .A(n9639), .B(n7354), .Z(n7278) );
  AND U7483 ( .A(n7279), .B(n7278), .Z(n7382) );
  NANDN U7484 ( .A(n9374), .B(n7280), .Z(n7282) );
  XOR U7485 ( .A(b[3]), .B(a[100]), .Z(n7357) );
  NANDN U7486 ( .A(n9375), .B(n7357), .Z(n7281) );
  NAND U7487 ( .A(n7282), .B(n7281), .Z(n7381) );
  XNOR U7488 ( .A(n7382), .B(n7381), .Z(n7383) );
  XOR U7489 ( .A(n7384), .B(n7383), .Z(n7361) );
  XOR U7490 ( .A(n7360), .B(n7361), .Z(n7363) );
  XOR U7491 ( .A(n7362), .B(n7363), .Z(n7334) );
  NANDN U7492 ( .A(n7284), .B(n7283), .Z(n7288) );
  OR U7493 ( .A(n7286), .B(n7285), .Z(n7287) );
  AND U7494 ( .A(n7288), .B(n7287), .Z(n7333) );
  XNOR U7495 ( .A(n7334), .B(n7333), .Z(n7336) );
  NAND U7496 ( .A(n7289), .B(n9883), .Z(n7291) );
  XOR U7497 ( .A(b[11]), .B(a[92]), .Z(n7366) );
  NANDN U7498 ( .A(n9856), .B(n7366), .Z(n7290) );
  AND U7499 ( .A(n7291), .B(n7290), .Z(n7377) );
  NANDN U7500 ( .A(n10005), .B(n7292), .Z(n7294) );
  XOR U7501 ( .A(b[15]), .B(a[88]), .Z(n7369) );
  NANDN U7502 ( .A(n10006), .B(n7369), .Z(n7293) );
  AND U7503 ( .A(n7294), .B(n7293), .Z(n7376) );
  NANDN U7504 ( .A(n9685), .B(n7295), .Z(n7297) );
  XOR U7505 ( .A(b[9]), .B(a[94]), .Z(n7372) );
  NANDN U7506 ( .A(n9758), .B(n7372), .Z(n7296) );
  NAND U7507 ( .A(n7297), .B(n7296), .Z(n7375) );
  XOR U7508 ( .A(n7376), .B(n7375), .Z(n7378) );
  XOR U7509 ( .A(n7377), .B(n7378), .Z(n7388) );
  NANDN U7510 ( .A(n7299), .B(n7298), .Z(n7303) );
  OR U7511 ( .A(n7301), .B(n7300), .Z(n7302) );
  AND U7512 ( .A(n7303), .B(n7302), .Z(n7387) );
  XNOR U7513 ( .A(n7388), .B(n7387), .Z(n7389) );
  NANDN U7514 ( .A(n7305), .B(n7304), .Z(n7309) );
  NANDN U7515 ( .A(n7307), .B(n7306), .Z(n7308) );
  NAND U7516 ( .A(n7309), .B(n7308), .Z(n7390) );
  XNOR U7517 ( .A(n7389), .B(n7390), .Z(n7335) );
  XOR U7518 ( .A(n7336), .B(n7335), .Z(n7394) );
  NANDN U7519 ( .A(n7311), .B(n7310), .Z(n7315) );
  NANDN U7520 ( .A(n7313), .B(n7312), .Z(n7314) );
  AND U7521 ( .A(n7315), .B(n7314), .Z(n7393) );
  XNOR U7522 ( .A(n7394), .B(n7393), .Z(n7395) );
  XOR U7523 ( .A(n7396), .B(n7395), .Z(n7328) );
  NANDN U7524 ( .A(n7317), .B(n7316), .Z(n7321) );
  NAND U7525 ( .A(n7319), .B(n7318), .Z(n7320) );
  AND U7526 ( .A(n7321), .B(n7320), .Z(n7327) );
  XNOR U7527 ( .A(n7328), .B(n7327), .Z(n7329) );
  XNOR U7528 ( .A(n7330), .B(n7329), .Z(n7399) );
  XNOR U7529 ( .A(sreg[214]), .B(n7399), .Z(n7401) );
  NANDN U7530 ( .A(sreg[213]), .B(n7322), .Z(n7326) );
  NAND U7531 ( .A(n7324), .B(n7323), .Z(n7325) );
  NAND U7532 ( .A(n7326), .B(n7325), .Z(n7400) );
  XNOR U7533 ( .A(n7401), .B(n7400), .Z(c[214]) );
  NANDN U7534 ( .A(n7328), .B(n7327), .Z(n7332) );
  NANDN U7535 ( .A(n7330), .B(n7329), .Z(n7331) );
  AND U7536 ( .A(n7332), .B(n7331), .Z(n7407) );
  NANDN U7537 ( .A(n7334), .B(n7333), .Z(n7338) );
  NAND U7538 ( .A(n7336), .B(n7335), .Z(n7337) );
  AND U7539 ( .A(n7338), .B(n7337), .Z(n7473) );
  NANDN U7540 ( .A(n7340), .B(n7339), .Z(n7344) );
  NANDN U7541 ( .A(n7342), .B(n7341), .Z(n7343) );
  AND U7542 ( .A(n7344), .B(n7343), .Z(n7439) );
  NAND U7543 ( .A(b[0]), .B(a[103]), .Z(n7345) );
  XNOR U7544 ( .A(b[1]), .B(n7345), .Z(n7347) );
  NANDN U7545 ( .A(b[0]), .B(a[102]), .Z(n7346) );
  NAND U7546 ( .A(n7347), .B(n7346), .Z(n7419) );
  NANDN U7547 ( .A(n9891), .B(n7348), .Z(n7350) );
  XOR U7548 ( .A(b[13]), .B(a[91]), .Z(n7422) );
  NANDN U7549 ( .A(n9935), .B(n7422), .Z(n7349) );
  AND U7550 ( .A(n7350), .B(n7349), .Z(n7417) );
  AND U7551 ( .A(b[15]), .B(a[87]), .Z(n7416) );
  XNOR U7552 ( .A(n7417), .B(n7416), .Z(n7418) );
  XNOR U7553 ( .A(n7419), .B(n7418), .Z(n7437) );
  NANDN U7554 ( .A(n9437), .B(n7351), .Z(n7353) );
  XOR U7555 ( .A(b[5]), .B(a[99]), .Z(n7428) );
  NANDN U7556 ( .A(n9503), .B(n7428), .Z(n7352) );
  AND U7557 ( .A(n7353), .B(n7352), .Z(n7461) );
  NANDN U7558 ( .A(n9588), .B(n7354), .Z(n7356) );
  XOR U7559 ( .A(b[7]), .B(a[97]), .Z(n7431) );
  NANDN U7560 ( .A(n9639), .B(n7431), .Z(n7355) );
  AND U7561 ( .A(n7356), .B(n7355), .Z(n7459) );
  NANDN U7562 ( .A(n9374), .B(n7357), .Z(n7359) );
  XOR U7563 ( .A(b[3]), .B(a[101]), .Z(n7434) );
  NANDN U7564 ( .A(n9375), .B(n7434), .Z(n7358) );
  NAND U7565 ( .A(n7359), .B(n7358), .Z(n7458) );
  XNOR U7566 ( .A(n7459), .B(n7458), .Z(n7460) );
  XOR U7567 ( .A(n7461), .B(n7460), .Z(n7438) );
  XOR U7568 ( .A(n7437), .B(n7438), .Z(n7440) );
  XOR U7569 ( .A(n7439), .B(n7440), .Z(n7411) );
  NANDN U7570 ( .A(n7361), .B(n7360), .Z(n7365) );
  OR U7571 ( .A(n7363), .B(n7362), .Z(n7364) );
  AND U7572 ( .A(n7365), .B(n7364), .Z(n7410) );
  XNOR U7573 ( .A(n7411), .B(n7410), .Z(n7413) );
  NAND U7574 ( .A(n7366), .B(n9883), .Z(n7368) );
  XOR U7575 ( .A(b[11]), .B(a[93]), .Z(n7443) );
  NANDN U7576 ( .A(n9856), .B(n7443), .Z(n7367) );
  AND U7577 ( .A(n7368), .B(n7367), .Z(n7454) );
  NANDN U7578 ( .A(n10005), .B(n7369), .Z(n7371) );
  XOR U7579 ( .A(b[15]), .B(a[89]), .Z(n7446) );
  NANDN U7580 ( .A(n10006), .B(n7446), .Z(n7370) );
  AND U7581 ( .A(n7371), .B(n7370), .Z(n7453) );
  NANDN U7582 ( .A(n9685), .B(n7372), .Z(n7374) );
  XOR U7583 ( .A(b[9]), .B(a[95]), .Z(n7449) );
  NANDN U7584 ( .A(n9758), .B(n7449), .Z(n7373) );
  NAND U7585 ( .A(n7374), .B(n7373), .Z(n7452) );
  XOR U7586 ( .A(n7453), .B(n7452), .Z(n7455) );
  XOR U7587 ( .A(n7454), .B(n7455), .Z(n7465) );
  NANDN U7588 ( .A(n7376), .B(n7375), .Z(n7380) );
  OR U7589 ( .A(n7378), .B(n7377), .Z(n7379) );
  AND U7590 ( .A(n7380), .B(n7379), .Z(n7464) );
  XNOR U7591 ( .A(n7465), .B(n7464), .Z(n7466) );
  NANDN U7592 ( .A(n7382), .B(n7381), .Z(n7386) );
  NANDN U7593 ( .A(n7384), .B(n7383), .Z(n7385) );
  NAND U7594 ( .A(n7386), .B(n7385), .Z(n7467) );
  XNOR U7595 ( .A(n7466), .B(n7467), .Z(n7412) );
  XOR U7596 ( .A(n7413), .B(n7412), .Z(n7471) );
  NANDN U7597 ( .A(n7388), .B(n7387), .Z(n7392) );
  NANDN U7598 ( .A(n7390), .B(n7389), .Z(n7391) );
  AND U7599 ( .A(n7392), .B(n7391), .Z(n7470) );
  XNOR U7600 ( .A(n7471), .B(n7470), .Z(n7472) );
  XOR U7601 ( .A(n7473), .B(n7472), .Z(n7405) );
  NANDN U7602 ( .A(n7394), .B(n7393), .Z(n7398) );
  NAND U7603 ( .A(n7396), .B(n7395), .Z(n7397) );
  AND U7604 ( .A(n7398), .B(n7397), .Z(n7404) );
  XNOR U7605 ( .A(n7405), .B(n7404), .Z(n7406) );
  XNOR U7606 ( .A(n7407), .B(n7406), .Z(n7476) );
  XNOR U7607 ( .A(sreg[215]), .B(n7476), .Z(n7478) );
  NANDN U7608 ( .A(sreg[214]), .B(n7399), .Z(n7403) );
  NAND U7609 ( .A(n7401), .B(n7400), .Z(n7402) );
  NAND U7610 ( .A(n7403), .B(n7402), .Z(n7477) );
  XNOR U7611 ( .A(n7478), .B(n7477), .Z(c[215]) );
  NANDN U7612 ( .A(n7405), .B(n7404), .Z(n7409) );
  NANDN U7613 ( .A(n7407), .B(n7406), .Z(n7408) );
  AND U7614 ( .A(n7409), .B(n7408), .Z(n7484) );
  NANDN U7615 ( .A(n7411), .B(n7410), .Z(n7415) );
  NAND U7616 ( .A(n7413), .B(n7412), .Z(n7414) );
  AND U7617 ( .A(n7415), .B(n7414), .Z(n7550) );
  NANDN U7618 ( .A(n7417), .B(n7416), .Z(n7421) );
  NANDN U7619 ( .A(n7419), .B(n7418), .Z(n7420) );
  AND U7620 ( .A(n7421), .B(n7420), .Z(n7516) );
  NANDN U7621 ( .A(n9891), .B(n7422), .Z(n7424) );
  XOR U7622 ( .A(b[13]), .B(a[92]), .Z(n7502) );
  NANDN U7623 ( .A(n9935), .B(n7502), .Z(n7423) );
  AND U7624 ( .A(n7424), .B(n7423), .Z(n7494) );
  AND U7625 ( .A(b[15]), .B(a[88]), .Z(n7493) );
  XNOR U7626 ( .A(n7494), .B(n7493), .Z(n7495) );
  NAND U7627 ( .A(b[0]), .B(a[104]), .Z(n7425) );
  XNOR U7628 ( .A(b[1]), .B(n7425), .Z(n7427) );
  NANDN U7629 ( .A(b[0]), .B(a[103]), .Z(n7426) );
  NAND U7630 ( .A(n7427), .B(n7426), .Z(n7496) );
  XNOR U7631 ( .A(n7495), .B(n7496), .Z(n7514) );
  NANDN U7632 ( .A(n9437), .B(n7428), .Z(n7430) );
  XOR U7633 ( .A(b[5]), .B(a[100]), .Z(n7505) );
  NANDN U7634 ( .A(n9503), .B(n7505), .Z(n7429) );
  AND U7635 ( .A(n7430), .B(n7429), .Z(n7538) );
  NANDN U7636 ( .A(n9588), .B(n7431), .Z(n7433) );
  XOR U7637 ( .A(b[7]), .B(a[98]), .Z(n7508) );
  NANDN U7638 ( .A(n9639), .B(n7508), .Z(n7432) );
  AND U7639 ( .A(n7433), .B(n7432), .Z(n7536) );
  NANDN U7640 ( .A(n9374), .B(n7434), .Z(n7436) );
  XOR U7641 ( .A(b[3]), .B(a[102]), .Z(n7511) );
  NANDN U7642 ( .A(n9375), .B(n7511), .Z(n7435) );
  NAND U7643 ( .A(n7436), .B(n7435), .Z(n7535) );
  XNOR U7644 ( .A(n7536), .B(n7535), .Z(n7537) );
  XOR U7645 ( .A(n7538), .B(n7537), .Z(n7515) );
  XOR U7646 ( .A(n7514), .B(n7515), .Z(n7517) );
  XOR U7647 ( .A(n7516), .B(n7517), .Z(n7488) );
  NANDN U7648 ( .A(n7438), .B(n7437), .Z(n7442) );
  OR U7649 ( .A(n7440), .B(n7439), .Z(n7441) );
  AND U7650 ( .A(n7442), .B(n7441), .Z(n7487) );
  XNOR U7651 ( .A(n7488), .B(n7487), .Z(n7490) );
  NAND U7652 ( .A(n7443), .B(n9883), .Z(n7445) );
  XOR U7653 ( .A(b[11]), .B(a[94]), .Z(n7520) );
  NANDN U7654 ( .A(n9856), .B(n7520), .Z(n7444) );
  AND U7655 ( .A(n7445), .B(n7444), .Z(n7531) );
  NANDN U7656 ( .A(n10005), .B(n7446), .Z(n7448) );
  XOR U7657 ( .A(b[15]), .B(a[90]), .Z(n7523) );
  NANDN U7658 ( .A(n10006), .B(n7523), .Z(n7447) );
  AND U7659 ( .A(n7448), .B(n7447), .Z(n7530) );
  NANDN U7660 ( .A(n9685), .B(n7449), .Z(n7451) );
  XOR U7661 ( .A(b[9]), .B(a[96]), .Z(n7526) );
  NANDN U7662 ( .A(n9758), .B(n7526), .Z(n7450) );
  NAND U7663 ( .A(n7451), .B(n7450), .Z(n7529) );
  XOR U7664 ( .A(n7530), .B(n7529), .Z(n7532) );
  XOR U7665 ( .A(n7531), .B(n7532), .Z(n7542) );
  NANDN U7666 ( .A(n7453), .B(n7452), .Z(n7457) );
  OR U7667 ( .A(n7455), .B(n7454), .Z(n7456) );
  AND U7668 ( .A(n7457), .B(n7456), .Z(n7541) );
  XNOR U7669 ( .A(n7542), .B(n7541), .Z(n7543) );
  NANDN U7670 ( .A(n7459), .B(n7458), .Z(n7463) );
  NANDN U7671 ( .A(n7461), .B(n7460), .Z(n7462) );
  NAND U7672 ( .A(n7463), .B(n7462), .Z(n7544) );
  XNOR U7673 ( .A(n7543), .B(n7544), .Z(n7489) );
  XOR U7674 ( .A(n7490), .B(n7489), .Z(n7548) );
  NANDN U7675 ( .A(n7465), .B(n7464), .Z(n7469) );
  NANDN U7676 ( .A(n7467), .B(n7466), .Z(n7468) );
  AND U7677 ( .A(n7469), .B(n7468), .Z(n7547) );
  XNOR U7678 ( .A(n7548), .B(n7547), .Z(n7549) );
  XOR U7679 ( .A(n7550), .B(n7549), .Z(n7482) );
  NANDN U7680 ( .A(n7471), .B(n7470), .Z(n7475) );
  NAND U7681 ( .A(n7473), .B(n7472), .Z(n7474) );
  AND U7682 ( .A(n7475), .B(n7474), .Z(n7481) );
  XNOR U7683 ( .A(n7482), .B(n7481), .Z(n7483) );
  XNOR U7684 ( .A(n7484), .B(n7483), .Z(n7553) );
  XNOR U7685 ( .A(sreg[216]), .B(n7553), .Z(n7555) );
  NANDN U7686 ( .A(sreg[215]), .B(n7476), .Z(n7480) );
  NAND U7687 ( .A(n7478), .B(n7477), .Z(n7479) );
  NAND U7688 ( .A(n7480), .B(n7479), .Z(n7554) );
  XNOR U7689 ( .A(n7555), .B(n7554), .Z(c[216]) );
  NANDN U7690 ( .A(n7482), .B(n7481), .Z(n7486) );
  NANDN U7691 ( .A(n7484), .B(n7483), .Z(n7485) );
  AND U7692 ( .A(n7486), .B(n7485), .Z(n7561) );
  NANDN U7693 ( .A(n7488), .B(n7487), .Z(n7492) );
  NAND U7694 ( .A(n7490), .B(n7489), .Z(n7491) );
  AND U7695 ( .A(n7492), .B(n7491), .Z(n7627) );
  NANDN U7696 ( .A(n7494), .B(n7493), .Z(n7498) );
  NANDN U7697 ( .A(n7496), .B(n7495), .Z(n7497) );
  AND U7698 ( .A(n7498), .B(n7497), .Z(n7593) );
  NAND U7699 ( .A(b[0]), .B(a[105]), .Z(n7499) );
  XNOR U7700 ( .A(b[1]), .B(n7499), .Z(n7501) );
  NANDN U7701 ( .A(b[0]), .B(a[104]), .Z(n7500) );
  NAND U7702 ( .A(n7501), .B(n7500), .Z(n7573) );
  NANDN U7703 ( .A(n9891), .B(n7502), .Z(n7504) );
  XOR U7704 ( .A(b[13]), .B(a[93]), .Z(n7576) );
  NANDN U7705 ( .A(n9935), .B(n7576), .Z(n7503) );
  AND U7706 ( .A(n7504), .B(n7503), .Z(n7571) );
  AND U7707 ( .A(b[15]), .B(a[89]), .Z(n7570) );
  XNOR U7708 ( .A(n7571), .B(n7570), .Z(n7572) );
  XNOR U7709 ( .A(n7573), .B(n7572), .Z(n7591) );
  NANDN U7710 ( .A(n9437), .B(n7505), .Z(n7507) );
  XOR U7711 ( .A(b[5]), .B(a[101]), .Z(n7582) );
  NANDN U7712 ( .A(n9503), .B(n7582), .Z(n7506) );
  AND U7713 ( .A(n7507), .B(n7506), .Z(n7615) );
  NANDN U7714 ( .A(n9588), .B(n7508), .Z(n7510) );
  XOR U7715 ( .A(b[7]), .B(a[99]), .Z(n7585) );
  NANDN U7716 ( .A(n9639), .B(n7585), .Z(n7509) );
  AND U7717 ( .A(n7510), .B(n7509), .Z(n7613) );
  NANDN U7718 ( .A(n9374), .B(n7511), .Z(n7513) );
  XOR U7719 ( .A(b[3]), .B(a[103]), .Z(n7588) );
  NANDN U7720 ( .A(n9375), .B(n7588), .Z(n7512) );
  NAND U7721 ( .A(n7513), .B(n7512), .Z(n7612) );
  XNOR U7722 ( .A(n7613), .B(n7612), .Z(n7614) );
  XOR U7723 ( .A(n7615), .B(n7614), .Z(n7592) );
  XOR U7724 ( .A(n7591), .B(n7592), .Z(n7594) );
  XOR U7725 ( .A(n7593), .B(n7594), .Z(n7565) );
  NANDN U7726 ( .A(n7515), .B(n7514), .Z(n7519) );
  OR U7727 ( .A(n7517), .B(n7516), .Z(n7518) );
  AND U7728 ( .A(n7519), .B(n7518), .Z(n7564) );
  XNOR U7729 ( .A(n7565), .B(n7564), .Z(n7567) );
  NAND U7730 ( .A(n7520), .B(n9883), .Z(n7522) );
  XOR U7731 ( .A(b[11]), .B(a[95]), .Z(n7597) );
  NANDN U7732 ( .A(n9856), .B(n7597), .Z(n7521) );
  AND U7733 ( .A(n7522), .B(n7521), .Z(n7608) );
  NANDN U7734 ( .A(n10005), .B(n7523), .Z(n7525) );
  XOR U7735 ( .A(b[15]), .B(a[91]), .Z(n7600) );
  NANDN U7736 ( .A(n10006), .B(n7600), .Z(n7524) );
  AND U7737 ( .A(n7525), .B(n7524), .Z(n7607) );
  NANDN U7738 ( .A(n9685), .B(n7526), .Z(n7528) );
  XOR U7739 ( .A(b[9]), .B(a[97]), .Z(n7603) );
  NANDN U7740 ( .A(n9758), .B(n7603), .Z(n7527) );
  NAND U7741 ( .A(n7528), .B(n7527), .Z(n7606) );
  XOR U7742 ( .A(n7607), .B(n7606), .Z(n7609) );
  XOR U7743 ( .A(n7608), .B(n7609), .Z(n7619) );
  NANDN U7744 ( .A(n7530), .B(n7529), .Z(n7534) );
  OR U7745 ( .A(n7532), .B(n7531), .Z(n7533) );
  AND U7746 ( .A(n7534), .B(n7533), .Z(n7618) );
  XNOR U7747 ( .A(n7619), .B(n7618), .Z(n7620) );
  NANDN U7748 ( .A(n7536), .B(n7535), .Z(n7540) );
  NANDN U7749 ( .A(n7538), .B(n7537), .Z(n7539) );
  NAND U7750 ( .A(n7540), .B(n7539), .Z(n7621) );
  XNOR U7751 ( .A(n7620), .B(n7621), .Z(n7566) );
  XOR U7752 ( .A(n7567), .B(n7566), .Z(n7625) );
  NANDN U7753 ( .A(n7542), .B(n7541), .Z(n7546) );
  NANDN U7754 ( .A(n7544), .B(n7543), .Z(n7545) );
  AND U7755 ( .A(n7546), .B(n7545), .Z(n7624) );
  XNOR U7756 ( .A(n7625), .B(n7624), .Z(n7626) );
  XOR U7757 ( .A(n7627), .B(n7626), .Z(n7559) );
  NANDN U7758 ( .A(n7548), .B(n7547), .Z(n7552) );
  NAND U7759 ( .A(n7550), .B(n7549), .Z(n7551) );
  AND U7760 ( .A(n7552), .B(n7551), .Z(n7558) );
  XNOR U7761 ( .A(n7559), .B(n7558), .Z(n7560) );
  XNOR U7762 ( .A(n7561), .B(n7560), .Z(n7630) );
  XNOR U7763 ( .A(sreg[217]), .B(n7630), .Z(n7632) );
  NANDN U7764 ( .A(sreg[216]), .B(n7553), .Z(n7557) );
  NAND U7765 ( .A(n7555), .B(n7554), .Z(n7556) );
  NAND U7766 ( .A(n7557), .B(n7556), .Z(n7631) );
  XNOR U7767 ( .A(n7632), .B(n7631), .Z(c[217]) );
  NANDN U7768 ( .A(n7559), .B(n7558), .Z(n7563) );
  NANDN U7769 ( .A(n7561), .B(n7560), .Z(n7562) );
  AND U7770 ( .A(n7563), .B(n7562), .Z(n7638) );
  NANDN U7771 ( .A(n7565), .B(n7564), .Z(n7569) );
  NAND U7772 ( .A(n7567), .B(n7566), .Z(n7568) );
  AND U7773 ( .A(n7569), .B(n7568), .Z(n7704) );
  NANDN U7774 ( .A(n7571), .B(n7570), .Z(n7575) );
  NANDN U7775 ( .A(n7573), .B(n7572), .Z(n7574) );
  AND U7776 ( .A(n7575), .B(n7574), .Z(n7670) );
  NANDN U7777 ( .A(n9891), .B(n7576), .Z(n7578) );
  XOR U7778 ( .A(b[13]), .B(a[94]), .Z(n7656) );
  NANDN U7779 ( .A(n9935), .B(n7656), .Z(n7577) );
  AND U7780 ( .A(n7578), .B(n7577), .Z(n7648) );
  AND U7781 ( .A(b[15]), .B(a[90]), .Z(n7647) );
  XNOR U7782 ( .A(n7648), .B(n7647), .Z(n7649) );
  NAND U7783 ( .A(b[0]), .B(a[106]), .Z(n7579) );
  XNOR U7784 ( .A(b[1]), .B(n7579), .Z(n7581) );
  NANDN U7785 ( .A(b[0]), .B(a[105]), .Z(n7580) );
  NAND U7786 ( .A(n7581), .B(n7580), .Z(n7650) );
  XNOR U7787 ( .A(n7649), .B(n7650), .Z(n7668) );
  NANDN U7788 ( .A(n9437), .B(n7582), .Z(n7584) );
  XOR U7789 ( .A(b[5]), .B(a[102]), .Z(n7659) );
  NANDN U7790 ( .A(n9503), .B(n7659), .Z(n7583) );
  AND U7791 ( .A(n7584), .B(n7583), .Z(n7692) );
  NANDN U7792 ( .A(n9588), .B(n7585), .Z(n7587) );
  XOR U7793 ( .A(b[7]), .B(a[100]), .Z(n7662) );
  NANDN U7794 ( .A(n9639), .B(n7662), .Z(n7586) );
  AND U7795 ( .A(n7587), .B(n7586), .Z(n7690) );
  NANDN U7796 ( .A(n9374), .B(n7588), .Z(n7590) );
  XOR U7797 ( .A(b[3]), .B(a[104]), .Z(n7665) );
  NANDN U7798 ( .A(n9375), .B(n7665), .Z(n7589) );
  NAND U7799 ( .A(n7590), .B(n7589), .Z(n7689) );
  XNOR U7800 ( .A(n7690), .B(n7689), .Z(n7691) );
  XOR U7801 ( .A(n7692), .B(n7691), .Z(n7669) );
  XOR U7802 ( .A(n7668), .B(n7669), .Z(n7671) );
  XOR U7803 ( .A(n7670), .B(n7671), .Z(n7642) );
  NANDN U7804 ( .A(n7592), .B(n7591), .Z(n7596) );
  OR U7805 ( .A(n7594), .B(n7593), .Z(n7595) );
  AND U7806 ( .A(n7596), .B(n7595), .Z(n7641) );
  XNOR U7807 ( .A(n7642), .B(n7641), .Z(n7644) );
  NAND U7808 ( .A(n7597), .B(n9883), .Z(n7599) );
  XOR U7809 ( .A(b[11]), .B(a[96]), .Z(n7674) );
  NANDN U7810 ( .A(n9856), .B(n7674), .Z(n7598) );
  AND U7811 ( .A(n7599), .B(n7598), .Z(n7685) );
  NANDN U7812 ( .A(n10005), .B(n7600), .Z(n7602) );
  XOR U7813 ( .A(b[15]), .B(a[92]), .Z(n7677) );
  NANDN U7814 ( .A(n10006), .B(n7677), .Z(n7601) );
  AND U7815 ( .A(n7602), .B(n7601), .Z(n7684) );
  NANDN U7816 ( .A(n9685), .B(n7603), .Z(n7605) );
  XOR U7817 ( .A(b[9]), .B(a[98]), .Z(n7680) );
  NANDN U7818 ( .A(n9758), .B(n7680), .Z(n7604) );
  NAND U7819 ( .A(n7605), .B(n7604), .Z(n7683) );
  XOR U7820 ( .A(n7684), .B(n7683), .Z(n7686) );
  XOR U7821 ( .A(n7685), .B(n7686), .Z(n7696) );
  NANDN U7822 ( .A(n7607), .B(n7606), .Z(n7611) );
  OR U7823 ( .A(n7609), .B(n7608), .Z(n7610) );
  AND U7824 ( .A(n7611), .B(n7610), .Z(n7695) );
  XNOR U7825 ( .A(n7696), .B(n7695), .Z(n7697) );
  NANDN U7826 ( .A(n7613), .B(n7612), .Z(n7617) );
  NANDN U7827 ( .A(n7615), .B(n7614), .Z(n7616) );
  NAND U7828 ( .A(n7617), .B(n7616), .Z(n7698) );
  XNOR U7829 ( .A(n7697), .B(n7698), .Z(n7643) );
  XOR U7830 ( .A(n7644), .B(n7643), .Z(n7702) );
  NANDN U7831 ( .A(n7619), .B(n7618), .Z(n7623) );
  NANDN U7832 ( .A(n7621), .B(n7620), .Z(n7622) );
  AND U7833 ( .A(n7623), .B(n7622), .Z(n7701) );
  XNOR U7834 ( .A(n7702), .B(n7701), .Z(n7703) );
  XOR U7835 ( .A(n7704), .B(n7703), .Z(n7636) );
  NANDN U7836 ( .A(n7625), .B(n7624), .Z(n7629) );
  NAND U7837 ( .A(n7627), .B(n7626), .Z(n7628) );
  AND U7838 ( .A(n7629), .B(n7628), .Z(n7635) );
  XNOR U7839 ( .A(n7636), .B(n7635), .Z(n7637) );
  XNOR U7840 ( .A(n7638), .B(n7637), .Z(n7707) );
  XNOR U7841 ( .A(sreg[218]), .B(n7707), .Z(n7709) );
  NANDN U7842 ( .A(sreg[217]), .B(n7630), .Z(n7634) );
  NAND U7843 ( .A(n7632), .B(n7631), .Z(n7633) );
  NAND U7844 ( .A(n7634), .B(n7633), .Z(n7708) );
  XNOR U7845 ( .A(n7709), .B(n7708), .Z(c[218]) );
  NANDN U7846 ( .A(n7636), .B(n7635), .Z(n7640) );
  NANDN U7847 ( .A(n7638), .B(n7637), .Z(n7639) );
  AND U7848 ( .A(n7640), .B(n7639), .Z(n7715) );
  NANDN U7849 ( .A(n7642), .B(n7641), .Z(n7646) );
  NAND U7850 ( .A(n7644), .B(n7643), .Z(n7645) );
  AND U7851 ( .A(n7646), .B(n7645), .Z(n7781) );
  NANDN U7852 ( .A(n7648), .B(n7647), .Z(n7652) );
  NANDN U7853 ( .A(n7650), .B(n7649), .Z(n7651) );
  AND U7854 ( .A(n7652), .B(n7651), .Z(n7747) );
  NAND U7855 ( .A(b[0]), .B(a[107]), .Z(n7653) );
  XNOR U7856 ( .A(b[1]), .B(n7653), .Z(n7655) );
  NANDN U7857 ( .A(b[0]), .B(a[106]), .Z(n7654) );
  NAND U7858 ( .A(n7655), .B(n7654), .Z(n7727) );
  NANDN U7859 ( .A(n9891), .B(n7656), .Z(n7658) );
  XOR U7860 ( .A(b[13]), .B(a[95]), .Z(n7733) );
  NANDN U7861 ( .A(n9935), .B(n7733), .Z(n7657) );
  AND U7862 ( .A(n7658), .B(n7657), .Z(n7725) );
  AND U7863 ( .A(b[15]), .B(a[91]), .Z(n7724) );
  XNOR U7864 ( .A(n7725), .B(n7724), .Z(n7726) );
  XNOR U7865 ( .A(n7727), .B(n7726), .Z(n7745) );
  NANDN U7866 ( .A(n9437), .B(n7659), .Z(n7661) );
  XOR U7867 ( .A(b[5]), .B(a[103]), .Z(n7736) );
  NANDN U7868 ( .A(n9503), .B(n7736), .Z(n7660) );
  AND U7869 ( .A(n7661), .B(n7660), .Z(n7769) );
  NANDN U7870 ( .A(n9588), .B(n7662), .Z(n7664) );
  XOR U7871 ( .A(b[7]), .B(a[101]), .Z(n7739) );
  NANDN U7872 ( .A(n9639), .B(n7739), .Z(n7663) );
  AND U7873 ( .A(n7664), .B(n7663), .Z(n7767) );
  NANDN U7874 ( .A(n9374), .B(n7665), .Z(n7667) );
  XOR U7875 ( .A(b[3]), .B(a[105]), .Z(n7742) );
  NANDN U7876 ( .A(n9375), .B(n7742), .Z(n7666) );
  NAND U7877 ( .A(n7667), .B(n7666), .Z(n7766) );
  XNOR U7878 ( .A(n7767), .B(n7766), .Z(n7768) );
  XOR U7879 ( .A(n7769), .B(n7768), .Z(n7746) );
  XOR U7880 ( .A(n7745), .B(n7746), .Z(n7748) );
  XOR U7881 ( .A(n7747), .B(n7748), .Z(n7719) );
  NANDN U7882 ( .A(n7669), .B(n7668), .Z(n7673) );
  OR U7883 ( .A(n7671), .B(n7670), .Z(n7672) );
  AND U7884 ( .A(n7673), .B(n7672), .Z(n7718) );
  XNOR U7885 ( .A(n7719), .B(n7718), .Z(n7721) );
  NAND U7886 ( .A(n7674), .B(n9883), .Z(n7676) );
  XOR U7887 ( .A(b[11]), .B(a[97]), .Z(n7751) );
  NANDN U7888 ( .A(n9856), .B(n7751), .Z(n7675) );
  AND U7889 ( .A(n7676), .B(n7675), .Z(n7762) );
  NANDN U7890 ( .A(n10005), .B(n7677), .Z(n7679) );
  XOR U7891 ( .A(b[15]), .B(a[93]), .Z(n7754) );
  NANDN U7892 ( .A(n10006), .B(n7754), .Z(n7678) );
  AND U7893 ( .A(n7679), .B(n7678), .Z(n7761) );
  NANDN U7894 ( .A(n9685), .B(n7680), .Z(n7682) );
  XOR U7895 ( .A(b[9]), .B(a[99]), .Z(n7757) );
  NANDN U7896 ( .A(n9758), .B(n7757), .Z(n7681) );
  NAND U7897 ( .A(n7682), .B(n7681), .Z(n7760) );
  XOR U7898 ( .A(n7761), .B(n7760), .Z(n7763) );
  XOR U7899 ( .A(n7762), .B(n7763), .Z(n7773) );
  NANDN U7900 ( .A(n7684), .B(n7683), .Z(n7688) );
  OR U7901 ( .A(n7686), .B(n7685), .Z(n7687) );
  AND U7902 ( .A(n7688), .B(n7687), .Z(n7772) );
  XNOR U7903 ( .A(n7773), .B(n7772), .Z(n7774) );
  NANDN U7904 ( .A(n7690), .B(n7689), .Z(n7694) );
  NANDN U7905 ( .A(n7692), .B(n7691), .Z(n7693) );
  NAND U7906 ( .A(n7694), .B(n7693), .Z(n7775) );
  XNOR U7907 ( .A(n7774), .B(n7775), .Z(n7720) );
  XOR U7908 ( .A(n7721), .B(n7720), .Z(n7779) );
  NANDN U7909 ( .A(n7696), .B(n7695), .Z(n7700) );
  NANDN U7910 ( .A(n7698), .B(n7697), .Z(n7699) );
  AND U7911 ( .A(n7700), .B(n7699), .Z(n7778) );
  XNOR U7912 ( .A(n7779), .B(n7778), .Z(n7780) );
  XOR U7913 ( .A(n7781), .B(n7780), .Z(n7713) );
  NANDN U7914 ( .A(n7702), .B(n7701), .Z(n7706) );
  NAND U7915 ( .A(n7704), .B(n7703), .Z(n7705) );
  AND U7916 ( .A(n7706), .B(n7705), .Z(n7712) );
  XNOR U7917 ( .A(n7713), .B(n7712), .Z(n7714) );
  XNOR U7918 ( .A(n7715), .B(n7714), .Z(n7784) );
  XNOR U7919 ( .A(sreg[219]), .B(n7784), .Z(n7786) );
  NANDN U7920 ( .A(sreg[218]), .B(n7707), .Z(n7711) );
  NAND U7921 ( .A(n7709), .B(n7708), .Z(n7710) );
  NAND U7922 ( .A(n7711), .B(n7710), .Z(n7785) );
  XNOR U7923 ( .A(n7786), .B(n7785), .Z(c[219]) );
  NANDN U7924 ( .A(n7713), .B(n7712), .Z(n7717) );
  NANDN U7925 ( .A(n7715), .B(n7714), .Z(n7716) );
  AND U7926 ( .A(n7717), .B(n7716), .Z(n7792) );
  NANDN U7927 ( .A(n7719), .B(n7718), .Z(n7723) );
  NAND U7928 ( .A(n7721), .B(n7720), .Z(n7722) );
  AND U7929 ( .A(n7723), .B(n7722), .Z(n7858) );
  NANDN U7930 ( .A(n7725), .B(n7724), .Z(n7729) );
  NANDN U7931 ( .A(n7727), .B(n7726), .Z(n7728) );
  AND U7932 ( .A(n7729), .B(n7728), .Z(n7824) );
  NAND U7933 ( .A(b[0]), .B(a[108]), .Z(n7730) );
  XNOR U7934 ( .A(b[1]), .B(n7730), .Z(n7732) );
  NANDN U7935 ( .A(b[0]), .B(a[107]), .Z(n7731) );
  NAND U7936 ( .A(n7732), .B(n7731), .Z(n7804) );
  NANDN U7937 ( .A(n9891), .B(n7733), .Z(n7735) );
  XOR U7938 ( .A(b[13]), .B(a[96]), .Z(n7807) );
  NANDN U7939 ( .A(n9935), .B(n7807), .Z(n7734) );
  AND U7940 ( .A(n7735), .B(n7734), .Z(n7802) );
  AND U7941 ( .A(b[15]), .B(a[92]), .Z(n7801) );
  XNOR U7942 ( .A(n7802), .B(n7801), .Z(n7803) );
  XNOR U7943 ( .A(n7804), .B(n7803), .Z(n7822) );
  NANDN U7944 ( .A(n9437), .B(n7736), .Z(n7738) );
  XOR U7945 ( .A(b[5]), .B(a[104]), .Z(n7813) );
  NANDN U7946 ( .A(n9503), .B(n7813), .Z(n7737) );
  AND U7947 ( .A(n7738), .B(n7737), .Z(n7846) );
  NANDN U7948 ( .A(n9588), .B(n7739), .Z(n7741) );
  XOR U7949 ( .A(b[7]), .B(a[102]), .Z(n7816) );
  NANDN U7950 ( .A(n9639), .B(n7816), .Z(n7740) );
  AND U7951 ( .A(n7741), .B(n7740), .Z(n7844) );
  NANDN U7952 ( .A(n9374), .B(n7742), .Z(n7744) );
  XOR U7953 ( .A(b[3]), .B(a[106]), .Z(n7819) );
  NANDN U7954 ( .A(n9375), .B(n7819), .Z(n7743) );
  NAND U7955 ( .A(n7744), .B(n7743), .Z(n7843) );
  XNOR U7956 ( .A(n7844), .B(n7843), .Z(n7845) );
  XOR U7957 ( .A(n7846), .B(n7845), .Z(n7823) );
  XOR U7958 ( .A(n7822), .B(n7823), .Z(n7825) );
  XOR U7959 ( .A(n7824), .B(n7825), .Z(n7796) );
  NANDN U7960 ( .A(n7746), .B(n7745), .Z(n7750) );
  OR U7961 ( .A(n7748), .B(n7747), .Z(n7749) );
  AND U7962 ( .A(n7750), .B(n7749), .Z(n7795) );
  XNOR U7963 ( .A(n7796), .B(n7795), .Z(n7798) );
  NAND U7964 ( .A(n7751), .B(n9883), .Z(n7753) );
  XOR U7965 ( .A(b[11]), .B(a[98]), .Z(n7828) );
  NANDN U7966 ( .A(n9856), .B(n7828), .Z(n7752) );
  AND U7967 ( .A(n7753), .B(n7752), .Z(n7839) );
  NANDN U7968 ( .A(n10005), .B(n7754), .Z(n7756) );
  XOR U7969 ( .A(b[15]), .B(a[94]), .Z(n7831) );
  NANDN U7970 ( .A(n10006), .B(n7831), .Z(n7755) );
  AND U7971 ( .A(n7756), .B(n7755), .Z(n7838) );
  NANDN U7972 ( .A(n9685), .B(n7757), .Z(n7759) );
  XOR U7973 ( .A(b[9]), .B(a[100]), .Z(n7834) );
  NANDN U7974 ( .A(n9758), .B(n7834), .Z(n7758) );
  NAND U7975 ( .A(n7759), .B(n7758), .Z(n7837) );
  XOR U7976 ( .A(n7838), .B(n7837), .Z(n7840) );
  XOR U7977 ( .A(n7839), .B(n7840), .Z(n7850) );
  NANDN U7978 ( .A(n7761), .B(n7760), .Z(n7765) );
  OR U7979 ( .A(n7763), .B(n7762), .Z(n7764) );
  AND U7980 ( .A(n7765), .B(n7764), .Z(n7849) );
  XNOR U7981 ( .A(n7850), .B(n7849), .Z(n7851) );
  NANDN U7982 ( .A(n7767), .B(n7766), .Z(n7771) );
  NANDN U7983 ( .A(n7769), .B(n7768), .Z(n7770) );
  NAND U7984 ( .A(n7771), .B(n7770), .Z(n7852) );
  XNOR U7985 ( .A(n7851), .B(n7852), .Z(n7797) );
  XOR U7986 ( .A(n7798), .B(n7797), .Z(n7856) );
  NANDN U7987 ( .A(n7773), .B(n7772), .Z(n7777) );
  NANDN U7988 ( .A(n7775), .B(n7774), .Z(n7776) );
  AND U7989 ( .A(n7777), .B(n7776), .Z(n7855) );
  XNOR U7990 ( .A(n7856), .B(n7855), .Z(n7857) );
  XOR U7991 ( .A(n7858), .B(n7857), .Z(n7790) );
  NANDN U7992 ( .A(n7779), .B(n7778), .Z(n7783) );
  NAND U7993 ( .A(n7781), .B(n7780), .Z(n7782) );
  AND U7994 ( .A(n7783), .B(n7782), .Z(n7789) );
  XNOR U7995 ( .A(n7790), .B(n7789), .Z(n7791) );
  XNOR U7996 ( .A(n7792), .B(n7791), .Z(n7861) );
  XNOR U7997 ( .A(sreg[220]), .B(n7861), .Z(n7863) );
  NANDN U7998 ( .A(sreg[219]), .B(n7784), .Z(n7788) );
  NAND U7999 ( .A(n7786), .B(n7785), .Z(n7787) );
  NAND U8000 ( .A(n7788), .B(n7787), .Z(n7862) );
  XNOR U8001 ( .A(n7863), .B(n7862), .Z(c[220]) );
  NANDN U8002 ( .A(n7790), .B(n7789), .Z(n7794) );
  NANDN U8003 ( .A(n7792), .B(n7791), .Z(n7793) );
  AND U8004 ( .A(n7794), .B(n7793), .Z(n7869) );
  NANDN U8005 ( .A(n7796), .B(n7795), .Z(n7800) );
  NAND U8006 ( .A(n7798), .B(n7797), .Z(n7799) );
  AND U8007 ( .A(n7800), .B(n7799), .Z(n7935) );
  NANDN U8008 ( .A(n7802), .B(n7801), .Z(n7806) );
  NANDN U8009 ( .A(n7804), .B(n7803), .Z(n7805) );
  AND U8010 ( .A(n7806), .B(n7805), .Z(n7901) );
  NANDN U8011 ( .A(n9891), .B(n7807), .Z(n7809) );
  XOR U8012 ( .A(b[13]), .B(a[97]), .Z(n7887) );
  NANDN U8013 ( .A(n9935), .B(n7887), .Z(n7808) );
  AND U8014 ( .A(n7809), .B(n7808), .Z(n7879) );
  AND U8015 ( .A(b[15]), .B(a[93]), .Z(n7878) );
  XNOR U8016 ( .A(n7879), .B(n7878), .Z(n7880) );
  NAND U8017 ( .A(b[0]), .B(a[109]), .Z(n7810) );
  XNOR U8018 ( .A(b[1]), .B(n7810), .Z(n7812) );
  NANDN U8019 ( .A(b[0]), .B(a[108]), .Z(n7811) );
  NAND U8020 ( .A(n7812), .B(n7811), .Z(n7881) );
  XNOR U8021 ( .A(n7880), .B(n7881), .Z(n7899) );
  NANDN U8022 ( .A(n9437), .B(n7813), .Z(n7815) );
  XOR U8023 ( .A(b[5]), .B(a[105]), .Z(n7890) );
  NANDN U8024 ( .A(n9503), .B(n7890), .Z(n7814) );
  AND U8025 ( .A(n7815), .B(n7814), .Z(n7923) );
  NANDN U8026 ( .A(n9588), .B(n7816), .Z(n7818) );
  XOR U8027 ( .A(b[7]), .B(a[103]), .Z(n7893) );
  NANDN U8028 ( .A(n9639), .B(n7893), .Z(n7817) );
  AND U8029 ( .A(n7818), .B(n7817), .Z(n7921) );
  NANDN U8030 ( .A(n9374), .B(n7819), .Z(n7821) );
  XOR U8031 ( .A(b[3]), .B(a[107]), .Z(n7896) );
  NANDN U8032 ( .A(n9375), .B(n7896), .Z(n7820) );
  NAND U8033 ( .A(n7821), .B(n7820), .Z(n7920) );
  XNOR U8034 ( .A(n7921), .B(n7920), .Z(n7922) );
  XOR U8035 ( .A(n7923), .B(n7922), .Z(n7900) );
  XOR U8036 ( .A(n7899), .B(n7900), .Z(n7902) );
  XOR U8037 ( .A(n7901), .B(n7902), .Z(n7873) );
  NANDN U8038 ( .A(n7823), .B(n7822), .Z(n7827) );
  OR U8039 ( .A(n7825), .B(n7824), .Z(n7826) );
  AND U8040 ( .A(n7827), .B(n7826), .Z(n7872) );
  XNOR U8041 ( .A(n7873), .B(n7872), .Z(n7875) );
  NAND U8042 ( .A(n7828), .B(n9883), .Z(n7830) );
  XOR U8043 ( .A(b[11]), .B(a[99]), .Z(n7905) );
  NANDN U8044 ( .A(n9856), .B(n7905), .Z(n7829) );
  AND U8045 ( .A(n7830), .B(n7829), .Z(n7916) );
  NANDN U8046 ( .A(n10005), .B(n7831), .Z(n7833) );
  XOR U8047 ( .A(b[15]), .B(a[95]), .Z(n7908) );
  NANDN U8048 ( .A(n10006), .B(n7908), .Z(n7832) );
  AND U8049 ( .A(n7833), .B(n7832), .Z(n7915) );
  NANDN U8050 ( .A(n9685), .B(n7834), .Z(n7836) );
  XOR U8051 ( .A(b[9]), .B(a[101]), .Z(n7911) );
  NANDN U8052 ( .A(n9758), .B(n7911), .Z(n7835) );
  NAND U8053 ( .A(n7836), .B(n7835), .Z(n7914) );
  XOR U8054 ( .A(n7915), .B(n7914), .Z(n7917) );
  XOR U8055 ( .A(n7916), .B(n7917), .Z(n7927) );
  NANDN U8056 ( .A(n7838), .B(n7837), .Z(n7842) );
  OR U8057 ( .A(n7840), .B(n7839), .Z(n7841) );
  AND U8058 ( .A(n7842), .B(n7841), .Z(n7926) );
  XNOR U8059 ( .A(n7927), .B(n7926), .Z(n7928) );
  NANDN U8060 ( .A(n7844), .B(n7843), .Z(n7848) );
  NANDN U8061 ( .A(n7846), .B(n7845), .Z(n7847) );
  NAND U8062 ( .A(n7848), .B(n7847), .Z(n7929) );
  XNOR U8063 ( .A(n7928), .B(n7929), .Z(n7874) );
  XOR U8064 ( .A(n7875), .B(n7874), .Z(n7933) );
  NANDN U8065 ( .A(n7850), .B(n7849), .Z(n7854) );
  NANDN U8066 ( .A(n7852), .B(n7851), .Z(n7853) );
  AND U8067 ( .A(n7854), .B(n7853), .Z(n7932) );
  XNOR U8068 ( .A(n7933), .B(n7932), .Z(n7934) );
  XOR U8069 ( .A(n7935), .B(n7934), .Z(n7867) );
  NANDN U8070 ( .A(n7856), .B(n7855), .Z(n7860) );
  NAND U8071 ( .A(n7858), .B(n7857), .Z(n7859) );
  AND U8072 ( .A(n7860), .B(n7859), .Z(n7866) );
  XNOR U8073 ( .A(n7867), .B(n7866), .Z(n7868) );
  XNOR U8074 ( .A(n7869), .B(n7868), .Z(n7938) );
  XNOR U8075 ( .A(sreg[221]), .B(n7938), .Z(n7940) );
  NANDN U8076 ( .A(sreg[220]), .B(n7861), .Z(n7865) );
  NAND U8077 ( .A(n7863), .B(n7862), .Z(n7864) );
  NAND U8078 ( .A(n7865), .B(n7864), .Z(n7939) );
  XNOR U8079 ( .A(n7940), .B(n7939), .Z(c[221]) );
  NANDN U8080 ( .A(n7867), .B(n7866), .Z(n7871) );
  NANDN U8081 ( .A(n7869), .B(n7868), .Z(n7870) );
  AND U8082 ( .A(n7871), .B(n7870), .Z(n7946) );
  NANDN U8083 ( .A(n7873), .B(n7872), .Z(n7877) );
  NAND U8084 ( .A(n7875), .B(n7874), .Z(n7876) );
  AND U8085 ( .A(n7877), .B(n7876), .Z(n8012) );
  NANDN U8086 ( .A(n7879), .B(n7878), .Z(n7883) );
  NANDN U8087 ( .A(n7881), .B(n7880), .Z(n7882) );
  AND U8088 ( .A(n7883), .B(n7882), .Z(n7978) );
  NAND U8089 ( .A(b[0]), .B(a[110]), .Z(n7884) );
  XNOR U8090 ( .A(b[1]), .B(n7884), .Z(n7886) );
  NANDN U8091 ( .A(b[0]), .B(a[109]), .Z(n7885) );
  NAND U8092 ( .A(n7886), .B(n7885), .Z(n7958) );
  NANDN U8093 ( .A(n9891), .B(n7887), .Z(n7889) );
  XOR U8094 ( .A(b[13]), .B(a[98]), .Z(n7964) );
  NANDN U8095 ( .A(n9935), .B(n7964), .Z(n7888) );
  AND U8096 ( .A(n7889), .B(n7888), .Z(n7956) );
  AND U8097 ( .A(b[15]), .B(a[94]), .Z(n7955) );
  XNOR U8098 ( .A(n7956), .B(n7955), .Z(n7957) );
  XNOR U8099 ( .A(n7958), .B(n7957), .Z(n7976) );
  NANDN U8100 ( .A(n9437), .B(n7890), .Z(n7892) );
  XOR U8101 ( .A(b[5]), .B(a[106]), .Z(n7967) );
  NANDN U8102 ( .A(n9503), .B(n7967), .Z(n7891) );
  AND U8103 ( .A(n7892), .B(n7891), .Z(n8000) );
  NANDN U8104 ( .A(n9588), .B(n7893), .Z(n7895) );
  XOR U8105 ( .A(b[7]), .B(a[104]), .Z(n7970) );
  NANDN U8106 ( .A(n9639), .B(n7970), .Z(n7894) );
  AND U8107 ( .A(n7895), .B(n7894), .Z(n7998) );
  NANDN U8108 ( .A(n9374), .B(n7896), .Z(n7898) );
  XOR U8109 ( .A(b[3]), .B(a[108]), .Z(n7973) );
  NANDN U8110 ( .A(n9375), .B(n7973), .Z(n7897) );
  NAND U8111 ( .A(n7898), .B(n7897), .Z(n7997) );
  XNOR U8112 ( .A(n7998), .B(n7997), .Z(n7999) );
  XOR U8113 ( .A(n8000), .B(n7999), .Z(n7977) );
  XOR U8114 ( .A(n7976), .B(n7977), .Z(n7979) );
  XOR U8115 ( .A(n7978), .B(n7979), .Z(n7950) );
  NANDN U8116 ( .A(n7900), .B(n7899), .Z(n7904) );
  OR U8117 ( .A(n7902), .B(n7901), .Z(n7903) );
  AND U8118 ( .A(n7904), .B(n7903), .Z(n7949) );
  XNOR U8119 ( .A(n7950), .B(n7949), .Z(n7952) );
  NAND U8120 ( .A(n7905), .B(n9883), .Z(n7907) );
  XOR U8121 ( .A(b[11]), .B(a[100]), .Z(n7982) );
  NANDN U8122 ( .A(n9856), .B(n7982), .Z(n7906) );
  AND U8123 ( .A(n7907), .B(n7906), .Z(n7993) );
  NANDN U8124 ( .A(n10005), .B(n7908), .Z(n7910) );
  XOR U8125 ( .A(b[15]), .B(a[96]), .Z(n7985) );
  NANDN U8126 ( .A(n10006), .B(n7985), .Z(n7909) );
  AND U8127 ( .A(n7910), .B(n7909), .Z(n7992) );
  NANDN U8128 ( .A(n9685), .B(n7911), .Z(n7913) );
  XOR U8129 ( .A(b[9]), .B(a[102]), .Z(n7988) );
  NANDN U8130 ( .A(n9758), .B(n7988), .Z(n7912) );
  NAND U8131 ( .A(n7913), .B(n7912), .Z(n7991) );
  XOR U8132 ( .A(n7992), .B(n7991), .Z(n7994) );
  XOR U8133 ( .A(n7993), .B(n7994), .Z(n8004) );
  NANDN U8134 ( .A(n7915), .B(n7914), .Z(n7919) );
  OR U8135 ( .A(n7917), .B(n7916), .Z(n7918) );
  AND U8136 ( .A(n7919), .B(n7918), .Z(n8003) );
  XNOR U8137 ( .A(n8004), .B(n8003), .Z(n8005) );
  NANDN U8138 ( .A(n7921), .B(n7920), .Z(n7925) );
  NANDN U8139 ( .A(n7923), .B(n7922), .Z(n7924) );
  NAND U8140 ( .A(n7925), .B(n7924), .Z(n8006) );
  XNOR U8141 ( .A(n8005), .B(n8006), .Z(n7951) );
  XOR U8142 ( .A(n7952), .B(n7951), .Z(n8010) );
  NANDN U8143 ( .A(n7927), .B(n7926), .Z(n7931) );
  NANDN U8144 ( .A(n7929), .B(n7928), .Z(n7930) );
  AND U8145 ( .A(n7931), .B(n7930), .Z(n8009) );
  XNOR U8146 ( .A(n8010), .B(n8009), .Z(n8011) );
  XOR U8147 ( .A(n8012), .B(n8011), .Z(n7944) );
  NANDN U8148 ( .A(n7933), .B(n7932), .Z(n7937) );
  NAND U8149 ( .A(n7935), .B(n7934), .Z(n7936) );
  AND U8150 ( .A(n7937), .B(n7936), .Z(n7943) );
  XNOR U8151 ( .A(n7944), .B(n7943), .Z(n7945) );
  XNOR U8152 ( .A(n7946), .B(n7945), .Z(n8015) );
  XNOR U8153 ( .A(sreg[222]), .B(n8015), .Z(n8017) );
  NANDN U8154 ( .A(sreg[221]), .B(n7938), .Z(n7942) );
  NAND U8155 ( .A(n7940), .B(n7939), .Z(n7941) );
  NAND U8156 ( .A(n7942), .B(n7941), .Z(n8016) );
  XNOR U8157 ( .A(n8017), .B(n8016), .Z(c[222]) );
  NANDN U8158 ( .A(n7944), .B(n7943), .Z(n7948) );
  NANDN U8159 ( .A(n7946), .B(n7945), .Z(n7947) );
  AND U8160 ( .A(n7948), .B(n7947), .Z(n8023) );
  NANDN U8161 ( .A(n7950), .B(n7949), .Z(n7954) );
  NAND U8162 ( .A(n7952), .B(n7951), .Z(n7953) );
  AND U8163 ( .A(n7954), .B(n7953), .Z(n8089) );
  NANDN U8164 ( .A(n7956), .B(n7955), .Z(n7960) );
  NANDN U8165 ( .A(n7958), .B(n7957), .Z(n7959) );
  AND U8166 ( .A(n7960), .B(n7959), .Z(n8055) );
  NAND U8167 ( .A(b[0]), .B(a[111]), .Z(n7961) );
  XNOR U8168 ( .A(b[1]), .B(n7961), .Z(n7963) );
  NANDN U8169 ( .A(b[0]), .B(a[110]), .Z(n7962) );
  NAND U8170 ( .A(n7963), .B(n7962), .Z(n8035) );
  NANDN U8171 ( .A(n9891), .B(n7964), .Z(n7966) );
  XOR U8172 ( .A(b[13]), .B(a[99]), .Z(n8041) );
  NANDN U8173 ( .A(n9935), .B(n8041), .Z(n7965) );
  AND U8174 ( .A(n7966), .B(n7965), .Z(n8033) );
  AND U8175 ( .A(b[15]), .B(a[95]), .Z(n8032) );
  XNOR U8176 ( .A(n8033), .B(n8032), .Z(n8034) );
  XNOR U8177 ( .A(n8035), .B(n8034), .Z(n8053) );
  NANDN U8178 ( .A(n9437), .B(n7967), .Z(n7969) );
  XOR U8179 ( .A(b[5]), .B(a[107]), .Z(n8044) );
  NANDN U8180 ( .A(n9503), .B(n8044), .Z(n7968) );
  AND U8181 ( .A(n7969), .B(n7968), .Z(n8077) );
  NANDN U8182 ( .A(n9588), .B(n7970), .Z(n7972) );
  XOR U8183 ( .A(b[7]), .B(a[105]), .Z(n8047) );
  NANDN U8184 ( .A(n9639), .B(n8047), .Z(n7971) );
  AND U8185 ( .A(n7972), .B(n7971), .Z(n8075) );
  NANDN U8186 ( .A(n9374), .B(n7973), .Z(n7975) );
  XOR U8187 ( .A(b[3]), .B(a[109]), .Z(n8050) );
  NANDN U8188 ( .A(n9375), .B(n8050), .Z(n7974) );
  NAND U8189 ( .A(n7975), .B(n7974), .Z(n8074) );
  XNOR U8190 ( .A(n8075), .B(n8074), .Z(n8076) );
  XOR U8191 ( .A(n8077), .B(n8076), .Z(n8054) );
  XOR U8192 ( .A(n8053), .B(n8054), .Z(n8056) );
  XOR U8193 ( .A(n8055), .B(n8056), .Z(n8027) );
  NANDN U8194 ( .A(n7977), .B(n7976), .Z(n7981) );
  OR U8195 ( .A(n7979), .B(n7978), .Z(n7980) );
  AND U8196 ( .A(n7981), .B(n7980), .Z(n8026) );
  XNOR U8197 ( .A(n8027), .B(n8026), .Z(n8029) );
  NAND U8198 ( .A(n7982), .B(n9883), .Z(n7984) );
  XOR U8199 ( .A(b[11]), .B(a[101]), .Z(n8059) );
  NANDN U8200 ( .A(n9856), .B(n8059), .Z(n7983) );
  AND U8201 ( .A(n7984), .B(n7983), .Z(n8070) );
  NANDN U8202 ( .A(n10005), .B(n7985), .Z(n7987) );
  XOR U8203 ( .A(b[15]), .B(a[97]), .Z(n8062) );
  NANDN U8204 ( .A(n10006), .B(n8062), .Z(n7986) );
  AND U8205 ( .A(n7987), .B(n7986), .Z(n8069) );
  NANDN U8206 ( .A(n9685), .B(n7988), .Z(n7990) );
  XOR U8207 ( .A(b[9]), .B(a[103]), .Z(n8065) );
  NANDN U8208 ( .A(n9758), .B(n8065), .Z(n7989) );
  NAND U8209 ( .A(n7990), .B(n7989), .Z(n8068) );
  XOR U8210 ( .A(n8069), .B(n8068), .Z(n8071) );
  XOR U8211 ( .A(n8070), .B(n8071), .Z(n8081) );
  NANDN U8212 ( .A(n7992), .B(n7991), .Z(n7996) );
  OR U8213 ( .A(n7994), .B(n7993), .Z(n7995) );
  AND U8214 ( .A(n7996), .B(n7995), .Z(n8080) );
  XNOR U8215 ( .A(n8081), .B(n8080), .Z(n8082) );
  NANDN U8216 ( .A(n7998), .B(n7997), .Z(n8002) );
  NANDN U8217 ( .A(n8000), .B(n7999), .Z(n8001) );
  NAND U8218 ( .A(n8002), .B(n8001), .Z(n8083) );
  XNOR U8219 ( .A(n8082), .B(n8083), .Z(n8028) );
  XOR U8220 ( .A(n8029), .B(n8028), .Z(n8087) );
  NANDN U8221 ( .A(n8004), .B(n8003), .Z(n8008) );
  NANDN U8222 ( .A(n8006), .B(n8005), .Z(n8007) );
  AND U8223 ( .A(n8008), .B(n8007), .Z(n8086) );
  XNOR U8224 ( .A(n8087), .B(n8086), .Z(n8088) );
  XOR U8225 ( .A(n8089), .B(n8088), .Z(n8021) );
  NANDN U8226 ( .A(n8010), .B(n8009), .Z(n8014) );
  NAND U8227 ( .A(n8012), .B(n8011), .Z(n8013) );
  AND U8228 ( .A(n8014), .B(n8013), .Z(n8020) );
  XNOR U8229 ( .A(n8021), .B(n8020), .Z(n8022) );
  XNOR U8230 ( .A(n8023), .B(n8022), .Z(n8092) );
  XNOR U8231 ( .A(sreg[223]), .B(n8092), .Z(n8094) );
  NANDN U8232 ( .A(sreg[222]), .B(n8015), .Z(n8019) );
  NAND U8233 ( .A(n8017), .B(n8016), .Z(n8018) );
  NAND U8234 ( .A(n8019), .B(n8018), .Z(n8093) );
  XNOR U8235 ( .A(n8094), .B(n8093), .Z(c[223]) );
  NANDN U8236 ( .A(n8021), .B(n8020), .Z(n8025) );
  NANDN U8237 ( .A(n8023), .B(n8022), .Z(n8024) );
  AND U8238 ( .A(n8025), .B(n8024), .Z(n8100) );
  NANDN U8239 ( .A(n8027), .B(n8026), .Z(n8031) );
  NAND U8240 ( .A(n8029), .B(n8028), .Z(n8030) );
  AND U8241 ( .A(n8031), .B(n8030), .Z(n8166) );
  NANDN U8242 ( .A(n8033), .B(n8032), .Z(n8037) );
  NANDN U8243 ( .A(n8035), .B(n8034), .Z(n8036) );
  AND U8244 ( .A(n8037), .B(n8036), .Z(n8132) );
  NAND U8245 ( .A(b[0]), .B(a[112]), .Z(n8038) );
  XNOR U8246 ( .A(b[1]), .B(n8038), .Z(n8040) );
  NANDN U8247 ( .A(b[0]), .B(a[111]), .Z(n8039) );
  NAND U8248 ( .A(n8040), .B(n8039), .Z(n8112) );
  NANDN U8249 ( .A(n9891), .B(n8041), .Z(n8043) );
  XOR U8250 ( .A(b[13]), .B(a[100]), .Z(n8118) );
  NANDN U8251 ( .A(n9935), .B(n8118), .Z(n8042) );
  AND U8252 ( .A(n8043), .B(n8042), .Z(n8110) );
  AND U8253 ( .A(b[15]), .B(a[96]), .Z(n8109) );
  XNOR U8254 ( .A(n8110), .B(n8109), .Z(n8111) );
  XNOR U8255 ( .A(n8112), .B(n8111), .Z(n8130) );
  NANDN U8256 ( .A(n9437), .B(n8044), .Z(n8046) );
  XOR U8257 ( .A(b[5]), .B(a[108]), .Z(n8121) );
  NANDN U8258 ( .A(n9503), .B(n8121), .Z(n8045) );
  AND U8259 ( .A(n8046), .B(n8045), .Z(n8154) );
  NANDN U8260 ( .A(n9588), .B(n8047), .Z(n8049) );
  XOR U8261 ( .A(b[7]), .B(a[106]), .Z(n8124) );
  NANDN U8262 ( .A(n9639), .B(n8124), .Z(n8048) );
  AND U8263 ( .A(n8049), .B(n8048), .Z(n8152) );
  NANDN U8264 ( .A(n9374), .B(n8050), .Z(n8052) );
  XOR U8265 ( .A(b[3]), .B(a[110]), .Z(n8127) );
  NANDN U8266 ( .A(n9375), .B(n8127), .Z(n8051) );
  NAND U8267 ( .A(n8052), .B(n8051), .Z(n8151) );
  XNOR U8268 ( .A(n8152), .B(n8151), .Z(n8153) );
  XOR U8269 ( .A(n8154), .B(n8153), .Z(n8131) );
  XOR U8270 ( .A(n8130), .B(n8131), .Z(n8133) );
  XOR U8271 ( .A(n8132), .B(n8133), .Z(n8104) );
  NANDN U8272 ( .A(n8054), .B(n8053), .Z(n8058) );
  OR U8273 ( .A(n8056), .B(n8055), .Z(n8057) );
  AND U8274 ( .A(n8058), .B(n8057), .Z(n8103) );
  XNOR U8275 ( .A(n8104), .B(n8103), .Z(n8106) );
  NAND U8276 ( .A(n8059), .B(n9883), .Z(n8061) );
  XOR U8277 ( .A(b[11]), .B(a[102]), .Z(n8136) );
  NANDN U8278 ( .A(n9856), .B(n8136), .Z(n8060) );
  AND U8279 ( .A(n8061), .B(n8060), .Z(n8147) );
  NANDN U8280 ( .A(n10005), .B(n8062), .Z(n8064) );
  XOR U8281 ( .A(b[15]), .B(a[98]), .Z(n8139) );
  NANDN U8282 ( .A(n10006), .B(n8139), .Z(n8063) );
  AND U8283 ( .A(n8064), .B(n8063), .Z(n8146) );
  NANDN U8284 ( .A(n9685), .B(n8065), .Z(n8067) );
  XOR U8285 ( .A(b[9]), .B(a[104]), .Z(n8142) );
  NANDN U8286 ( .A(n9758), .B(n8142), .Z(n8066) );
  NAND U8287 ( .A(n8067), .B(n8066), .Z(n8145) );
  XOR U8288 ( .A(n8146), .B(n8145), .Z(n8148) );
  XOR U8289 ( .A(n8147), .B(n8148), .Z(n8158) );
  NANDN U8290 ( .A(n8069), .B(n8068), .Z(n8073) );
  OR U8291 ( .A(n8071), .B(n8070), .Z(n8072) );
  AND U8292 ( .A(n8073), .B(n8072), .Z(n8157) );
  XNOR U8293 ( .A(n8158), .B(n8157), .Z(n8159) );
  NANDN U8294 ( .A(n8075), .B(n8074), .Z(n8079) );
  NANDN U8295 ( .A(n8077), .B(n8076), .Z(n8078) );
  NAND U8296 ( .A(n8079), .B(n8078), .Z(n8160) );
  XNOR U8297 ( .A(n8159), .B(n8160), .Z(n8105) );
  XOR U8298 ( .A(n8106), .B(n8105), .Z(n8164) );
  NANDN U8299 ( .A(n8081), .B(n8080), .Z(n8085) );
  NANDN U8300 ( .A(n8083), .B(n8082), .Z(n8084) );
  AND U8301 ( .A(n8085), .B(n8084), .Z(n8163) );
  XNOR U8302 ( .A(n8164), .B(n8163), .Z(n8165) );
  XOR U8303 ( .A(n8166), .B(n8165), .Z(n8098) );
  NANDN U8304 ( .A(n8087), .B(n8086), .Z(n8091) );
  NAND U8305 ( .A(n8089), .B(n8088), .Z(n8090) );
  AND U8306 ( .A(n8091), .B(n8090), .Z(n8097) );
  XNOR U8307 ( .A(n8098), .B(n8097), .Z(n8099) );
  XNOR U8308 ( .A(n8100), .B(n8099), .Z(n8169) );
  XNOR U8309 ( .A(sreg[224]), .B(n8169), .Z(n8171) );
  NANDN U8310 ( .A(sreg[223]), .B(n8092), .Z(n8096) );
  NAND U8311 ( .A(n8094), .B(n8093), .Z(n8095) );
  NAND U8312 ( .A(n8096), .B(n8095), .Z(n8170) );
  XNOR U8313 ( .A(n8171), .B(n8170), .Z(c[224]) );
  NANDN U8314 ( .A(n8098), .B(n8097), .Z(n8102) );
  NANDN U8315 ( .A(n8100), .B(n8099), .Z(n8101) );
  AND U8316 ( .A(n8102), .B(n8101), .Z(n8177) );
  NANDN U8317 ( .A(n8104), .B(n8103), .Z(n8108) );
  NAND U8318 ( .A(n8106), .B(n8105), .Z(n8107) );
  AND U8319 ( .A(n8108), .B(n8107), .Z(n8243) );
  NANDN U8320 ( .A(n8110), .B(n8109), .Z(n8114) );
  NANDN U8321 ( .A(n8112), .B(n8111), .Z(n8113) );
  AND U8322 ( .A(n8114), .B(n8113), .Z(n8230) );
  NAND U8323 ( .A(b[0]), .B(a[113]), .Z(n8115) );
  XNOR U8324 ( .A(b[1]), .B(n8115), .Z(n8117) );
  NANDN U8325 ( .A(b[0]), .B(a[112]), .Z(n8116) );
  NAND U8326 ( .A(n8117), .B(n8116), .Z(n8210) );
  NANDN U8327 ( .A(n9891), .B(n8118), .Z(n8120) );
  XOR U8328 ( .A(b[13]), .B(a[101]), .Z(n8216) );
  NANDN U8329 ( .A(n9935), .B(n8216), .Z(n8119) );
  AND U8330 ( .A(n8120), .B(n8119), .Z(n8208) );
  AND U8331 ( .A(b[15]), .B(a[97]), .Z(n8207) );
  XNOR U8332 ( .A(n8208), .B(n8207), .Z(n8209) );
  XNOR U8333 ( .A(n8210), .B(n8209), .Z(n8228) );
  NANDN U8334 ( .A(n9437), .B(n8121), .Z(n8123) );
  XOR U8335 ( .A(b[5]), .B(a[109]), .Z(n8219) );
  NANDN U8336 ( .A(n9503), .B(n8219), .Z(n8122) );
  AND U8337 ( .A(n8123), .B(n8122), .Z(n8204) );
  NANDN U8338 ( .A(n9588), .B(n8124), .Z(n8126) );
  XOR U8339 ( .A(b[7]), .B(a[107]), .Z(n8222) );
  NANDN U8340 ( .A(n9639), .B(n8222), .Z(n8125) );
  AND U8341 ( .A(n8126), .B(n8125), .Z(n8202) );
  NANDN U8342 ( .A(n9374), .B(n8127), .Z(n8129) );
  XOR U8343 ( .A(b[3]), .B(a[111]), .Z(n8225) );
  NANDN U8344 ( .A(n9375), .B(n8225), .Z(n8128) );
  NAND U8345 ( .A(n8129), .B(n8128), .Z(n8201) );
  XNOR U8346 ( .A(n8202), .B(n8201), .Z(n8203) );
  XOR U8347 ( .A(n8204), .B(n8203), .Z(n8229) );
  XOR U8348 ( .A(n8228), .B(n8229), .Z(n8231) );
  XOR U8349 ( .A(n8230), .B(n8231), .Z(n8181) );
  NANDN U8350 ( .A(n8131), .B(n8130), .Z(n8135) );
  OR U8351 ( .A(n8133), .B(n8132), .Z(n8134) );
  AND U8352 ( .A(n8135), .B(n8134), .Z(n8180) );
  XNOR U8353 ( .A(n8181), .B(n8180), .Z(n8183) );
  NAND U8354 ( .A(n8136), .B(n9883), .Z(n8138) );
  XOR U8355 ( .A(b[11]), .B(a[103]), .Z(n8186) );
  NANDN U8356 ( .A(n9856), .B(n8186), .Z(n8137) );
  AND U8357 ( .A(n8138), .B(n8137), .Z(n8197) );
  NANDN U8358 ( .A(n10005), .B(n8139), .Z(n8141) );
  XOR U8359 ( .A(b[15]), .B(a[99]), .Z(n8189) );
  NANDN U8360 ( .A(n10006), .B(n8189), .Z(n8140) );
  AND U8361 ( .A(n8141), .B(n8140), .Z(n8196) );
  NANDN U8362 ( .A(n9685), .B(n8142), .Z(n8144) );
  XOR U8363 ( .A(b[9]), .B(a[105]), .Z(n8192) );
  NANDN U8364 ( .A(n9758), .B(n8192), .Z(n8143) );
  NAND U8365 ( .A(n8144), .B(n8143), .Z(n8195) );
  XOR U8366 ( .A(n8196), .B(n8195), .Z(n8198) );
  XOR U8367 ( .A(n8197), .B(n8198), .Z(n8235) );
  NANDN U8368 ( .A(n8146), .B(n8145), .Z(n8150) );
  OR U8369 ( .A(n8148), .B(n8147), .Z(n8149) );
  AND U8370 ( .A(n8150), .B(n8149), .Z(n8234) );
  XNOR U8371 ( .A(n8235), .B(n8234), .Z(n8236) );
  NANDN U8372 ( .A(n8152), .B(n8151), .Z(n8156) );
  NANDN U8373 ( .A(n8154), .B(n8153), .Z(n8155) );
  NAND U8374 ( .A(n8156), .B(n8155), .Z(n8237) );
  XNOR U8375 ( .A(n8236), .B(n8237), .Z(n8182) );
  XOR U8376 ( .A(n8183), .B(n8182), .Z(n8241) );
  NANDN U8377 ( .A(n8158), .B(n8157), .Z(n8162) );
  NANDN U8378 ( .A(n8160), .B(n8159), .Z(n8161) );
  AND U8379 ( .A(n8162), .B(n8161), .Z(n8240) );
  XNOR U8380 ( .A(n8241), .B(n8240), .Z(n8242) );
  XOR U8381 ( .A(n8243), .B(n8242), .Z(n8175) );
  NANDN U8382 ( .A(n8164), .B(n8163), .Z(n8168) );
  NAND U8383 ( .A(n8166), .B(n8165), .Z(n8167) );
  AND U8384 ( .A(n8168), .B(n8167), .Z(n8174) );
  XNOR U8385 ( .A(n8175), .B(n8174), .Z(n8176) );
  XNOR U8386 ( .A(n8177), .B(n8176), .Z(n8246) );
  XNOR U8387 ( .A(sreg[225]), .B(n8246), .Z(n8248) );
  NANDN U8388 ( .A(sreg[224]), .B(n8169), .Z(n8173) );
  NAND U8389 ( .A(n8171), .B(n8170), .Z(n8172) );
  NAND U8390 ( .A(n8173), .B(n8172), .Z(n8247) );
  XNOR U8391 ( .A(n8248), .B(n8247), .Z(c[225]) );
  NANDN U8392 ( .A(n8175), .B(n8174), .Z(n8179) );
  NANDN U8393 ( .A(n8177), .B(n8176), .Z(n8178) );
  AND U8394 ( .A(n8179), .B(n8178), .Z(n8254) );
  NANDN U8395 ( .A(n8181), .B(n8180), .Z(n8185) );
  NAND U8396 ( .A(n8183), .B(n8182), .Z(n8184) );
  AND U8397 ( .A(n8185), .B(n8184), .Z(n8320) );
  NAND U8398 ( .A(n8186), .B(n9883), .Z(n8188) );
  XOR U8399 ( .A(b[11]), .B(a[104]), .Z(n8290) );
  NANDN U8400 ( .A(n9856), .B(n8290), .Z(n8187) );
  AND U8401 ( .A(n8188), .B(n8187), .Z(n8301) );
  NANDN U8402 ( .A(n10005), .B(n8189), .Z(n8191) );
  XOR U8403 ( .A(b[15]), .B(a[100]), .Z(n8293) );
  NANDN U8404 ( .A(n10006), .B(n8293), .Z(n8190) );
  AND U8405 ( .A(n8191), .B(n8190), .Z(n8300) );
  NANDN U8406 ( .A(n9685), .B(n8192), .Z(n8194) );
  XOR U8407 ( .A(b[9]), .B(a[106]), .Z(n8296) );
  NANDN U8408 ( .A(n9758), .B(n8296), .Z(n8193) );
  NAND U8409 ( .A(n8194), .B(n8193), .Z(n8299) );
  XOR U8410 ( .A(n8300), .B(n8299), .Z(n8302) );
  XOR U8411 ( .A(n8301), .B(n8302), .Z(n8312) );
  NANDN U8412 ( .A(n8196), .B(n8195), .Z(n8200) );
  OR U8413 ( .A(n8198), .B(n8197), .Z(n8199) );
  AND U8414 ( .A(n8200), .B(n8199), .Z(n8311) );
  XNOR U8415 ( .A(n8312), .B(n8311), .Z(n8313) );
  NANDN U8416 ( .A(n8202), .B(n8201), .Z(n8206) );
  NANDN U8417 ( .A(n8204), .B(n8203), .Z(n8205) );
  NAND U8418 ( .A(n8206), .B(n8205), .Z(n8314) );
  XNOR U8419 ( .A(n8313), .B(n8314), .Z(n8260) );
  NANDN U8420 ( .A(n8208), .B(n8207), .Z(n8212) );
  NANDN U8421 ( .A(n8210), .B(n8209), .Z(n8211) );
  AND U8422 ( .A(n8212), .B(n8211), .Z(n8286) );
  NAND U8423 ( .A(b[0]), .B(a[114]), .Z(n8213) );
  XNOR U8424 ( .A(b[1]), .B(n8213), .Z(n8215) );
  NANDN U8425 ( .A(b[0]), .B(a[113]), .Z(n8214) );
  NAND U8426 ( .A(n8215), .B(n8214), .Z(n8266) );
  NANDN U8427 ( .A(n9891), .B(n8216), .Z(n8218) );
  XOR U8428 ( .A(b[13]), .B(a[102]), .Z(n8269) );
  NANDN U8429 ( .A(n9935), .B(n8269), .Z(n8217) );
  AND U8430 ( .A(n8218), .B(n8217), .Z(n8264) );
  AND U8431 ( .A(b[15]), .B(a[98]), .Z(n8263) );
  XNOR U8432 ( .A(n8264), .B(n8263), .Z(n8265) );
  XNOR U8433 ( .A(n8266), .B(n8265), .Z(n8284) );
  NANDN U8434 ( .A(n9437), .B(n8219), .Z(n8221) );
  XOR U8435 ( .A(b[5]), .B(a[110]), .Z(n8275) );
  NANDN U8436 ( .A(n9503), .B(n8275), .Z(n8220) );
  AND U8437 ( .A(n8221), .B(n8220), .Z(n8308) );
  NANDN U8438 ( .A(n9588), .B(n8222), .Z(n8224) );
  XOR U8439 ( .A(b[7]), .B(a[108]), .Z(n8278) );
  NANDN U8440 ( .A(n9639), .B(n8278), .Z(n8223) );
  AND U8441 ( .A(n8224), .B(n8223), .Z(n8306) );
  NANDN U8442 ( .A(n9374), .B(n8225), .Z(n8227) );
  XOR U8443 ( .A(b[3]), .B(a[112]), .Z(n8281) );
  NANDN U8444 ( .A(n9375), .B(n8281), .Z(n8226) );
  NAND U8445 ( .A(n8227), .B(n8226), .Z(n8305) );
  XNOR U8446 ( .A(n8306), .B(n8305), .Z(n8307) );
  XOR U8447 ( .A(n8308), .B(n8307), .Z(n8285) );
  XOR U8448 ( .A(n8284), .B(n8285), .Z(n8287) );
  XOR U8449 ( .A(n8286), .B(n8287), .Z(n8258) );
  NANDN U8450 ( .A(n8229), .B(n8228), .Z(n8233) );
  OR U8451 ( .A(n8231), .B(n8230), .Z(n8232) );
  AND U8452 ( .A(n8233), .B(n8232), .Z(n8257) );
  XNOR U8453 ( .A(n8258), .B(n8257), .Z(n8259) );
  XOR U8454 ( .A(n8260), .B(n8259), .Z(n8318) );
  NANDN U8455 ( .A(n8235), .B(n8234), .Z(n8239) );
  NANDN U8456 ( .A(n8237), .B(n8236), .Z(n8238) );
  AND U8457 ( .A(n8239), .B(n8238), .Z(n8317) );
  XNOR U8458 ( .A(n8318), .B(n8317), .Z(n8319) );
  XOR U8459 ( .A(n8320), .B(n8319), .Z(n8252) );
  NANDN U8460 ( .A(n8241), .B(n8240), .Z(n8245) );
  NAND U8461 ( .A(n8243), .B(n8242), .Z(n8244) );
  AND U8462 ( .A(n8245), .B(n8244), .Z(n8251) );
  XNOR U8463 ( .A(n8252), .B(n8251), .Z(n8253) );
  XNOR U8464 ( .A(n8254), .B(n8253), .Z(n8323) );
  XNOR U8465 ( .A(sreg[226]), .B(n8323), .Z(n8325) );
  NANDN U8466 ( .A(sreg[225]), .B(n8246), .Z(n8250) );
  NAND U8467 ( .A(n8248), .B(n8247), .Z(n8249) );
  NAND U8468 ( .A(n8250), .B(n8249), .Z(n8324) );
  XNOR U8469 ( .A(n8325), .B(n8324), .Z(c[226]) );
  NANDN U8470 ( .A(n8252), .B(n8251), .Z(n8256) );
  NANDN U8471 ( .A(n8254), .B(n8253), .Z(n8255) );
  AND U8472 ( .A(n8256), .B(n8255), .Z(n8331) );
  NANDN U8473 ( .A(n8258), .B(n8257), .Z(n8262) );
  NAND U8474 ( .A(n8260), .B(n8259), .Z(n8261) );
  AND U8475 ( .A(n8262), .B(n8261), .Z(n8397) );
  NANDN U8476 ( .A(n8264), .B(n8263), .Z(n8268) );
  NANDN U8477 ( .A(n8266), .B(n8265), .Z(n8267) );
  AND U8478 ( .A(n8268), .B(n8267), .Z(n8363) );
  NANDN U8479 ( .A(n9891), .B(n8269), .Z(n8271) );
  XOR U8480 ( .A(b[13]), .B(a[103]), .Z(n8349) );
  NANDN U8481 ( .A(n9935), .B(n8349), .Z(n8270) );
  AND U8482 ( .A(n8271), .B(n8270), .Z(n8341) );
  AND U8483 ( .A(b[15]), .B(a[99]), .Z(n8340) );
  XNOR U8484 ( .A(n8341), .B(n8340), .Z(n8342) );
  NAND U8485 ( .A(b[0]), .B(a[115]), .Z(n8272) );
  XNOR U8486 ( .A(b[1]), .B(n8272), .Z(n8274) );
  NANDN U8487 ( .A(b[0]), .B(a[114]), .Z(n8273) );
  NAND U8488 ( .A(n8274), .B(n8273), .Z(n8343) );
  XNOR U8489 ( .A(n8342), .B(n8343), .Z(n8361) );
  NANDN U8490 ( .A(n9437), .B(n8275), .Z(n8277) );
  XOR U8491 ( .A(b[5]), .B(a[111]), .Z(n8352) );
  NANDN U8492 ( .A(n9503), .B(n8352), .Z(n8276) );
  AND U8493 ( .A(n8277), .B(n8276), .Z(n8385) );
  NANDN U8494 ( .A(n9588), .B(n8278), .Z(n8280) );
  XOR U8495 ( .A(b[7]), .B(a[109]), .Z(n8355) );
  NANDN U8496 ( .A(n9639), .B(n8355), .Z(n8279) );
  AND U8497 ( .A(n8280), .B(n8279), .Z(n8383) );
  NANDN U8498 ( .A(n9374), .B(n8281), .Z(n8283) );
  XOR U8499 ( .A(b[3]), .B(a[113]), .Z(n8358) );
  NANDN U8500 ( .A(n9375), .B(n8358), .Z(n8282) );
  NAND U8501 ( .A(n8283), .B(n8282), .Z(n8382) );
  XNOR U8502 ( .A(n8383), .B(n8382), .Z(n8384) );
  XOR U8503 ( .A(n8385), .B(n8384), .Z(n8362) );
  XOR U8504 ( .A(n8361), .B(n8362), .Z(n8364) );
  XOR U8505 ( .A(n8363), .B(n8364), .Z(n8335) );
  NANDN U8506 ( .A(n8285), .B(n8284), .Z(n8289) );
  OR U8507 ( .A(n8287), .B(n8286), .Z(n8288) );
  AND U8508 ( .A(n8289), .B(n8288), .Z(n8334) );
  XNOR U8509 ( .A(n8335), .B(n8334), .Z(n8337) );
  NAND U8510 ( .A(n8290), .B(n9883), .Z(n8292) );
  XOR U8511 ( .A(b[11]), .B(a[105]), .Z(n8367) );
  NANDN U8512 ( .A(n9856), .B(n8367), .Z(n8291) );
  AND U8513 ( .A(n8292), .B(n8291), .Z(n8378) );
  NANDN U8514 ( .A(n10005), .B(n8293), .Z(n8295) );
  XOR U8515 ( .A(b[15]), .B(a[101]), .Z(n8370) );
  NANDN U8516 ( .A(n10006), .B(n8370), .Z(n8294) );
  AND U8517 ( .A(n8295), .B(n8294), .Z(n8377) );
  NANDN U8518 ( .A(n9685), .B(n8296), .Z(n8298) );
  XOR U8519 ( .A(b[9]), .B(a[107]), .Z(n8373) );
  NANDN U8520 ( .A(n9758), .B(n8373), .Z(n8297) );
  NAND U8521 ( .A(n8298), .B(n8297), .Z(n8376) );
  XOR U8522 ( .A(n8377), .B(n8376), .Z(n8379) );
  XOR U8523 ( .A(n8378), .B(n8379), .Z(n8389) );
  NANDN U8524 ( .A(n8300), .B(n8299), .Z(n8304) );
  OR U8525 ( .A(n8302), .B(n8301), .Z(n8303) );
  AND U8526 ( .A(n8304), .B(n8303), .Z(n8388) );
  XNOR U8527 ( .A(n8389), .B(n8388), .Z(n8390) );
  NANDN U8528 ( .A(n8306), .B(n8305), .Z(n8310) );
  NANDN U8529 ( .A(n8308), .B(n8307), .Z(n8309) );
  NAND U8530 ( .A(n8310), .B(n8309), .Z(n8391) );
  XNOR U8531 ( .A(n8390), .B(n8391), .Z(n8336) );
  XOR U8532 ( .A(n8337), .B(n8336), .Z(n8395) );
  NANDN U8533 ( .A(n8312), .B(n8311), .Z(n8316) );
  NANDN U8534 ( .A(n8314), .B(n8313), .Z(n8315) );
  AND U8535 ( .A(n8316), .B(n8315), .Z(n8394) );
  XNOR U8536 ( .A(n8395), .B(n8394), .Z(n8396) );
  XOR U8537 ( .A(n8397), .B(n8396), .Z(n8329) );
  NANDN U8538 ( .A(n8318), .B(n8317), .Z(n8322) );
  NAND U8539 ( .A(n8320), .B(n8319), .Z(n8321) );
  AND U8540 ( .A(n8322), .B(n8321), .Z(n8328) );
  XNOR U8541 ( .A(n8329), .B(n8328), .Z(n8330) );
  XNOR U8542 ( .A(n8331), .B(n8330), .Z(n8400) );
  XNOR U8543 ( .A(sreg[227]), .B(n8400), .Z(n8402) );
  NANDN U8544 ( .A(sreg[226]), .B(n8323), .Z(n8327) );
  NAND U8545 ( .A(n8325), .B(n8324), .Z(n8326) );
  NAND U8546 ( .A(n8327), .B(n8326), .Z(n8401) );
  XNOR U8547 ( .A(n8402), .B(n8401), .Z(c[227]) );
  NANDN U8548 ( .A(n8329), .B(n8328), .Z(n8333) );
  NANDN U8549 ( .A(n8331), .B(n8330), .Z(n8332) );
  AND U8550 ( .A(n8333), .B(n8332), .Z(n8408) );
  NANDN U8551 ( .A(n8335), .B(n8334), .Z(n8339) );
  NAND U8552 ( .A(n8337), .B(n8336), .Z(n8338) );
  AND U8553 ( .A(n8339), .B(n8338), .Z(n8474) );
  NANDN U8554 ( .A(n8341), .B(n8340), .Z(n8345) );
  NANDN U8555 ( .A(n8343), .B(n8342), .Z(n8344) );
  AND U8556 ( .A(n8345), .B(n8344), .Z(n8440) );
  NAND U8557 ( .A(b[0]), .B(a[116]), .Z(n8346) );
  XNOR U8558 ( .A(b[1]), .B(n8346), .Z(n8348) );
  NANDN U8559 ( .A(b[0]), .B(a[115]), .Z(n8347) );
  NAND U8560 ( .A(n8348), .B(n8347), .Z(n8420) );
  NANDN U8561 ( .A(n9891), .B(n8349), .Z(n8351) );
  XOR U8562 ( .A(b[13]), .B(a[104]), .Z(n8426) );
  NANDN U8563 ( .A(n9935), .B(n8426), .Z(n8350) );
  AND U8564 ( .A(n8351), .B(n8350), .Z(n8418) );
  AND U8565 ( .A(b[15]), .B(a[100]), .Z(n8417) );
  XNOR U8566 ( .A(n8418), .B(n8417), .Z(n8419) );
  XNOR U8567 ( .A(n8420), .B(n8419), .Z(n8438) );
  NANDN U8568 ( .A(n9437), .B(n8352), .Z(n8354) );
  XOR U8569 ( .A(b[5]), .B(a[112]), .Z(n8429) );
  NANDN U8570 ( .A(n9503), .B(n8429), .Z(n8353) );
  AND U8571 ( .A(n8354), .B(n8353), .Z(n8462) );
  NANDN U8572 ( .A(n9588), .B(n8355), .Z(n8357) );
  XOR U8573 ( .A(b[7]), .B(a[110]), .Z(n8432) );
  NANDN U8574 ( .A(n9639), .B(n8432), .Z(n8356) );
  AND U8575 ( .A(n8357), .B(n8356), .Z(n8460) );
  NANDN U8576 ( .A(n9374), .B(n8358), .Z(n8360) );
  XOR U8577 ( .A(b[3]), .B(a[114]), .Z(n8435) );
  NANDN U8578 ( .A(n9375), .B(n8435), .Z(n8359) );
  NAND U8579 ( .A(n8360), .B(n8359), .Z(n8459) );
  XNOR U8580 ( .A(n8460), .B(n8459), .Z(n8461) );
  XOR U8581 ( .A(n8462), .B(n8461), .Z(n8439) );
  XOR U8582 ( .A(n8438), .B(n8439), .Z(n8441) );
  XOR U8583 ( .A(n8440), .B(n8441), .Z(n8412) );
  NANDN U8584 ( .A(n8362), .B(n8361), .Z(n8366) );
  OR U8585 ( .A(n8364), .B(n8363), .Z(n8365) );
  AND U8586 ( .A(n8366), .B(n8365), .Z(n8411) );
  XNOR U8587 ( .A(n8412), .B(n8411), .Z(n8414) );
  NAND U8588 ( .A(n8367), .B(n9883), .Z(n8369) );
  XOR U8589 ( .A(b[11]), .B(a[106]), .Z(n8444) );
  NANDN U8590 ( .A(n9856), .B(n8444), .Z(n8368) );
  AND U8591 ( .A(n8369), .B(n8368), .Z(n8455) );
  NANDN U8592 ( .A(n10005), .B(n8370), .Z(n8372) );
  XOR U8593 ( .A(b[15]), .B(a[102]), .Z(n8447) );
  NANDN U8594 ( .A(n10006), .B(n8447), .Z(n8371) );
  AND U8595 ( .A(n8372), .B(n8371), .Z(n8454) );
  NANDN U8596 ( .A(n9685), .B(n8373), .Z(n8375) );
  XOR U8597 ( .A(b[9]), .B(a[108]), .Z(n8450) );
  NANDN U8598 ( .A(n9758), .B(n8450), .Z(n8374) );
  NAND U8599 ( .A(n8375), .B(n8374), .Z(n8453) );
  XOR U8600 ( .A(n8454), .B(n8453), .Z(n8456) );
  XOR U8601 ( .A(n8455), .B(n8456), .Z(n8466) );
  NANDN U8602 ( .A(n8377), .B(n8376), .Z(n8381) );
  OR U8603 ( .A(n8379), .B(n8378), .Z(n8380) );
  AND U8604 ( .A(n8381), .B(n8380), .Z(n8465) );
  XNOR U8605 ( .A(n8466), .B(n8465), .Z(n8467) );
  NANDN U8606 ( .A(n8383), .B(n8382), .Z(n8387) );
  NANDN U8607 ( .A(n8385), .B(n8384), .Z(n8386) );
  NAND U8608 ( .A(n8387), .B(n8386), .Z(n8468) );
  XNOR U8609 ( .A(n8467), .B(n8468), .Z(n8413) );
  XOR U8610 ( .A(n8414), .B(n8413), .Z(n8472) );
  NANDN U8611 ( .A(n8389), .B(n8388), .Z(n8393) );
  NANDN U8612 ( .A(n8391), .B(n8390), .Z(n8392) );
  AND U8613 ( .A(n8393), .B(n8392), .Z(n8471) );
  XNOR U8614 ( .A(n8472), .B(n8471), .Z(n8473) );
  XOR U8615 ( .A(n8474), .B(n8473), .Z(n8406) );
  NANDN U8616 ( .A(n8395), .B(n8394), .Z(n8399) );
  NAND U8617 ( .A(n8397), .B(n8396), .Z(n8398) );
  AND U8618 ( .A(n8399), .B(n8398), .Z(n8405) );
  XNOR U8619 ( .A(n8406), .B(n8405), .Z(n8407) );
  XNOR U8620 ( .A(n8408), .B(n8407), .Z(n8477) );
  XNOR U8621 ( .A(sreg[228]), .B(n8477), .Z(n8479) );
  NANDN U8622 ( .A(sreg[227]), .B(n8400), .Z(n8404) );
  NAND U8623 ( .A(n8402), .B(n8401), .Z(n8403) );
  NAND U8624 ( .A(n8404), .B(n8403), .Z(n8478) );
  XNOR U8625 ( .A(n8479), .B(n8478), .Z(c[228]) );
  NANDN U8626 ( .A(n8406), .B(n8405), .Z(n8410) );
  NANDN U8627 ( .A(n8408), .B(n8407), .Z(n8409) );
  AND U8628 ( .A(n8410), .B(n8409), .Z(n8485) );
  NANDN U8629 ( .A(n8412), .B(n8411), .Z(n8416) );
  NAND U8630 ( .A(n8414), .B(n8413), .Z(n8415) );
  AND U8631 ( .A(n8416), .B(n8415), .Z(n8551) );
  NANDN U8632 ( .A(n8418), .B(n8417), .Z(n8422) );
  NANDN U8633 ( .A(n8420), .B(n8419), .Z(n8421) );
  AND U8634 ( .A(n8422), .B(n8421), .Z(n8517) );
  NAND U8635 ( .A(b[0]), .B(a[117]), .Z(n8423) );
  XNOR U8636 ( .A(b[1]), .B(n8423), .Z(n8425) );
  NANDN U8637 ( .A(b[0]), .B(a[116]), .Z(n8424) );
  NAND U8638 ( .A(n8425), .B(n8424), .Z(n8497) );
  NANDN U8639 ( .A(n9891), .B(n8426), .Z(n8428) );
  XOR U8640 ( .A(b[13]), .B(a[105]), .Z(n8503) );
  NANDN U8641 ( .A(n9935), .B(n8503), .Z(n8427) );
  AND U8642 ( .A(n8428), .B(n8427), .Z(n8495) );
  AND U8643 ( .A(b[15]), .B(a[101]), .Z(n8494) );
  XNOR U8644 ( .A(n8495), .B(n8494), .Z(n8496) );
  XNOR U8645 ( .A(n8497), .B(n8496), .Z(n8515) );
  NANDN U8646 ( .A(n9437), .B(n8429), .Z(n8431) );
  XOR U8647 ( .A(b[5]), .B(a[113]), .Z(n8506) );
  NANDN U8648 ( .A(n9503), .B(n8506), .Z(n8430) );
  AND U8649 ( .A(n8431), .B(n8430), .Z(n8539) );
  NANDN U8650 ( .A(n9588), .B(n8432), .Z(n8434) );
  XOR U8651 ( .A(b[7]), .B(a[111]), .Z(n8509) );
  NANDN U8652 ( .A(n9639), .B(n8509), .Z(n8433) );
  AND U8653 ( .A(n8434), .B(n8433), .Z(n8537) );
  NANDN U8654 ( .A(n9374), .B(n8435), .Z(n8437) );
  XOR U8655 ( .A(b[3]), .B(a[115]), .Z(n8512) );
  NANDN U8656 ( .A(n9375), .B(n8512), .Z(n8436) );
  NAND U8657 ( .A(n8437), .B(n8436), .Z(n8536) );
  XNOR U8658 ( .A(n8537), .B(n8536), .Z(n8538) );
  XOR U8659 ( .A(n8539), .B(n8538), .Z(n8516) );
  XOR U8660 ( .A(n8515), .B(n8516), .Z(n8518) );
  XOR U8661 ( .A(n8517), .B(n8518), .Z(n8489) );
  NANDN U8662 ( .A(n8439), .B(n8438), .Z(n8443) );
  OR U8663 ( .A(n8441), .B(n8440), .Z(n8442) );
  AND U8664 ( .A(n8443), .B(n8442), .Z(n8488) );
  XNOR U8665 ( .A(n8489), .B(n8488), .Z(n8491) );
  NAND U8666 ( .A(n8444), .B(n9883), .Z(n8446) );
  XOR U8667 ( .A(b[11]), .B(a[107]), .Z(n8521) );
  NANDN U8668 ( .A(n9856), .B(n8521), .Z(n8445) );
  AND U8669 ( .A(n8446), .B(n8445), .Z(n8532) );
  NANDN U8670 ( .A(n10005), .B(n8447), .Z(n8449) );
  XOR U8671 ( .A(b[15]), .B(a[103]), .Z(n8524) );
  NANDN U8672 ( .A(n10006), .B(n8524), .Z(n8448) );
  AND U8673 ( .A(n8449), .B(n8448), .Z(n8531) );
  NANDN U8674 ( .A(n9685), .B(n8450), .Z(n8452) );
  XOR U8675 ( .A(b[9]), .B(a[109]), .Z(n8527) );
  NANDN U8676 ( .A(n9758), .B(n8527), .Z(n8451) );
  NAND U8677 ( .A(n8452), .B(n8451), .Z(n8530) );
  XOR U8678 ( .A(n8531), .B(n8530), .Z(n8533) );
  XOR U8679 ( .A(n8532), .B(n8533), .Z(n8543) );
  NANDN U8680 ( .A(n8454), .B(n8453), .Z(n8458) );
  OR U8681 ( .A(n8456), .B(n8455), .Z(n8457) );
  AND U8682 ( .A(n8458), .B(n8457), .Z(n8542) );
  XNOR U8683 ( .A(n8543), .B(n8542), .Z(n8544) );
  NANDN U8684 ( .A(n8460), .B(n8459), .Z(n8464) );
  NANDN U8685 ( .A(n8462), .B(n8461), .Z(n8463) );
  NAND U8686 ( .A(n8464), .B(n8463), .Z(n8545) );
  XNOR U8687 ( .A(n8544), .B(n8545), .Z(n8490) );
  XOR U8688 ( .A(n8491), .B(n8490), .Z(n8549) );
  NANDN U8689 ( .A(n8466), .B(n8465), .Z(n8470) );
  NANDN U8690 ( .A(n8468), .B(n8467), .Z(n8469) );
  AND U8691 ( .A(n8470), .B(n8469), .Z(n8548) );
  XNOR U8692 ( .A(n8549), .B(n8548), .Z(n8550) );
  XOR U8693 ( .A(n8551), .B(n8550), .Z(n8483) );
  NANDN U8694 ( .A(n8472), .B(n8471), .Z(n8476) );
  NAND U8695 ( .A(n8474), .B(n8473), .Z(n8475) );
  AND U8696 ( .A(n8476), .B(n8475), .Z(n8482) );
  XNOR U8697 ( .A(n8483), .B(n8482), .Z(n8484) );
  XNOR U8698 ( .A(n8485), .B(n8484), .Z(n8554) );
  XNOR U8699 ( .A(sreg[229]), .B(n8554), .Z(n8556) );
  NANDN U8700 ( .A(sreg[228]), .B(n8477), .Z(n8481) );
  NAND U8701 ( .A(n8479), .B(n8478), .Z(n8480) );
  NAND U8702 ( .A(n8481), .B(n8480), .Z(n8555) );
  XNOR U8703 ( .A(n8556), .B(n8555), .Z(c[229]) );
  NANDN U8704 ( .A(n8483), .B(n8482), .Z(n8487) );
  NANDN U8705 ( .A(n8485), .B(n8484), .Z(n8486) );
  AND U8706 ( .A(n8487), .B(n8486), .Z(n8562) );
  NANDN U8707 ( .A(n8489), .B(n8488), .Z(n8493) );
  NAND U8708 ( .A(n8491), .B(n8490), .Z(n8492) );
  AND U8709 ( .A(n8493), .B(n8492), .Z(n8628) );
  NANDN U8710 ( .A(n8495), .B(n8494), .Z(n8499) );
  NANDN U8711 ( .A(n8497), .B(n8496), .Z(n8498) );
  AND U8712 ( .A(n8499), .B(n8498), .Z(n8594) );
  NAND U8713 ( .A(b[0]), .B(a[118]), .Z(n8500) );
  XNOR U8714 ( .A(b[1]), .B(n8500), .Z(n8502) );
  NANDN U8715 ( .A(b[0]), .B(a[117]), .Z(n8501) );
  NAND U8716 ( .A(n8502), .B(n8501), .Z(n8574) );
  NANDN U8717 ( .A(n9891), .B(n8503), .Z(n8505) );
  XOR U8718 ( .A(b[13]), .B(a[106]), .Z(n8580) );
  NANDN U8719 ( .A(n9935), .B(n8580), .Z(n8504) );
  AND U8720 ( .A(n8505), .B(n8504), .Z(n8572) );
  AND U8721 ( .A(b[15]), .B(a[102]), .Z(n8571) );
  XNOR U8722 ( .A(n8572), .B(n8571), .Z(n8573) );
  XNOR U8723 ( .A(n8574), .B(n8573), .Z(n8592) );
  NANDN U8724 ( .A(n9437), .B(n8506), .Z(n8508) );
  XOR U8725 ( .A(b[5]), .B(a[114]), .Z(n8583) );
  NANDN U8726 ( .A(n9503), .B(n8583), .Z(n8507) );
  AND U8727 ( .A(n8508), .B(n8507), .Z(n8616) );
  NANDN U8728 ( .A(n9588), .B(n8509), .Z(n8511) );
  XOR U8729 ( .A(b[7]), .B(a[112]), .Z(n8586) );
  NANDN U8730 ( .A(n9639), .B(n8586), .Z(n8510) );
  AND U8731 ( .A(n8511), .B(n8510), .Z(n8614) );
  NANDN U8732 ( .A(n9374), .B(n8512), .Z(n8514) );
  XOR U8733 ( .A(b[3]), .B(a[116]), .Z(n8589) );
  NANDN U8734 ( .A(n9375), .B(n8589), .Z(n8513) );
  NAND U8735 ( .A(n8514), .B(n8513), .Z(n8613) );
  XNOR U8736 ( .A(n8614), .B(n8613), .Z(n8615) );
  XOR U8737 ( .A(n8616), .B(n8615), .Z(n8593) );
  XOR U8738 ( .A(n8592), .B(n8593), .Z(n8595) );
  XOR U8739 ( .A(n8594), .B(n8595), .Z(n8566) );
  NANDN U8740 ( .A(n8516), .B(n8515), .Z(n8520) );
  OR U8741 ( .A(n8518), .B(n8517), .Z(n8519) );
  AND U8742 ( .A(n8520), .B(n8519), .Z(n8565) );
  XNOR U8743 ( .A(n8566), .B(n8565), .Z(n8568) );
  NAND U8744 ( .A(n8521), .B(n9883), .Z(n8523) );
  XOR U8745 ( .A(b[11]), .B(a[108]), .Z(n8598) );
  NANDN U8746 ( .A(n9856), .B(n8598), .Z(n8522) );
  AND U8747 ( .A(n8523), .B(n8522), .Z(n8609) );
  NANDN U8748 ( .A(n10005), .B(n8524), .Z(n8526) );
  XOR U8749 ( .A(b[15]), .B(a[104]), .Z(n8601) );
  NANDN U8750 ( .A(n10006), .B(n8601), .Z(n8525) );
  AND U8751 ( .A(n8526), .B(n8525), .Z(n8608) );
  NANDN U8752 ( .A(n9685), .B(n8527), .Z(n8529) );
  XOR U8753 ( .A(b[9]), .B(a[110]), .Z(n8604) );
  NANDN U8754 ( .A(n9758), .B(n8604), .Z(n8528) );
  NAND U8755 ( .A(n8529), .B(n8528), .Z(n8607) );
  XOR U8756 ( .A(n8608), .B(n8607), .Z(n8610) );
  XOR U8757 ( .A(n8609), .B(n8610), .Z(n8620) );
  NANDN U8758 ( .A(n8531), .B(n8530), .Z(n8535) );
  OR U8759 ( .A(n8533), .B(n8532), .Z(n8534) );
  AND U8760 ( .A(n8535), .B(n8534), .Z(n8619) );
  XNOR U8761 ( .A(n8620), .B(n8619), .Z(n8621) );
  NANDN U8762 ( .A(n8537), .B(n8536), .Z(n8541) );
  NANDN U8763 ( .A(n8539), .B(n8538), .Z(n8540) );
  NAND U8764 ( .A(n8541), .B(n8540), .Z(n8622) );
  XNOR U8765 ( .A(n8621), .B(n8622), .Z(n8567) );
  XOR U8766 ( .A(n8568), .B(n8567), .Z(n8626) );
  NANDN U8767 ( .A(n8543), .B(n8542), .Z(n8547) );
  NANDN U8768 ( .A(n8545), .B(n8544), .Z(n8546) );
  AND U8769 ( .A(n8547), .B(n8546), .Z(n8625) );
  XNOR U8770 ( .A(n8626), .B(n8625), .Z(n8627) );
  XOR U8771 ( .A(n8628), .B(n8627), .Z(n8560) );
  NANDN U8772 ( .A(n8549), .B(n8548), .Z(n8553) );
  NAND U8773 ( .A(n8551), .B(n8550), .Z(n8552) );
  AND U8774 ( .A(n8553), .B(n8552), .Z(n8559) );
  XNOR U8775 ( .A(n8560), .B(n8559), .Z(n8561) );
  XNOR U8776 ( .A(n8562), .B(n8561), .Z(n8631) );
  XNOR U8777 ( .A(sreg[230]), .B(n8631), .Z(n8633) );
  NANDN U8778 ( .A(sreg[229]), .B(n8554), .Z(n8558) );
  NAND U8779 ( .A(n8556), .B(n8555), .Z(n8557) );
  NAND U8780 ( .A(n8558), .B(n8557), .Z(n8632) );
  XNOR U8781 ( .A(n8633), .B(n8632), .Z(c[230]) );
  NANDN U8782 ( .A(n8560), .B(n8559), .Z(n8564) );
  NANDN U8783 ( .A(n8562), .B(n8561), .Z(n8563) );
  AND U8784 ( .A(n8564), .B(n8563), .Z(n8639) );
  NANDN U8785 ( .A(n8566), .B(n8565), .Z(n8570) );
  NAND U8786 ( .A(n8568), .B(n8567), .Z(n8569) );
  AND U8787 ( .A(n8570), .B(n8569), .Z(n8705) );
  NANDN U8788 ( .A(n8572), .B(n8571), .Z(n8576) );
  NANDN U8789 ( .A(n8574), .B(n8573), .Z(n8575) );
  AND U8790 ( .A(n8576), .B(n8575), .Z(n8671) );
  NAND U8791 ( .A(b[0]), .B(a[119]), .Z(n8577) );
  XNOR U8792 ( .A(b[1]), .B(n8577), .Z(n8579) );
  NANDN U8793 ( .A(b[0]), .B(a[118]), .Z(n8578) );
  NAND U8794 ( .A(n8579), .B(n8578), .Z(n8651) );
  NANDN U8795 ( .A(n9891), .B(n8580), .Z(n8582) );
  XOR U8796 ( .A(b[13]), .B(a[107]), .Z(n8657) );
  NANDN U8797 ( .A(n9935), .B(n8657), .Z(n8581) );
  AND U8798 ( .A(n8582), .B(n8581), .Z(n8649) );
  AND U8799 ( .A(b[15]), .B(a[103]), .Z(n8648) );
  XNOR U8800 ( .A(n8649), .B(n8648), .Z(n8650) );
  XNOR U8801 ( .A(n8651), .B(n8650), .Z(n8669) );
  NANDN U8802 ( .A(n9437), .B(n8583), .Z(n8585) );
  XOR U8803 ( .A(b[5]), .B(a[115]), .Z(n8660) );
  NANDN U8804 ( .A(n9503), .B(n8660), .Z(n8584) );
  AND U8805 ( .A(n8585), .B(n8584), .Z(n8693) );
  NANDN U8806 ( .A(n9588), .B(n8586), .Z(n8588) );
  XOR U8807 ( .A(b[7]), .B(a[113]), .Z(n8663) );
  NANDN U8808 ( .A(n9639), .B(n8663), .Z(n8587) );
  AND U8809 ( .A(n8588), .B(n8587), .Z(n8691) );
  NANDN U8810 ( .A(n9374), .B(n8589), .Z(n8591) );
  XOR U8811 ( .A(b[3]), .B(a[117]), .Z(n8666) );
  NANDN U8812 ( .A(n9375), .B(n8666), .Z(n8590) );
  NAND U8813 ( .A(n8591), .B(n8590), .Z(n8690) );
  XNOR U8814 ( .A(n8691), .B(n8690), .Z(n8692) );
  XOR U8815 ( .A(n8693), .B(n8692), .Z(n8670) );
  XOR U8816 ( .A(n8669), .B(n8670), .Z(n8672) );
  XOR U8817 ( .A(n8671), .B(n8672), .Z(n8643) );
  NANDN U8818 ( .A(n8593), .B(n8592), .Z(n8597) );
  OR U8819 ( .A(n8595), .B(n8594), .Z(n8596) );
  AND U8820 ( .A(n8597), .B(n8596), .Z(n8642) );
  XNOR U8821 ( .A(n8643), .B(n8642), .Z(n8645) );
  NAND U8822 ( .A(n8598), .B(n9883), .Z(n8600) );
  XOR U8823 ( .A(b[11]), .B(a[109]), .Z(n8675) );
  NANDN U8824 ( .A(n9856), .B(n8675), .Z(n8599) );
  AND U8825 ( .A(n8600), .B(n8599), .Z(n8686) );
  NANDN U8826 ( .A(n10005), .B(n8601), .Z(n8603) );
  XOR U8827 ( .A(b[15]), .B(a[105]), .Z(n8678) );
  NANDN U8828 ( .A(n10006), .B(n8678), .Z(n8602) );
  AND U8829 ( .A(n8603), .B(n8602), .Z(n8685) );
  NANDN U8830 ( .A(n9685), .B(n8604), .Z(n8606) );
  XOR U8831 ( .A(b[9]), .B(a[111]), .Z(n8681) );
  NANDN U8832 ( .A(n9758), .B(n8681), .Z(n8605) );
  NAND U8833 ( .A(n8606), .B(n8605), .Z(n8684) );
  XOR U8834 ( .A(n8685), .B(n8684), .Z(n8687) );
  XOR U8835 ( .A(n8686), .B(n8687), .Z(n8697) );
  NANDN U8836 ( .A(n8608), .B(n8607), .Z(n8612) );
  OR U8837 ( .A(n8610), .B(n8609), .Z(n8611) );
  AND U8838 ( .A(n8612), .B(n8611), .Z(n8696) );
  XNOR U8839 ( .A(n8697), .B(n8696), .Z(n8698) );
  NANDN U8840 ( .A(n8614), .B(n8613), .Z(n8618) );
  NANDN U8841 ( .A(n8616), .B(n8615), .Z(n8617) );
  NAND U8842 ( .A(n8618), .B(n8617), .Z(n8699) );
  XNOR U8843 ( .A(n8698), .B(n8699), .Z(n8644) );
  XOR U8844 ( .A(n8645), .B(n8644), .Z(n8703) );
  NANDN U8845 ( .A(n8620), .B(n8619), .Z(n8624) );
  NANDN U8846 ( .A(n8622), .B(n8621), .Z(n8623) );
  AND U8847 ( .A(n8624), .B(n8623), .Z(n8702) );
  XNOR U8848 ( .A(n8703), .B(n8702), .Z(n8704) );
  XOR U8849 ( .A(n8705), .B(n8704), .Z(n8637) );
  NANDN U8850 ( .A(n8626), .B(n8625), .Z(n8630) );
  NAND U8851 ( .A(n8628), .B(n8627), .Z(n8629) );
  AND U8852 ( .A(n8630), .B(n8629), .Z(n8636) );
  XNOR U8853 ( .A(n8637), .B(n8636), .Z(n8638) );
  XNOR U8854 ( .A(n8639), .B(n8638), .Z(n8708) );
  XNOR U8855 ( .A(sreg[231]), .B(n8708), .Z(n8710) );
  NANDN U8856 ( .A(sreg[230]), .B(n8631), .Z(n8635) );
  NAND U8857 ( .A(n8633), .B(n8632), .Z(n8634) );
  NAND U8858 ( .A(n8635), .B(n8634), .Z(n8709) );
  XNOR U8859 ( .A(n8710), .B(n8709), .Z(c[231]) );
  NANDN U8860 ( .A(n8637), .B(n8636), .Z(n8641) );
  NANDN U8861 ( .A(n8639), .B(n8638), .Z(n8640) );
  AND U8862 ( .A(n8641), .B(n8640), .Z(n8716) );
  NANDN U8863 ( .A(n8643), .B(n8642), .Z(n8647) );
  NAND U8864 ( .A(n8645), .B(n8644), .Z(n8646) );
  AND U8865 ( .A(n8647), .B(n8646), .Z(n8782) );
  NANDN U8866 ( .A(n8649), .B(n8648), .Z(n8653) );
  NANDN U8867 ( .A(n8651), .B(n8650), .Z(n8652) );
  AND U8868 ( .A(n8653), .B(n8652), .Z(n8748) );
  NAND U8869 ( .A(b[0]), .B(a[120]), .Z(n8654) );
  XNOR U8870 ( .A(b[1]), .B(n8654), .Z(n8656) );
  NANDN U8871 ( .A(b[0]), .B(a[119]), .Z(n8655) );
  NAND U8872 ( .A(n8656), .B(n8655), .Z(n8728) );
  NANDN U8873 ( .A(n9891), .B(n8657), .Z(n8659) );
  XOR U8874 ( .A(b[13]), .B(a[108]), .Z(n8734) );
  NANDN U8875 ( .A(n9935), .B(n8734), .Z(n8658) );
  AND U8876 ( .A(n8659), .B(n8658), .Z(n8726) );
  AND U8877 ( .A(b[15]), .B(a[104]), .Z(n8725) );
  XNOR U8878 ( .A(n8726), .B(n8725), .Z(n8727) );
  XNOR U8879 ( .A(n8728), .B(n8727), .Z(n8746) );
  NANDN U8880 ( .A(n9437), .B(n8660), .Z(n8662) );
  XOR U8881 ( .A(b[5]), .B(a[116]), .Z(n8737) );
  NANDN U8882 ( .A(n9503), .B(n8737), .Z(n8661) );
  AND U8883 ( .A(n8662), .B(n8661), .Z(n8770) );
  NANDN U8884 ( .A(n9588), .B(n8663), .Z(n8665) );
  XOR U8885 ( .A(b[7]), .B(a[114]), .Z(n8740) );
  NANDN U8886 ( .A(n9639), .B(n8740), .Z(n8664) );
  AND U8887 ( .A(n8665), .B(n8664), .Z(n8768) );
  NANDN U8888 ( .A(n9374), .B(n8666), .Z(n8668) );
  XOR U8889 ( .A(a[118]), .B(b[3]), .Z(n8743) );
  NANDN U8890 ( .A(n9375), .B(n8743), .Z(n8667) );
  NAND U8891 ( .A(n8668), .B(n8667), .Z(n8767) );
  XNOR U8892 ( .A(n8768), .B(n8767), .Z(n8769) );
  XOR U8893 ( .A(n8770), .B(n8769), .Z(n8747) );
  XOR U8894 ( .A(n8746), .B(n8747), .Z(n8749) );
  XOR U8895 ( .A(n8748), .B(n8749), .Z(n8720) );
  NANDN U8896 ( .A(n8670), .B(n8669), .Z(n8674) );
  OR U8897 ( .A(n8672), .B(n8671), .Z(n8673) );
  AND U8898 ( .A(n8674), .B(n8673), .Z(n8719) );
  XNOR U8899 ( .A(n8720), .B(n8719), .Z(n8722) );
  NAND U8900 ( .A(n8675), .B(n9883), .Z(n8677) );
  XOR U8901 ( .A(b[11]), .B(a[110]), .Z(n8752) );
  NANDN U8902 ( .A(n9856), .B(n8752), .Z(n8676) );
  AND U8903 ( .A(n8677), .B(n8676), .Z(n8763) );
  NANDN U8904 ( .A(n10005), .B(n8678), .Z(n8680) );
  XOR U8905 ( .A(b[15]), .B(a[106]), .Z(n8755) );
  NANDN U8906 ( .A(n10006), .B(n8755), .Z(n8679) );
  AND U8907 ( .A(n8680), .B(n8679), .Z(n8762) );
  NANDN U8908 ( .A(n9685), .B(n8681), .Z(n8683) );
  XOR U8909 ( .A(b[9]), .B(a[112]), .Z(n8758) );
  NANDN U8910 ( .A(n9758), .B(n8758), .Z(n8682) );
  NAND U8911 ( .A(n8683), .B(n8682), .Z(n8761) );
  XOR U8912 ( .A(n8762), .B(n8761), .Z(n8764) );
  XOR U8913 ( .A(n8763), .B(n8764), .Z(n8774) );
  NANDN U8914 ( .A(n8685), .B(n8684), .Z(n8689) );
  OR U8915 ( .A(n8687), .B(n8686), .Z(n8688) );
  AND U8916 ( .A(n8689), .B(n8688), .Z(n8773) );
  XNOR U8917 ( .A(n8774), .B(n8773), .Z(n8775) );
  NANDN U8918 ( .A(n8691), .B(n8690), .Z(n8695) );
  NANDN U8919 ( .A(n8693), .B(n8692), .Z(n8694) );
  NAND U8920 ( .A(n8695), .B(n8694), .Z(n8776) );
  XNOR U8921 ( .A(n8775), .B(n8776), .Z(n8721) );
  XOR U8922 ( .A(n8722), .B(n8721), .Z(n8780) );
  NANDN U8923 ( .A(n8697), .B(n8696), .Z(n8701) );
  NANDN U8924 ( .A(n8699), .B(n8698), .Z(n8700) );
  AND U8925 ( .A(n8701), .B(n8700), .Z(n8779) );
  XNOR U8926 ( .A(n8780), .B(n8779), .Z(n8781) );
  XOR U8927 ( .A(n8782), .B(n8781), .Z(n8714) );
  NANDN U8928 ( .A(n8703), .B(n8702), .Z(n8707) );
  NAND U8929 ( .A(n8705), .B(n8704), .Z(n8706) );
  AND U8930 ( .A(n8707), .B(n8706), .Z(n8713) );
  XNOR U8931 ( .A(n8714), .B(n8713), .Z(n8715) );
  XNOR U8932 ( .A(n8716), .B(n8715), .Z(n8785) );
  XNOR U8933 ( .A(sreg[232]), .B(n8785), .Z(n8787) );
  NANDN U8934 ( .A(sreg[231]), .B(n8708), .Z(n8712) );
  NAND U8935 ( .A(n8710), .B(n8709), .Z(n8711) );
  NAND U8936 ( .A(n8712), .B(n8711), .Z(n8786) );
  XNOR U8937 ( .A(n8787), .B(n8786), .Z(c[232]) );
  NANDN U8938 ( .A(n8714), .B(n8713), .Z(n8718) );
  NANDN U8939 ( .A(n8716), .B(n8715), .Z(n8717) );
  AND U8940 ( .A(n8718), .B(n8717), .Z(n8793) );
  NANDN U8941 ( .A(n8720), .B(n8719), .Z(n8724) );
  NAND U8942 ( .A(n8722), .B(n8721), .Z(n8723) );
  AND U8943 ( .A(n8724), .B(n8723), .Z(n8859) );
  NANDN U8944 ( .A(n8726), .B(n8725), .Z(n8730) );
  NANDN U8945 ( .A(n8728), .B(n8727), .Z(n8729) );
  AND U8946 ( .A(n8730), .B(n8729), .Z(n8825) );
  NAND U8947 ( .A(b[0]), .B(a[121]), .Z(n8731) );
  XNOR U8948 ( .A(b[1]), .B(n8731), .Z(n8733) );
  NANDN U8949 ( .A(b[0]), .B(a[120]), .Z(n8732) );
  NAND U8950 ( .A(n8733), .B(n8732), .Z(n8805) );
  NANDN U8951 ( .A(n9891), .B(n8734), .Z(n8736) );
  XOR U8952 ( .A(b[13]), .B(a[109]), .Z(n8811) );
  NANDN U8953 ( .A(n9935), .B(n8811), .Z(n8735) );
  AND U8954 ( .A(n8736), .B(n8735), .Z(n8803) );
  AND U8955 ( .A(b[15]), .B(a[105]), .Z(n8802) );
  XNOR U8956 ( .A(n8803), .B(n8802), .Z(n8804) );
  XNOR U8957 ( .A(n8805), .B(n8804), .Z(n8823) );
  NANDN U8958 ( .A(n9437), .B(n8737), .Z(n8739) );
  XOR U8959 ( .A(b[5]), .B(a[117]), .Z(n8814) );
  NANDN U8960 ( .A(n9503), .B(n8814), .Z(n8738) );
  AND U8961 ( .A(n8739), .B(n8738), .Z(n8847) );
  NANDN U8962 ( .A(n9588), .B(n8740), .Z(n8742) );
  XOR U8963 ( .A(b[7]), .B(a[115]), .Z(n8817) );
  NANDN U8964 ( .A(n9639), .B(n8817), .Z(n8741) );
  AND U8965 ( .A(n8742), .B(n8741), .Z(n8845) );
  NANDN U8966 ( .A(n9374), .B(n8743), .Z(n8745) );
  XOR U8967 ( .A(a[119]), .B(b[3]), .Z(n8820) );
  NANDN U8968 ( .A(n9375), .B(n8820), .Z(n8744) );
  NAND U8969 ( .A(n8745), .B(n8744), .Z(n8844) );
  XNOR U8970 ( .A(n8845), .B(n8844), .Z(n8846) );
  XOR U8971 ( .A(n8847), .B(n8846), .Z(n8824) );
  XOR U8972 ( .A(n8823), .B(n8824), .Z(n8826) );
  XOR U8973 ( .A(n8825), .B(n8826), .Z(n8797) );
  NANDN U8974 ( .A(n8747), .B(n8746), .Z(n8751) );
  OR U8975 ( .A(n8749), .B(n8748), .Z(n8750) );
  AND U8976 ( .A(n8751), .B(n8750), .Z(n8796) );
  XNOR U8977 ( .A(n8797), .B(n8796), .Z(n8799) );
  NAND U8978 ( .A(n8752), .B(n9883), .Z(n8754) );
  XOR U8979 ( .A(b[11]), .B(a[111]), .Z(n8829) );
  NANDN U8980 ( .A(n9856), .B(n8829), .Z(n8753) );
  AND U8981 ( .A(n8754), .B(n8753), .Z(n8840) );
  NANDN U8982 ( .A(n10005), .B(n8755), .Z(n8757) );
  XOR U8983 ( .A(b[15]), .B(a[107]), .Z(n8832) );
  NANDN U8984 ( .A(n10006), .B(n8832), .Z(n8756) );
  AND U8985 ( .A(n8757), .B(n8756), .Z(n8839) );
  NANDN U8986 ( .A(n9685), .B(n8758), .Z(n8760) );
  XOR U8987 ( .A(b[9]), .B(a[113]), .Z(n8835) );
  NANDN U8988 ( .A(n9758), .B(n8835), .Z(n8759) );
  NAND U8989 ( .A(n8760), .B(n8759), .Z(n8838) );
  XOR U8990 ( .A(n8839), .B(n8838), .Z(n8841) );
  XOR U8991 ( .A(n8840), .B(n8841), .Z(n8851) );
  NANDN U8992 ( .A(n8762), .B(n8761), .Z(n8766) );
  OR U8993 ( .A(n8764), .B(n8763), .Z(n8765) );
  AND U8994 ( .A(n8766), .B(n8765), .Z(n8850) );
  XNOR U8995 ( .A(n8851), .B(n8850), .Z(n8852) );
  NANDN U8996 ( .A(n8768), .B(n8767), .Z(n8772) );
  NANDN U8997 ( .A(n8770), .B(n8769), .Z(n8771) );
  NAND U8998 ( .A(n8772), .B(n8771), .Z(n8853) );
  XNOR U8999 ( .A(n8852), .B(n8853), .Z(n8798) );
  XOR U9000 ( .A(n8799), .B(n8798), .Z(n8857) );
  NANDN U9001 ( .A(n8774), .B(n8773), .Z(n8778) );
  NANDN U9002 ( .A(n8776), .B(n8775), .Z(n8777) );
  AND U9003 ( .A(n8778), .B(n8777), .Z(n8856) );
  XNOR U9004 ( .A(n8857), .B(n8856), .Z(n8858) );
  XOR U9005 ( .A(n8859), .B(n8858), .Z(n8791) );
  NANDN U9006 ( .A(n8780), .B(n8779), .Z(n8784) );
  NAND U9007 ( .A(n8782), .B(n8781), .Z(n8783) );
  AND U9008 ( .A(n8784), .B(n8783), .Z(n8790) );
  XNOR U9009 ( .A(n8791), .B(n8790), .Z(n8792) );
  XNOR U9010 ( .A(n8793), .B(n8792), .Z(n8862) );
  XNOR U9011 ( .A(sreg[233]), .B(n8862), .Z(n8864) );
  NANDN U9012 ( .A(sreg[232]), .B(n8785), .Z(n8789) );
  NAND U9013 ( .A(n8787), .B(n8786), .Z(n8788) );
  NAND U9014 ( .A(n8789), .B(n8788), .Z(n8863) );
  XNOR U9015 ( .A(n8864), .B(n8863), .Z(c[233]) );
  NANDN U9016 ( .A(n8791), .B(n8790), .Z(n8795) );
  NANDN U9017 ( .A(n8793), .B(n8792), .Z(n8794) );
  AND U9018 ( .A(n8795), .B(n8794), .Z(n8870) );
  NANDN U9019 ( .A(n8797), .B(n8796), .Z(n8801) );
  NAND U9020 ( .A(n8799), .B(n8798), .Z(n8800) );
  AND U9021 ( .A(n8801), .B(n8800), .Z(n8936) );
  NANDN U9022 ( .A(n8803), .B(n8802), .Z(n8807) );
  NANDN U9023 ( .A(n8805), .B(n8804), .Z(n8806) );
  AND U9024 ( .A(n8807), .B(n8806), .Z(n8923) );
  NAND U9025 ( .A(b[0]), .B(a[122]), .Z(n8808) );
  XNOR U9026 ( .A(b[1]), .B(n8808), .Z(n8810) );
  NANDN U9027 ( .A(b[0]), .B(a[121]), .Z(n8809) );
  NAND U9028 ( .A(n8810), .B(n8809), .Z(n8903) );
  NANDN U9029 ( .A(n9891), .B(n8811), .Z(n8813) );
  XOR U9030 ( .A(b[13]), .B(a[110]), .Z(n8909) );
  NANDN U9031 ( .A(n9935), .B(n8909), .Z(n8812) );
  AND U9032 ( .A(n8813), .B(n8812), .Z(n8901) );
  AND U9033 ( .A(b[15]), .B(a[106]), .Z(n8900) );
  XNOR U9034 ( .A(n8901), .B(n8900), .Z(n8902) );
  XNOR U9035 ( .A(n8903), .B(n8902), .Z(n8921) );
  NANDN U9036 ( .A(n9437), .B(n8814), .Z(n8816) );
  XOR U9037 ( .A(b[5]), .B(a[118]), .Z(n8912) );
  NANDN U9038 ( .A(n9503), .B(n8912), .Z(n8815) );
  AND U9039 ( .A(n8816), .B(n8815), .Z(n8897) );
  NANDN U9040 ( .A(n9588), .B(n8817), .Z(n8819) );
  XOR U9041 ( .A(b[7]), .B(a[116]), .Z(n8915) );
  NANDN U9042 ( .A(n9639), .B(n8915), .Z(n8818) );
  AND U9043 ( .A(n8819), .B(n8818), .Z(n8895) );
  NANDN U9044 ( .A(n9374), .B(n8820), .Z(n8822) );
  XOR U9045 ( .A(a[120]), .B(b[3]), .Z(n8918) );
  NANDN U9046 ( .A(n9375), .B(n8918), .Z(n8821) );
  NAND U9047 ( .A(n8822), .B(n8821), .Z(n8894) );
  XNOR U9048 ( .A(n8895), .B(n8894), .Z(n8896) );
  XOR U9049 ( .A(n8897), .B(n8896), .Z(n8922) );
  XOR U9050 ( .A(n8921), .B(n8922), .Z(n8924) );
  XOR U9051 ( .A(n8923), .B(n8924), .Z(n8874) );
  NANDN U9052 ( .A(n8824), .B(n8823), .Z(n8828) );
  OR U9053 ( .A(n8826), .B(n8825), .Z(n8827) );
  AND U9054 ( .A(n8828), .B(n8827), .Z(n8873) );
  XNOR U9055 ( .A(n8874), .B(n8873), .Z(n8876) );
  NAND U9056 ( .A(n8829), .B(n9883), .Z(n8831) );
  XOR U9057 ( .A(b[11]), .B(a[112]), .Z(n8879) );
  NANDN U9058 ( .A(n9856), .B(n8879), .Z(n8830) );
  AND U9059 ( .A(n8831), .B(n8830), .Z(n8890) );
  NANDN U9060 ( .A(n10005), .B(n8832), .Z(n8834) );
  XOR U9061 ( .A(b[15]), .B(a[108]), .Z(n8882) );
  NANDN U9062 ( .A(n10006), .B(n8882), .Z(n8833) );
  AND U9063 ( .A(n8834), .B(n8833), .Z(n8889) );
  NANDN U9064 ( .A(n9685), .B(n8835), .Z(n8837) );
  XOR U9065 ( .A(b[9]), .B(a[114]), .Z(n8885) );
  NANDN U9066 ( .A(n9758), .B(n8885), .Z(n8836) );
  NAND U9067 ( .A(n8837), .B(n8836), .Z(n8888) );
  XOR U9068 ( .A(n8889), .B(n8888), .Z(n8891) );
  XOR U9069 ( .A(n8890), .B(n8891), .Z(n8928) );
  NANDN U9070 ( .A(n8839), .B(n8838), .Z(n8843) );
  OR U9071 ( .A(n8841), .B(n8840), .Z(n8842) );
  AND U9072 ( .A(n8843), .B(n8842), .Z(n8927) );
  XNOR U9073 ( .A(n8928), .B(n8927), .Z(n8929) );
  NANDN U9074 ( .A(n8845), .B(n8844), .Z(n8849) );
  NANDN U9075 ( .A(n8847), .B(n8846), .Z(n8848) );
  NAND U9076 ( .A(n8849), .B(n8848), .Z(n8930) );
  XNOR U9077 ( .A(n8929), .B(n8930), .Z(n8875) );
  XOR U9078 ( .A(n8876), .B(n8875), .Z(n8934) );
  NANDN U9079 ( .A(n8851), .B(n8850), .Z(n8855) );
  NANDN U9080 ( .A(n8853), .B(n8852), .Z(n8854) );
  AND U9081 ( .A(n8855), .B(n8854), .Z(n8933) );
  XNOR U9082 ( .A(n8934), .B(n8933), .Z(n8935) );
  XOR U9083 ( .A(n8936), .B(n8935), .Z(n8868) );
  NANDN U9084 ( .A(n8857), .B(n8856), .Z(n8861) );
  NAND U9085 ( .A(n8859), .B(n8858), .Z(n8860) );
  AND U9086 ( .A(n8861), .B(n8860), .Z(n8867) );
  XNOR U9087 ( .A(n8868), .B(n8867), .Z(n8869) );
  XNOR U9088 ( .A(n8870), .B(n8869), .Z(n8939) );
  XNOR U9089 ( .A(sreg[234]), .B(n8939), .Z(n8941) );
  NANDN U9090 ( .A(sreg[233]), .B(n8862), .Z(n8866) );
  NAND U9091 ( .A(n8864), .B(n8863), .Z(n8865) );
  NAND U9092 ( .A(n8866), .B(n8865), .Z(n8940) );
  XNOR U9093 ( .A(n8941), .B(n8940), .Z(c[234]) );
  NANDN U9094 ( .A(n8868), .B(n8867), .Z(n8872) );
  NANDN U9095 ( .A(n8870), .B(n8869), .Z(n8871) );
  AND U9096 ( .A(n8872), .B(n8871), .Z(n8947) );
  NANDN U9097 ( .A(n8874), .B(n8873), .Z(n8878) );
  NAND U9098 ( .A(n8876), .B(n8875), .Z(n8877) );
  AND U9099 ( .A(n8878), .B(n8877), .Z(n9013) );
  NAND U9100 ( .A(n8879), .B(n9883), .Z(n8881) );
  XOR U9101 ( .A(b[11]), .B(a[113]), .Z(n8956) );
  NANDN U9102 ( .A(n9856), .B(n8956), .Z(n8880) );
  AND U9103 ( .A(n8881), .B(n8880), .Z(n8967) );
  NANDN U9104 ( .A(n10005), .B(n8882), .Z(n8884) );
  XOR U9105 ( .A(b[15]), .B(a[109]), .Z(n8959) );
  NANDN U9106 ( .A(n10006), .B(n8959), .Z(n8883) );
  AND U9107 ( .A(n8884), .B(n8883), .Z(n8966) );
  NANDN U9108 ( .A(n9685), .B(n8885), .Z(n8887) );
  XOR U9109 ( .A(b[9]), .B(a[115]), .Z(n8962) );
  NANDN U9110 ( .A(n9758), .B(n8962), .Z(n8886) );
  NAND U9111 ( .A(n8887), .B(n8886), .Z(n8965) );
  XOR U9112 ( .A(n8966), .B(n8965), .Z(n8968) );
  XOR U9113 ( .A(n8967), .B(n8968), .Z(n9005) );
  NANDN U9114 ( .A(n8889), .B(n8888), .Z(n8893) );
  OR U9115 ( .A(n8891), .B(n8890), .Z(n8892) );
  AND U9116 ( .A(n8893), .B(n8892), .Z(n9004) );
  XNOR U9117 ( .A(n9005), .B(n9004), .Z(n9006) );
  NANDN U9118 ( .A(n8895), .B(n8894), .Z(n8899) );
  NANDN U9119 ( .A(n8897), .B(n8896), .Z(n8898) );
  NAND U9120 ( .A(n8899), .B(n8898), .Z(n9007) );
  XNOR U9121 ( .A(n9006), .B(n9007), .Z(n8953) );
  NANDN U9122 ( .A(n8901), .B(n8900), .Z(n8905) );
  NANDN U9123 ( .A(n8903), .B(n8902), .Z(n8904) );
  AND U9124 ( .A(n8905), .B(n8904), .Z(n9000) );
  NAND U9125 ( .A(b[0]), .B(a[123]), .Z(n8906) );
  XNOR U9126 ( .A(b[1]), .B(n8906), .Z(n8908) );
  NANDN U9127 ( .A(b[0]), .B(a[122]), .Z(n8907) );
  NAND U9128 ( .A(n8908), .B(n8907), .Z(n8980) );
  NANDN U9129 ( .A(n9891), .B(n8909), .Z(n8911) );
  XOR U9130 ( .A(b[13]), .B(a[111]), .Z(n8986) );
  NANDN U9131 ( .A(n9935), .B(n8986), .Z(n8910) );
  AND U9132 ( .A(n8911), .B(n8910), .Z(n8978) );
  AND U9133 ( .A(b[15]), .B(a[107]), .Z(n8977) );
  XNOR U9134 ( .A(n8978), .B(n8977), .Z(n8979) );
  XNOR U9135 ( .A(n8980), .B(n8979), .Z(n8998) );
  NANDN U9136 ( .A(n9437), .B(n8912), .Z(n8914) );
  XOR U9137 ( .A(b[5]), .B(a[119]), .Z(n8989) );
  NANDN U9138 ( .A(n9503), .B(n8989), .Z(n8913) );
  AND U9139 ( .A(n8914), .B(n8913), .Z(n8974) );
  NANDN U9140 ( .A(n9588), .B(n8915), .Z(n8917) );
  XOR U9141 ( .A(b[7]), .B(a[117]), .Z(n8992) );
  NANDN U9142 ( .A(n9639), .B(n8992), .Z(n8916) );
  AND U9143 ( .A(n8917), .B(n8916), .Z(n8972) );
  NANDN U9144 ( .A(n9374), .B(n8918), .Z(n8920) );
  XOR U9145 ( .A(a[121]), .B(b[3]), .Z(n8995) );
  NANDN U9146 ( .A(n9375), .B(n8995), .Z(n8919) );
  NAND U9147 ( .A(n8920), .B(n8919), .Z(n8971) );
  XNOR U9148 ( .A(n8972), .B(n8971), .Z(n8973) );
  XOR U9149 ( .A(n8974), .B(n8973), .Z(n8999) );
  XOR U9150 ( .A(n8998), .B(n8999), .Z(n9001) );
  XOR U9151 ( .A(n9000), .B(n9001), .Z(n8951) );
  NANDN U9152 ( .A(n8922), .B(n8921), .Z(n8926) );
  OR U9153 ( .A(n8924), .B(n8923), .Z(n8925) );
  AND U9154 ( .A(n8926), .B(n8925), .Z(n8950) );
  XNOR U9155 ( .A(n8951), .B(n8950), .Z(n8952) );
  XOR U9156 ( .A(n8953), .B(n8952), .Z(n9011) );
  NANDN U9157 ( .A(n8928), .B(n8927), .Z(n8932) );
  NANDN U9158 ( .A(n8930), .B(n8929), .Z(n8931) );
  AND U9159 ( .A(n8932), .B(n8931), .Z(n9010) );
  XNOR U9160 ( .A(n9011), .B(n9010), .Z(n9012) );
  XOR U9161 ( .A(n9013), .B(n9012), .Z(n8945) );
  NANDN U9162 ( .A(n8934), .B(n8933), .Z(n8938) );
  NAND U9163 ( .A(n8936), .B(n8935), .Z(n8937) );
  AND U9164 ( .A(n8938), .B(n8937), .Z(n8944) );
  XNOR U9165 ( .A(n8945), .B(n8944), .Z(n8946) );
  XNOR U9166 ( .A(n8947), .B(n8946), .Z(n9016) );
  XNOR U9167 ( .A(sreg[235]), .B(n9016), .Z(n9018) );
  NANDN U9168 ( .A(sreg[234]), .B(n8939), .Z(n8943) );
  NAND U9169 ( .A(n8941), .B(n8940), .Z(n8942) );
  NAND U9170 ( .A(n8943), .B(n8942), .Z(n9017) );
  XNOR U9171 ( .A(n9018), .B(n9017), .Z(c[235]) );
  NANDN U9172 ( .A(n8945), .B(n8944), .Z(n8949) );
  NANDN U9173 ( .A(n8947), .B(n8946), .Z(n8948) );
  AND U9174 ( .A(n8949), .B(n8948), .Z(n9024) );
  NANDN U9175 ( .A(n8951), .B(n8950), .Z(n8955) );
  NAND U9176 ( .A(n8953), .B(n8952), .Z(n8954) );
  AND U9177 ( .A(n8955), .B(n8954), .Z(n9090) );
  NAND U9178 ( .A(n8956), .B(n9883), .Z(n8958) );
  XOR U9179 ( .A(b[11]), .B(a[114]), .Z(n9060) );
  NANDN U9180 ( .A(n9856), .B(n9060), .Z(n8957) );
  AND U9181 ( .A(n8958), .B(n8957), .Z(n9071) );
  NANDN U9182 ( .A(n10005), .B(n8959), .Z(n8961) );
  XOR U9183 ( .A(b[15]), .B(a[110]), .Z(n9063) );
  NANDN U9184 ( .A(n10006), .B(n9063), .Z(n8960) );
  AND U9185 ( .A(n8961), .B(n8960), .Z(n9070) );
  NANDN U9186 ( .A(n9685), .B(n8962), .Z(n8964) );
  XOR U9187 ( .A(b[9]), .B(a[116]), .Z(n9066) );
  NANDN U9188 ( .A(n9758), .B(n9066), .Z(n8963) );
  NAND U9189 ( .A(n8964), .B(n8963), .Z(n9069) );
  XOR U9190 ( .A(n9070), .B(n9069), .Z(n9072) );
  XOR U9191 ( .A(n9071), .B(n9072), .Z(n9082) );
  NANDN U9192 ( .A(n8966), .B(n8965), .Z(n8970) );
  OR U9193 ( .A(n8968), .B(n8967), .Z(n8969) );
  AND U9194 ( .A(n8970), .B(n8969), .Z(n9081) );
  XNOR U9195 ( .A(n9082), .B(n9081), .Z(n9083) );
  NANDN U9196 ( .A(n8972), .B(n8971), .Z(n8976) );
  NANDN U9197 ( .A(n8974), .B(n8973), .Z(n8975) );
  NAND U9198 ( .A(n8976), .B(n8975), .Z(n9084) );
  XNOR U9199 ( .A(n9083), .B(n9084), .Z(n9030) );
  NANDN U9200 ( .A(n8978), .B(n8977), .Z(n8982) );
  NANDN U9201 ( .A(n8980), .B(n8979), .Z(n8981) );
  AND U9202 ( .A(n8982), .B(n8981), .Z(n9056) );
  NAND U9203 ( .A(b[0]), .B(a[124]), .Z(n8983) );
  XNOR U9204 ( .A(b[1]), .B(n8983), .Z(n8985) );
  NANDN U9205 ( .A(b[0]), .B(a[123]), .Z(n8984) );
  NAND U9206 ( .A(n8985), .B(n8984), .Z(n9036) );
  NANDN U9207 ( .A(n9891), .B(n8986), .Z(n8988) );
  XOR U9208 ( .A(b[13]), .B(a[112]), .Z(n9042) );
  NANDN U9209 ( .A(n9935), .B(n9042), .Z(n8987) );
  AND U9210 ( .A(n8988), .B(n8987), .Z(n9034) );
  AND U9211 ( .A(b[15]), .B(a[108]), .Z(n9033) );
  XNOR U9212 ( .A(n9034), .B(n9033), .Z(n9035) );
  XNOR U9213 ( .A(n9036), .B(n9035), .Z(n9054) );
  NANDN U9214 ( .A(n9437), .B(n8989), .Z(n8991) );
  XOR U9215 ( .A(a[120]), .B(b[5]), .Z(n9045) );
  NANDN U9216 ( .A(n9503), .B(n9045), .Z(n8990) );
  AND U9217 ( .A(n8991), .B(n8990), .Z(n9078) );
  NANDN U9218 ( .A(n9588), .B(n8992), .Z(n8994) );
  XOR U9219 ( .A(b[7]), .B(a[118]), .Z(n9048) );
  NANDN U9220 ( .A(n9639), .B(n9048), .Z(n8993) );
  AND U9221 ( .A(n8994), .B(n8993), .Z(n9076) );
  NANDN U9222 ( .A(n9374), .B(n8995), .Z(n8997) );
  XOR U9223 ( .A(a[122]), .B(b[3]), .Z(n9051) );
  NANDN U9224 ( .A(n9375), .B(n9051), .Z(n8996) );
  NAND U9225 ( .A(n8997), .B(n8996), .Z(n9075) );
  XNOR U9226 ( .A(n9076), .B(n9075), .Z(n9077) );
  XOR U9227 ( .A(n9078), .B(n9077), .Z(n9055) );
  XOR U9228 ( .A(n9054), .B(n9055), .Z(n9057) );
  XOR U9229 ( .A(n9056), .B(n9057), .Z(n9028) );
  NANDN U9230 ( .A(n8999), .B(n8998), .Z(n9003) );
  OR U9231 ( .A(n9001), .B(n9000), .Z(n9002) );
  AND U9232 ( .A(n9003), .B(n9002), .Z(n9027) );
  XNOR U9233 ( .A(n9028), .B(n9027), .Z(n9029) );
  XOR U9234 ( .A(n9030), .B(n9029), .Z(n9088) );
  NANDN U9235 ( .A(n9005), .B(n9004), .Z(n9009) );
  NANDN U9236 ( .A(n9007), .B(n9006), .Z(n9008) );
  AND U9237 ( .A(n9009), .B(n9008), .Z(n9087) );
  XNOR U9238 ( .A(n9088), .B(n9087), .Z(n9089) );
  XOR U9239 ( .A(n9090), .B(n9089), .Z(n9022) );
  NANDN U9240 ( .A(n9011), .B(n9010), .Z(n9015) );
  NAND U9241 ( .A(n9013), .B(n9012), .Z(n9014) );
  AND U9242 ( .A(n9015), .B(n9014), .Z(n9021) );
  XNOR U9243 ( .A(n9022), .B(n9021), .Z(n9023) );
  XNOR U9244 ( .A(n9024), .B(n9023), .Z(n9093) );
  XNOR U9245 ( .A(sreg[236]), .B(n9093), .Z(n9095) );
  NANDN U9246 ( .A(sreg[235]), .B(n9016), .Z(n9020) );
  NAND U9247 ( .A(n9018), .B(n9017), .Z(n9019) );
  NAND U9248 ( .A(n9020), .B(n9019), .Z(n9094) );
  XNOR U9249 ( .A(n9095), .B(n9094), .Z(c[236]) );
  NANDN U9250 ( .A(n9022), .B(n9021), .Z(n9026) );
  NANDN U9251 ( .A(n9024), .B(n9023), .Z(n9025) );
  AND U9252 ( .A(n9026), .B(n9025), .Z(n9101) );
  NANDN U9253 ( .A(n9028), .B(n9027), .Z(n9032) );
  NAND U9254 ( .A(n9030), .B(n9029), .Z(n9031) );
  AND U9255 ( .A(n9032), .B(n9031), .Z(n9167) );
  NANDN U9256 ( .A(n9034), .B(n9033), .Z(n9038) );
  NANDN U9257 ( .A(n9036), .B(n9035), .Z(n9037) );
  AND U9258 ( .A(n9038), .B(n9037), .Z(n9133) );
  NAND U9259 ( .A(b[0]), .B(a[125]), .Z(n9039) );
  XNOR U9260 ( .A(b[1]), .B(n9039), .Z(n9041) );
  NANDN U9261 ( .A(b[0]), .B(a[124]), .Z(n9040) );
  NAND U9262 ( .A(n9041), .B(n9040), .Z(n9113) );
  NANDN U9263 ( .A(n9891), .B(n9042), .Z(n9044) );
  XOR U9264 ( .A(b[13]), .B(a[113]), .Z(n9116) );
  NANDN U9265 ( .A(n9935), .B(n9116), .Z(n9043) );
  AND U9266 ( .A(n9044), .B(n9043), .Z(n9111) );
  AND U9267 ( .A(b[15]), .B(a[109]), .Z(n9110) );
  XNOR U9268 ( .A(n9111), .B(n9110), .Z(n9112) );
  XNOR U9269 ( .A(n9113), .B(n9112), .Z(n9131) );
  NANDN U9270 ( .A(n9437), .B(n9045), .Z(n9047) );
  XOR U9271 ( .A(a[121]), .B(b[5]), .Z(n9122) );
  NANDN U9272 ( .A(n9503), .B(n9122), .Z(n9046) );
  AND U9273 ( .A(n9047), .B(n9046), .Z(n9155) );
  NANDN U9274 ( .A(n9588), .B(n9048), .Z(n9050) );
  XOR U9275 ( .A(b[7]), .B(a[119]), .Z(n9125) );
  NANDN U9276 ( .A(n9639), .B(n9125), .Z(n9049) );
  AND U9277 ( .A(n9050), .B(n9049), .Z(n9153) );
  NANDN U9278 ( .A(n9374), .B(n9051), .Z(n9053) );
  XOR U9279 ( .A(a[123]), .B(b[3]), .Z(n9128) );
  NANDN U9280 ( .A(n9375), .B(n9128), .Z(n9052) );
  NAND U9281 ( .A(n9053), .B(n9052), .Z(n9152) );
  XNOR U9282 ( .A(n9153), .B(n9152), .Z(n9154) );
  XOR U9283 ( .A(n9155), .B(n9154), .Z(n9132) );
  XOR U9284 ( .A(n9131), .B(n9132), .Z(n9134) );
  XOR U9285 ( .A(n9133), .B(n9134), .Z(n9105) );
  NANDN U9286 ( .A(n9055), .B(n9054), .Z(n9059) );
  OR U9287 ( .A(n9057), .B(n9056), .Z(n9058) );
  AND U9288 ( .A(n9059), .B(n9058), .Z(n9104) );
  XNOR U9289 ( .A(n9105), .B(n9104), .Z(n9107) );
  NAND U9290 ( .A(n9060), .B(n9883), .Z(n9062) );
  XOR U9291 ( .A(b[11]), .B(a[115]), .Z(n9137) );
  NANDN U9292 ( .A(n9856), .B(n9137), .Z(n9061) );
  AND U9293 ( .A(n9062), .B(n9061), .Z(n9148) );
  NANDN U9294 ( .A(n10005), .B(n9063), .Z(n9065) );
  XOR U9295 ( .A(b[15]), .B(a[111]), .Z(n9140) );
  NANDN U9296 ( .A(n10006), .B(n9140), .Z(n9064) );
  AND U9297 ( .A(n9065), .B(n9064), .Z(n9147) );
  NANDN U9298 ( .A(n9685), .B(n9066), .Z(n9068) );
  XOR U9299 ( .A(b[9]), .B(a[117]), .Z(n9143) );
  NANDN U9300 ( .A(n9758), .B(n9143), .Z(n9067) );
  NAND U9301 ( .A(n9068), .B(n9067), .Z(n9146) );
  XOR U9302 ( .A(n9147), .B(n9146), .Z(n9149) );
  XOR U9303 ( .A(n9148), .B(n9149), .Z(n9159) );
  NANDN U9304 ( .A(n9070), .B(n9069), .Z(n9074) );
  OR U9305 ( .A(n9072), .B(n9071), .Z(n9073) );
  AND U9306 ( .A(n9074), .B(n9073), .Z(n9158) );
  XNOR U9307 ( .A(n9159), .B(n9158), .Z(n9160) );
  NANDN U9308 ( .A(n9076), .B(n9075), .Z(n9080) );
  NANDN U9309 ( .A(n9078), .B(n9077), .Z(n9079) );
  NAND U9310 ( .A(n9080), .B(n9079), .Z(n9161) );
  XNOR U9311 ( .A(n9160), .B(n9161), .Z(n9106) );
  XOR U9312 ( .A(n9107), .B(n9106), .Z(n9165) );
  NANDN U9313 ( .A(n9082), .B(n9081), .Z(n9086) );
  NANDN U9314 ( .A(n9084), .B(n9083), .Z(n9085) );
  AND U9315 ( .A(n9086), .B(n9085), .Z(n9164) );
  XNOR U9316 ( .A(n9165), .B(n9164), .Z(n9166) );
  XOR U9317 ( .A(n9167), .B(n9166), .Z(n9099) );
  NANDN U9318 ( .A(n9088), .B(n9087), .Z(n9092) );
  NAND U9319 ( .A(n9090), .B(n9089), .Z(n9091) );
  AND U9320 ( .A(n9092), .B(n9091), .Z(n9098) );
  XNOR U9321 ( .A(n9099), .B(n9098), .Z(n9100) );
  XNOR U9322 ( .A(n9101), .B(n9100), .Z(n9170) );
  XNOR U9323 ( .A(sreg[237]), .B(n9170), .Z(n9172) );
  NANDN U9324 ( .A(sreg[236]), .B(n9093), .Z(n9097) );
  NAND U9325 ( .A(n9095), .B(n9094), .Z(n9096) );
  NAND U9326 ( .A(n9097), .B(n9096), .Z(n9171) );
  XNOR U9327 ( .A(n9172), .B(n9171), .Z(c[237]) );
  NANDN U9328 ( .A(n9099), .B(n9098), .Z(n9103) );
  NANDN U9329 ( .A(n9101), .B(n9100), .Z(n9102) );
  AND U9330 ( .A(n9103), .B(n9102), .Z(n9178) );
  NANDN U9331 ( .A(n9105), .B(n9104), .Z(n9109) );
  NAND U9332 ( .A(n9107), .B(n9106), .Z(n9108) );
  AND U9333 ( .A(n9109), .B(n9108), .Z(n9244) );
  NANDN U9334 ( .A(n9111), .B(n9110), .Z(n9115) );
  NANDN U9335 ( .A(n9113), .B(n9112), .Z(n9114) );
  AND U9336 ( .A(n9115), .B(n9114), .Z(n9210) );
  NANDN U9337 ( .A(n9891), .B(n9116), .Z(n9118) );
  XOR U9338 ( .A(b[13]), .B(a[114]), .Z(n9196) );
  NANDN U9339 ( .A(n9935), .B(n9196), .Z(n9117) );
  AND U9340 ( .A(n9118), .B(n9117), .Z(n9188) );
  AND U9341 ( .A(b[15]), .B(a[110]), .Z(n9187) );
  XNOR U9342 ( .A(n9188), .B(n9187), .Z(n9189) );
  NAND U9343 ( .A(b[0]), .B(a[126]), .Z(n9119) );
  XNOR U9344 ( .A(b[1]), .B(n9119), .Z(n9121) );
  NANDN U9345 ( .A(b[0]), .B(a[125]), .Z(n9120) );
  NAND U9346 ( .A(n9121), .B(n9120), .Z(n9190) );
  XNOR U9347 ( .A(n9189), .B(n9190), .Z(n9208) );
  NANDN U9348 ( .A(n9437), .B(n9122), .Z(n9124) );
  XOR U9349 ( .A(a[122]), .B(b[5]), .Z(n9199) );
  NANDN U9350 ( .A(n9503), .B(n9199), .Z(n9123) );
  AND U9351 ( .A(n9124), .B(n9123), .Z(n9232) );
  NANDN U9352 ( .A(n9588), .B(n9125), .Z(n9127) );
  XOR U9353 ( .A(b[7]), .B(a[120]), .Z(n9202) );
  NANDN U9354 ( .A(n9639), .B(n9202), .Z(n9126) );
  AND U9355 ( .A(n9127), .B(n9126), .Z(n9230) );
  NANDN U9356 ( .A(n9374), .B(n9128), .Z(n9130) );
  XOR U9357 ( .A(a[124]), .B(b[3]), .Z(n9205) );
  NANDN U9358 ( .A(n9375), .B(n9205), .Z(n9129) );
  NAND U9359 ( .A(n9130), .B(n9129), .Z(n9229) );
  XNOR U9360 ( .A(n9230), .B(n9229), .Z(n9231) );
  XOR U9361 ( .A(n9232), .B(n9231), .Z(n9209) );
  XOR U9362 ( .A(n9208), .B(n9209), .Z(n9211) );
  XOR U9363 ( .A(n9210), .B(n9211), .Z(n9182) );
  NANDN U9364 ( .A(n9132), .B(n9131), .Z(n9136) );
  OR U9365 ( .A(n9134), .B(n9133), .Z(n9135) );
  AND U9366 ( .A(n9136), .B(n9135), .Z(n9181) );
  XNOR U9367 ( .A(n9182), .B(n9181), .Z(n9184) );
  NAND U9368 ( .A(n9137), .B(n9883), .Z(n9139) );
  XOR U9369 ( .A(b[11]), .B(a[116]), .Z(n9214) );
  NANDN U9370 ( .A(n9856), .B(n9214), .Z(n9138) );
  AND U9371 ( .A(n9139), .B(n9138), .Z(n9225) );
  NANDN U9372 ( .A(n10005), .B(n9140), .Z(n9142) );
  XOR U9373 ( .A(b[15]), .B(a[112]), .Z(n9217) );
  NANDN U9374 ( .A(n10006), .B(n9217), .Z(n9141) );
  AND U9375 ( .A(n9142), .B(n9141), .Z(n9224) );
  NANDN U9376 ( .A(n9685), .B(n9143), .Z(n9145) );
  XOR U9377 ( .A(b[9]), .B(a[118]), .Z(n9220) );
  NANDN U9378 ( .A(n9758), .B(n9220), .Z(n9144) );
  NAND U9379 ( .A(n9145), .B(n9144), .Z(n9223) );
  XOR U9380 ( .A(n9224), .B(n9223), .Z(n9226) );
  XOR U9381 ( .A(n9225), .B(n9226), .Z(n9236) );
  NANDN U9382 ( .A(n9147), .B(n9146), .Z(n9151) );
  OR U9383 ( .A(n9149), .B(n9148), .Z(n9150) );
  AND U9384 ( .A(n9151), .B(n9150), .Z(n9235) );
  XNOR U9385 ( .A(n9236), .B(n9235), .Z(n9237) );
  NANDN U9386 ( .A(n9153), .B(n9152), .Z(n9157) );
  NANDN U9387 ( .A(n9155), .B(n9154), .Z(n9156) );
  NAND U9388 ( .A(n9157), .B(n9156), .Z(n9238) );
  XNOR U9389 ( .A(n9237), .B(n9238), .Z(n9183) );
  XOR U9390 ( .A(n9184), .B(n9183), .Z(n9242) );
  NANDN U9391 ( .A(n9159), .B(n9158), .Z(n9163) );
  NANDN U9392 ( .A(n9161), .B(n9160), .Z(n9162) );
  AND U9393 ( .A(n9163), .B(n9162), .Z(n9241) );
  XNOR U9394 ( .A(n9242), .B(n9241), .Z(n9243) );
  XOR U9395 ( .A(n9244), .B(n9243), .Z(n9176) );
  NANDN U9396 ( .A(n9165), .B(n9164), .Z(n9169) );
  NAND U9397 ( .A(n9167), .B(n9166), .Z(n9168) );
  AND U9398 ( .A(n9169), .B(n9168), .Z(n9175) );
  XNOR U9399 ( .A(n9176), .B(n9175), .Z(n9177) );
  XNOR U9400 ( .A(n9178), .B(n9177), .Z(n9247) );
  XNOR U9401 ( .A(sreg[238]), .B(n9247), .Z(n9249) );
  NANDN U9402 ( .A(sreg[237]), .B(n9170), .Z(n9174) );
  NAND U9403 ( .A(n9172), .B(n9171), .Z(n9173) );
  NAND U9404 ( .A(n9174), .B(n9173), .Z(n9248) );
  XNOR U9405 ( .A(n9249), .B(n9248), .Z(c[238]) );
  NANDN U9406 ( .A(n9176), .B(n9175), .Z(n9180) );
  NANDN U9407 ( .A(n9178), .B(n9177), .Z(n9179) );
  AND U9408 ( .A(n9180), .B(n9179), .Z(n9260) );
  NANDN U9409 ( .A(n9182), .B(n9181), .Z(n9186) );
  NAND U9410 ( .A(n9184), .B(n9183), .Z(n9185) );
  AND U9411 ( .A(n9186), .B(n9185), .Z(n9323) );
  NANDN U9412 ( .A(n9188), .B(n9187), .Z(n9192) );
  NANDN U9413 ( .A(n9190), .B(n9189), .Z(n9191) );
  AND U9414 ( .A(n9192), .B(n9191), .Z(n9310) );
  NAND U9415 ( .A(b[0]), .B(a[127]), .Z(n9193) );
  XNOR U9416 ( .A(b[1]), .B(n9193), .Z(n9195) );
  NANDN U9417 ( .A(b[0]), .B(a[126]), .Z(n9194) );
  NAND U9418 ( .A(n9195), .B(n9194), .Z(n9293) );
  NANDN U9419 ( .A(n9891), .B(n9196), .Z(n9198) );
  XOR U9420 ( .A(b[13]), .B(a[115]), .Z(n9296) );
  NANDN U9421 ( .A(n9935), .B(n9296), .Z(n9197) );
  AND U9422 ( .A(n9198), .B(n9197), .Z(n9291) );
  AND U9423 ( .A(b[15]), .B(a[111]), .Z(n9290) );
  XNOR U9424 ( .A(n9291), .B(n9290), .Z(n9292) );
  XNOR U9425 ( .A(n9293), .B(n9292), .Z(n9308) );
  NANDN U9426 ( .A(n9437), .B(n9199), .Z(n9201) );
  XOR U9427 ( .A(a[123]), .B(b[5]), .Z(n9299) );
  NANDN U9428 ( .A(n9503), .B(n9299), .Z(n9200) );
  AND U9429 ( .A(n9201), .B(n9200), .Z(n9287) );
  NANDN U9430 ( .A(n9588), .B(n9202), .Z(n9204) );
  XOR U9431 ( .A(b[7]), .B(a[121]), .Z(n9302) );
  NANDN U9432 ( .A(n9639), .B(n9302), .Z(n9203) );
  AND U9433 ( .A(n9204), .B(n9203), .Z(n9285) );
  NANDN U9434 ( .A(n9374), .B(n9205), .Z(n9207) );
  XOR U9435 ( .A(a[125]), .B(b[3]), .Z(n9305) );
  NANDN U9436 ( .A(n9375), .B(n9305), .Z(n9206) );
  NAND U9437 ( .A(n9207), .B(n9206), .Z(n9284) );
  XNOR U9438 ( .A(n9285), .B(n9284), .Z(n9286) );
  XOR U9439 ( .A(n9287), .B(n9286), .Z(n9309) );
  XOR U9440 ( .A(n9308), .B(n9309), .Z(n9311) );
  XOR U9441 ( .A(n9310), .B(n9311), .Z(n9264) );
  NANDN U9442 ( .A(n9209), .B(n9208), .Z(n9213) );
  OR U9443 ( .A(n9211), .B(n9210), .Z(n9212) );
  AND U9444 ( .A(n9213), .B(n9212), .Z(n9263) );
  XNOR U9445 ( .A(n9264), .B(n9263), .Z(n9266) );
  NAND U9446 ( .A(n9214), .B(n9883), .Z(n9216) );
  XOR U9447 ( .A(b[11]), .B(a[117]), .Z(n9269) );
  NANDN U9448 ( .A(n9856), .B(n9269), .Z(n9215) );
  AND U9449 ( .A(n9216), .B(n9215), .Z(n9280) );
  NANDN U9450 ( .A(n10005), .B(n9217), .Z(n9219) );
  XOR U9451 ( .A(b[15]), .B(a[113]), .Z(n9272) );
  NANDN U9452 ( .A(n10006), .B(n9272), .Z(n9218) );
  AND U9453 ( .A(n9219), .B(n9218), .Z(n9279) );
  NANDN U9454 ( .A(n9685), .B(n9220), .Z(n9222) );
  XOR U9455 ( .A(b[9]), .B(a[119]), .Z(n9275) );
  NANDN U9456 ( .A(n9758), .B(n9275), .Z(n9221) );
  NAND U9457 ( .A(n9222), .B(n9221), .Z(n9278) );
  XOR U9458 ( .A(n9279), .B(n9278), .Z(n9281) );
  XOR U9459 ( .A(n9280), .B(n9281), .Z(n9315) );
  NANDN U9460 ( .A(n9224), .B(n9223), .Z(n9228) );
  OR U9461 ( .A(n9226), .B(n9225), .Z(n9227) );
  AND U9462 ( .A(n9228), .B(n9227), .Z(n9314) );
  XNOR U9463 ( .A(n9315), .B(n9314), .Z(n9316) );
  NANDN U9464 ( .A(n9230), .B(n9229), .Z(n9234) );
  NANDN U9465 ( .A(n9232), .B(n9231), .Z(n9233) );
  NAND U9466 ( .A(n9234), .B(n9233), .Z(n9317) );
  XNOR U9467 ( .A(n9316), .B(n9317), .Z(n9265) );
  XOR U9468 ( .A(n9266), .B(n9265), .Z(n9321) );
  NANDN U9469 ( .A(n9236), .B(n9235), .Z(n9240) );
  NANDN U9470 ( .A(n9238), .B(n9237), .Z(n9239) );
  AND U9471 ( .A(n9240), .B(n9239), .Z(n9320) );
  XNOR U9472 ( .A(n9321), .B(n9320), .Z(n9322) );
  XOR U9473 ( .A(n9323), .B(n9322), .Z(n9258) );
  NANDN U9474 ( .A(n9242), .B(n9241), .Z(n9246) );
  NAND U9475 ( .A(n9244), .B(n9243), .Z(n9245) );
  AND U9476 ( .A(n9246), .B(n9245), .Z(n9257) );
  XNOR U9477 ( .A(n9258), .B(n9257), .Z(n9259) );
  XNOR U9478 ( .A(n9260), .B(n9259), .Z(n9252) );
  XNOR U9479 ( .A(sreg[239]), .B(n9252), .Z(n9254) );
  NANDN U9480 ( .A(sreg[238]), .B(n9247), .Z(n9251) );
  NAND U9481 ( .A(n9249), .B(n9248), .Z(n9250) );
  NAND U9482 ( .A(n9251), .B(n9250), .Z(n9253) );
  XNOR U9483 ( .A(n9254), .B(n9253), .Z(c[239]) );
  NANDN U9484 ( .A(sreg[239]), .B(n9252), .Z(n9256) );
  NAND U9485 ( .A(n9254), .B(n9253), .Z(n9255) );
  AND U9486 ( .A(n9256), .B(n9255), .Z(n9327) );
  NANDN U9487 ( .A(n9258), .B(n9257), .Z(n9262) );
  NANDN U9488 ( .A(n9260), .B(n9259), .Z(n9261) );
  AND U9489 ( .A(n9262), .B(n9261), .Z(n9330) );
  NANDN U9490 ( .A(n9264), .B(n9263), .Z(n9268) );
  NAND U9491 ( .A(n9266), .B(n9265), .Z(n9267) );
  AND U9492 ( .A(n9268), .B(n9267), .Z(n9396) );
  NAND U9493 ( .A(n9269), .B(n9883), .Z(n9271) );
  XOR U9494 ( .A(b[11]), .B(a[118]), .Z(n9343) );
  NANDN U9495 ( .A(n9856), .B(n9343), .Z(n9270) );
  AND U9496 ( .A(n9271), .B(n9270), .Z(n9351) );
  NANDN U9497 ( .A(n10005), .B(n9272), .Z(n9274) );
  XOR U9498 ( .A(b[15]), .B(a[114]), .Z(n9367) );
  NANDN U9499 ( .A(n10006), .B(n9367), .Z(n9273) );
  AND U9500 ( .A(n9274), .B(n9273), .Z(n9350) );
  NANDN U9501 ( .A(n9685), .B(n9275), .Z(n9277) );
  XOR U9502 ( .A(b[9]), .B(a[120]), .Z(n9340) );
  NANDN U9503 ( .A(n9758), .B(n9340), .Z(n9276) );
  NAND U9504 ( .A(n9277), .B(n9276), .Z(n9349) );
  XOR U9505 ( .A(n9350), .B(n9349), .Z(n9352) );
  XOR U9506 ( .A(n9351), .B(n9352), .Z(n9388) );
  NANDN U9507 ( .A(n9279), .B(n9278), .Z(n9283) );
  OR U9508 ( .A(n9281), .B(n9280), .Z(n9282) );
  AND U9509 ( .A(n9283), .B(n9282), .Z(n9387) );
  XNOR U9510 ( .A(n9388), .B(n9387), .Z(n9389) );
  NANDN U9511 ( .A(n9285), .B(n9284), .Z(n9289) );
  NANDN U9512 ( .A(n9287), .B(n9286), .Z(n9288) );
  NAND U9513 ( .A(n9289), .B(n9288), .Z(n9390) );
  XNOR U9514 ( .A(n9389), .B(n9390), .Z(n9337) );
  NANDN U9515 ( .A(n9291), .B(n9290), .Z(n9295) );
  NANDN U9516 ( .A(n9293), .B(n9292), .Z(n9294) );
  AND U9517 ( .A(n9295), .B(n9294), .Z(n9383) );
  NANDN U9518 ( .A(n9891), .B(n9296), .Z(n9298) );
  XOR U9519 ( .A(b[13]), .B(a[116]), .Z(n9370) );
  NANDN U9520 ( .A(n9935), .B(n9370), .Z(n9297) );
  AND U9521 ( .A(n9298), .B(n9297), .Z(n9364) );
  AND U9522 ( .A(b[15]), .B(a[112]), .Z(n9361) );
  XNOR U9523 ( .A(n9362), .B(n9361), .Z(n9363) );
  XNOR U9524 ( .A(n9364), .B(n9363), .Z(n9381) );
  NANDN U9525 ( .A(n9437), .B(n9299), .Z(n9301) );
  XOR U9526 ( .A(a[124]), .B(b[5]), .Z(n9378) );
  NANDN U9527 ( .A(n9503), .B(n9378), .Z(n9300) );
  AND U9528 ( .A(n9301), .B(n9300), .Z(n9358) );
  NANDN U9529 ( .A(n9588), .B(n9302), .Z(n9304) );
  XOR U9530 ( .A(a[122]), .B(b[7]), .Z(n9346) );
  NANDN U9531 ( .A(n9639), .B(n9346), .Z(n9303) );
  AND U9532 ( .A(n9304), .B(n9303), .Z(n9356) );
  NANDN U9533 ( .A(n9374), .B(n9305), .Z(n9307) );
  XOR U9534 ( .A(a[126]), .B(b[3]), .Z(n9373) );
  NANDN U9535 ( .A(n9375), .B(n9373), .Z(n9306) );
  NAND U9536 ( .A(n9307), .B(n9306), .Z(n9355) );
  XNOR U9537 ( .A(n9356), .B(n9355), .Z(n9357) );
  XOR U9538 ( .A(n9358), .B(n9357), .Z(n9382) );
  XOR U9539 ( .A(n9381), .B(n9382), .Z(n9384) );
  XOR U9540 ( .A(n9383), .B(n9384), .Z(n9335) );
  NANDN U9541 ( .A(n9309), .B(n9308), .Z(n9313) );
  OR U9542 ( .A(n9311), .B(n9310), .Z(n9312) );
  AND U9543 ( .A(n9313), .B(n9312), .Z(n9334) );
  XNOR U9544 ( .A(n9335), .B(n9334), .Z(n9336) );
  XOR U9545 ( .A(n9337), .B(n9336), .Z(n9394) );
  NANDN U9546 ( .A(n9315), .B(n9314), .Z(n9319) );
  NANDN U9547 ( .A(n9317), .B(n9316), .Z(n9318) );
  AND U9548 ( .A(n9319), .B(n9318), .Z(n9393) );
  XNOR U9549 ( .A(n9394), .B(n9393), .Z(n9395) );
  XOR U9550 ( .A(n9396), .B(n9395), .Z(n9329) );
  NANDN U9551 ( .A(n9321), .B(n9320), .Z(n9325) );
  NAND U9552 ( .A(n9323), .B(n9322), .Z(n9324) );
  AND U9553 ( .A(n9325), .B(n9324), .Z(n9328) );
  XOR U9554 ( .A(n9329), .B(n9328), .Z(n9331) );
  XNOR U9555 ( .A(n9330), .B(n9331), .Z(n9326) );
  XOR U9556 ( .A(n9327), .B(n9326), .Z(c[240]) );
  AND U9557 ( .A(n9327), .B(n9326), .Z(n9400) );
  NANDN U9558 ( .A(n9329), .B(n9328), .Z(n9333) );
  OR U9559 ( .A(n9331), .B(n9330), .Z(n9332) );
  AND U9560 ( .A(n9333), .B(n9332), .Z(n9403) );
  NANDN U9561 ( .A(n9335), .B(n9334), .Z(n9339) );
  NAND U9562 ( .A(n9337), .B(n9336), .Z(n9338) );
  AND U9563 ( .A(n9339), .B(n9338), .Z(n9468) );
  NANDN U9564 ( .A(n9685), .B(n9340), .Z(n9342) );
  XOR U9565 ( .A(b[9]), .B(a[121]), .Z(n9440) );
  NANDN U9566 ( .A(n9758), .B(n9440), .Z(n9341) );
  AND U9567 ( .A(n9342), .B(n9341), .Z(n9445) );
  NAND U9568 ( .A(n9343), .B(n9883), .Z(n9345) );
  XOR U9569 ( .A(b[11]), .B(a[119]), .Z(n9427) );
  NANDN U9570 ( .A(n9856), .B(n9427), .Z(n9344) );
  AND U9571 ( .A(n9345), .B(n9344), .Z(n9444) );
  NANDN U9572 ( .A(n9588), .B(n9346), .Z(n9348) );
  XOR U9573 ( .A(a[123]), .B(b[7]), .Z(n9433) );
  NANDN U9574 ( .A(n9639), .B(n9433), .Z(n9347) );
  NAND U9575 ( .A(n9348), .B(n9347), .Z(n9443) );
  XOR U9576 ( .A(n9444), .B(n9443), .Z(n9446) );
  XOR U9577 ( .A(n9445), .B(n9446), .Z(n9414) );
  NANDN U9578 ( .A(n9350), .B(n9349), .Z(n9354) );
  OR U9579 ( .A(n9352), .B(n9351), .Z(n9353) );
  AND U9580 ( .A(n9354), .B(n9353), .Z(n9413) );
  XNOR U9581 ( .A(n9414), .B(n9413), .Z(n9415) );
  NANDN U9582 ( .A(n9356), .B(n9355), .Z(n9360) );
  NANDN U9583 ( .A(n9358), .B(n9357), .Z(n9359) );
  NAND U9584 ( .A(n9360), .B(n9359), .Z(n9416) );
  XNOR U9585 ( .A(n9415), .B(n9416), .Z(n9410) );
  NANDN U9586 ( .A(n9362), .B(n9361), .Z(n9366) );
  NANDN U9587 ( .A(n9364), .B(n9363), .Z(n9365) );
  AND U9588 ( .A(n9366), .B(n9365), .Z(n9461) );
  NANDN U9589 ( .A(n10005), .B(n9367), .Z(n9369) );
  XOR U9590 ( .A(b[15]), .B(a[115]), .Z(n9424) );
  NANDN U9591 ( .A(n10006), .B(n9424), .Z(n9368) );
  AND U9592 ( .A(n9369), .B(n9368), .Z(n9456) );
  NAND U9593 ( .A(b[15]), .B(a[113]), .Z(n9510) );
  NANDN U9594 ( .A(n9891), .B(n9370), .Z(n9372) );
  XOR U9595 ( .A(b[13]), .B(a[117]), .Z(n9430) );
  NANDN U9596 ( .A(n9935), .B(n9430), .Z(n9371) );
  NAND U9597 ( .A(n9372), .B(n9371), .Z(n9454) );
  XOR U9598 ( .A(n9510), .B(n9454), .Z(n9455) );
  XNOR U9599 ( .A(n9456), .B(n9455), .Z(n9459) );
  NANDN U9600 ( .A(n9374), .B(n9373), .Z(n9377) );
  XOR U9601 ( .A(a[127]), .B(b[3]), .Z(n9419) );
  NANDN U9602 ( .A(n9375), .B(n9419), .Z(n9376) );
  AND U9603 ( .A(n9377), .B(n9376), .Z(n9451) );
  NANDN U9604 ( .A(n9437), .B(n9378), .Z(n9380) );
  XOR U9605 ( .A(a[125]), .B(b[5]), .Z(n9436) );
  NANDN U9606 ( .A(n9503), .B(n9436), .Z(n9379) );
  NAND U9607 ( .A(n9380), .B(n9379), .Z(n9449) );
  XNOR U9608 ( .A(b[1]), .B(n9449), .Z(n9450) );
  XOR U9609 ( .A(n9451), .B(n9450), .Z(n9460) );
  XOR U9610 ( .A(n9459), .B(n9460), .Z(n9462) );
  XOR U9611 ( .A(n9461), .B(n9462), .Z(n9408) );
  NANDN U9612 ( .A(n9382), .B(n9381), .Z(n9386) );
  OR U9613 ( .A(n9384), .B(n9383), .Z(n9385) );
  AND U9614 ( .A(n9386), .B(n9385), .Z(n9407) );
  XNOR U9615 ( .A(n9408), .B(n9407), .Z(n9409) );
  XOR U9616 ( .A(n9410), .B(n9409), .Z(n9466) );
  NANDN U9617 ( .A(n9388), .B(n9387), .Z(n9392) );
  NANDN U9618 ( .A(n9390), .B(n9389), .Z(n9391) );
  AND U9619 ( .A(n9392), .B(n9391), .Z(n9465) );
  XNOR U9620 ( .A(n9466), .B(n9465), .Z(n9467) );
  XOR U9621 ( .A(n9468), .B(n9467), .Z(n9402) );
  NANDN U9622 ( .A(n9394), .B(n9393), .Z(n9398) );
  NAND U9623 ( .A(n9396), .B(n9395), .Z(n9397) );
  AND U9624 ( .A(n9398), .B(n9397), .Z(n9401) );
  XOR U9625 ( .A(n9402), .B(n9401), .Z(n9404) );
  XNOR U9626 ( .A(n9403), .B(n9404), .Z(n9399) );
  XOR U9627 ( .A(n9400), .B(n9399), .Z(c[241]) );
  AND U9628 ( .A(n9400), .B(n9399), .Z(n9472) );
  NANDN U9629 ( .A(n9402), .B(n9401), .Z(n9406) );
  OR U9630 ( .A(n9404), .B(n9403), .Z(n9405) );
  AND U9631 ( .A(n9406), .B(n9405), .Z(n9475) );
  NANDN U9632 ( .A(n9408), .B(n9407), .Z(n9412) );
  NAND U9633 ( .A(n9410), .B(n9409), .Z(n9411) );
  AND U9634 ( .A(n9412), .B(n9411), .Z(n9537) );
  NANDN U9635 ( .A(n9414), .B(n9413), .Z(n9418) );
  NANDN U9636 ( .A(n9416), .B(n9415), .Z(n9417) );
  AND U9637 ( .A(n9418), .B(n9417), .Z(n9535) );
  NAND U9638 ( .A(n9420), .B(n9419), .Z(n9423) );
  NAND U9639 ( .A(n9421), .B(b[3]), .Z(n9422) );
  NAND U9640 ( .A(n9423), .B(n9422), .Z(n9523) );
  AND U9641 ( .A(b[15]), .B(a[114]), .Z(n9524) );
  XOR U9642 ( .A(n9523), .B(n9524), .Z(n9525) );
  XOR U9643 ( .A(n9510), .B(n9525), .Z(n9519) );
  NANDN U9644 ( .A(n10005), .B(n9424), .Z(n9426) );
  XOR U9645 ( .A(b[15]), .B(a[116]), .Z(n9491) );
  NANDN U9646 ( .A(n10006), .B(n9491), .Z(n9425) );
  AND U9647 ( .A(n9426), .B(n9425), .Z(n9518) );
  NAND U9648 ( .A(n9427), .B(n9883), .Z(n9429) );
  XOR U9649 ( .A(b[11]), .B(a[120]), .Z(n9507) );
  NANDN U9650 ( .A(n9856), .B(n9507), .Z(n9428) );
  NAND U9651 ( .A(n9429), .B(n9428), .Z(n9517) );
  XOR U9652 ( .A(n9518), .B(n9517), .Z(n9520) );
  XNOR U9653 ( .A(n9519), .B(n9520), .Z(n9487) );
  NANDN U9654 ( .A(n9891), .B(n9430), .Z(n9432) );
  XOR U9655 ( .A(b[13]), .B(a[118]), .Z(n9500) );
  NANDN U9656 ( .A(n9935), .B(n9500), .Z(n9431) );
  AND U9657 ( .A(n9432), .B(n9431), .Z(n9486) );
  NANDN U9658 ( .A(n9588), .B(n9433), .Z(n9435) );
  XOR U9659 ( .A(a[124]), .B(b[7]), .Z(n9497) );
  NANDN U9660 ( .A(n9639), .B(n9497), .Z(n9434) );
  AND U9661 ( .A(n9435), .B(n9434), .Z(n9514) );
  NANDN U9662 ( .A(n9437), .B(n9436), .Z(n9439) );
  XOR U9663 ( .A(a[126]), .B(b[5]), .Z(n9504) );
  NANDN U9664 ( .A(n9503), .B(n9504), .Z(n9438) );
  AND U9665 ( .A(n9439), .B(n9438), .Z(n9512) );
  NANDN U9666 ( .A(n9685), .B(n9440), .Z(n9442) );
  XOR U9667 ( .A(b[9]), .B(a[122]), .Z(n9494) );
  NANDN U9668 ( .A(n9758), .B(n9494), .Z(n9441) );
  NAND U9669 ( .A(n9442), .B(n9441), .Z(n9511) );
  XNOR U9670 ( .A(n9512), .B(n9511), .Z(n9513) );
  XNOR U9671 ( .A(n9514), .B(n9513), .Z(n9485) );
  XOR U9672 ( .A(n9486), .B(n9485), .Z(n9488) );
  XNOR U9673 ( .A(n9487), .B(n9488), .Z(n9482) );
  NANDN U9674 ( .A(n9444), .B(n9443), .Z(n9448) );
  OR U9675 ( .A(n9446), .B(n9445), .Z(n9447) );
  AND U9676 ( .A(n9448), .B(n9447), .Z(n9480) );
  NANDN U9677 ( .A(b[1]), .B(n9449), .Z(n9453) );
  NANDN U9678 ( .A(n9451), .B(n9450), .Z(n9452) );
  NAND U9679 ( .A(n9453), .B(n9452), .Z(n9479) );
  XNOR U9680 ( .A(n9480), .B(n9479), .Z(n9481) );
  XOR U9681 ( .A(n9482), .B(n9481), .Z(n9531) );
  IV U9682 ( .A(n9510), .Z(n9568) );
  NANDN U9683 ( .A(n9568), .B(n9454), .Z(n9458) );
  NANDN U9684 ( .A(n9456), .B(n9455), .Z(n9457) );
  AND U9685 ( .A(n9458), .B(n9457), .Z(n9528) );
  NANDN U9686 ( .A(n9460), .B(n9459), .Z(n9464) );
  OR U9687 ( .A(n9462), .B(n9461), .Z(n9463) );
  NAND U9688 ( .A(n9464), .B(n9463), .Z(n9529) );
  XNOR U9689 ( .A(n9528), .B(n9529), .Z(n9530) );
  XNOR U9690 ( .A(n9531), .B(n9530), .Z(n9534) );
  XNOR U9691 ( .A(n9535), .B(n9534), .Z(n9536) );
  XNOR U9692 ( .A(n9537), .B(n9536), .Z(n9473) );
  NANDN U9693 ( .A(n9466), .B(n9465), .Z(n9470) );
  NAND U9694 ( .A(n9468), .B(n9467), .Z(n9469) );
  NAND U9695 ( .A(n9470), .B(n9469), .Z(n9474) );
  XOR U9696 ( .A(n9473), .B(n9474), .Z(n9476) );
  XNOR U9697 ( .A(n9475), .B(n9476), .Z(n9471) );
  XOR U9698 ( .A(n9472), .B(n9471), .Z(c[242]) );
  AND U9699 ( .A(n9472), .B(n9471), .Z(n9541) );
  NANDN U9700 ( .A(n9474), .B(n9473), .Z(n9478) );
  OR U9701 ( .A(n9476), .B(n9475), .Z(n9477) );
  AND U9702 ( .A(n9478), .B(n9477), .Z(n9544) );
  NANDN U9703 ( .A(n9480), .B(n9479), .Z(n9484) );
  NAND U9704 ( .A(n9482), .B(n9481), .Z(n9483) );
  AND U9705 ( .A(n9484), .B(n9483), .Z(n9549) );
  NANDN U9706 ( .A(n9486), .B(n9485), .Z(n9490) );
  NANDN U9707 ( .A(n9488), .B(n9487), .Z(n9489) );
  AND U9708 ( .A(n9490), .B(n9489), .Z(n9555) );
  NANDN U9709 ( .A(n10005), .B(n9491), .Z(n9493) );
  XOR U9710 ( .A(b[15]), .B(a[117]), .Z(n9576) );
  NANDN U9711 ( .A(n10006), .B(n9576), .Z(n9492) );
  AND U9712 ( .A(n9493), .B(n9492), .Z(n9598) );
  NANDN U9713 ( .A(n9685), .B(n9494), .Z(n9496) );
  XOR U9714 ( .A(b[9]), .B(a[123]), .Z(n9584) );
  NANDN U9715 ( .A(n9758), .B(n9584), .Z(n9495) );
  AND U9716 ( .A(n9496), .B(n9495), .Z(n9563) );
  NANDN U9717 ( .A(n9588), .B(n9497), .Z(n9499) );
  XOR U9718 ( .A(a[125]), .B(b[7]), .Z(n9587) );
  NANDN U9719 ( .A(n9639), .B(n9587), .Z(n9498) );
  AND U9720 ( .A(n9499), .B(n9498), .Z(n9561) );
  NANDN U9721 ( .A(n9891), .B(n9500), .Z(n9502) );
  XOR U9722 ( .A(b[13]), .B(a[119]), .Z(n9594) );
  NANDN U9723 ( .A(n9935), .B(n9594), .Z(n9501) );
  NAND U9724 ( .A(n9502), .B(n9501), .Z(n9560) );
  XNOR U9725 ( .A(n9561), .B(n9560), .Z(n9562) );
  XNOR U9726 ( .A(n9563), .B(n9562), .Z(n9597) );
  XNOR U9727 ( .A(n9598), .B(n9597), .Z(n9600) );
  XNOR U9728 ( .A(a[127]), .B(b[5]), .Z(n9579) );
  OR U9729 ( .A(n9579), .B(n9503), .Z(n9506) );
  NAND U9730 ( .A(n9580), .B(n9504), .Z(n9505) );
  AND U9731 ( .A(n9506), .B(n9505), .Z(n9573) );
  NAND U9732 ( .A(n9507), .B(n9883), .Z(n9509) );
  XOR U9733 ( .A(b[11]), .B(a[121]), .Z(n9591) );
  NANDN U9734 ( .A(n9856), .B(n9591), .Z(n9508) );
  NAND U9735 ( .A(n9509), .B(n9508), .Z(n9572) );
  XNOR U9736 ( .A(n9573), .B(n9572), .Z(n9575) );
  AND U9737 ( .A(b[15]), .B(a[115]), .Z(n9566) );
  XOR U9738 ( .A(n9567), .B(n9566), .Z(n9569) );
  XOR U9739 ( .A(n9510), .B(n9569), .Z(n9574) );
  XOR U9740 ( .A(n9575), .B(n9574), .Z(n9599) );
  XOR U9741 ( .A(n9600), .B(n9599), .Z(n9554) );
  XNOR U9742 ( .A(n9555), .B(n9554), .Z(n9556) );
  NANDN U9743 ( .A(n9512), .B(n9511), .Z(n9516) );
  NANDN U9744 ( .A(n9514), .B(n9513), .Z(n9515) );
  AND U9745 ( .A(n9516), .B(n9515), .Z(n9604) );
  NANDN U9746 ( .A(n9518), .B(n9517), .Z(n9522) );
  NANDN U9747 ( .A(n9520), .B(n9519), .Z(n9521) );
  AND U9748 ( .A(n9522), .B(n9521), .Z(n9602) );
  NAND U9749 ( .A(n9524), .B(n9523), .Z(n9527) );
  NANDN U9750 ( .A(n9568), .B(n9525), .Z(n9526) );
  NAND U9751 ( .A(n9527), .B(n9526), .Z(n9601) );
  XNOR U9752 ( .A(n9602), .B(n9601), .Z(n9603) );
  XOR U9753 ( .A(n9604), .B(n9603), .Z(n9557) );
  XNOR U9754 ( .A(n9556), .B(n9557), .Z(n9548) );
  XNOR U9755 ( .A(n9549), .B(n9548), .Z(n9551) );
  NANDN U9756 ( .A(n9529), .B(n9528), .Z(n9533) );
  NANDN U9757 ( .A(n9531), .B(n9530), .Z(n9532) );
  AND U9758 ( .A(n9533), .B(n9532), .Z(n9550) );
  XOR U9759 ( .A(n9551), .B(n9550), .Z(n9543) );
  NANDN U9760 ( .A(n9535), .B(n9534), .Z(n9539) );
  NANDN U9761 ( .A(n9537), .B(n9536), .Z(n9538) );
  NAND U9762 ( .A(n9539), .B(n9538), .Z(n9542) );
  XOR U9763 ( .A(n9543), .B(n9542), .Z(n9545) );
  XNOR U9764 ( .A(n9544), .B(n9545), .Z(n9540) );
  XOR U9765 ( .A(n9541), .B(n9540), .Z(c[243]) );
  AND U9766 ( .A(n9541), .B(n9540), .Z(n9608) );
  NANDN U9767 ( .A(n9543), .B(n9542), .Z(n9547) );
  OR U9768 ( .A(n9545), .B(n9544), .Z(n9546) );
  AND U9769 ( .A(n9547), .B(n9546), .Z(n9612) );
  NANDN U9770 ( .A(n9549), .B(n9548), .Z(n9553) );
  NAND U9771 ( .A(n9551), .B(n9550), .Z(n9552) );
  AND U9772 ( .A(n9553), .B(n9552), .Z(n9610) );
  NANDN U9773 ( .A(n9555), .B(n9554), .Z(n9559) );
  NANDN U9774 ( .A(n9557), .B(n9556), .Z(n9558) );
  AND U9775 ( .A(n9559), .B(n9558), .Z(n9616) );
  NANDN U9776 ( .A(n9561), .B(n9560), .Z(n9565) );
  NANDN U9777 ( .A(n9563), .B(n9562), .Z(n9564) );
  AND U9778 ( .A(n9565), .B(n9564), .Z(n9624) );
  NANDN U9779 ( .A(n9567), .B(n9566), .Z(n9571) );
  NANDN U9780 ( .A(n9569), .B(n9568), .Z(n9570) );
  AND U9781 ( .A(n9571), .B(n9570), .Z(n9621) );
  XNOR U9782 ( .A(n9621), .B(n9622), .Z(n9623) );
  XOR U9783 ( .A(n9624), .B(n9623), .Z(n9620) );
  NANDN U9784 ( .A(n10005), .B(n9576), .Z(n9578) );
  XOR U9785 ( .A(b[15]), .B(a[118]), .Z(n9652) );
  NANDN U9786 ( .A(n10006), .B(n9652), .Z(n9577) );
  AND U9787 ( .A(n9578), .B(n9577), .Z(n9658) );
  NAND U9788 ( .A(b[15]), .B(a[116]), .Z(n9655) );
  ANDN U9789 ( .B(n9580), .A(n9579), .Z(n9583) );
  NAND U9790 ( .A(b[5]), .B(n9581), .Z(n9582) );
  NANDN U9791 ( .A(n9583), .B(n9582), .Z(n9656) );
  XOR U9792 ( .A(n9655), .B(n9656), .Z(n9657) );
  XOR U9793 ( .A(n9658), .B(n9657), .Z(n9629) );
  NANDN U9794 ( .A(n9685), .B(n9584), .Z(n9586) );
  XOR U9795 ( .A(a[124]), .B(b[9]), .Z(n9646) );
  NANDN U9796 ( .A(n9758), .B(n9646), .Z(n9585) );
  AND U9797 ( .A(n9586), .B(n9585), .Z(n9635) );
  NANDN U9798 ( .A(n9588), .B(n9587), .Z(n9590) );
  XOR U9799 ( .A(a[126]), .B(b[7]), .Z(n9640) );
  NANDN U9800 ( .A(n9639), .B(n9640), .Z(n9589) );
  AND U9801 ( .A(n9590), .B(n9589), .Z(n9634) );
  NAND U9802 ( .A(n9591), .B(n9883), .Z(n9593) );
  XOR U9803 ( .A(b[11]), .B(a[122]), .Z(n9643) );
  NANDN U9804 ( .A(n9856), .B(n9643), .Z(n9592) );
  NAND U9805 ( .A(n9593), .B(n9592), .Z(n9633) );
  XOR U9806 ( .A(n9634), .B(n9633), .Z(n9636) );
  XOR U9807 ( .A(n9635), .B(n9636), .Z(n9628) );
  NAND U9808 ( .A(n9972), .B(n9594), .Z(n9596) );
  XNOR U9809 ( .A(b[13]), .B(a[120]), .Z(n9649) );
  NANDN U9810 ( .A(n9649), .B(n9973), .Z(n9595) );
  AND U9811 ( .A(n9596), .B(n9595), .Z(n9627) );
  XOR U9812 ( .A(n9628), .B(n9627), .Z(n9630) );
  XOR U9813 ( .A(n9629), .B(n9630), .Z(n9617) );
  XOR U9814 ( .A(n9617), .B(n9618), .Z(n9619) );
  XOR U9815 ( .A(n9620), .B(n9619), .Z(n9613) );
  NANDN U9816 ( .A(n9602), .B(n9601), .Z(n9606) );
  NANDN U9817 ( .A(n9604), .B(n9603), .Z(n9605) );
  AND U9818 ( .A(n9606), .B(n9605), .Z(n9614) );
  XOR U9819 ( .A(n9613), .B(n9614), .Z(n9615) );
  XOR U9820 ( .A(n9616), .B(n9615), .Z(n9609) );
  XOR U9821 ( .A(n9610), .B(n9609), .Z(n9611) );
  XOR U9822 ( .A(n9612), .B(n9611), .Z(n9607) );
  XOR U9823 ( .A(n9608), .B(n9607), .Z(c[244]) );
  AND U9824 ( .A(n9608), .B(n9607), .Z(n9662) );
  NANDN U9825 ( .A(n9622), .B(n9621), .Z(n9626) );
  NAND U9826 ( .A(n9624), .B(n9623), .Z(n9625) );
  AND U9827 ( .A(n9626), .B(n9625), .Z(n9670) );
  NANDN U9828 ( .A(n9628), .B(n9627), .Z(n9632) );
  NANDN U9829 ( .A(n9630), .B(n9629), .Z(n9631) );
  AND U9830 ( .A(n9632), .B(n9631), .Z(n9678) );
  NANDN U9831 ( .A(n9634), .B(n9633), .Z(n9638) );
  OR U9832 ( .A(n9636), .B(n9635), .Z(n9637) );
  AND U9833 ( .A(n9638), .B(n9637), .Z(n9720) );
  XNOR U9834 ( .A(a[127]), .B(b[7]), .Z(n9694) );
  OR U9835 ( .A(n9694), .B(n9639), .Z(n9642) );
  NAND U9836 ( .A(n9695), .B(n9640), .Z(n9641) );
  AND U9837 ( .A(n9642), .B(n9641), .Z(n9712) );
  NAND U9838 ( .A(n9643), .B(n9883), .Z(n9645) );
  XOR U9839 ( .A(b[11]), .B(a[123]), .Z(n9681) );
  NANDN U9840 ( .A(n9856), .B(n9681), .Z(n9644) );
  NAND U9841 ( .A(n9645), .B(n9644), .Z(n9711) );
  XNOR U9842 ( .A(n9712), .B(n9711), .Z(n9713) );
  XOR U9843 ( .A(n9706), .B(n9655), .Z(n9707) );
  NAND U9844 ( .A(b[15]), .B(a[117]), .Z(n9708) );
  XOR U9845 ( .A(n9707), .B(n9708), .Z(n9714) );
  XNOR U9846 ( .A(n9713), .B(n9714), .Z(n9718) );
  NANDN U9847 ( .A(n9685), .B(n9646), .Z(n9648) );
  XOR U9848 ( .A(a[125]), .B(b[9]), .Z(n9684) );
  NANDN U9849 ( .A(n9758), .B(n9684), .Z(n9647) );
  AND U9850 ( .A(n9648), .B(n9647), .Z(n9702) );
  NANDN U9851 ( .A(n9649), .B(n9972), .Z(n9651) );
  XOR U9852 ( .A(b[13]), .B(a[121]), .Z(n9688) );
  NANDN U9853 ( .A(n9935), .B(n9688), .Z(n9650) );
  AND U9854 ( .A(n9651), .B(n9650), .Z(n9700) );
  NANDN U9855 ( .A(n10005), .B(n9652), .Z(n9654) );
  XOR U9856 ( .A(b[15]), .B(a[119]), .Z(n9691) );
  NANDN U9857 ( .A(n10006), .B(n9691), .Z(n9653) );
  NAND U9858 ( .A(n9654), .B(n9653), .Z(n9699) );
  XNOR U9859 ( .A(n9700), .B(n9699), .Z(n9701) );
  XOR U9860 ( .A(n9702), .B(n9701), .Z(n9719) );
  XOR U9861 ( .A(n9718), .B(n9719), .Z(n9721) );
  XOR U9862 ( .A(n9720), .B(n9721), .Z(n9676) );
  IV U9863 ( .A(n9655), .Z(n9705) );
  NANDN U9864 ( .A(n9705), .B(n9656), .Z(n9660) );
  NANDN U9865 ( .A(n9658), .B(n9657), .Z(n9659) );
  AND U9866 ( .A(n9660), .B(n9659), .Z(n9675) );
  XNOR U9867 ( .A(n9676), .B(n9675), .Z(n9677) );
  XNOR U9868 ( .A(n9678), .B(n9677), .Z(n9669) );
  XOR U9869 ( .A(n9670), .B(n9669), .Z(n9672) );
  XNOR U9870 ( .A(n9671), .B(n9672), .Z(n9663) );
  XOR U9871 ( .A(n9664), .B(n9663), .Z(n9666) );
  XNOR U9872 ( .A(n9665), .B(n9666), .Z(n9661) );
  XOR U9873 ( .A(n9662), .B(n9661), .Z(c[245]) );
  AND U9874 ( .A(n9662), .B(n9661), .Z(n9725) );
  NANDN U9875 ( .A(n9664), .B(n9663), .Z(n9668) );
  OR U9876 ( .A(n9666), .B(n9665), .Z(n9667) );
  AND U9877 ( .A(n9668), .B(n9667), .Z(n9728) );
  NANDN U9878 ( .A(n9670), .B(n9669), .Z(n9674) );
  NANDN U9879 ( .A(n9672), .B(n9671), .Z(n9673) );
  AND U9880 ( .A(n9674), .B(n9673), .Z(n9727) );
  NANDN U9881 ( .A(n9676), .B(n9675), .Z(n9680) );
  NANDN U9882 ( .A(n9678), .B(n9677), .Z(n9679) );
  AND U9883 ( .A(n9680), .B(n9679), .Z(n9735) );
  NAND U9884 ( .A(n9681), .B(n9883), .Z(n9683) );
  XOR U9885 ( .A(b[11]), .B(a[124]), .Z(n9755) );
  NANDN U9886 ( .A(n9856), .B(n9755), .Z(n9682) );
  AND U9887 ( .A(n9683), .B(n9682), .Z(n9743) );
  NANDN U9888 ( .A(n9685), .B(n9684), .Z(n9687) );
  XOR U9889 ( .A(a[126]), .B(b[9]), .Z(n9759) );
  NANDN U9890 ( .A(n9758), .B(n9759), .Z(n9686) );
  AND U9891 ( .A(n9687), .B(n9686), .Z(n9742) );
  NANDN U9892 ( .A(n9891), .B(n9688), .Z(n9690) );
  XOR U9893 ( .A(b[13]), .B(a[122]), .Z(n9762) );
  NANDN U9894 ( .A(n9935), .B(n9762), .Z(n9689) );
  NAND U9895 ( .A(n9690), .B(n9689), .Z(n9741) );
  XOR U9896 ( .A(n9742), .B(n9741), .Z(n9744) );
  XOR U9897 ( .A(n9743), .B(n9744), .Z(n9768) );
  NANDN U9898 ( .A(n10005), .B(n9691), .Z(n9693) );
  XOR U9899 ( .A(b[15]), .B(a[120]), .Z(n9752) );
  NANDN U9900 ( .A(n10006), .B(n9752), .Z(n9692) );
  AND U9901 ( .A(n9693), .B(n9692), .Z(n9749) );
  NAND U9902 ( .A(b[15]), .B(a[118]), .Z(n9766) );
  ANDN U9903 ( .B(n9695), .A(n9694), .Z(n9698) );
  NAND U9904 ( .A(b[7]), .B(n9696), .Z(n9697) );
  NANDN U9905 ( .A(n9698), .B(n9697), .Z(n9747) );
  XOR U9906 ( .A(n9766), .B(n9747), .Z(n9748) );
  XOR U9907 ( .A(n9749), .B(n9748), .Z(n9767) );
  XNOR U9908 ( .A(n9768), .B(n9767), .Z(n9769) );
  NANDN U9909 ( .A(n9700), .B(n9699), .Z(n9704) );
  NANDN U9910 ( .A(n9702), .B(n9701), .Z(n9703) );
  NAND U9911 ( .A(n9704), .B(n9703), .Z(n9770) );
  XNOR U9912 ( .A(n9769), .B(n9770), .Z(n9738) );
  NANDN U9913 ( .A(n9706), .B(n9705), .Z(n9710) );
  NANDN U9914 ( .A(n9708), .B(n9707), .Z(n9709) );
  AND U9915 ( .A(n9710), .B(n9709), .Z(n9740) );
  NANDN U9916 ( .A(n9712), .B(n9711), .Z(n9716) );
  NANDN U9917 ( .A(n9714), .B(n9713), .Z(n9715) );
  AND U9918 ( .A(n9716), .B(n9715), .Z(n9739) );
  XNOR U9919 ( .A(n9740), .B(n9739), .Z(n9717) );
  XNOR U9920 ( .A(n9738), .B(n9717), .Z(n9732) );
  NANDN U9921 ( .A(n9719), .B(n9718), .Z(n9723) );
  OR U9922 ( .A(n9721), .B(n9720), .Z(n9722) );
  NAND U9923 ( .A(n9723), .B(n9722), .Z(n9733) );
  XNOR U9924 ( .A(n9732), .B(n9733), .Z(n9734) );
  XNOR U9925 ( .A(n9735), .B(n9734), .Z(n9726) );
  XOR U9926 ( .A(n9727), .B(n9726), .Z(n9729) );
  XNOR U9927 ( .A(n9728), .B(n9729), .Z(n9724) );
  XOR U9928 ( .A(n9725), .B(n9724), .Z(c[246]) );
  AND U9929 ( .A(n9725), .B(n9724), .Z(n9774) );
  NANDN U9930 ( .A(n9727), .B(n9726), .Z(n9731) );
  OR U9931 ( .A(n9729), .B(n9728), .Z(n9730) );
  AND U9932 ( .A(n9731), .B(n9730), .Z(n9777) );
  NANDN U9933 ( .A(n9733), .B(n9732), .Z(n9737) );
  NANDN U9934 ( .A(n9735), .B(n9734), .Z(n9736) );
  AND U9935 ( .A(n9737), .B(n9736), .Z(n9776) );
  NANDN U9936 ( .A(n9742), .B(n9741), .Z(n9746) );
  OR U9937 ( .A(n9744), .B(n9743), .Z(n9745) );
  AND U9938 ( .A(n9746), .B(n9745), .Z(n9789) );
  IV U9939 ( .A(n9766), .Z(n9810) );
  NANDN U9940 ( .A(n9810), .B(n9747), .Z(n9751) );
  NANDN U9941 ( .A(n9749), .B(n9748), .Z(n9750) );
  AND U9942 ( .A(n9751), .B(n9750), .Z(n9788) );
  NANDN U9943 ( .A(n10005), .B(n9752), .Z(n9754) );
  XOR U9944 ( .A(b[15]), .B(a[121]), .Z(n9799) );
  NANDN U9945 ( .A(n10006), .B(n9799), .Z(n9753) );
  AND U9946 ( .A(n9754), .B(n9753), .Z(n9822) );
  NAND U9947 ( .A(n9755), .B(n9883), .Z(n9757) );
  XOR U9948 ( .A(b[11]), .B(a[125]), .Z(n9816) );
  NANDN U9949 ( .A(n9856), .B(n9816), .Z(n9756) );
  AND U9950 ( .A(n9757), .B(n9756), .Z(n9820) );
  XNOR U9951 ( .A(a[127]), .B(b[9]), .Z(n9802) );
  OR U9952 ( .A(n9802), .B(n9758), .Z(n9761) );
  NAND U9953 ( .A(n9803), .B(n9759), .Z(n9760) );
  AND U9954 ( .A(n9761), .B(n9760), .Z(n9794) );
  NANDN U9955 ( .A(n9891), .B(n9762), .Z(n9764) );
  XOR U9956 ( .A(b[13]), .B(a[123]), .Z(n9813) );
  NANDN U9957 ( .A(n9935), .B(n9813), .Z(n9763) );
  NAND U9958 ( .A(n9764), .B(n9763), .Z(n9793) );
  XNOR U9959 ( .A(n9794), .B(n9793), .Z(n9795) );
  IV U9960 ( .A(n9765), .Z(n9808) );
  AND U9961 ( .A(b[15]), .B(a[119]), .Z(n9807) );
  XOR U9962 ( .A(n9808), .B(n9807), .Z(n9809) );
  XOR U9963 ( .A(n9766), .B(n9809), .Z(n9796) );
  XOR U9964 ( .A(n9795), .B(n9796), .Z(n9819) );
  XNOR U9965 ( .A(n9820), .B(n9819), .Z(n9821) );
  XNOR U9966 ( .A(n9822), .B(n9821), .Z(n9787) );
  XOR U9967 ( .A(n9788), .B(n9787), .Z(n9790) );
  XOR U9968 ( .A(n9789), .B(n9790), .Z(n9782) );
  NANDN U9969 ( .A(n9768), .B(n9767), .Z(n9772) );
  NANDN U9970 ( .A(n9770), .B(n9769), .Z(n9771) );
  NAND U9971 ( .A(n9772), .B(n9771), .Z(n9781) );
  XNOR U9972 ( .A(n9782), .B(n9781), .Z(n9783) );
  XNOR U9973 ( .A(n9784), .B(n9783), .Z(n9775) );
  XOR U9974 ( .A(n9776), .B(n9775), .Z(n9778) );
  XNOR U9975 ( .A(n9777), .B(n9778), .Z(n9773) );
  XOR U9976 ( .A(n9774), .B(n9773), .Z(c[247]) );
  AND U9977 ( .A(n9774), .B(n9773), .Z(n9826) );
  NANDN U9978 ( .A(n9776), .B(n9775), .Z(n9780) );
  OR U9979 ( .A(n9778), .B(n9777), .Z(n9779) );
  AND U9980 ( .A(n9780), .B(n9779), .Z(n9829) );
  NANDN U9981 ( .A(n9782), .B(n9781), .Z(n9786) );
  NANDN U9982 ( .A(n9784), .B(n9783), .Z(n9785) );
  AND U9983 ( .A(n9786), .B(n9785), .Z(n9828) );
  NANDN U9984 ( .A(n9788), .B(n9787), .Z(n9792) );
  OR U9985 ( .A(n9790), .B(n9789), .Z(n9791) );
  AND U9986 ( .A(n9792), .B(n9791), .Z(n9835) );
  NANDN U9987 ( .A(n9794), .B(n9793), .Z(n9798) );
  NAND U9988 ( .A(n9796), .B(n9795), .Z(n9797) );
  AND U9989 ( .A(n9798), .B(n9797), .Z(n9840) );
  NANDN U9990 ( .A(n10005), .B(n9799), .Z(n9801) );
  XOR U9991 ( .A(b[15]), .B(a[122]), .Z(n9863) );
  NANDN U9992 ( .A(n10006), .B(n9863), .Z(n9800) );
  AND U9993 ( .A(n9801), .B(n9800), .Z(n9853) );
  NAND U9994 ( .A(b[15]), .B(a[120]), .Z(n9867) );
  ANDN U9995 ( .B(n9803), .A(n9802), .Z(n9806) );
  NAND U9996 ( .A(b[9]), .B(n9804), .Z(n9805) );
  NANDN U9997 ( .A(n9806), .B(n9805), .Z(n9851) );
  XOR U9998 ( .A(n9867), .B(n9851), .Z(n9852) );
  XNOR U9999 ( .A(n9853), .B(n9852), .Z(n9839) );
  XNOR U10000 ( .A(n9840), .B(n9839), .Z(n9842) );
  NANDN U10001 ( .A(n9808), .B(n9807), .Z(n9812) );
  ANDN U10002 ( .B(n9810), .A(n9809), .Z(n9811) );
  ANDN U10003 ( .B(n9812), .A(n9811), .Z(n9848) );
  NANDN U10004 ( .A(n9891), .B(n9813), .Z(n9815) );
  XOR U10005 ( .A(b[13]), .B(a[124]), .Z(n9860) );
  NANDN U10006 ( .A(n9935), .B(n9860), .Z(n9814) );
  AND U10007 ( .A(n9815), .B(n9814), .Z(n9846) );
  NAND U10008 ( .A(n9816), .B(n9883), .Z(n9818) );
  XOR U10009 ( .A(a[126]), .B(b[11]), .Z(n9857) );
  NANDN U10010 ( .A(n9856), .B(n9857), .Z(n9817) );
  NAND U10011 ( .A(n9818), .B(n9817), .Z(n9845) );
  XNOR U10012 ( .A(n9846), .B(n9845), .Z(n9847) );
  XNOR U10013 ( .A(n9848), .B(n9847), .Z(n9841) );
  XOR U10014 ( .A(n9842), .B(n9841), .Z(n9834) );
  NANDN U10015 ( .A(n9820), .B(n9819), .Z(n9824) );
  NANDN U10016 ( .A(n9822), .B(n9821), .Z(n9823) );
  AND U10017 ( .A(n9824), .B(n9823), .Z(n9833) );
  XOR U10018 ( .A(n9834), .B(n9833), .Z(n9836) );
  XNOR U10019 ( .A(n9835), .B(n9836), .Z(n9827) );
  XOR U10020 ( .A(n9828), .B(n9827), .Z(n9830) );
  XNOR U10021 ( .A(n9829), .B(n9830), .Z(n9825) );
  XOR U10022 ( .A(n9826), .B(n9825), .Z(c[248]) );
  AND U10023 ( .A(n9826), .B(n9825), .Z(n9869) );
  NANDN U10024 ( .A(n9828), .B(n9827), .Z(n9832) );
  OR U10025 ( .A(n9830), .B(n9829), .Z(n9831) );
  AND U10026 ( .A(n9832), .B(n9831), .Z(n9872) );
  NANDN U10027 ( .A(n9834), .B(n9833), .Z(n9838) );
  NANDN U10028 ( .A(n9836), .B(n9835), .Z(n9837) );
  AND U10029 ( .A(n9838), .B(n9837), .Z(n9871) );
  NANDN U10030 ( .A(n9840), .B(n9839), .Z(n9844) );
  NAND U10031 ( .A(n9842), .B(n9841), .Z(n9843) );
  AND U10032 ( .A(n9844), .B(n9843), .Z(n9908) );
  NANDN U10033 ( .A(n9846), .B(n9845), .Z(n9850) );
  NANDN U10034 ( .A(n9848), .B(n9847), .Z(n9849) );
  AND U10035 ( .A(n9850), .B(n9849), .Z(n9907) );
  IV U10036 ( .A(n9867), .Z(n9895) );
  NANDN U10037 ( .A(n9895), .B(n9851), .Z(n9855) );
  NANDN U10038 ( .A(n9853), .B(n9852), .Z(n9854) );
  AND U10039 ( .A(n9855), .B(n9854), .Z(n9879) );
  XNOR U10040 ( .A(a[127]), .B(b[11]), .Z(n9884) );
  OR U10041 ( .A(n9884), .B(n9856), .Z(n9859) );
  NAND U10042 ( .A(n9883), .B(n9857), .Z(n9858) );
  AND U10043 ( .A(n9859), .B(n9858), .Z(n9877) );
  NANDN U10044 ( .A(n9891), .B(n9860), .Z(n9862) );
  XOR U10045 ( .A(b[13]), .B(a[125]), .Z(n9890) );
  NANDN U10046 ( .A(n9935), .B(n9890), .Z(n9861) );
  AND U10047 ( .A(n9862), .B(n9861), .Z(n9901) );
  NANDN U10048 ( .A(n10005), .B(n9863), .Z(n9865) );
  XOR U10049 ( .A(b[15]), .B(a[123]), .Z(n9887) );
  NANDN U10050 ( .A(n10006), .B(n9887), .Z(n9864) );
  NAND U10051 ( .A(n9865), .B(n9864), .Z(n9900) );
  XNOR U10052 ( .A(n9901), .B(n9900), .Z(n9902) );
  IV U10053 ( .A(n9866), .Z(n9897) );
  AND U10054 ( .A(b[15]), .B(a[121]), .Z(n9896) );
  XOR U10055 ( .A(n9897), .B(n9896), .Z(n9894) );
  XOR U10056 ( .A(n9867), .B(n9894), .Z(n9903) );
  XOR U10057 ( .A(n9902), .B(n9903), .Z(n9876) );
  XNOR U10058 ( .A(n9877), .B(n9876), .Z(n9878) );
  XNOR U10059 ( .A(n9879), .B(n9878), .Z(n9906) );
  XOR U10060 ( .A(n9907), .B(n9906), .Z(n9909) );
  XNOR U10061 ( .A(n9908), .B(n9909), .Z(n9870) );
  XOR U10062 ( .A(n9871), .B(n9870), .Z(n9873) );
  XNOR U10063 ( .A(n9872), .B(n9873), .Z(n9868) );
  XOR U10064 ( .A(n9869), .B(n9868), .Z(c[249]) );
  AND U10065 ( .A(n9869), .B(n9868), .Z(n9913) );
  NANDN U10066 ( .A(n9871), .B(n9870), .Z(n9875) );
  OR U10067 ( .A(n9873), .B(n9872), .Z(n9874) );
  AND U10068 ( .A(n9875), .B(n9874), .Z(n9916) );
  NANDN U10069 ( .A(n9877), .B(n9876), .Z(n9881) );
  NANDN U10070 ( .A(n9879), .B(n9878), .Z(n9880) );
  AND U10071 ( .A(n9881), .B(n9880), .Z(n9922) );
  AND U10072 ( .A(b[15]), .B(a[122]), .Z(n9967) );
  XOR U10073 ( .A(b[9]), .B(b[10]), .Z(n9882) );
  AND U10074 ( .A(b[11]), .B(n9882), .Z(n9886) );
  NANDN U10075 ( .A(n9884), .B(n9883), .Z(n9885) );
  NANDN U10076 ( .A(n9886), .B(n9885), .Z(n9939) );
  XNOR U10077 ( .A(n9967), .B(n9939), .Z(n9941) );
  NAND U10078 ( .A(n9987), .B(n9887), .Z(n9889) );
  XNOR U10079 ( .A(b[15]), .B(a[124]), .Z(n9932) );
  NANDN U10080 ( .A(n9932), .B(n9989), .Z(n9888) );
  AND U10081 ( .A(n9889), .B(n9888), .Z(n9940) );
  XOR U10082 ( .A(n9941), .B(n9940), .Z(n9928) );
  NANDN U10083 ( .A(n9891), .B(n9890), .Z(n9893) );
  XOR U10084 ( .A(b[13]), .B(a[126]), .Z(n9936) );
  NANDN U10085 ( .A(n9935), .B(n9936), .Z(n9892) );
  AND U10086 ( .A(n9893), .B(n9892), .Z(n9927) );
  ANDN U10087 ( .B(n9895), .A(n9894), .Z(n9899) );
  NANDN U10088 ( .A(n9897), .B(n9896), .Z(n9898) );
  NANDN U10089 ( .A(n9899), .B(n9898), .Z(n9926) );
  XOR U10090 ( .A(n9927), .B(n9926), .Z(n9929) );
  XOR U10091 ( .A(n9928), .B(n9929), .Z(n9921) );
  NANDN U10092 ( .A(n9901), .B(n9900), .Z(n9905) );
  NAND U10093 ( .A(n9903), .B(n9902), .Z(n9904) );
  AND U10094 ( .A(n9905), .B(n9904), .Z(n9920) );
  XOR U10095 ( .A(n9921), .B(n9920), .Z(n9923) );
  XNOR U10096 ( .A(n9922), .B(n9923), .Z(n9914) );
  NANDN U10097 ( .A(n9907), .B(n9906), .Z(n9911) );
  OR U10098 ( .A(n9909), .B(n9908), .Z(n9910) );
  NAND U10099 ( .A(n9911), .B(n9910), .Z(n9915) );
  XOR U10100 ( .A(n9914), .B(n9915), .Z(n9917) );
  XNOR U10101 ( .A(n9916), .B(n9917), .Z(n9912) );
  XOR U10102 ( .A(n9913), .B(n9912), .Z(c[250]) );
  AND U10103 ( .A(n9913), .B(n9912), .Z(n9945) );
  NANDN U10104 ( .A(n9915), .B(n9914), .Z(n9919) );
  OR U10105 ( .A(n9917), .B(n9916), .Z(n9918) );
  AND U10106 ( .A(n9919), .B(n9918), .Z(n9948) );
  NANDN U10107 ( .A(n9921), .B(n9920), .Z(n9925) );
  NANDN U10108 ( .A(n9923), .B(n9922), .Z(n9924) );
  AND U10109 ( .A(n9925), .B(n9924), .Z(n9947) );
  NANDN U10110 ( .A(n9927), .B(n9926), .Z(n9931) );
  OR U10111 ( .A(n9929), .B(n9928), .Z(n9930) );
  AND U10112 ( .A(n9931), .B(n9930), .Z(n9954) );
  NANDN U10113 ( .A(n9932), .B(n9987), .Z(n9934) );
  XOR U10114 ( .A(b[15]), .B(a[125]), .Z(n9968) );
  NANDN U10115 ( .A(n10006), .B(n9968), .Z(n9933) );
  AND U10116 ( .A(n9934), .B(n9933), .Z(n9959) );
  XNOR U10117 ( .A(a[127]), .B(b[13]), .Z(n9971) );
  OR U10118 ( .A(n9971), .B(n9935), .Z(n9938) );
  NAND U10119 ( .A(n9972), .B(n9936), .Z(n9937) );
  NAND U10120 ( .A(n9938), .B(n9937), .Z(n9958) );
  XNOR U10121 ( .A(n9959), .B(n9958), .Z(n9961) );
  AND U10122 ( .A(b[15]), .B(a[123]), .Z(n9964) );
  XNOR U10123 ( .A(n9965), .B(n9964), .Z(n9966) );
  XOR U10124 ( .A(n9967), .B(n9966), .Z(n9960) );
  XOR U10125 ( .A(n9961), .B(n9960), .Z(n9953) );
  NANDN U10126 ( .A(n9939), .B(n9967), .Z(n9943) );
  NAND U10127 ( .A(n9941), .B(n9940), .Z(n9942) );
  NAND U10128 ( .A(n9943), .B(n9942), .Z(n9952) );
  XOR U10129 ( .A(n9953), .B(n9952), .Z(n9955) );
  XNOR U10130 ( .A(n9954), .B(n9955), .Z(n9946) );
  XOR U10131 ( .A(n9947), .B(n9946), .Z(n9949) );
  XNOR U10132 ( .A(n9948), .B(n9949), .Z(n9944) );
  XOR U10133 ( .A(n9945), .B(n9944), .Z(c[251]) );
  AND U10134 ( .A(n9945), .B(n9944), .Z(n9977) );
  NANDN U10135 ( .A(n9947), .B(n9946), .Z(n9951) );
  OR U10136 ( .A(n9949), .B(n9948), .Z(n9950) );
  AND U10137 ( .A(n9951), .B(n9950), .Z(n9980) );
  NANDN U10138 ( .A(n9953), .B(n9952), .Z(n9957) );
  NANDN U10139 ( .A(n9955), .B(n9954), .Z(n9956) );
  AND U10140 ( .A(n9957), .B(n9956), .Z(n9979) );
  NANDN U10141 ( .A(n9959), .B(n9958), .Z(n9963) );
  NAND U10142 ( .A(n9961), .B(n9960), .Z(n9962) );
  AND U10143 ( .A(n9963), .B(n9962), .Z(n9994) );
  NAND U10144 ( .A(n9987), .B(n9968), .Z(n9970) );
  XNOR U10145 ( .A(b[15]), .B(a[126]), .Z(n9988) );
  NANDN U10146 ( .A(n9988), .B(n9989), .Z(n9969) );
  NAND U10147 ( .A(n9970), .B(n9969), .Z(n9985) );
  NAND U10148 ( .A(b[15]), .B(a[124]), .Z(n10000) );
  ANDN U10149 ( .B(n9972), .A(n9971), .Z(n9975) );
  NAND U10150 ( .A(b[13]), .B(n9973), .Z(n9974) );
  NANDN U10151 ( .A(n9975), .B(n9974), .Z(n9984) );
  XOR U10152 ( .A(n10000), .B(n9984), .Z(n9986) );
  XOR U10153 ( .A(n9985), .B(n9986), .Z(n9992) );
  XOR U10154 ( .A(n9993), .B(n9992), .Z(n9995) );
  XNOR U10155 ( .A(n9994), .B(n9995), .Z(n9978) );
  XOR U10156 ( .A(n9979), .B(n9978), .Z(n9981) );
  XNOR U10157 ( .A(n9980), .B(n9981), .Z(n9976) );
  XOR U10158 ( .A(n9977), .B(n9976), .Z(c[252]) );
  AND U10159 ( .A(n9977), .B(n9976), .Z(n10010) );
  NANDN U10160 ( .A(n9979), .B(n9978), .Z(n9983) );
  OR U10161 ( .A(n9981), .B(n9980), .Z(n9982) );
  AND U10162 ( .A(n9983), .B(n9982), .Z(n10020) );
  NANDN U10163 ( .A(n9988), .B(n9987), .Z(n9991) );
  XOR U10164 ( .A(a[127]), .B(b[15]), .Z(n10004) );
  NAND U10165 ( .A(n9989), .B(n10004), .Z(n9990) );
  NAND U10166 ( .A(n9991), .B(n9990), .Z(n10011) );
  AND U10167 ( .A(b[15]), .B(a[125]), .Z(n9998) );
  XNOR U10168 ( .A(n9999), .B(n9998), .Z(n10001) );
  XOR U10169 ( .A(n10001), .B(n10000), .Z(n10012) );
  XOR U10170 ( .A(n10011), .B(n10012), .Z(n10014) );
  XOR U10171 ( .A(n10013), .B(n10014), .Z(n10017) );
  NANDN U10172 ( .A(n9993), .B(n9992), .Z(n9997) );
  OR U10173 ( .A(n9995), .B(n9994), .Z(n9996) );
  AND U10174 ( .A(n9997), .B(n9996), .Z(n10018) );
  XOR U10175 ( .A(n10017), .B(n10018), .Z(n10019) );
  XOR U10176 ( .A(n10020), .B(n10019), .Z(n10009) );
  XOR U10177 ( .A(n10010), .B(n10009), .Z(c[253]) );
  NANDN U10178 ( .A(n9999), .B(n9998), .Z(n10003) );
  ANDN U10179 ( .B(n10001), .A(n10000), .Z(n10002) );
  ANDN U10180 ( .B(n10003), .A(n10002), .Z(n10026) );
  AND U10181 ( .A(b[15]), .B(a[126]), .Z(n10024) );
  NANDN U10182 ( .A(n10005), .B(n10004), .Z(n10008) );
  NANDN U10183 ( .A(n10006), .B(b[15]), .Z(n10007) );
  NAND U10184 ( .A(n10008), .B(n10007), .Z(n10025) );
  XNOR U10185 ( .A(n10024), .B(n10025), .Z(n10027) );
  XOR U10186 ( .A(n10026), .B(n10027), .Z(n10030) );
  AND U10187 ( .A(n10010), .B(n10009), .Z(n10029) );
  XNOR U10188 ( .A(n10030), .B(n10029), .Z(n10022) );
  NANDN U10189 ( .A(n10012), .B(n10011), .Z(n10016) );
  NANDN U10190 ( .A(n10014), .B(n10013), .Z(n10015) );
  AND U10191 ( .A(n10016), .B(n10015), .Z(n10031) );
  IV U10192 ( .A(n10032), .Z(n10028) );
  XOR U10193 ( .A(n10031), .B(n10028), .Z(n10021) );
  XNOR U10194 ( .A(n10022), .B(n10021), .Z(c[254]) );
endmodule

